module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251;
  assign n65 = ~x29 & x61;
  assign n66 = ~x28 & x60;
  assign n67 = ~n65 & ~n66;
  assign n68 = ~x30 & x62;
  assign n69 = ~x31 & x63;
  assign n70 = ~n68 & ~n69;
  assign n71 = n67 & n70;
  assign n72 = x59 ^ x27;
  assign n74 = x58 ^ x26;
  assign n73 = ~x27 & x59;
  assign n75 = n74 ^ n73;
  assign n76 = x57 ^ x25;
  assign n77 = ~x57 & ~n76;
  assign n78 = n77 ^ x26;
  assign n79 = n78 ^ x57;
  assign n80 = n75 & ~n79;
  assign n81 = n80 ^ n77;
  assign n82 = n81 ^ x57;
  assign n83 = n82 ^ x59;
  assign n84 = ~n72 & n83;
  assign n85 = n84 ^ x59;
  assign n86 = ~x26 & x58;
  assign n87 = ~n73 & ~n86;
  assign n88 = n77 ^ x25;
  assign n89 = n87 & n88;
  assign n90 = ~x56 & n89;
  assign n91 = x24 & n89;
  assign n92 = ~n90 & ~n91;
  assign n93 = n92 ^ n90;
  assign n94 = n93 ^ n91;
  assign n95 = n85 & n94;
  assign n96 = n71 & ~n95;
  assign n97 = n71 & ~n92;
  assign n98 = ~x22 & x54;
  assign n99 = ~x23 & x55;
  assign n100 = ~n98 & ~n99;
  assign n101 = x53 ^ x21;
  assign n103 = x52 ^ x20;
  assign n102 = ~x20 & x52;
  assign n104 = n103 ^ n102;
  assign n105 = n104 ^ x53;
  assign n106 = ~n101 & n105;
  assign n107 = n106 ^ x21;
  assign n108 = n100 & n107;
  assign n109 = ~x21 & x53;
  assign n110 = ~n102 & ~n109;
  assign n111 = n100 & n110;
  assign n112 = x51 ^ x19;
  assign n113 = x50 ^ x18;
  assign n122 = x51 ^ x50;
  assign n114 = x49 ^ x17;
  assign n116 = x48 ^ x16;
  assign n115 = ~x16 & x48;
  assign n117 = n116 ^ n115;
  assign n118 = n117 ^ x49;
  assign n119 = ~n114 & n118;
  assign n120 = n119 ^ x17;
  assign n121 = n120 ^ x51;
  assign n123 = n122 ^ n121;
  assign n124 = ~n113 & ~n123;
  assign n125 = n124 ^ x51;
  assign n126 = n125 ^ x50;
  assign n127 = ~n112 & ~n126;
  assign n128 = n127 ^ x19;
  assign n129 = n111 & n128;
  assign n130 = ~n108 & ~n129;
  assign n131 = x55 ^ x23;
  assign n132 = x54 ^ x22;
  assign n133 = n132 ^ n98;
  assign n134 = n133 ^ x55;
  assign n135 = ~n131 & n134;
  assign n136 = n135 ^ x23;
  assign n137 = n130 & ~n136;
  assign n138 = n97 & ~n137;
  assign n139 = ~n96 & ~n138;
  assign n140 = ~x17 & x49;
  assign n141 = ~x18 & x50;
  assign n142 = ~x19 & x51;
  assign n143 = ~n141 & ~n142;
  assign n144 = ~x15 & x47;
  assign n145 = ~x14 & x46;
  assign n146 = ~n144 & ~n145;
  assign n147 = x45 ^ x13;
  assign n148 = ~x45 & ~n147;
  assign n149 = n148 ^ x13;
  assign n150 = n146 & n149;
  assign n151 = ~x12 & x44;
  assign n152 = x43 ^ x11;
  assign n153 = x42 ^ x10;
  assign n154 = x9 & ~x41;
  assign n155 = n154 ^ x42;
  assign n156 = ~n153 & ~n155;
  assign n157 = n156 ^ x42;
  assign n158 = n157 ^ x43;
  assign n159 = ~n152 & n158;
  assign n160 = n159 ^ x43;
  assign n161 = ~x11 & x43;
  assign n162 = ~x10 & x42;
  assign n163 = ~n161 & ~n162;
  assign n164 = x41 ^ x9;
  assign n165 = n164 ^ n154;
  assign n168 = ~x40 & ~n165;
  assign n169 = n163 & n168;
  assign n166 = x8 & ~n165;
  assign n167 = n163 & n166;
  assign n170 = n169 ^ n167;
  assign n171 = x39 ^ x7;
  assign n173 = x38 ^ x6;
  assign n172 = ~x6 & x38;
  assign n174 = n173 ^ n172;
  assign n175 = n174 ^ x39;
  assign n176 = ~n171 & n175;
  assign n177 = n176 ^ x7;
  assign n178 = ~x7 & x39;
  assign n179 = ~n172 & ~n178;
  assign n180 = x37 ^ x5;
  assign n181 = x36 ^ x4;
  assign n182 = x35 ^ x3;
  assign n183 = x34 ^ x2;
  assign n185 = x33 ^ x1;
  assign n184 = ~x2 & x34;
  assign n186 = n185 ^ n184;
  assign n187 = x32 ^ x0;
  assign n188 = x32 & ~n187;
  assign n189 = n188 ^ x1;
  assign n190 = n189 ^ x32;
  assign n191 = n186 & ~n190;
  assign n192 = n191 ^ n188;
  assign n193 = n192 ^ x32;
  assign n194 = n193 ^ x34;
  assign n195 = ~n183 & n194;
  assign n196 = n195 ^ x34;
  assign n197 = n196 ^ x35;
  assign n198 = ~n182 & n197;
  assign n199 = n198 ^ x35;
  assign n200 = n199 ^ x36;
  assign n201 = ~n181 & n200;
  assign n202 = n201 ^ x36;
  assign n203 = n202 ^ x37;
  assign n204 = ~n180 & n203;
  assign n205 = n204 ^ x37;
  assign n206 = n179 & ~n205;
  assign n207 = ~n177 & ~n206;
  assign n208 = n207 ^ n167;
  assign n209 = n170 & ~n208;
  assign n210 = n209 ^ n167;
  assign n211 = n160 & ~n210;
  assign n212 = ~n151 & ~n211;
  assign n213 = n150 & n212;
  assign n214 = x12 & n150;
  assign n215 = ~x44 & n214;
  assign n216 = x47 ^ x15;
  assign n217 = x46 ^ x14;
  assign n218 = n217 ^ n144;
  assign n219 = n148 ^ x14;
  assign n220 = n219 ^ x45;
  assign n221 = n218 & ~n220;
  assign n222 = n221 ^ n148;
  assign n223 = n222 ^ x45;
  assign n224 = n223 ^ x47;
  assign n225 = ~n216 & n224;
  assign n226 = n225 ^ x47;
  assign n227 = ~n215 & n226;
  assign n228 = ~n213 & n227;
  assign n229 = ~n115 & ~n228;
  assign n230 = n143 & n229;
  assign n231 = ~n140 & n230;
  assign n232 = n111 & n231;
  assign n233 = n97 & n232;
  assign n234 = x63 ^ x31;
  assign n235 = x62 ^ x30;
  assign n243 = x63 ^ x62;
  assign n236 = x61 ^ x29;
  assign n237 = x60 ^ x28;
  assign n238 = n237 ^ n66;
  assign n239 = n238 ^ x61;
  assign n240 = ~n236 & n239;
  assign n241 = n240 ^ x29;
  assign n242 = n241 ^ x63;
  assign n244 = n243 ^ n242;
  assign n245 = ~n235 & ~n244;
  assign n246 = n245 ^ x63;
  assign n247 = n246 ^ x62;
  assign n248 = ~n234 & ~n247;
  assign n249 = n248 ^ x31;
  assign n250 = ~n233 & ~n249;
  assign n251 = n139 & n250;
  assign y0 = n251;
endmodule
