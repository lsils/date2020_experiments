module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, y0, y1, y2, y3, y4, y5, y6);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10;
  output y0, y1, y2, y3, y4, y5, y6;
  wire n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184;
  assign n40 = x7 ^ x6;
  assign n34 = x6 & x7;
  assign n36 = ~x8 & ~n34;
  assign n35 = n34 ^ x8;
  assign n37 = n36 ^ n35;
  assign n38 = ~x9 & ~n37;
  assign n39 = n38 ^ n37;
  assign n41 = n40 ^ n39;
  assign n27 = x5 ^ x4;
  assign n20 = x3 ^ x2;
  assign n15 = x1 & x4;
  assign n16 = n15 ^ x0;
  assign n14 = x2 ^ x1;
  assign n17 = n16 ^ n14;
  assign n18 = x5 & n17;
  assign n19 = n18 ^ n16;
  assign n21 = n20 ^ n19;
  assign n22 = ~x6 & n21;
  assign n23 = n22 ^ n20;
  assign n13 = x4 ^ x3;
  assign n24 = n23 ^ n13;
  assign n25 = x7 & n24;
  assign n26 = n25 ^ n23;
  assign n28 = n27 ^ n26;
  assign n29 = ~x8 & n28;
  assign n30 = n29 ^ n27;
  assign n12 = x6 ^ x5;
  assign n31 = n30 ^ n12;
  assign n32 = x9 & n31;
  assign n33 = n32 ^ n30;
  assign n42 = n41 ^ n33;
  assign n43 = x10 & ~n42;
  assign n44 = n43 ^ n33;
  assign n45 = ~x7 & ~x8;
  assign n53 = x1 & x2;
  assign n54 = n53 ^ x3;
  assign n50 = ~x0 & n15;
  assign n51 = n50 ^ x1;
  assign n49 = x2 & x4;
  assign n52 = n51 ^ n49;
  assign n55 = n54 ^ n52;
  assign n56 = x5 & n55;
  assign n57 = n56 ^ n52;
  assign n46 = ~x2 & ~x3;
  assign n47 = n46 ^ n20;
  assign n48 = n47 ^ x4;
  assign n58 = n57 ^ n48;
  assign n59 = n58 ^ n57;
  assign n60 = ~x9 & n59;
  assign n61 = n60 ^ n57;
  assign n62 = x6 & ~n61;
  assign n63 = n62 ^ n57;
  assign n64 = n45 & ~n63;
  assign n72 = x4 & x5;
  assign n73 = n72 ^ x6;
  assign n68 = x3 & x4;
  assign n69 = n68 ^ x5;
  assign n70 = n69 ^ x7;
  assign n71 = x7 & ~n70;
  assign n74 = n73 ^ n71;
  assign n75 = n74 ^ x7;
  assign n76 = x9 ^ x8;
  assign n77 = ~n75 & n76;
  assign n78 = n77 ^ n71;
  assign n79 = n78 ^ x7;
  assign n65 = ~x5 & ~x6;
  assign n66 = n65 ^ n12;
  assign n67 = n66 ^ x7;
  assign n80 = n79 ^ n67;
  assign n81 = ~x9 & n80;
  assign n82 = n81 ^ n67;
  assign n83 = ~x10 & ~n82;
  assign n84 = ~n64 & n83;
  assign n85 = x10 & ~n36;
  assign n86 = ~n38 & n85;
  assign n87 = ~n84 & ~n86;
  assign n88 = x5 & n34;
  assign n89 = n88 ^ x8;
  assign n90 = n89 ^ n37;
  assign n91 = ~x10 & n90;
  assign n92 = n91 ^ n37;
  assign n93 = n92 ^ x9;
  assign n94 = n93 ^ x10;
  assign n95 = n94 ^ n92;
  assign n96 = x6 & n72;
  assign n97 = ~n47 & n96;
  assign n98 = ~x7 & ~n97;
  assign n101 = x6 ^ x2;
  assign n102 = n101 ^ x4;
  assign n103 = ~n101 & ~n102;
  assign n99 = x5 ^ x2;
  assign n100 = n99 ^ x6;
  assign n104 = n103 ^ n100;
  assign n105 = n104 ^ n101;
  assign n106 = x6 ^ x3;
  assign n107 = n103 ^ n101;
  assign n108 = ~n106 & ~n107;
  assign n109 = n108 ^ x6;
  assign n110 = ~n105 & ~n109;
  assign n111 = n110 ^ x6;
  assign n112 = n111 ^ x5;
  assign n113 = n112 ^ x6;
  assign n114 = n98 & n113;
  assign n117 = ~x3 & x5;
  assign n118 = n117 ^ x3;
  assign n119 = n118 ^ n12;
  assign n120 = x4 & ~n119;
  assign n121 = n120 ^ n12;
  assign n115 = x3 & ~x6;
  assign n116 = n49 & n115;
  assign n122 = n121 ^ n116;
  assign n123 = x3 ^ x0;
  assign n124 = x5 & n123;
  assign n125 = n124 ^ x0;
  assign n126 = x1 & n125;
  assign n127 = n122 & n126;
  assign n128 = n127 ^ n121;
  assign n129 = n114 & ~n128;
  assign n130 = ~x3 & n34;
  assign n131 = ~n129 & ~n130;
  assign n132 = ~x8 & ~n131;
  assign n133 = x7 & ~n96;
  assign n134 = ~n36 & n133;
  assign n135 = n72 ^ n40;
  assign n136 = x8 ^ x3;
  assign n137 = x7 & n136;
  assign n138 = n137 ^ x8;
  assign n139 = n138 ^ n40;
  assign n140 = n135 & n139;
  assign n141 = n140 ^ n137;
  assign n142 = n141 ^ x8;
  assign n143 = n142 ^ n72;
  assign n144 = n40 & n143;
  assign n145 = n144 ^ n40;
  assign n146 = ~n134 & ~n145;
  assign n147 = ~n132 & n146;
  assign n148 = n147 ^ n92;
  assign n149 = n148 ^ n92;
  assign n150 = ~x10 & ~n149;
  assign n151 = n150 ^ n92;
  assign n152 = ~n95 & ~n151;
  assign n153 = n152 ^ n93;
  assign n154 = ~x9 & ~x10;
  assign n155 = ~x3 & n154;
  assign n159 = ~x2 & ~n37;
  assign n160 = n72 & n159;
  assign n156 = x4 & n65;
  assign n157 = n156 ^ n65;
  assign n158 = n45 & n157;
  assign n161 = n160 ^ n158;
  assign n162 = n155 & n161;
  assign n164 = n156 ^ x6;
  assign n163 = n116 & n126;
  assign n165 = n164 ^ n163;
  assign n166 = n98 & n165;
  assign n167 = ~x8 & ~n166;
  assign n168 = ~n46 & n72;
  assign n169 = n34 & n168;
  assign n170 = ~x9 & ~n169;
  assign n171 = ~n167 & n170;
  assign n172 = ~x9 & ~n68;
  assign n173 = ~n76 & n172;
  assign n174 = n173 ^ n76;
  assign n175 = n88 & ~n174;
  assign n176 = ~x10 & ~n175;
  assign n177 = ~n171 & n176;
  assign n178 = n65 & ~n163;
  assign n179 = n45 & ~n97;
  assign n180 = ~n178 & n179;
  assign n181 = x8 & n169;
  assign n182 = n154 & ~n181;
  assign n183 = ~n180 & n182;
  assign n184 = n154 & n179;
  assign y0 = n44;
  assign y1 = ~n87;
  assign y2 = ~n153;
  assign y3 = ~n162;
  assign y4 = ~n177;
  assign y5 = ~n183;
  assign y6 = ~n184;
endmodule
