module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 ;
  wire n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 ;
  assign n597 = x527 ^ x495 ;
  assign n596 = x526 ^ x494 ;
  assign n598 = n597 ^ n596 ;
  assign n595 = x528 ^ x496 ;
  assign n599 = n598 ^ n595 ;
  assign n594 = x522 ^ x490 ;
  assign n600 = n599 ^ n594 ;
  assign n591 = x524 ^ x492 ;
  assign n590 = x523 ^ x491 ;
  assign n592 = n591 ^ n590 ;
  assign n589 = x525 ^ x493 ;
  assign n593 = n592 ^ n589 ;
  assign n656 = n599 ^ n593 ;
  assign n657 = ~n600 & n656 ;
  assign n658 = n657 ^ n593 ;
  assign n653 = n596 ^ n595 ;
  assign n654 = n598 & ~n653 ;
  assign n655 = n654 ^ n597 ;
  assign n659 = n658 ^ n655 ;
  assign n650 = n590 ^ n589 ;
  assign n651 = n592 & ~n650 ;
  assign n652 = n651 ^ n591 ;
  assign n660 = n659 ^ n652 ;
  assign n584 = x520 ^ x488 ;
  assign n583 = x519 ^ x487 ;
  assign n585 = n584 ^ n583 ;
  assign n582 = x521 ^ x489 ;
  assign n645 = n583 ^ n582 ;
  assign n646 = n585 & ~n645 ;
  assign n647 = n646 ^ n584 ;
  assign n586 = n585 ^ n582 ;
  assign n581 = x515 ^ x483 ;
  assign n587 = n586 ^ n581 ;
  assign n578 = x517 ^ x485 ;
  assign n577 = x516 ^ x484 ;
  assign n579 = n578 ^ n577 ;
  assign n576 = x518 ^ x486 ;
  assign n580 = n579 ^ n576 ;
  assign n642 = n586 ^ n580 ;
  assign n643 = ~n587 & n642 ;
  assign n644 = n643 ^ n580 ;
  assign n648 = n647 ^ n644 ;
  assign n639 = n577 ^ n576 ;
  assign n640 = n579 & ~n639 ;
  assign n641 = n640 ^ n578 ;
  assign n649 = n648 ^ n641 ;
  assign n661 = n660 ^ n649 ;
  assign n602 = x514 ^ x482 ;
  assign n601 = n600 ^ n593 ;
  assign n603 = n602 ^ n601 ;
  assign n588 = n587 ^ n580 ;
  assign n636 = n601 ^ n588 ;
  assign n637 = n603 & ~n636 ;
  assign n638 = n637 ^ n602 ;
  assign n684 = n660 ^ n638 ;
  assign n685 = ~n661 & n684 ;
  assign n686 = n685 ^ n638 ;
  assign n681 = n655 ^ n652 ;
  assign n682 = n659 & ~n681 ;
  assign n683 = n682 ^ n658 ;
  assign n687 = n686 ^ n683 ;
  assign n678 = n644 ^ n641 ;
  assign n679 = n648 & n678 ;
  assign n680 = n679 ^ n644 ;
  assign n688 = n687 ^ n680 ;
  assign n565 = x541 ^ x509 ;
  assign n564 = x542 ^ x510 ;
  assign n566 = n565 ^ n564 ;
  assign n563 = x543 ^ x511 ;
  assign n628 = n564 ^ n563 ;
  assign n629 = n566 & ~n628 ;
  assign n630 = n629 ^ n565 ;
  assign n568 = x537 ^ x505 ;
  assign n567 = n566 ^ n563 ;
  assign n569 = n568 ^ n567 ;
  assign n560 = x539 ^ x507 ;
  assign n559 = x538 ^ x506 ;
  assign n561 = n560 ^ n559 ;
  assign n558 = x540 ^ x508 ;
  assign n562 = n561 ^ n558 ;
  assign n625 = n568 ^ n562 ;
  assign n626 = ~n569 & n625 ;
  assign n627 = n626 ^ n562 ;
  assign n631 = n630 ^ n627 ;
  assign n622 = n559 ^ n558 ;
  assign n623 = n561 & ~n622 ;
  assign n624 = n623 ^ n560 ;
  assign n632 = n631 ^ n624 ;
  assign n571 = x529 ^ x497 ;
  assign n570 = n569 ^ n562 ;
  assign n572 = n571 ^ n570 ;
  assign n555 = x530 ^ x498 ;
  assign n553 = x536 ^ x504 ;
  assign n551 = x534 ^ x502 ;
  assign n550 = x535 ^ x503 ;
  assign n552 = n551 ^ n550 ;
  assign n554 = n553 ^ n552 ;
  assign n556 = n555 ^ n554 ;
  assign n547 = x532 ^ x500 ;
  assign n546 = x531 ^ x499 ;
  assign n548 = n547 ^ n546 ;
  assign n545 = x533 ^ x501 ;
  assign n549 = n548 ^ n545 ;
  assign n557 = n556 ^ n549 ;
  assign n619 = n571 ^ n557 ;
  assign n620 = ~n572 & n619 ;
  assign n621 = n620 ^ n557 ;
  assign n633 = n632 ^ n621 ;
  assign n614 = n553 ^ n550 ;
  assign n615 = n552 & ~n614 ;
  assign n616 = n615 ^ n551 ;
  assign n611 = n554 ^ n549 ;
  assign n612 = n556 & ~n611 ;
  assign n613 = n612 ^ n555 ;
  assign n617 = n616 ^ n613 ;
  assign n608 = n546 ^ n545 ;
  assign n609 = n548 & ~n608 ;
  assign n610 = n609 ^ n547 ;
  assign n618 = n617 ^ n610 ;
  assign n672 = n632 ^ n618 ;
  assign n673 = ~n633 & n672 ;
  assign n674 = n673 ^ n618 ;
  assign n669 = n630 ^ n624 ;
  assign n670 = n631 & n669 ;
  assign n671 = n670 ^ n630 ;
  assign n675 = n674 ^ n671 ;
  assign n666 = n613 ^ n610 ;
  assign n667 = n617 & n666 ;
  assign n668 = n667 ^ n613 ;
  assign n676 = n675 ^ n668 ;
  assign n634 = n633 ^ n618 ;
  assign n574 = x513 ^ x481 ;
  assign n573 = n572 ^ n557 ;
  assign n575 = n574 ^ n573 ;
  assign n604 = n603 ^ n588 ;
  assign n605 = n604 ^ n573 ;
  assign n606 = n575 & ~n605 ;
  assign n607 = n606 ^ n574 ;
  assign n635 = n634 ^ n607 ;
  assign n662 = n661 ^ n638 ;
  assign n663 = n662 ^ n634 ;
  assign n664 = n635 & ~n663 ;
  assign n665 = n664 ^ n607 ;
  assign n677 = n676 ^ n665 ;
  assign n689 = n688 ^ n677 ;
  assign n690 = n662 ^ n635 ;
  assign n691 = x512 ^ x480 ;
  assign n692 = n604 ^ n575 ;
  assign n693 = n691 & n692 ;
  assign n694 = n690 & n693 ;
  assign n695 = n689 & n694 ;
  assign n702 = n688 ^ n676 ;
  assign n703 = ~n677 & n702 ;
  assign n704 = n703 ^ n688 ;
  assign n699 = n671 ^ n668 ;
  assign n700 = n675 & ~n699 ;
  assign n701 = n700 ^ n674 ;
  assign n705 = n704 ^ n701 ;
  assign n696 = n683 ^ n680 ;
  assign n697 = n687 & ~n696 ;
  assign n698 = n697 ^ n686 ;
  assign n706 = n705 ^ n698 ;
  assign n707 = n695 & n706 ;
  assign n708 = n701 ^ n698 ;
  assign n709 = n705 & ~n708 ;
  assign n710 = n709 ^ n704 ;
  assign n711 = n707 & n710 ;
  assign n747 = x534 ^ x470 ;
  assign n746 = x535 ^ x471 ;
  assign n748 = n747 ^ n746 ;
  assign n745 = x536 ^ x472 ;
  assign n764 = n746 ^ n745 ;
  assign n765 = n748 & ~n764 ;
  assign n766 = n765 ^ n747 ;
  assign n750 = x530 ^ x466 ;
  assign n749 = n748 ^ n745 ;
  assign n751 = n750 ^ n749 ;
  assign n742 = x532 ^ x468 ;
  assign n741 = x531 ^ x467 ;
  assign n743 = n742 ^ n741 ;
  assign n740 = x533 ^ x469 ;
  assign n744 = n743 ^ n740 ;
  assign n761 = n749 ^ n744 ;
  assign n762 = n751 & ~n761 ;
  assign n763 = n762 ^ n750 ;
  assign n767 = n766 ^ n763 ;
  assign n758 = n741 ^ n740 ;
  assign n759 = n743 & ~n758 ;
  assign n760 = n759 ^ n742 ;
  assign n773 = n763 ^ n760 ;
  assign n774 = n767 & n773 ;
  assign n775 = n774 ^ n763 ;
  assign n721 = x539 ^ x475 ;
  assign n720 = x538 ^ x474 ;
  assign n722 = n721 ^ n720 ;
  assign n719 = x540 ^ x476 ;
  assign n731 = n720 ^ n719 ;
  assign n732 = n722 & ~n731 ;
  assign n733 = n732 ^ n721 ;
  assign n714 = x541 ^ x477 ;
  assign n713 = x542 ^ x478 ;
  assign n715 = n714 ^ n713 ;
  assign n712 = x543 ^ x479 ;
  assign n727 = n713 ^ n712 ;
  assign n728 = n715 & ~n727 ;
  assign n729 = n728 ^ n714 ;
  assign n717 = x537 ^ x473 ;
  assign n716 = n715 ^ n712 ;
  assign n718 = n717 ^ n716 ;
  assign n723 = n722 ^ n719 ;
  assign n724 = n723 ^ n717 ;
  assign n725 = ~n718 & n724 ;
  assign n726 = n725 ^ n723 ;
  assign n730 = n729 ^ n726 ;
  assign n756 = n733 ^ n730 ;
  assign n738 = x529 ^ x465 ;
  assign n737 = n723 ^ n718 ;
  assign n739 = n738 ^ n737 ;
  assign n752 = n751 ^ n744 ;
  assign n753 = n752 ^ n738 ;
  assign n754 = ~n739 & n753 ;
  assign n755 = n754 ^ n752 ;
  assign n757 = n756 ^ n755 ;
  assign n768 = n767 ^ n760 ;
  assign n769 = n768 ^ n756 ;
  assign n770 = ~n757 & n769 ;
  assign n771 = n770 ^ n768 ;
  assign n734 = n733 ^ n729 ;
  assign n735 = n730 & n734 ;
  assign n736 = n735 ^ n729 ;
  assign n772 = n771 ^ n736 ;
  assign n846 = n775 ^ n772 ;
  assign n814 = n768 ^ n757 ;
  assign n780 = x513 ^ x449 ;
  assign n779 = n752 ^ n739 ;
  assign n781 = n780 ^ n779 ;
  assign n806 = x517 ^ x453 ;
  assign n805 = x516 ^ x452 ;
  assign n807 = n806 ^ n805 ;
  assign n804 = x518 ^ x454 ;
  assign n808 = n807 ^ n804 ;
  assign n800 = x520 ^ x456 ;
  assign n799 = x519 ^ x455 ;
  assign n801 = n800 ^ n799 ;
  assign n798 = x521 ^ x457 ;
  assign n802 = n801 ^ n798 ;
  assign n797 = x515 ^ x451 ;
  assign n803 = n802 ^ n797 ;
  assign n809 = n808 ^ n803 ;
  assign n795 = x514 ^ x450 ;
  assign n791 = x524 ^ x460 ;
  assign n790 = x523 ^ x459 ;
  assign n792 = n791 ^ n790 ;
  assign n789 = x525 ^ x461 ;
  assign n793 = n792 ^ n789 ;
  assign n786 = x528 ^ x464 ;
  assign n784 = x527 ^ x463 ;
  assign n783 = x526 ^ x462 ;
  assign n785 = n784 ^ n783 ;
  assign n787 = n786 ^ n785 ;
  assign n782 = x522 ^ x458 ;
  assign n788 = n787 ^ n782 ;
  assign n794 = n793 ^ n788 ;
  assign n796 = n795 ^ n794 ;
  assign n810 = n809 ^ n796 ;
  assign n811 = n810 ^ n779 ;
  assign n812 = n781 & ~n811 ;
  assign n813 = n812 ^ n780 ;
  assign n815 = n814 ^ n813 ;
  assign n839 = n809 ^ n794 ;
  assign n840 = n796 & ~n839 ;
  assign n841 = n840 ^ n795 ;
  assign n834 = n790 ^ n789 ;
  assign n835 = n792 & ~n834 ;
  assign n836 = n835 ^ n791 ;
  assign n830 = n793 ^ n787 ;
  assign n831 = ~n788 & n830 ;
  assign n832 = n831 ^ n793 ;
  assign n827 = n786 ^ n783 ;
  assign n828 = n785 & ~n827 ;
  assign n829 = n828 ^ n784 ;
  assign n833 = n832 ^ n829 ;
  assign n837 = n836 ^ n833 ;
  assign n823 = n805 ^ n804 ;
  assign n824 = n807 & ~n823 ;
  assign n825 = n824 ^ n806 ;
  assign n819 = n799 ^ n798 ;
  assign n820 = n801 & ~n819 ;
  assign n821 = n820 ^ n800 ;
  assign n816 = n808 ^ n802 ;
  assign n817 = ~n803 & n816 ;
  assign n818 = n817 ^ n808 ;
  assign n822 = n821 ^ n818 ;
  assign n826 = n825 ^ n822 ;
  assign n838 = n837 ^ n826 ;
  assign n842 = n841 ^ n838 ;
  assign n843 = n842 ^ n814 ;
  assign n844 = n815 & ~n843 ;
  assign n845 = n844 ^ n813 ;
  assign n847 = n846 ^ n845 ;
  assign n854 = n841 ^ n837 ;
  assign n855 = ~n838 & n854 ;
  assign n856 = n855 ^ n841 ;
  assign n851 = n836 ^ n829 ;
  assign n852 = n833 & ~n851 ;
  assign n853 = n852 ^ n832 ;
  assign n857 = n856 ^ n853 ;
  assign n848 = n825 ^ n818 ;
  assign n849 = n822 & n848 ;
  assign n850 = n849 ^ n818 ;
  assign n858 = n857 ^ n850 ;
  assign n859 = n858 ^ n846 ;
  assign n860 = ~n847 & n859 ;
  assign n861 = n860 ^ n858 ;
  assign n776 = n775 ^ n736 ;
  assign n777 = n772 & ~n776 ;
  assign n778 = n777 ^ n771 ;
  assign n862 = n861 ^ n778 ;
  assign n863 = n853 ^ n850 ;
  assign n864 = n857 & ~n863 ;
  assign n865 = n864 ^ n856 ;
  assign n866 = n865 ^ n778 ;
  assign n867 = n862 & ~n866 ;
  assign n868 = n867 ^ n861 ;
  assign n869 = n858 ^ n847 ;
  assign n870 = n842 ^ n815 ;
  assign n871 = x512 ^ x448 ;
  assign n872 = n810 ^ n781 ;
  assign n873 = n871 & n872 ;
  assign n874 = n870 & n873 ;
  assign n875 = n869 & n874 ;
  assign n876 = n865 ^ n862 ;
  assign n877 = n875 & n876 ;
  assign n879 = ~n868 & ~n877 ;
  assign n878 = n877 ^ n868 ;
  assign n880 = n879 ^ n878 ;
  assign n881 = ~n711 & ~n880 ;
  assign n882 = n881 ^ n711 ;
  assign n973 = x543 ^ x447 ;
  assign n971 = x542 ^ x446 ;
  assign n970 = x541 ^ x445 ;
  assign n972 = n971 ^ n970 ;
  assign n974 = n973 ^ n972 ;
  assign n969 = x537 ^ x441 ;
  assign n975 = n974 ^ n969 ;
  assign n967 = x540 ^ x444 ;
  assign n965 = x539 ^ x443 ;
  assign n964 = x538 ^ x442 ;
  assign n966 = n965 ^ n964 ;
  assign n968 = n967 ^ n966 ;
  assign n1005 = n969 ^ n968 ;
  assign n1006 = n975 & ~n1005 ;
  assign n1007 = n1006 ^ n974 ;
  assign n1002 = n973 ^ n971 ;
  assign n1003 = ~n972 & n1002 ;
  assign n1004 = n1003 ^ n973 ;
  assign n1008 = n1007 ^ n1004 ;
  assign n999 = n967 ^ n965 ;
  assign n1000 = ~n966 & n999 ;
  assign n1001 = n1000 ^ n967 ;
  assign n1009 = n1008 ^ n1001 ;
  assign n977 = x529 ^ x433 ;
  assign n976 = n975 ^ n968 ;
  assign n978 = n977 ^ n976 ;
  assign n959 = x535 ^ x439 ;
  assign n958 = x534 ^ x438 ;
  assign n960 = n959 ^ n958 ;
  assign n957 = x536 ^ x440 ;
  assign n961 = n960 ^ n957 ;
  assign n956 = x530 ^ x434 ;
  assign n962 = n961 ^ n956 ;
  assign n953 = x532 ^ x436 ;
  assign n952 = x531 ^ x435 ;
  assign n954 = n953 ^ n952 ;
  assign n951 = x533 ^ x437 ;
  assign n955 = n954 ^ n951 ;
  assign n963 = n962 ^ n955 ;
  assign n996 = n976 ^ n963 ;
  assign n997 = n978 & ~n996 ;
  assign n998 = n997 ^ n977 ;
  assign n1010 = n1009 ^ n998 ;
  assign n991 = n956 ^ n955 ;
  assign n992 = n962 & ~n991 ;
  assign n993 = n992 ^ n961 ;
  assign n988 = n958 ^ n957 ;
  assign n989 = n960 & ~n988 ;
  assign n990 = n989 ^ n959 ;
  assign n994 = n993 ^ n990 ;
  assign n985 = n952 ^ n951 ;
  assign n986 = n954 & ~n985 ;
  assign n987 = n986 ^ n953 ;
  assign n995 = n994 ^ n987 ;
  assign n1023 = n998 ^ n995 ;
  assign n1024 = n1010 & ~n1023 ;
  assign n1025 = n1024 ^ n1009 ;
  assign n1020 = n1004 ^ n1001 ;
  assign n1021 = n1008 & ~n1020 ;
  assign n1022 = n1021 ^ n1007 ;
  assign n1026 = n1025 ^ n1022 ;
  assign n1017 = n990 ^ n987 ;
  assign n1018 = n994 & ~n1017 ;
  assign n1019 = n1018 ^ n993 ;
  assign n1033 = n1022 ^ n1019 ;
  assign n1034 = n1026 & ~n1033 ;
  assign n1035 = n1034 ^ n1025 ;
  assign n1027 = n1026 ^ n1019 ;
  assign n1011 = n1010 ^ n995 ;
  assign n979 = n978 ^ n963 ;
  assign n950 = x513 ^ x417 ;
  assign n980 = n979 ^ n950 ;
  assign n907 = x517 ^ x421 ;
  assign n906 = x516 ^ x420 ;
  assign n908 = n907 ^ n906 ;
  assign n905 = x518 ^ x422 ;
  assign n909 = n908 ^ n905 ;
  assign n901 = x520 ^ x424 ;
  assign n900 = x519 ^ x423 ;
  assign n902 = n901 ^ n900 ;
  assign n899 = x521 ^ x425 ;
  assign n903 = n902 ^ n899 ;
  assign n898 = x515 ^ x419 ;
  assign n904 = n903 ^ n898 ;
  assign n910 = n909 ^ n904 ;
  assign n893 = x524 ^ x428 ;
  assign n892 = x523 ^ x427 ;
  assign n894 = n893 ^ n892 ;
  assign n891 = x525 ^ x429 ;
  assign n895 = n894 ^ n891 ;
  assign n887 = x527 ^ x431 ;
  assign n886 = x526 ^ x430 ;
  assign n888 = n887 ^ n886 ;
  assign n885 = x528 ^ x432 ;
  assign n889 = n888 ^ n885 ;
  assign n884 = x522 ^ x426 ;
  assign n890 = n889 ^ n884 ;
  assign n896 = n895 ^ n890 ;
  assign n883 = x514 ^ x418 ;
  assign n897 = n896 ^ n883 ;
  assign n981 = n910 ^ n897 ;
  assign n982 = n981 ^ n950 ;
  assign n983 = n980 & ~n982 ;
  assign n984 = n983 ^ n979 ;
  assign n1012 = n1011 ^ n984 ;
  assign n932 = n900 ^ n899 ;
  assign n933 = n902 & ~n932 ;
  assign n934 = n933 ^ n901 ;
  assign n929 = n909 ^ n903 ;
  assign n930 = ~n904 & n929 ;
  assign n931 = n930 ^ n909 ;
  assign n935 = n934 ^ n931 ;
  assign n926 = n906 ^ n905 ;
  assign n927 = n908 & ~n926 ;
  assign n928 = n927 ^ n907 ;
  assign n936 = n935 ^ n928 ;
  assign n920 = n895 ^ n889 ;
  assign n921 = ~n890 & n920 ;
  assign n922 = n921 ^ n895 ;
  assign n917 = n886 ^ n885 ;
  assign n918 = n888 & ~n917 ;
  assign n919 = n918 ^ n887 ;
  assign n923 = n922 ^ n919 ;
  assign n914 = n892 ^ n891 ;
  assign n915 = n894 & ~n914 ;
  assign n916 = n915 ^ n893 ;
  assign n924 = n923 ^ n916 ;
  assign n911 = n910 ^ n883 ;
  assign n912 = n897 & ~n911 ;
  assign n913 = n912 ^ n896 ;
  assign n925 = n924 ^ n913 ;
  assign n1013 = n936 ^ n925 ;
  assign n1014 = n1013 ^ n1011 ;
  assign n1015 = n1012 & ~n1014 ;
  assign n1016 = n1015 ^ n984 ;
  assign n1028 = n1027 ^ n1016 ;
  assign n944 = n931 ^ n928 ;
  assign n945 = n935 & ~n944 ;
  assign n946 = n945 ^ n934 ;
  assign n940 = n919 ^ n916 ;
  assign n941 = n923 & ~n940 ;
  assign n942 = n941 ^ n922 ;
  assign n937 = n936 ^ n913 ;
  assign n938 = n925 & ~n937 ;
  assign n939 = n938 ^ n924 ;
  assign n943 = n942 ^ n939 ;
  assign n1029 = n946 ^ n943 ;
  assign n1030 = n1029 ^ n1016 ;
  assign n1031 = n1028 & ~n1030 ;
  assign n1032 = n1031 ^ n1027 ;
  assign n1036 = n1035 ^ n1032 ;
  assign n947 = n946 ^ n942 ;
  assign n948 = ~n943 & n947 ;
  assign n949 = n948 ^ n946 ;
  assign n1037 = n1036 ^ n949 ;
  assign n1038 = n1013 ^ n1012 ;
  assign n1039 = n981 ^ n980 ;
  assign n1040 = x512 ^ x416 ;
  assign n1041 = n1039 & n1040 ;
  assign n1042 = n1038 & n1041 ;
  assign n1043 = n1029 ^ n1028 ;
  assign n1044 = n1042 & n1043 ;
  assign n1045 = n1037 & n1044 ;
  assign n1046 = n1032 ^ n949 ;
  assign n1047 = n1036 & ~n1046 ;
  assign n1048 = n1047 ^ n1035 ;
  assign n1049 = n1045 & n1048 ;
  assign n1050 = n882 & n1049 ;
  assign n1051 = n882 ^ n880 ;
  assign n1052 = n1051 ^ n711 ;
  assign n1053 = n1050 & n1052 ;
  assign n1054 = n1053 ^ n1050 ;
  assign n1055 = n1054 ^ n1052 ;
  assign n1056 = n1055 ^ n1050 ;
  assign n1057 = n1049 ^ n882 ;
  assign n1058 = n1057 ^ n1050 ;
  assign n1149 = x543 ^ x415 ;
  assign n1147 = x542 ^ x414 ;
  assign n1146 = x541 ^ x413 ;
  assign n1148 = n1147 ^ n1146 ;
  assign n1150 = n1149 ^ n1148 ;
  assign n1145 = x537 ^ x409 ;
  assign n1151 = n1150 ^ n1145 ;
  assign n1143 = x540 ^ x412 ;
  assign n1141 = x539 ^ x411 ;
  assign n1140 = x538 ^ x410 ;
  assign n1142 = n1141 ^ n1140 ;
  assign n1144 = n1143 ^ n1142 ;
  assign n1181 = n1145 ^ n1144 ;
  assign n1182 = n1151 & ~n1181 ;
  assign n1183 = n1182 ^ n1150 ;
  assign n1178 = n1149 ^ n1147 ;
  assign n1179 = ~n1148 & n1178 ;
  assign n1180 = n1179 ^ n1149 ;
  assign n1184 = n1183 ^ n1180 ;
  assign n1175 = n1143 ^ n1141 ;
  assign n1176 = ~n1142 & n1175 ;
  assign n1177 = n1176 ^ n1143 ;
  assign n1185 = n1184 ^ n1177 ;
  assign n1153 = x529 ^ x401 ;
  assign n1152 = n1151 ^ n1144 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n1135 = x535 ^ x407 ;
  assign n1134 = x534 ^ x406 ;
  assign n1136 = n1135 ^ n1134 ;
  assign n1133 = x536 ^ x408 ;
  assign n1137 = n1136 ^ n1133 ;
  assign n1132 = x530 ^ x402 ;
  assign n1138 = n1137 ^ n1132 ;
  assign n1129 = x532 ^ x404 ;
  assign n1128 = x531 ^ x403 ;
  assign n1130 = n1129 ^ n1128 ;
  assign n1127 = x533 ^ x405 ;
  assign n1131 = n1130 ^ n1127 ;
  assign n1139 = n1138 ^ n1131 ;
  assign n1172 = n1152 ^ n1139 ;
  assign n1173 = n1154 & ~n1172 ;
  assign n1174 = n1173 ^ n1153 ;
  assign n1186 = n1185 ^ n1174 ;
  assign n1167 = n1132 ^ n1131 ;
  assign n1168 = n1138 & ~n1167 ;
  assign n1169 = n1168 ^ n1137 ;
  assign n1164 = n1134 ^ n1133 ;
  assign n1165 = n1136 & ~n1164 ;
  assign n1166 = n1165 ^ n1135 ;
  assign n1170 = n1169 ^ n1166 ;
  assign n1161 = n1128 ^ n1127 ;
  assign n1162 = n1130 & ~n1161 ;
  assign n1163 = n1162 ^ n1129 ;
  assign n1171 = n1170 ^ n1163 ;
  assign n1199 = n1174 ^ n1171 ;
  assign n1200 = n1186 & ~n1199 ;
  assign n1201 = n1200 ^ n1185 ;
  assign n1196 = n1180 ^ n1177 ;
  assign n1197 = n1184 & ~n1196 ;
  assign n1198 = n1197 ^ n1183 ;
  assign n1202 = n1201 ^ n1198 ;
  assign n1193 = n1166 ^ n1163 ;
  assign n1194 = n1170 & ~n1193 ;
  assign n1195 = n1194 ^ n1169 ;
  assign n1209 = n1198 ^ n1195 ;
  assign n1210 = n1202 & ~n1209 ;
  assign n1211 = n1210 ^ n1201 ;
  assign n1203 = n1202 ^ n1195 ;
  assign n1187 = n1186 ^ n1171 ;
  assign n1155 = n1154 ^ n1139 ;
  assign n1126 = x513 ^ x385 ;
  assign n1156 = n1155 ^ n1126 ;
  assign n1083 = x517 ^ x389 ;
  assign n1082 = x516 ^ x388 ;
  assign n1084 = n1083 ^ n1082 ;
  assign n1081 = x518 ^ x390 ;
  assign n1085 = n1084 ^ n1081 ;
  assign n1077 = x520 ^ x392 ;
  assign n1076 = x519 ^ x391 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1075 = x521 ^ x393 ;
  assign n1079 = n1078 ^ n1075 ;
  assign n1074 = x515 ^ x387 ;
  assign n1080 = n1079 ^ n1074 ;
  assign n1086 = n1085 ^ n1080 ;
  assign n1069 = x524 ^ x396 ;
  assign n1068 = x523 ^ x395 ;
  assign n1070 = n1069 ^ n1068 ;
  assign n1067 = x525 ^ x397 ;
  assign n1071 = n1070 ^ n1067 ;
  assign n1063 = x527 ^ x399 ;
  assign n1062 = x526 ^ x398 ;
  assign n1064 = n1063 ^ n1062 ;
  assign n1061 = x528 ^ x400 ;
  assign n1065 = n1064 ^ n1061 ;
  assign n1060 = x522 ^ x394 ;
  assign n1066 = n1065 ^ n1060 ;
  assign n1072 = n1071 ^ n1066 ;
  assign n1059 = x514 ^ x386 ;
  assign n1073 = n1072 ^ n1059 ;
  assign n1157 = n1086 ^ n1073 ;
  assign n1158 = n1157 ^ n1126 ;
  assign n1159 = n1156 & ~n1158 ;
  assign n1160 = n1159 ^ n1155 ;
  assign n1188 = n1187 ^ n1160 ;
  assign n1108 = n1076 ^ n1075 ;
  assign n1109 = n1078 & ~n1108 ;
  assign n1110 = n1109 ^ n1077 ;
  assign n1105 = n1085 ^ n1079 ;
  assign n1106 = ~n1080 & n1105 ;
  assign n1107 = n1106 ^ n1085 ;
  assign n1111 = n1110 ^ n1107 ;
  assign n1102 = n1082 ^ n1081 ;
  assign n1103 = n1084 & ~n1102 ;
  assign n1104 = n1103 ^ n1083 ;
  assign n1112 = n1111 ^ n1104 ;
  assign n1096 = n1071 ^ n1065 ;
  assign n1097 = ~n1066 & n1096 ;
  assign n1098 = n1097 ^ n1071 ;
  assign n1093 = n1062 ^ n1061 ;
  assign n1094 = n1064 & ~n1093 ;
  assign n1095 = n1094 ^ n1063 ;
  assign n1099 = n1098 ^ n1095 ;
  assign n1090 = n1068 ^ n1067 ;
  assign n1091 = n1070 & ~n1090 ;
  assign n1092 = n1091 ^ n1069 ;
  assign n1100 = n1099 ^ n1092 ;
  assign n1087 = n1086 ^ n1059 ;
  assign n1088 = n1073 & ~n1087 ;
  assign n1089 = n1088 ^ n1072 ;
  assign n1101 = n1100 ^ n1089 ;
  assign n1189 = n1112 ^ n1101 ;
  assign n1190 = n1189 ^ n1187 ;
  assign n1191 = n1188 & ~n1190 ;
  assign n1192 = n1191 ^ n1160 ;
  assign n1204 = n1203 ^ n1192 ;
  assign n1120 = n1107 ^ n1104 ;
  assign n1121 = n1111 & ~n1120 ;
  assign n1122 = n1121 ^ n1110 ;
  assign n1116 = n1095 ^ n1092 ;
  assign n1117 = n1099 & ~n1116 ;
  assign n1118 = n1117 ^ n1098 ;
  assign n1113 = n1112 ^ n1089 ;
  assign n1114 = n1101 & ~n1113 ;
  assign n1115 = n1114 ^ n1100 ;
  assign n1119 = n1118 ^ n1115 ;
  assign n1205 = n1122 ^ n1119 ;
  assign n1206 = n1205 ^ n1192 ;
  assign n1207 = n1204 & ~n1206 ;
  assign n1208 = n1207 ^ n1203 ;
  assign n1212 = n1211 ^ n1208 ;
  assign n1123 = n1122 ^ n1118 ;
  assign n1124 = ~n1119 & n1123 ;
  assign n1125 = n1124 ^ n1122 ;
  assign n1213 = n1212 ^ n1125 ;
  assign n1214 = n1189 ^ n1188 ;
  assign n1215 = n1157 ^ n1156 ;
  assign n1216 = x512 ^ x384 ;
  assign n1217 = n1215 & n1216 ;
  assign n1218 = n1214 & n1217 ;
  assign n1219 = n1205 ^ n1204 ;
  assign n1220 = n1218 & n1219 ;
  assign n1221 = n1213 & n1220 ;
  assign n1222 = n1208 ^ n1125 ;
  assign n1223 = n1212 & ~n1222 ;
  assign n1224 = n1223 ^ n1211 ;
  assign n1225 = n1221 & n1224 ;
  assign n1226 = n1058 & ~n1225 ;
  assign n1227 = n1226 ^ n1058 ;
  assign n1228 = ~n1056 & n1227 ;
  assign n1400 = ~n1054 & n1228 ;
  assign n1401 = n1400 ^ n1228 ;
  assign n1402 = n1401 ^ n1054 ;
  assign n1403 = n1402 ^ n1228 ;
  assign n1229 = n1227 ^ n1056 ;
  assign n1230 = n1229 ^ n1228 ;
  assign n1321 = x543 ^ x383 ;
  assign n1319 = x542 ^ x382 ;
  assign n1318 = x541 ^ x381 ;
  assign n1320 = n1319 ^ n1318 ;
  assign n1322 = n1321 ^ n1320 ;
  assign n1317 = x537 ^ x377 ;
  assign n1323 = n1322 ^ n1317 ;
  assign n1315 = x540 ^ x380 ;
  assign n1313 = x539 ^ x379 ;
  assign n1312 = x538 ^ x378 ;
  assign n1314 = n1313 ^ n1312 ;
  assign n1316 = n1315 ^ n1314 ;
  assign n1353 = n1317 ^ n1316 ;
  assign n1354 = n1323 & ~n1353 ;
  assign n1355 = n1354 ^ n1322 ;
  assign n1350 = n1321 ^ n1319 ;
  assign n1351 = ~n1320 & n1350 ;
  assign n1352 = n1351 ^ n1321 ;
  assign n1356 = n1355 ^ n1352 ;
  assign n1347 = n1315 ^ n1313 ;
  assign n1348 = ~n1314 & n1347 ;
  assign n1349 = n1348 ^ n1315 ;
  assign n1357 = n1356 ^ n1349 ;
  assign n1325 = x529 ^ x369 ;
  assign n1324 = n1323 ^ n1316 ;
  assign n1326 = n1325 ^ n1324 ;
  assign n1307 = x535 ^ x375 ;
  assign n1306 = x534 ^ x374 ;
  assign n1308 = n1307 ^ n1306 ;
  assign n1305 = x536 ^ x376 ;
  assign n1309 = n1308 ^ n1305 ;
  assign n1304 = x530 ^ x370 ;
  assign n1310 = n1309 ^ n1304 ;
  assign n1301 = x532 ^ x372 ;
  assign n1300 = x531 ^ x371 ;
  assign n1302 = n1301 ^ n1300 ;
  assign n1299 = x533 ^ x373 ;
  assign n1303 = n1302 ^ n1299 ;
  assign n1311 = n1310 ^ n1303 ;
  assign n1344 = n1324 ^ n1311 ;
  assign n1345 = n1326 & ~n1344 ;
  assign n1346 = n1345 ^ n1325 ;
  assign n1358 = n1357 ^ n1346 ;
  assign n1339 = n1304 ^ n1303 ;
  assign n1340 = n1310 & ~n1339 ;
  assign n1341 = n1340 ^ n1309 ;
  assign n1336 = n1306 ^ n1305 ;
  assign n1337 = n1308 & ~n1336 ;
  assign n1338 = n1337 ^ n1307 ;
  assign n1342 = n1341 ^ n1338 ;
  assign n1333 = n1300 ^ n1299 ;
  assign n1334 = n1302 & ~n1333 ;
  assign n1335 = n1334 ^ n1301 ;
  assign n1343 = n1342 ^ n1335 ;
  assign n1371 = n1346 ^ n1343 ;
  assign n1372 = n1358 & ~n1371 ;
  assign n1373 = n1372 ^ n1357 ;
  assign n1368 = n1352 ^ n1349 ;
  assign n1369 = n1356 & ~n1368 ;
  assign n1370 = n1369 ^ n1355 ;
  assign n1374 = n1373 ^ n1370 ;
  assign n1365 = n1338 ^ n1335 ;
  assign n1366 = n1342 & ~n1365 ;
  assign n1367 = n1366 ^ n1341 ;
  assign n1381 = n1370 ^ n1367 ;
  assign n1382 = n1374 & ~n1381 ;
  assign n1383 = n1382 ^ n1373 ;
  assign n1375 = n1374 ^ n1367 ;
  assign n1359 = n1358 ^ n1343 ;
  assign n1327 = n1326 ^ n1311 ;
  assign n1298 = x513 ^ x353 ;
  assign n1328 = n1327 ^ n1298 ;
  assign n1255 = x517 ^ x357 ;
  assign n1254 = x516 ^ x356 ;
  assign n1256 = n1255 ^ n1254 ;
  assign n1253 = x518 ^ x358 ;
  assign n1257 = n1256 ^ n1253 ;
  assign n1249 = x520 ^ x360 ;
  assign n1248 = x519 ^ x359 ;
  assign n1250 = n1249 ^ n1248 ;
  assign n1247 = x521 ^ x361 ;
  assign n1251 = n1250 ^ n1247 ;
  assign n1246 = x515 ^ x355 ;
  assign n1252 = n1251 ^ n1246 ;
  assign n1258 = n1257 ^ n1252 ;
  assign n1241 = x524 ^ x364 ;
  assign n1240 = x523 ^ x363 ;
  assign n1242 = n1241 ^ n1240 ;
  assign n1239 = x525 ^ x365 ;
  assign n1243 = n1242 ^ n1239 ;
  assign n1235 = x527 ^ x367 ;
  assign n1234 = x526 ^ x366 ;
  assign n1236 = n1235 ^ n1234 ;
  assign n1233 = x528 ^ x368 ;
  assign n1237 = n1236 ^ n1233 ;
  assign n1232 = x522 ^ x362 ;
  assign n1238 = n1237 ^ n1232 ;
  assign n1244 = n1243 ^ n1238 ;
  assign n1231 = x514 ^ x354 ;
  assign n1245 = n1244 ^ n1231 ;
  assign n1329 = n1258 ^ n1245 ;
  assign n1330 = n1329 ^ n1298 ;
  assign n1331 = n1328 & ~n1330 ;
  assign n1332 = n1331 ^ n1327 ;
  assign n1360 = n1359 ^ n1332 ;
  assign n1280 = n1248 ^ n1247 ;
  assign n1281 = n1250 & ~n1280 ;
  assign n1282 = n1281 ^ n1249 ;
  assign n1277 = n1257 ^ n1251 ;
  assign n1278 = ~n1252 & n1277 ;
  assign n1279 = n1278 ^ n1257 ;
  assign n1283 = n1282 ^ n1279 ;
  assign n1274 = n1254 ^ n1253 ;
  assign n1275 = n1256 & ~n1274 ;
  assign n1276 = n1275 ^ n1255 ;
  assign n1284 = n1283 ^ n1276 ;
  assign n1268 = n1243 ^ n1237 ;
  assign n1269 = ~n1238 & n1268 ;
  assign n1270 = n1269 ^ n1243 ;
  assign n1265 = n1234 ^ n1233 ;
  assign n1266 = n1236 & ~n1265 ;
  assign n1267 = n1266 ^ n1235 ;
  assign n1271 = n1270 ^ n1267 ;
  assign n1262 = n1240 ^ n1239 ;
  assign n1263 = n1242 & ~n1262 ;
  assign n1264 = n1263 ^ n1241 ;
  assign n1272 = n1271 ^ n1264 ;
  assign n1259 = n1258 ^ n1231 ;
  assign n1260 = n1245 & ~n1259 ;
  assign n1261 = n1260 ^ n1244 ;
  assign n1273 = n1272 ^ n1261 ;
  assign n1361 = n1284 ^ n1273 ;
  assign n1362 = n1361 ^ n1359 ;
  assign n1363 = n1360 & ~n1362 ;
  assign n1364 = n1363 ^ n1332 ;
  assign n1376 = n1375 ^ n1364 ;
  assign n1292 = n1279 ^ n1276 ;
  assign n1293 = n1283 & ~n1292 ;
  assign n1294 = n1293 ^ n1282 ;
  assign n1288 = n1267 ^ n1264 ;
  assign n1289 = n1271 & ~n1288 ;
  assign n1290 = n1289 ^ n1270 ;
  assign n1285 = n1284 ^ n1261 ;
  assign n1286 = n1273 & ~n1285 ;
  assign n1287 = n1286 ^ n1272 ;
  assign n1291 = n1290 ^ n1287 ;
  assign n1377 = n1294 ^ n1291 ;
  assign n1378 = n1377 ^ n1364 ;
  assign n1379 = n1376 & ~n1378 ;
  assign n1380 = n1379 ^ n1375 ;
  assign n1384 = n1383 ^ n1380 ;
  assign n1295 = n1294 ^ n1290 ;
  assign n1296 = ~n1291 & n1295 ;
  assign n1297 = n1296 ^ n1294 ;
  assign n1385 = n1384 ^ n1297 ;
  assign n1386 = n1361 ^ n1360 ;
  assign n1387 = n1329 ^ n1328 ;
  assign n1388 = x512 ^ x352 ;
  assign n1389 = n1387 & n1388 ;
  assign n1390 = n1386 & n1389 ;
  assign n1391 = n1377 ^ n1376 ;
  assign n1392 = n1390 & n1391 ;
  assign n1393 = n1385 & n1392 ;
  assign n1394 = n1380 ^ n1297 ;
  assign n1395 = n1384 & ~n1394 ;
  assign n1396 = n1395 ^ n1383 ;
  assign n1397 = n1393 & n1396 ;
  assign n1398 = ~n1230 & ~n1397 ;
  assign n1399 = n1398 ^ n1230 ;
  assign n1405 = n1403 ^ n1399 ;
  assign n1404 = ~n1399 & n1403 ;
  assign n1406 = n1405 ^ n1404 ;
  assign n1497 = x543 ^ x351 ;
  assign n1495 = x542 ^ x350 ;
  assign n1494 = x541 ^ x349 ;
  assign n1496 = n1495 ^ n1494 ;
  assign n1498 = n1497 ^ n1496 ;
  assign n1493 = x537 ^ x345 ;
  assign n1499 = n1498 ^ n1493 ;
  assign n1491 = x540 ^ x348 ;
  assign n1489 = x539 ^ x347 ;
  assign n1488 = x538 ^ x346 ;
  assign n1490 = n1489 ^ n1488 ;
  assign n1492 = n1491 ^ n1490 ;
  assign n1529 = n1493 ^ n1492 ;
  assign n1530 = n1499 & ~n1529 ;
  assign n1531 = n1530 ^ n1498 ;
  assign n1526 = n1497 ^ n1495 ;
  assign n1527 = ~n1496 & n1526 ;
  assign n1528 = n1527 ^ n1497 ;
  assign n1532 = n1531 ^ n1528 ;
  assign n1523 = n1491 ^ n1489 ;
  assign n1524 = ~n1490 & n1523 ;
  assign n1525 = n1524 ^ n1491 ;
  assign n1533 = n1532 ^ n1525 ;
  assign n1501 = x529 ^ x337 ;
  assign n1500 = n1499 ^ n1492 ;
  assign n1502 = n1501 ^ n1500 ;
  assign n1483 = x535 ^ x343 ;
  assign n1482 = x534 ^ x342 ;
  assign n1484 = n1483 ^ n1482 ;
  assign n1481 = x536 ^ x344 ;
  assign n1485 = n1484 ^ n1481 ;
  assign n1480 = x530 ^ x338 ;
  assign n1486 = n1485 ^ n1480 ;
  assign n1477 = x532 ^ x340 ;
  assign n1476 = x531 ^ x339 ;
  assign n1478 = n1477 ^ n1476 ;
  assign n1475 = x533 ^ x341 ;
  assign n1479 = n1478 ^ n1475 ;
  assign n1487 = n1486 ^ n1479 ;
  assign n1520 = n1500 ^ n1487 ;
  assign n1521 = n1502 & ~n1520 ;
  assign n1522 = n1521 ^ n1501 ;
  assign n1534 = n1533 ^ n1522 ;
  assign n1515 = n1480 ^ n1479 ;
  assign n1516 = n1486 & ~n1515 ;
  assign n1517 = n1516 ^ n1485 ;
  assign n1512 = n1482 ^ n1481 ;
  assign n1513 = n1484 & ~n1512 ;
  assign n1514 = n1513 ^ n1483 ;
  assign n1518 = n1517 ^ n1514 ;
  assign n1509 = n1476 ^ n1475 ;
  assign n1510 = n1478 & ~n1509 ;
  assign n1511 = n1510 ^ n1477 ;
  assign n1519 = n1518 ^ n1511 ;
  assign n1547 = n1522 ^ n1519 ;
  assign n1548 = n1534 & ~n1547 ;
  assign n1549 = n1548 ^ n1533 ;
  assign n1544 = n1528 ^ n1525 ;
  assign n1545 = n1532 & ~n1544 ;
  assign n1546 = n1545 ^ n1531 ;
  assign n1550 = n1549 ^ n1546 ;
  assign n1541 = n1514 ^ n1511 ;
  assign n1542 = n1518 & ~n1541 ;
  assign n1543 = n1542 ^ n1517 ;
  assign n1557 = n1546 ^ n1543 ;
  assign n1558 = n1550 & ~n1557 ;
  assign n1559 = n1558 ^ n1549 ;
  assign n1551 = n1550 ^ n1543 ;
  assign n1535 = n1534 ^ n1519 ;
  assign n1503 = n1502 ^ n1487 ;
  assign n1474 = x513 ^ x321 ;
  assign n1504 = n1503 ^ n1474 ;
  assign n1431 = x517 ^ x325 ;
  assign n1430 = x516 ^ x324 ;
  assign n1432 = n1431 ^ n1430 ;
  assign n1429 = x518 ^ x326 ;
  assign n1433 = n1432 ^ n1429 ;
  assign n1425 = x520 ^ x328 ;
  assign n1424 = x519 ^ x327 ;
  assign n1426 = n1425 ^ n1424 ;
  assign n1423 = x521 ^ x329 ;
  assign n1427 = n1426 ^ n1423 ;
  assign n1422 = x515 ^ x323 ;
  assign n1428 = n1427 ^ n1422 ;
  assign n1434 = n1433 ^ n1428 ;
  assign n1417 = x524 ^ x332 ;
  assign n1416 = x523 ^ x331 ;
  assign n1418 = n1417 ^ n1416 ;
  assign n1415 = x525 ^ x333 ;
  assign n1419 = n1418 ^ n1415 ;
  assign n1411 = x527 ^ x335 ;
  assign n1410 = x526 ^ x334 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1409 = x528 ^ x336 ;
  assign n1413 = n1412 ^ n1409 ;
  assign n1408 = x522 ^ x330 ;
  assign n1414 = n1413 ^ n1408 ;
  assign n1420 = n1419 ^ n1414 ;
  assign n1407 = x514 ^ x322 ;
  assign n1421 = n1420 ^ n1407 ;
  assign n1505 = n1434 ^ n1421 ;
  assign n1506 = n1505 ^ n1474 ;
  assign n1507 = n1504 & ~n1506 ;
  assign n1508 = n1507 ^ n1503 ;
  assign n1536 = n1535 ^ n1508 ;
  assign n1456 = n1424 ^ n1423 ;
  assign n1457 = n1426 & ~n1456 ;
  assign n1458 = n1457 ^ n1425 ;
  assign n1453 = n1433 ^ n1427 ;
  assign n1454 = ~n1428 & n1453 ;
  assign n1455 = n1454 ^ n1433 ;
  assign n1459 = n1458 ^ n1455 ;
  assign n1450 = n1430 ^ n1429 ;
  assign n1451 = n1432 & ~n1450 ;
  assign n1452 = n1451 ^ n1431 ;
  assign n1460 = n1459 ^ n1452 ;
  assign n1444 = n1419 ^ n1413 ;
  assign n1445 = ~n1414 & n1444 ;
  assign n1446 = n1445 ^ n1419 ;
  assign n1441 = n1410 ^ n1409 ;
  assign n1442 = n1412 & ~n1441 ;
  assign n1443 = n1442 ^ n1411 ;
  assign n1447 = n1446 ^ n1443 ;
  assign n1438 = n1416 ^ n1415 ;
  assign n1439 = n1418 & ~n1438 ;
  assign n1440 = n1439 ^ n1417 ;
  assign n1448 = n1447 ^ n1440 ;
  assign n1435 = n1434 ^ n1407 ;
  assign n1436 = n1421 & ~n1435 ;
  assign n1437 = n1436 ^ n1420 ;
  assign n1449 = n1448 ^ n1437 ;
  assign n1537 = n1460 ^ n1449 ;
  assign n1538 = n1537 ^ n1535 ;
  assign n1539 = n1536 & ~n1538 ;
  assign n1540 = n1539 ^ n1508 ;
  assign n1552 = n1551 ^ n1540 ;
  assign n1468 = n1455 ^ n1452 ;
  assign n1469 = n1459 & ~n1468 ;
  assign n1470 = n1469 ^ n1458 ;
  assign n1464 = n1443 ^ n1440 ;
  assign n1465 = n1447 & ~n1464 ;
  assign n1466 = n1465 ^ n1446 ;
  assign n1461 = n1460 ^ n1437 ;
  assign n1462 = n1449 & ~n1461 ;
  assign n1463 = n1462 ^ n1448 ;
  assign n1467 = n1466 ^ n1463 ;
  assign n1553 = n1470 ^ n1467 ;
  assign n1554 = n1553 ^ n1540 ;
  assign n1555 = n1552 & ~n1554 ;
  assign n1556 = n1555 ^ n1551 ;
  assign n1560 = n1559 ^ n1556 ;
  assign n1471 = n1470 ^ n1466 ;
  assign n1472 = ~n1467 & n1471 ;
  assign n1473 = n1472 ^ n1470 ;
  assign n1561 = n1560 ^ n1473 ;
  assign n1562 = n1537 ^ n1536 ;
  assign n1563 = n1505 ^ n1504 ;
  assign n1564 = x512 ^ x320 ;
  assign n1565 = n1563 & n1564 ;
  assign n1566 = n1562 & n1565 ;
  assign n1567 = n1553 ^ n1552 ;
  assign n1568 = n1566 & n1567 ;
  assign n1569 = n1561 & n1568 ;
  assign n1570 = n1556 ^ n1473 ;
  assign n1571 = n1560 & ~n1570 ;
  assign n1572 = n1571 ^ n1559 ;
  assign n1573 = n1569 & n1572 ;
  assign n1574 = ~n1406 & ~n1573 ;
  assign n1575 = n1574 ^ n1406 ;
  assign n1576 = n1401 & ~n1404 ;
  assign n1577 = n1576 ^ n1404 ;
  assign n1578 = ~n1575 & n1577 ;
  assign n1579 = n1576 ^ n1401 ;
  assign n1580 = n1578 & ~n1579 ;
  assign n1581 = n1580 ^ n1578 ;
  assign n1582 = n1581 ^ n1579 ;
  assign n1583 = n1582 ^ n1578 ;
  assign n1584 = n1577 ^ n1575 ;
  assign n1585 = n1584 ^ n1578 ;
  assign n1676 = x543 ^ x319 ;
  assign n1674 = x542 ^ x318 ;
  assign n1673 = x541 ^ x317 ;
  assign n1675 = n1674 ^ n1673 ;
  assign n1677 = n1676 ^ n1675 ;
  assign n1672 = x537 ^ x313 ;
  assign n1678 = n1677 ^ n1672 ;
  assign n1670 = x540 ^ x316 ;
  assign n1668 = x539 ^ x315 ;
  assign n1667 = x538 ^ x314 ;
  assign n1669 = n1668 ^ n1667 ;
  assign n1671 = n1670 ^ n1669 ;
  assign n1708 = n1672 ^ n1671 ;
  assign n1709 = n1678 & ~n1708 ;
  assign n1710 = n1709 ^ n1677 ;
  assign n1705 = n1676 ^ n1674 ;
  assign n1706 = ~n1675 & n1705 ;
  assign n1707 = n1706 ^ n1676 ;
  assign n1711 = n1710 ^ n1707 ;
  assign n1702 = n1670 ^ n1668 ;
  assign n1703 = ~n1669 & n1702 ;
  assign n1704 = n1703 ^ n1670 ;
  assign n1712 = n1711 ^ n1704 ;
  assign n1680 = x529 ^ x305 ;
  assign n1679 = n1678 ^ n1671 ;
  assign n1681 = n1680 ^ n1679 ;
  assign n1662 = x535 ^ x311 ;
  assign n1661 = x534 ^ x310 ;
  assign n1663 = n1662 ^ n1661 ;
  assign n1660 = x536 ^ x312 ;
  assign n1664 = n1663 ^ n1660 ;
  assign n1659 = x530 ^ x306 ;
  assign n1665 = n1664 ^ n1659 ;
  assign n1656 = x532 ^ x308 ;
  assign n1655 = x531 ^ x307 ;
  assign n1657 = n1656 ^ n1655 ;
  assign n1654 = x533 ^ x309 ;
  assign n1658 = n1657 ^ n1654 ;
  assign n1666 = n1665 ^ n1658 ;
  assign n1699 = n1679 ^ n1666 ;
  assign n1700 = n1681 & ~n1699 ;
  assign n1701 = n1700 ^ n1680 ;
  assign n1713 = n1712 ^ n1701 ;
  assign n1694 = n1659 ^ n1658 ;
  assign n1695 = n1665 & ~n1694 ;
  assign n1696 = n1695 ^ n1664 ;
  assign n1691 = n1661 ^ n1660 ;
  assign n1692 = n1663 & ~n1691 ;
  assign n1693 = n1692 ^ n1662 ;
  assign n1697 = n1696 ^ n1693 ;
  assign n1688 = n1655 ^ n1654 ;
  assign n1689 = n1657 & ~n1688 ;
  assign n1690 = n1689 ^ n1656 ;
  assign n1698 = n1697 ^ n1690 ;
  assign n1726 = n1701 ^ n1698 ;
  assign n1727 = n1713 & ~n1726 ;
  assign n1728 = n1727 ^ n1712 ;
  assign n1723 = n1707 ^ n1704 ;
  assign n1724 = n1711 & ~n1723 ;
  assign n1725 = n1724 ^ n1710 ;
  assign n1729 = n1728 ^ n1725 ;
  assign n1720 = n1693 ^ n1690 ;
  assign n1721 = n1697 & ~n1720 ;
  assign n1722 = n1721 ^ n1696 ;
  assign n1736 = n1725 ^ n1722 ;
  assign n1737 = n1729 & ~n1736 ;
  assign n1738 = n1737 ^ n1728 ;
  assign n1730 = n1729 ^ n1722 ;
  assign n1714 = n1713 ^ n1698 ;
  assign n1682 = n1681 ^ n1666 ;
  assign n1653 = x513 ^ x289 ;
  assign n1683 = n1682 ^ n1653 ;
  assign n1610 = x517 ^ x293 ;
  assign n1609 = x516 ^ x292 ;
  assign n1611 = n1610 ^ n1609 ;
  assign n1608 = x518 ^ x294 ;
  assign n1612 = n1611 ^ n1608 ;
  assign n1604 = x520 ^ x296 ;
  assign n1603 = x519 ^ x295 ;
  assign n1605 = n1604 ^ n1603 ;
  assign n1602 = x521 ^ x297 ;
  assign n1606 = n1605 ^ n1602 ;
  assign n1601 = x515 ^ x291 ;
  assign n1607 = n1606 ^ n1601 ;
  assign n1613 = n1612 ^ n1607 ;
  assign n1596 = x524 ^ x300 ;
  assign n1595 = x523 ^ x299 ;
  assign n1597 = n1596 ^ n1595 ;
  assign n1594 = x525 ^ x301 ;
  assign n1598 = n1597 ^ n1594 ;
  assign n1590 = x527 ^ x303 ;
  assign n1589 = x526 ^ x302 ;
  assign n1591 = n1590 ^ n1589 ;
  assign n1588 = x528 ^ x304 ;
  assign n1592 = n1591 ^ n1588 ;
  assign n1587 = x522 ^ x298 ;
  assign n1593 = n1592 ^ n1587 ;
  assign n1599 = n1598 ^ n1593 ;
  assign n1586 = x514 ^ x290 ;
  assign n1600 = n1599 ^ n1586 ;
  assign n1684 = n1613 ^ n1600 ;
  assign n1685 = n1684 ^ n1653 ;
  assign n1686 = n1683 & ~n1685 ;
  assign n1687 = n1686 ^ n1682 ;
  assign n1715 = n1714 ^ n1687 ;
  assign n1635 = n1603 ^ n1602 ;
  assign n1636 = n1605 & ~n1635 ;
  assign n1637 = n1636 ^ n1604 ;
  assign n1632 = n1612 ^ n1606 ;
  assign n1633 = ~n1607 & n1632 ;
  assign n1634 = n1633 ^ n1612 ;
  assign n1638 = n1637 ^ n1634 ;
  assign n1629 = n1609 ^ n1608 ;
  assign n1630 = n1611 & ~n1629 ;
  assign n1631 = n1630 ^ n1610 ;
  assign n1639 = n1638 ^ n1631 ;
  assign n1623 = n1598 ^ n1592 ;
  assign n1624 = ~n1593 & n1623 ;
  assign n1625 = n1624 ^ n1598 ;
  assign n1620 = n1589 ^ n1588 ;
  assign n1621 = n1591 & ~n1620 ;
  assign n1622 = n1621 ^ n1590 ;
  assign n1626 = n1625 ^ n1622 ;
  assign n1617 = n1595 ^ n1594 ;
  assign n1618 = n1597 & ~n1617 ;
  assign n1619 = n1618 ^ n1596 ;
  assign n1627 = n1626 ^ n1619 ;
  assign n1614 = n1613 ^ n1586 ;
  assign n1615 = n1600 & ~n1614 ;
  assign n1616 = n1615 ^ n1599 ;
  assign n1628 = n1627 ^ n1616 ;
  assign n1716 = n1639 ^ n1628 ;
  assign n1717 = n1716 ^ n1714 ;
  assign n1718 = n1715 & ~n1717 ;
  assign n1719 = n1718 ^ n1687 ;
  assign n1731 = n1730 ^ n1719 ;
  assign n1647 = n1634 ^ n1631 ;
  assign n1648 = n1638 & ~n1647 ;
  assign n1649 = n1648 ^ n1637 ;
  assign n1643 = n1622 ^ n1619 ;
  assign n1644 = n1626 & ~n1643 ;
  assign n1645 = n1644 ^ n1625 ;
  assign n1640 = n1639 ^ n1616 ;
  assign n1641 = n1628 & ~n1640 ;
  assign n1642 = n1641 ^ n1627 ;
  assign n1646 = n1645 ^ n1642 ;
  assign n1732 = n1649 ^ n1646 ;
  assign n1733 = n1732 ^ n1719 ;
  assign n1734 = n1731 & ~n1733 ;
  assign n1735 = n1734 ^ n1730 ;
  assign n1739 = n1738 ^ n1735 ;
  assign n1650 = n1649 ^ n1645 ;
  assign n1651 = ~n1646 & n1650 ;
  assign n1652 = n1651 ^ n1649 ;
  assign n1740 = n1739 ^ n1652 ;
  assign n1741 = n1716 ^ n1715 ;
  assign n1742 = n1684 ^ n1683 ;
  assign n1743 = x512 ^ x288 ;
  assign n1744 = n1742 & n1743 ;
  assign n1745 = n1741 & n1744 ;
  assign n1746 = n1732 ^ n1731 ;
  assign n1747 = n1745 & n1746 ;
  assign n1748 = n1740 & n1747 ;
  assign n1749 = n1735 ^ n1652 ;
  assign n1750 = n1739 & ~n1749 ;
  assign n1751 = n1750 ^ n1738 ;
  assign n1752 = n1748 & n1751 ;
  assign n1753 = ~n1585 & ~n1752 ;
  assign n1754 = n1753 ^ n1585 ;
  assign n1755 = n1583 & ~n1754 ;
  assign n1756 = ~n1581 & n1755 ;
  assign n1757 = n1756 ^ n1755 ;
  assign n1758 = n1757 ^ n1581 ;
  assign n1759 = n1758 ^ n1755 ;
  assign n1760 = n1754 ^ n1583 ;
  assign n1761 = n1760 ^ n1755 ;
  assign n1852 = x543 ^ x287 ;
  assign n1850 = x542 ^ x286 ;
  assign n1849 = x541 ^ x285 ;
  assign n1851 = n1850 ^ n1849 ;
  assign n1853 = n1852 ^ n1851 ;
  assign n1848 = x537 ^ x281 ;
  assign n1854 = n1853 ^ n1848 ;
  assign n1846 = x540 ^ x284 ;
  assign n1844 = x539 ^ x283 ;
  assign n1843 = x538 ^ x282 ;
  assign n1845 = n1844 ^ n1843 ;
  assign n1847 = n1846 ^ n1845 ;
  assign n1884 = n1848 ^ n1847 ;
  assign n1885 = n1854 & ~n1884 ;
  assign n1886 = n1885 ^ n1853 ;
  assign n1881 = n1852 ^ n1850 ;
  assign n1882 = ~n1851 & n1881 ;
  assign n1883 = n1882 ^ n1852 ;
  assign n1887 = n1886 ^ n1883 ;
  assign n1878 = n1846 ^ n1844 ;
  assign n1879 = ~n1845 & n1878 ;
  assign n1880 = n1879 ^ n1846 ;
  assign n1888 = n1887 ^ n1880 ;
  assign n1856 = x529 ^ x273 ;
  assign n1855 = n1854 ^ n1847 ;
  assign n1857 = n1856 ^ n1855 ;
  assign n1838 = x535 ^ x279 ;
  assign n1837 = x534 ^ x278 ;
  assign n1839 = n1838 ^ n1837 ;
  assign n1836 = x536 ^ x280 ;
  assign n1840 = n1839 ^ n1836 ;
  assign n1835 = x530 ^ x274 ;
  assign n1841 = n1840 ^ n1835 ;
  assign n1832 = x532 ^ x276 ;
  assign n1831 = x531 ^ x275 ;
  assign n1833 = n1832 ^ n1831 ;
  assign n1830 = x533 ^ x277 ;
  assign n1834 = n1833 ^ n1830 ;
  assign n1842 = n1841 ^ n1834 ;
  assign n1875 = n1855 ^ n1842 ;
  assign n1876 = n1857 & ~n1875 ;
  assign n1877 = n1876 ^ n1856 ;
  assign n1889 = n1888 ^ n1877 ;
  assign n1870 = n1835 ^ n1834 ;
  assign n1871 = n1841 & ~n1870 ;
  assign n1872 = n1871 ^ n1840 ;
  assign n1867 = n1837 ^ n1836 ;
  assign n1868 = n1839 & ~n1867 ;
  assign n1869 = n1868 ^ n1838 ;
  assign n1873 = n1872 ^ n1869 ;
  assign n1864 = n1831 ^ n1830 ;
  assign n1865 = n1833 & ~n1864 ;
  assign n1866 = n1865 ^ n1832 ;
  assign n1874 = n1873 ^ n1866 ;
  assign n1902 = n1877 ^ n1874 ;
  assign n1903 = n1889 & ~n1902 ;
  assign n1904 = n1903 ^ n1888 ;
  assign n1899 = n1883 ^ n1880 ;
  assign n1900 = n1887 & ~n1899 ;
  assign n1901 = n1900 ^ n1886 ;
  assign n1905 = n1904 ^ n1901 ;
  assign n1896 = n1869 ^ n1866 ;
  assign n1897 = n1873 & ~n1896 ;
  assign n1898 = n1897 ^ n1872 ;
  assign n1912 = n1901 ^ n1898 ;
  assign n1913 = n1905 & ~n1912 ;
  assign n1914 = n1913 ^ n1904 ;
  assign n1906 = n1905 ^ n1898 ;
  assign n1890 = n1889 ^ n1874 ;
  assign n1858 = n1857 ^ n1842 ;
  assign n1829 = x513 ^ x257 ;
  assign n1859 = n1858 ^ n1829 ;
  assign n1786 = x517 ^ x261 ;
  assign n1785 = x516 ^ x260 ;
  assign n1787 = n1786 ^ n1785 ;
  assign n1784 = x518 ^ x262 ;
  assign n1788 = n1787 ^ n1784 ;
  assign n1780 = x520 ^ x264 ;
  assign n1779 = x519 ^ x263 ;
  assign n1781 = n1780 ^ n1779 ;
  assign n1778 = x521 ^ x265 ;
  assign n1782 = n1781 ^ n1778 ;
  assign n1777 = x515 ^ x259 ;
  assign n1783 = n1782 ^ n1777 ;
  assign n1789 = n1788 ^ n1783 ;
  assign n1772 = x524 ^ x268 ;
  assign n1771 = x523 ^ x267 ;
  assign n1773 = n1772 ^ n1771 ;
  assign n1770 = x525 ^ x269 ;
  assign n1774 = n1773 ^ n1770 ;
  assign n1766 = x527 ^ x271 ;
  assign n1765 = x526 ^ x270 ;
  assign n1767 = n1766 ^ n1765 ;
  assign n1764 = x528 ^ x272 ;
  assign n1768 = n1767 ^ n1764 ;
  assign n1763 = x522 ^ x266 ;
  assign n1769 = n1768 ^ n1763 ;
  assign n1775 = n1774 ^ n1769 ;
  assign n1762 = x514 ^ x258 ;
  assign n1776 = n1775 ^ n1762 ;
  assign n1860 = n1789 ^ n1776 ;
  assign n1861 = n1860 ^ n1829 ;
  assign n1862 = n1859 & ~n1861 ;
  assign n1863 = n1862 ^ n1858 ;
  assign n1891 = n1890 ^ n1863 ;
  assign n1811 = n1779 ^ n1778 ;
  assign n1812 = n1781 & ~n1811 ;
  assign n1813 = n1812 ^ n1780 ;
  assign n1808 = n1788 ^ n1782 ;
  assign n1809 = ~n1783 & n1808 ;
  assign n1810 = n1809 ^ n1788 ;
  assign n1814 = n1813 ^ n1810 ;
  assign n1805 = n1785 ^ n1784 ;
  assign n1806 = n1787 & ~n1805 ;
  assign n1807 = n1806 ^ n1786 ;
  assign n1815 = n1814 ^ n1807 ;
  assign n1799 = n1774 ^ n1768 ;
  assign n1800 = ~n1769 & n1799 ;
  assign n1801 = n1800 ^ n1774 ;
  assign n1796 = n1765 ^ n1764 ;
  assign n1797 = n1767 & ~n1796 ;
  assign n1798 = n1797 ^ n1766 ;
  assign n1802 = n1801 ^ n1798 ;
  assign n1793 = n1771 ^ n1770 ;
  assign n1794 = n1773 & ~n1793 ;
  assign n1795 = n1794 ^ n1772 ;
  assign n1803 = n1802 ^ n1795 ;
  assign n1790 = n1789 ^ n1762 ;
  assign n1791 = n1776 & ~n1790 ;
  assign n1792 = n1791 ^ n1775 ;
  assign n1804 = n1803 ^ n1792 ;
  assign n1892 = n1815 ^ n1804 ;
  assign n1893 = n1892 ^ n1890 ;
  assign n1894 = n1891 & ~n1893 ;
  assign n1895 = n1894 ^ n1863 ;
  assign n1907 = n1906 ^ n1895 ;
  assign n1823 = n1810 ^ n1807 ;
  assign n1824 = n1814 & ~n1823 ;
  assign n1825 = n1824 ^ n1813 ;
  assign n1819 = n1798 ^ n1795 ;
  assign n1820 = n1802 & ~n1819 ;
  assign n1821 = n1820 ^ n1801 ;
  assign n1816 = n1815 ^ n1792 ;
  assign n1817 = n1804 & ~n1816 ;
  assign n1818 = n1817 ^ n1803 ;
  assign n1822 = n1821 ^ n1818 ;
  assign n1908 = n1825 ^ n1822 ;
  assign n1909 = n1908 ^ n1895 ;
  assign n1910 = n1907 & ~n1909 ;
  assign n1911 = n1910 ^ n1906 ;
  assign n1915 = n1914 ^ n1911 ;
  assign n1826 = n1825 ^ n1821 ;
  assign n1827 = ~n1822 & n1826 ;
  assign n1828 = n1827 ^ n1825 ;
  assign n1916 = n1915 ^ n1828 ;
  assign n1917 = n1892 ^ n1891 ;
  assign n1918 = n1860 ^ n1859 ;
  assign n1919 = x512 ^ x256 ;
  assign n1920 = n1918 & n1919 ;
  assign n1921 = n1917 & n1920 ;
  assign n1922 = n1908 ^ n1907 ;
  assign n1923 = n1921 & n1922 ;
  assign n1924 = n1916 & n1923 ;
  assign n1925 = n1911 ^ n1828 ;
  assign n1926 = n1915 & ~n1925 ;
  assign n1927 = n1926 ^ n1914 ;
  assign n1928 = n1924 & n1927 ;
  assign n1929 = ~n1761 & ~n1928 ;
  assign n1930 = n1929 ^ n1761 ;
  assign n1931 = n1759 & ~n1930 ;
  assign n1932 = n1757 & ~n1931 ;
  assign n1933 = n1932 ^ n1931 ;
  assign n1934 = n1930 ^ n1759 ;
  assign n1935 = n1934 ^ n1931 ;
  assign n2026 = x543 ^ x255 ;
  assign n2024 = x542 ^ x254 ;
  assign n2023 = x541 ^ x253 ;
  assign n2025 = n2024 ^ n2023 ;
  assign n2027 = n2026 ^ n2025 ;
  assign n2022 = x537 ^ x249 ;
  assign n2028 = n2027 ^ n2022 ;
  assign n2020 = x540 ^ x252 ;
  assign n2018 = x539 ^ x251 ;
  assign n2017 = x538 ^ x250 ;
  assign n2019 = n2018 ^ n2017 ;
  assign n2021 = n2020 ^ n2019 ;
  assign n2058 = n2022 ^ n2021 ;
  assign n2059 = n2028 & ~n2058 ;
  assign n2060 = n2059 ^ n2027 ;
  assign n2055 = n2026 ^ n2024 ;
  assign n2056 = ~n2025 & n2055 ;
  assign n2057 = n2056 ^ n2026 ;
  assign n2061 = n2060 ^ n2057 ;
  assign n2052 = n2020 ^ n2018 ;
  assign n2053 = ~n2019 & n2052 ;
  assign n2054 = n2053 ^ n2020 ;
  assign n2062 = n2061 ^ n2054 ;
  assign n2030 = x529 ^ x241 ;
  assign n2029 = n2028 ^ n2021 ;
  assign n2031 = n2030 ^ n2029 ;
  assign n2012 = x535 ^ x247 ;
  assign n2011 = x534 ^ x246 ;
  assign n2013 = n2012 ^ n2011 ;
  assign n2010 = x536 ^ x248 ;
  assign n2014 = n2013 ^ n2010 ;
  assign n2009 = x530 ^ x242 ;
  assign n2015 = n2014 ^ n2009 ;
  assign n2006 = x532 ^ x244 ;
  assign n2005 = x531 ^ x243 ;
  assign n2007 = n2006 ^ n2005 ;
  assign n2004 = x533 ^ x245 ;
  assign n2008 = n2007 ^ n2004 ;
  assign n2016 = n2015 ^ n2008 ;
  assign n2049 = n2029 ^ n2016 ;
  assign n2050 = n2031 & ~n2049 ;
  assign n2051 = n2050 ^ n2030 ;
  assign n2063 = n2062 ^ n2051 ;
  assign n2044 = n2009 ^ n2008 ;
  assign n2045 = n2015 & ~n2044 ;
  assign n2046 = n2045 ^ n2014 ;
  assign n2041 = n2011 ^ n2010 ;
  assign n2042 = n2013 & ~n2041 ;
  assign n2043 = n2042 ^ n2012 ;
  assign n2047 = n2046 ^ n2043 ;
  assign n2038 = n2005 ^ n2004 ;
  assign n2039 = n2007 & ~n2038 ;
  assign n2040 = n2039 ^ n2006 ;
  assign n2048 = n2047 ^ n2040 ;
  assign n2076 = n2051 ^ n2048 ;
  assign n2077 = n2063 & ~n2076 ;
  assign n2078 = n2077 ^ n2062 ;
  assign n2073 = n2057 ^ n2054 ;
  assign n2074 = n2061 & ~n2073 ;
  assign n2075 = n2074 ^ n2060 ;
  assign n2079 = n2078 ^ n2075 ;
  assign n2070 = n2043 ^ n2040 ;
  assign n2071 = n2047 & ~n2070 ;
  assign n2072 = n2071 ^ n2046 ;
  assign n2086 = n2075 ^ n2072 ;
  assign n2087 = n2079 & ~n2086 ;
  assign n2088 = n2087 ^ n2078 ;
  assign n2080 = n2079 ^ n2072 ;
  assign n2064 = n2063 ^ n2048 ;
  assign n2032 = n2031 ^ n2016 ;
  assign n2003 = x513 ^ x225 ;
  assign n2033 = n2032 ^ n2003 ;
  assign n1960 = x517 ^ x229 ;
  assign n1959 = x516 ^ x228 ;
  assign n1961 = n1960 ^ n1959 ;
  assign n1958 = x518 ^ x230 ;
  assign n1962 = n1961 ^ n1958 ;
  assign n1954 = x520 ^ x232 ;
  assign n1953 = x519 ^ x231 ;
  assign n1955 = n1954 ^ n1953 ;
  assign n1952 = x521 ^ x233 ;
  assign n1956 = n1955 ^ n1952 ;
  assign n1951 = x515 ^ x227 ;
  assign n1957 = n1956 ^ n1951 ;
  assign n1963 = n1962 ^ n1957 ;
  assign n1946 = x524 ^ x236 ;
  assign n1945 = x523 ^ x235 ;
  assign n1947 = n1946 ^ n1945 ;
  assign n1944 = x525 ^ x237 ;
  assign n1948 = n1947 ^ n1944 ;
  assign n1940 = x527 ^ x239 ;
  assign n1939 = x526 ^ x238 ;
  assign n1941 = n1940 ^ n1939 ;
  assign n1938 = x528 ^ x240 ;
  assign n1942 = n1941 ^ n1938 ;
  assign n1937 = x522 ^ x234 ;
  assign n1943 = n1942 ^ n1937 ;
  assign n1949 = n1948 ^ n1943 ;
  assign n1936 = x514 ^ x226 ;
  assign n1950 = n1949 ^ n1936 ;
  assign n2034 = n1963 ^ n1950 ;
  assign n2035 = n2034 ^ n2003 ;
  assign n2036 = n2033 & ~n2035 ;
  assign n2037 = n2036 ^ n2032 ;
  assign n2065 = n2064 ^ n2037 ;
  assign n1985 = n1953 ^ n1952 ;
  assign n1986 = n1955 & ~n1985 ;
  assign n1987 = n1986 ^ n1954 ;
  assign n1982 = n1962 ^ n1956 ;
  assign n1983 = ~n1957 & n1982 ;
  assign n1984 = n1983 ^ n1962 ;
  assign n1988 = n1987 ^ n1984 ;
  assign n1979 = n1959 ^ n1958 ;
  assign n1980 = n1961 & ~n1979 ;
  assign n1981 = n1980 ^ n1960 ;
  assign n1989 = n1988 ^ n1981 ;
  assign n1973 = n1948 ^ n1942 ;
  assign n1974 = ~n1943 & n1973 ;
  assign n1975 = n1974 ^ n1948 ;
  assign n1970 = n1939 ^ n1938 ;
  assign n1971 = n1941 & ~n1970 ;
  assign n1972 = n1971 ^ n1940 ;
  assign n1976 = n1975 ^ n1972 ;
  assign n1967 = n1945 ^ n1944 ;
  assign n1968 = n1947 & ~n1967 ;
  assign n1969 = n1968 ^ n1946 ;
  assign n1977 = n1976 ^ n1969 ;
  assign n1964 = n1963 ^ n1936 ;
  assign n1965 = n1950 & ~n1964 ;
  assign n1966 = n1965 ^ n1949 ;
  assign n1978 = n1977 ^ n1966 ;
  assign n2066 = n1989 ^ n1978 ;
  assign n2067 = n2066 ^ n2064 ;
  assign n2068 = n2065 & ~n2067 ;
  assign n2069 = n2068 ^ n2037 ;
  assign n2081 = n2080 ^ n2069 ;
  assign n1997 = n1984 ^ n1981 ;
  assign n1998 = n1988 & ~n1997 ;
  assign n1999 = n1998 ^ n1987 ;
  assign n1993 = n1972 ^ n1969 ;
  assign n1994 = n1976 & ~n1993 ;
  assign n1995 = n1994 ^ n1975 ;
  assign n1990 = n1989 ^ n1966 ;
  assign n1991 = n1978 & ~n1990 ;
  assign n1992 = n1991 ^ n1977 ;
  assign n1996 = n1995 ^ n1992 ;
  assign n2082 = n1999 ^ n1996 ;
  assign n2083 = n2082 ^ n2069 ;
  assign n2084 = n2081 & ~n2083 ;
  assign n2085 = n2084 ^ n2080 ;
  assign n2089 = n2088 ^ n2085 ;
  assign n2000 = n1999 ^ n1995 ;
  assign n2001 = ~n1996 & n2000 ;
  assign n2002 = n2001 ^ n1999 ;
  assign n2090 = n2089 ^ n2002 ;
  assign n2091 = n2066 ^ n2065 ;
  assign n2092 = n2034 ^ n2033 ;
  assign n2093 = x512 ^ x224 ;
  assign n2094 = n2092 & n2093 ;
  assign n2095 = n2091 & n2094 ;
  assign n2096 = n2082 ^ n2081 ;
  assign n2097 = n2095 & n2096 ;
  assign n2098 = n2090 & n2097 ;
  assign n2099 = n2085 ^ n2002 ;
  assign n2100 = n2089 & ~n2099 ;
  assign n2101 = n2100 ^ n2088 ;
  assign n2102 = n2098 & n2101 ;
  assign n2103 = ~n1935 & ~n2102 ;
  assign n2104 = n2103 ^ n1935 ;
  assign n2105 = n1933 & ~n2104 ;
  assign n2106 = n1932 ^ n1757 ;
  assign n2107 = n2105 & ~n2106 ;
  assign n2108 = n2107 ^ n2105 ;
  assign n2109 = n2104 ^ n1933 ;
  assign n2110 = n2109 ^ n2105 ;
  assign n2201 = x543 ^ x223 ;
  assign n2199 = x542 ^ x222 ;
  assign n2198 = x541 ^ x221 ;
  assign n2200 = n2199 ^ n2198 ;
  assign n2202 = n2201 ^ n2200 ;
  assign n2197 = x537 ^ x217 ;
  assign n2203 = n2202 ^ n2197 ;
  assign n2195 = x540 ^ x220 ;
  assign n2193 = x539 ^ x219 ;
  assign n2192 = x538 ^ x218 ;
  assign n2194 = n2193 ^ n2192 ;
  assign n2196 = n2195 ^ n2194 ;
  assign n2233 = n2197 ^ n2196 ;
  assign n2234 = n2203 & ~n2233 ;
  assign n2235 = n2234 ^ n2202 ;
  assign n2230 = n2201 ^ n2199 ;
  assign n2231 = ~n2200 & n2230 ;
  assign n2232 = n2231 ^ n2201 ;
  assign n2236 = n2235 ^ n2232 ;
  assign n2227 = n2195 ^ n2193 ;
  assign n2228 = ~n2194 & n2227 ;
  assign n2229 = n2228 ^ n2195 ;
  assign n2237 = n2236 ^ n2229 ;
  assign n2205 = x529 ^ x209 ;
  assign n2204 = n2203 ^ n2196 ;
  assign n2206 = n2205 ^ n2204 ;
  assign n2187 = x535 ^ x215 ;
  assign n2186 = x534 ^ x214 ;
  assign n2188 = n2187 ^ n2186 ;
  assign n2185 = x536 ^ x216 ;
  assign n2189 = n2188 ^ n2185 ;
  assign n2184 = x530 ^ x210 ;
  assign n2190 = n2189 ^ n2184 ;
  assign n2181 = x532 ^ x212 ;
  assign n2180 = x531 ^ x211 ;
  assign n2182 = n2181 ^ n2180 ;
  assign n2179 = x533 ^ x213 ;
  assign n2183 = n2182 ^ n2179 ;
  assign n2191 = n2190 ^ n2183 ;
  assign n2224 = n2204 ^ n2191 ;
  assign n2225 = n2206 & ~n2224 ;
  assign n2226 = n2225 ^ n2205 ;
  assign n2238 = n2237 ^ n2226 ;
  assign n2219 = n2184 ^ n2183 ;
  assign n2220 = n2190 & ~n2219 ;
  assign n2221 = n2220 ^ n2189 ;
  assign n2216 = n2186 ^ n2185 ;
  assign n2217 = n2188 & ~n2216 ;
  assign n2218 = n2217 ^ n2187 ;
  assign n2222 = n2221 ^ n2218 ;
  assign n2213 = n2180 ^ n2179 ;
  assign n2214 = n2182 & ~n2213 ;
  assign n2215 = n2214 ^ n2181 ;
  assign n2223 = n2222 ^ n2215 ;
  assign n2251 = n2226 ^ n2223 ;
  assign n2252 = n2238 & ~n2251 ;
  assign n2253 = n2252 ^ n2237 ;
  assign n2248 = n2232 ^ n2229 ;
  assign n2249 = n2236 & ~n2248 ;
  assign n2250 = n2249 ^ n2235 ;
  assign n2254 = n2253 ^ n2250 ;
  assign n2245 = n2218 ^ n2215 ;
  assign n2246 = n2222 & ~n2245 ;
  assign n2247 = n2246 ^ n2221 ;
  assign n2261 = n2250 ^ n2247 ;
  assign n2262 = n2254 & ~n2261 ;
  assign n2263 = n2262 ^ n2253 ;
  assign n2255 = n2254 ^ n2247 ;
  assign n2239 = n2238 ^ n2223 ;
  assign n2207 = n2206 ^ n2191 ;
  assign n2178 = x513 ^ x193 ;
  assign n2208 = n2207 ^ n2178 ;
  assign n2135 = x517 ^ x197 ;
  assign n2134 = x516 ^ x196 ;
  assign n2136 = n2135 ^ n2134 ;
  assign n2133 = x518 ^ x198 ;
  assign n2137 = n2136 ^ n2133 ;
  assign n2129 = x520 ^ x200 ;
  assign n2128 = x519 ^ x199 ;
  assign n2130 = n2129 ^ n2128 ;
  assign n2127 = x521 ^ x201 ;
  assign n2131 = n2130 ^ n2127 ;
  assign n2126 = x515 ^ x195 ;
  assign n2132 = n2131 ^ n2126 ;
  assign n2138 = n2137 ^ n2132 ;
  assign n2121 = x524 ^ x204 ;
  assign n2120 = x523 ^ x203 ;
  assign n2122 = n2121 ^ n2120 ;
  assign n2119 = x525 ^ x205 ;
  assign n2123 = n2122 ^ n2119 ;
  assign n2115 = x527 ^ x207 ;
  assign n2114 = x526 ^ x206 ;
  assign n2116 = n2115 ^ n2114 ;
  assign n2113 = x528 ^ x208 ;
  assign n2117 = n2116 ^ n2113 ;
  assign n2112 = x522 ^ x202 ;
  assign n2118 = n2117 ^ n2112 ;
  assign n2124 = n2123 ^ n2118 ;
  assign n2111 = x514 ^ x194 ;
  assign n2125 = n2124 ^ n2111 ;
  assign n2209 = n2138 ^ n2125 ;
  assign n2210 = n2209 ^ n2178 ;
  assign n2211 = n2208 & ~n2210 ;
  assign n2212 = n2211 ^ n2207 ;
  assign n2240 = n2239 ^ n2212 ;
  assign n2160 = n2128 ^ n2127 ;
  assign n2161 = n2130 & ~n2160 ;
  assign n2162 = n2161 ^ n2129 ;
  assign n2157 = n2137 ^ n2131 ;
  assign n2158 = ~n2132 & n2157 ;
  assign n2159 = n2158 ^ n2137 ;
  assign n2163 = n2162 ^ n2159 ;
  assign n2154 = n2134 ^ n2133 ;
  assign n2155 = n2136 & ~n2154 ;
  assign n2156 = n2155 ^ n2135 ;
  assign n2164 = n2163 ^ n2156 ;
  assign n2148 = n2123 ^ n2117 ;
  assign n2149 = ~n2118 & n2148 ;
  assign n2150 = n2149 ^ n2123 ;
  assign n2145 = n2114 ^ n2113 ;
  assign n2146 = n2116 & ~n2145 ;
  assign n2147 = n2146 ^ n2115 ;
  assign n2151 = n2150 ^ n2147 ;
  assign n2142 = n2120 ^ n2119 ;
  assign n2143 = n2122 & ~n2142 ;
  assign n2144 = n2143 ^ n2121 ;
  assign n2152 = n2151 ^ n2144 ;
  assign n2139 = n2138 ^ n2111 ;
  assign n2140 = n2125 & ~n2139 ;
  assign n2141 = n2140 ^ n2124 ;
  assign n2153 = n2152 ^ n2141 ;
  assign n2241 = n2164 ^ n2153 ;
  assign n2242 = n2241 ^ n2239 ;
  assign n2243 = n2240 & ~n2242 ;
  assign n2244 = n2243 ^ n2212 ;
  assign n2256 = n2255 ^ n2244 ;
  assign n2172 = n2159 ^ n2156 ;
  assign n2173 = n2163 & ~n2172 ;
  assign n2174 = n2173 ^ n2162 ;
  assign n2168 = n2147 ^ n2144 ;
  assign n2169 = n2151 & ~n2168 ;
  assign n2170 = n2169 ^ n2150 ;
  assign n2165 = n2164 ^ n2141 ;
  assign n2166 = n2153 & ~n2165 ;
  assign n2167 = n2166 ^ n2152 ;
  assign n2171 = n2170 ^ n2167 ;
  assign n2257 = n2174 ^ n2171 ;
  assign n2258 = n2257 ^ n2244 ;
  assign n2259 = n2256 & ~n2258 ;
  assign n2260 = n2259 ^ n2255 ;
  assign n2264 = n2263 ^ n2260 ;
  assign n2175 = n2174 ^ n2170 ;
  assign n2176 = ~n2171 & n2175 ;
  assign n2177 = n2176 ^ n2174 ;
  assign n2265 = n2264 ^ n2177 ;
  assign n2266 = n2241 ^ n2240 ;
  assign n2267 = n2209 ^ n2208 ;
  assign n2268 = x512 ^ x192 ;
  assign n2269 = n2267 & n2268 ;
  assign n2270 = n2266 & n2269 ;
  assign n2271 = n2257 ^ n2256 ;
  assign n2272 = n2270 & n2271 ;
  assign n2273 = n2265 & n2272 ;
  assign n2274 = n2260 ^ n2177 ;
  assign n2275 = n2264 & ~n2274 ;
  assign n2276 = n2275 ^ n2263 ;
  assign n2277 = n2273 & n2276 ;
  assign n2278 = ~n2110 & ~n2277 ;
  assign n2279 = n2278 ^ n2110 ;
  assign n2280 = n2108 ^ n2106 ;
  assign n2281 = n2280 ^ n2105 ;
  assign n2282 = ~n2279 & n2281 ;
  assign n2283 = ~n2108 & n2282 ;
  assign n2284 = n2283 ^ n2282 ;
  assign n2285 = n2281 ^ n2279 ;
  assign n2286 = n2285 ^ n2282 ;
  assign n2377 = x543 ^ x191 ;
  assign n2375 = x542 ^ x190 ;
  assign n2374 = x541 ^ x189 ;
  assign n2376 = n2375 ^ n2374 ;
  assign n2378 = n2377 ^ n2376 ;
  assign n2373 = x537 ^ x185 ;
  assign n2379 = n2378 ^ n2373 ;
  assign n2371 = x540 ^ x188 ;
  assign n2369 = x539 ^ x187 ;
  assign n2368 = x538 ^ x186 ;
  assign n2370 = n2369 ^ n2368 ;
  assign n2372 = n2371 ^ n2370 ;
  assign n2409 = n2373 ^ n2372 ;
  assign n2410 = n2379 & ~n2409 ;
  assign n2411 = n2410 ^ n2378 ;
  assign n2406 = n2377 ^ n2375 ;
  assign n2407 = ~n2376 & n2406 ;
  assign n2408 = n2407 ^ n2377 ;
  assign n2412 = n2411 ^ n2408 ;
  assign n2403 = n2371 ^ n2369 ;
  assign n2404 = ~n2370 & n2403 ;
  assign n2405 = n2404 ^ n2371 ;
  assign n2413 = n2412 ^ n2405 ;
  assign n2381 = x529 ^ x177 ;
  assign n2380 = n2379 ^ n2372 ;
  assign n2382 = n2381 ^ n2380 ;
  assign n2363 = x535 ^ x183 ;
  assign n2362 = x534 ^ x182 ;
  assign n2364 = n2363 ^ n2362 ;
  assign n2361 = x536 ^ x184 ;
  assign n2365 = n2364 ^ n2361 ;
  assign n2360 = x530 ^ x178 ;
  assign n2366 = n2365 ^ n2360 ;
  assign n2357 = x532 ^ x180 ;
  assign n2356 = x531 ^ x179 ;
  assign n2358 = n2357 ^ n2356 ;
  assign n2355 = x533 ^ x181 ;
  assign n2359 = n2358 ^ n2355 ;
  assign n2367 = n2366 ^ n2359 ;
  assign n2400 = n2380 ^ n2367 ;
  assign n2401 = n2382 & ~n2400 ;
  assign n2402 = n2401 ^ n2381 ;
  assign n2414 = n2413 ^ n2402 ;
  assign n2395 = n2360 ^ n2359 ;
  assign n2396 = n2366 & ~n2395 ;
  assign n2397 = n2396 ^ n2365 ;
  assign n2392 = n2362 ^ n2361 ;
  assign n2393 = n2364 & ~n2392 ;
  assign n2394 = n2393 ^ n2363 ;
  assign n2398 = n2397 ^ n2394 ;
  assign n2389 = n2356 ^ n2355 ;
  assign n2390 = n2358 & ~n2389 ;
  assign n2391 = n2390 ^ n2357 ;
  assign n2399 = n2398 ^ n2391 ;
  assign n2427 = n2402 ^ n2399 ;
  assign n2428 = n2414 & ~n2427 ;
  assign n2429 = n2428 ^ n2413 ;
  assign n2424 = n2408 ^ n2405 ;
  assign n2425 = n2412 & ~n2424 ;
  assign n2426 = n2425 ^ n2411 ;
  assign n2430 = n2429 ^ n2426 ;
  assign n2421 = n2394 ^ n2391 ;
  assign n2422 = n2398 & ~n2421 ;
  assign n2423 = n2422 ^ n2397 ;
  assign n2437 = n2426 ^ n2423 ;
  assign n2438 = n2430 & ~n2437 ;
  assign n2439 = n2438 ^ n2429 ;
  assign n2431 = n2430 ^ n2423 ;
  assign n2415 = n2414 ^ n2399 ;
  assign n2383 = n2382 ^ n2367 ;
  assign n2354 = x513 ^ x161 ;
  assign n2384 = n2383 ^ n2354 ;
  assign n2311 = x517 ^ x165 ;
  assign n2310 = x516 ^ x164 ;
  assign n2312 = n2311 ^ n2310 ;
  assign n2309 = x518 ^ x166 ;
  assign n2313 = n2312 ^ n2309 ;
  assign n2305 = x520 ^ x168 ;
  assign n2304 = x519 ^ x167 ;
  assign n2306 = n2305 ^ n2304 ;
  assign n2303 = x521 ^ x169 ;
  assign n2307 = n2306 ^ n2303 ;
  assign n2302 = x515 ^ x163 ;
  assign n2308 = n2307 ^ n2302 ;
  assign n2314 = n2313 ^ n2308 ;
  assign n2297 = x524 ^ x172 ;
  assign n2296 = x523 ^ x171 ;
  assign n2298 = n2297 ^ n2296 ;
  assign n2295 = x525 ^ x173 ;
  assign n2299 = n2298 ^ n2295 ;
  assign n2291 = x527 ^ x175 ;
  assign n2290 = x526 ^ x174 ;
  assign n2292 = n2291 ^ n2290 ;
  assign n2289 = x528 ^ x176 ;
  assign n2293 = n2292 ^ n2289 ;
  assign n2288 = x522 ^ x170 ;
  assign n2294 = n2293 ^ n2288 ;
  assign n2300 = n2299 ^ n2294 ;
  assign n2287 = x514 ^ x162 ;
  assign n2301 = n2300 ^ n2287 ;
  assign n2385 = n2314 ^ n2301 ;
  assign n2386 = n2385 ^ n2354 ;
  assign n2387 = n2384 & ~n2386 ;
  assign n2388 = n2387 ^ n2383 ;
  assign n2416 = n2415 ^ n2388 ;
  assign n2336 = n2304 ^ n2303 ;
  assign n2337 = n2306 & ~n2336 ;
  assign n2338 = n2337 ^ n2305 ;
  assign n2333 = n2313 ^ n2307 ;
  assign n2334 = ~n2308 & n2333 ;
  assign n2335 = n2334 ^ n2313 ;
  assign n2339 = n2338 ^ n2335 ;
  assign n2330 = n2310 ^ n2309 ;
  assign n2331 = n2312 & ~n2330 ;
  assign n2332 = n2331 ^ n2311 ;
  assign n2340 = n2339 ^ n2332 ;
  assign n2324 = n2299 ^ n2293 ;
  assign n2325 = ~n2294 & n2324 ;
  assign n2326 = n2325 ^ n2299 ;
  assign n2321 = n2290 ^ n2289 ;
  assign n2322 = n2292 & ~n2321 ;
  assign n2323 = n2322 ^ n2291 ;
  assign n2327 = n2326 ^ n2323 ;
  assign n2318 = n2296 ^ n2295 ;
  assign n2319 = n2298 & ~n2318 ;
  assign n2320 = n2319 ^ n2297 ;
  assign n2328 = n2327 ^ n2320 ;
  assign n2315 = n2314 ^ n2287 ;
  assign n2316 = n2301 & ~n2315 ;
  assign n2317 = n2316 ^ n2300 ;
  assign n2329 = n2328 ^ n2317 ;
  assign n2417 = n2340 ^ n2329 ;
  assign n2418 = n2417 ^ n2415 ;
  assign n2419 = n2416 & ~n2418 ;
  assign n2420 = n2419 ^ n2388 ;
  assign n2432 = n2431 ^ n2420 ;
  assign n2348 = n2335 ^ n2332 ;
  assign n2349 = n2339 & ~n2348 ;
  assign n2350 = n2349 ^ n2338 ;
  assign n2344 = n2323 ^ n2320 ;
  assign n2345 = n2327 & ~n2344 ;
  assign n2346 = n2345 ^ n2326 ;
  assign n2341 = n2340 ^ n2317 ;
  assign n2342 = n2329 & ~n2341 ;
  assign n2343 = n2342 ^ n2328 ;
  assign n2347 = n2346 ^ n2343 ;
  assign n2433 = n2350 ^ n2347 ;
  assign n2434 = n2433 ^ n2420 ;
  assign n2435 = n2432 & ~n2434 ;
  assign n2436 = n2435 ^ n2431 ;
  assign n2440 = n2439 ^ n2436 ;
  assign n2351 = n2350 ^ n2346 ;
  assign n2352 = ~n2347 & n2351 ;
  assign n2353 = n2352 ^ n2350 ;
  assign n2441 = n2440 ^ n2353 ;
  assign n2442 = n2417 ^ n2416 ;
  assign n2443 = n2385 ^ n2384 ;
  assign n2444 = x512 ^ x160 ;
  assign n2445 = n2443 & n2444 ;
  assign n2446 = n2442 & n2445 ;
  assign n2447 = n2433 ^ n2432 ;
  assign n2448 = n2446 & n2447 ;
  assign n2449 = n2441 & n2448 ;
  assign n2450 = n2436 ^ n2353 ;
  assign n2451 = n2440 & ~n2450 ;
  assign n2452 = n2451 ^ n2439 ;
  assign n2453 = n2449 & n2452 ;
  assign n2454 = ~n2286 & ~n2453 ;
  assign n2455 = n2454 ^ n2286 ;
  assign n2456 = n2284 ^ n2108 ;
  assign n2457 = n2456 ^ n2282 ;
  assign n2458 = ~n2455 & n2457 ;
  assign n2459 = n2284 & ~n2458 ;
  assign n2460 = n2459 ^ n2458 ;
  assign n2461 = n2457 ^ n2455 ;
  assign n2462 = n2461 ^ n2458 ;
  assign n2553 = x543 ^ x159 ;
  assign n2551 = x542 ^ x158 ;
  assign n2550 = x541 ^ x157 ;
  assign n2552 = n2551 ^ n2550 ;
  assign n2554 = n2553 ^ n2552 ;
  assign n2549 = x537 ^ x153 ;
  assign n2555 = n2554 ^ n2549 ;
  assign n2547 = x540 ^ x156 ;
  assign n2545 = x539 ^ x155 ;
  assign n2544 = x538 ^ x154 ;
  assign n2546 = n2545 ^ n2544 ;
  assign n2548 = n2547 ^ n2546 ;
  assign n2585 = n2549 ^ n2548 ;
  assign n2586 = n2555 & ~n2585 ;
  assign n2587 = n2586 ^ n2554 ;
  assign n2582 = n2553 ^ n2551 ;
  assign n2583 = ~n2552 & n2582 ;
  assign n2584 = n2583 ^ n2553 ;
  assign n2588 = n2587 ^ n2584 ;
  assign n2579 = n2547 ^ n2545 ;
  assign n2580 = ~n2546 & n2579 ;
  assign n2581 = n2580 ^ n2547 ;
  assign n2589 = n2588 ^ n2581 ;
  assign n2557 = x529 ^ x145 ;
  assign n2556 = n2555 ^ n2548 ;
  assign n2558 = n2557 ^ n2556 ;
  assign n2539 = x535 ^ x151 ;
  assign n2538 = x534 ^ x150 ;
  assign n2540 = n2539 ^ n2538 ;
  assign n2537 = x536 ^ x152 ;
  assign n2541 = n2540 ^ n2537 ;
  assign n2536 = x530 ^ x146 ;
  assign n2542 = n2541 ^ n2536 ;
  assign n2533 = x532 ^ x148 ;
  assign n2532 = x531 ^ x147 ;
  assign n2534 = n2533 ^ n2532 ;
  assign n2531 = x533 ^ x149 ;
  assign n2535 = n2534 ^ n2531 ;
  assign n2543 = n2542 ^ n2535 ;
  assign n2576 = n2556 ^ n2543 ;
  assign n2577 = n2558 & ~n2576 ;
  assign n2578 = n2577 ^ n2557 ;
  assign n2590 = n2589 ^ n2578 ;
  assign n2571 = n2536 ^ n2535 ;
  assign n2572 = n2542 & ~n2571 ;
  assign n2573 = n2572 ^ n2541 ;
  assign n2568 = n2538 ^ n2537 ;
  assign n2569 = n2540 & ~n2568 ;
  assign n2570 = n2569 ^ n2539 ;
  assign n2574 = n2573 ^ n2570 ;
  assign n2565 = n2532 ^ n2531 ;
  assign n2566 = n2534 & ~n2565 ;
  assign n2567 = n2566 ^ n2533 ;
  assign n2575 = n2574 ^ n2567 ;
  assign n2603 = n2578 ^ n2575 ;
  assign n2604 = n2590 & ~n2603 ;
  assign n2605 = n2604 ^ n2589 ;
  assign n2600 = n2584 ^ n2581 ;
  assign n2601 = n2588 & ~n2600 ;
  assign n2602 = n2601 ^ n2587 ;
  assign n2606 = n2605 ^ n2602 ;
  assign n2597 = n2570 ^ n2567 ;
  assign n2598 = n2574 & ~n2597 ;
  assign n2599 = n2598 ^ n2573 ;
  assign n2613 = n2602 ^ n2599 ;
  assign n2614 = n2606 & ~n2613 ;
  assign n2615 = n2614 ^ n2605 ;
  assign n2607 = n2606 ^ n2599 ;
  assign n2591 = n2590 ^ n2575 ;
  assign n2559 = n2558 ^ n2543 ;
  assign n2530 = x513 ^ x129 ;
  assign n2560 = n2559 ^ n2530 ;
  assign n2487 = x517 ^ x133 ;
  assign n2486 = x516 ^ x132 ;
  assign n2488 = n2487 ^ n2486 ;
  assign n2485 = x518 ^ x134 ;
  assign n2489 = n2488 ^ n2485 ;
  assign n2481 = x520 ^ x136 ;
  assign n2480 = x519 ^ x135 ;
  assign n2482 = n2481 ^ n2480 ;
  assign n2479 = x521 ^ x137 ;
  assign n2483 = n2482 ^ n2479 ;
  assign n2478 = x515 ^ x131 ;
  assign n2484 = n2483 ^ n2478 ;
  assign n2490 = n2489 ^ n2484 ;
  assign n2473 = x524 ^ x140 ;
  assign n2472 = x523 ^ x139 ;
  assign n2474 = n2473 ^ n2472 ;
  assign n2471 = x525 ^ x141 ;
  assign n2475 = n2474 ^ n2471 ;
  assign n2467 = x527 ^ x143 ;
  assign n2466 = x526 ^ x142 ;
  assign n2468 = n2467 ^ n2466 ;
  assign n2465 = x528 ^ x144 ;
  assign n2469 = n2468 ^ n2465 ;
  assign n2464 = x522 ^ x138 ;
  assign n2470 = n2469 ^ n2464 ;
  assign n2476 = n2475 ^ n2470 ;
  assign n2463 = x514 ^ x130 ;
  assign n2477 = n2476 ^ n2463 ;
  assign n2561 = n2490 ^ n2477 ;
  assign n2562 = n2561 ^ n2530 ;
  assign n2563 = n2560 & ~n2562 ;
  assign n2564 = n2563 ^ n2559 ;
  assign n2592 = n2591 ^ n2564 ;
  assign n2512 = n2480 ^ n2479 ;
  assign n2513 = n2482 & ~n2512 ;
  assign n2514 = n2513 ^ n2481 ;
  assign n2509 = n2489 ^ n2483 ;
  assign n2510 = ~n2484 & n2509 ;
  assign n2511 = n2510 ^ n2489 ;
  assign n2515 = n2514 ^ n2511 ;
  assign n2506 = n2486 ^ n2485 ;
  assign n2507 = n2488 & ~n2506 ;
  assign n2508 = n2507 ^ n2487 ;
  assign n2516 = n2515 ^ n2508 ;
  assign n2500 = n2475 ^ n2469 ;
  assign n2501 = ~n2470 & n2500 ;
  assign n2502 = n2501 ^ n2475 ;
  assign n2497 = n2466 ^ n2465 ;
  assign n2498 = n2468 & ~n2497 ;
  assign n2499 = n2498 ^ n2467 ;
  assign n2503 = n2502 ^ n2499 ;
  assign n2494 = n2472 ^ n2471 ;
  assign n2495 = n2474 & ~n2494 ;
  assign n2496 = n2495 ^ n2473 ;
  assign n2504 = n2503 ^ n2496 ;
  assign n2491 = n2490 ^ n2463 ;
  assign n2492 = n2477 & ~n2491 ;
  assign n2493 = n2492 ^ n2476 ;
  assign n2505 = n2504 ^ n2493 ;
  assign n2593 = n2516 ^ n2505 ;
  assign n2594 = n2593 ^ n2591 ;
  assign n2595 = n2592 & ~n2594 ;
  assign n2596 = n2595 ^ n2564 ;
  assign n2608 = n2607 ^ n2596 ;
  assign n2524 = n2511 ^ n2508 ;
  assign n2525 = n2515 & ~n2524 ;
  assign n2526 = n2525 ^ n2514 ;
  assign n2520 = n2499 ^ n2496 ;
  assign n2521 = n2503 & ~n2520 ;
  assign n2522 = n2521 ^ n2502 ;
  assign n2517 = n2516 ^ n2493 ;
  assign n2518 = n2505 & ~n2517 ;
  assign n2519 = n2518 ^ n2504 ;
  assign n2523 = n2522 ^ n2519 ;
  assign n2609 = n2526 ^ n2523 ;
  assign n2610 = n2609 ^ n2596 ;
  assign n2611 = n2608 & ~n2610 ;
  assign n2612 = n2611 ^ n2607 ;
  assign n2616 = n2615 ^ n2612 ;
  assign n2527 = n2526 ^ n2522 ;
  assign n2528 = ~n2523 & n2527 ;
  assign n2529 = n2528 ^ n2526 ;
  assign n2617 = n2616 ^ n2529 ;
  assign n2618 = n2593 ^ n2592 ;
  assign n2619 = n2561 ^ n2560 ;
  assign n2620 = x512 ^ x128 ;
  assign n2621 = n2619 & n2620 ;
  assign n2622 = n2618 & n2621 ;
  assign n2623 = n2609 ^ n2608 ;
  assign n2624 = n2622 & n2623 ;
  assign n2625 = n2617 & n2624 ;
  assign n2626 = n2612 ^ n2529 ;
  assign n2627 = n2616 & ~n2626 ;
  assign n2628 = n2627 ^ n2615 ;
  assign n2629 = n2625 & n2628 ;
  assign n2630 = ~n2462 & ~n2629 ;
  assign n2631 = n2630 ^ n2462 ;
  assign n2632 = n2460 & ~n2631 ;
  assign n2633 = n2459 ^ n2284 ;
  assign n2634 = n2632 & ~n2633 ;
  assign n2635 = n2634 ^ n2632 ;
  assign n2636 = n2631 ^ n2460 ;
  assign n2637 = n2636 ^ n2632 ;
  assign n2728 = x543 ^ x127 ;
  assign n2726 = x542 ^ x126 ;
  assign n2725 = x541 ^ x125 ;
  assign n2727 = n2726 ^ n2725 ;
  assign n2729 = n2728 ^ n2727 ;
  assign n2724 = x537 ^ x121 ;
  assign n2730 = n2729 ^ n2724 ;
  assign n2722 = x540 ^ x124 ;
  assign n2720 = x539 ^ x123 ;
  assign n2719 = x538 ^ x122 ;
  assign n2721 = n2720 ^ n2719 ;
  assign n2723 = n2722 ^ n2721 ;
  assign n2760 = n2724 ^ n2723 ;
  assign n2761 = n2730 & ~n2760 ;
  assign n2762 = n2761 ^ n2729 ;
  assign n2757 = n2728 ^ n2726 ;
  assign n2758 = ~n2727 & n2757 ;
  assign n2759 = n2758 ^ n2728 ;
  assign n2763 = n2762 ^ n2759 ;
  assign n2754 = n2722 ^ n2720 ;
  assign n2755 = ~n2721 & n2754 ;
  assign n2756 = n2755 ^ n2722 ;
  assign n2764 = n2763 ^ n2756 ;
  assign n2732 = x529 ^ x113 ;
  assign n2731 = n2730 ^ n2723 ;
  assign n2733 = n2732 ^ n2731 ;
  assign n2714 = x535 ^ x119 ;
  assign n2713 = x534 ^ x118 ;
  assign n2715 = n2714 ^ n2713 ;
  assign n2712 = x536 ^ x120 ;
  assign n2716 = n2715 ^ n2712 ;
  assign n2711 = x530 ^ x114 ;
  assign n2717 = n2716 ^ n2711 ;
  assign n2708 = x532 ^ x116 ;
  assign n2707 = x531 ^ x115 ;
  assign n2709 = n2708 ^ n2707 ;
  assign n2706 = x533 ^ x117 ;
  assign n2710 = n2709 ^ n2706 ;
  assign n2718 = n2717 ^ n2710 ;
  assign n2751 = n2731 ^ n2718 ;
  assign n2752 = n2733 & ~n2751 ;
  assign n2753 = n2752 ^ n2732 ;
  assign n2765 = n2764 ^ n2753 ;
  assign n2746 = n2711 ^ n2710 ;
  assign n2747 = n2717 & ~n2746 ;
  assign n2748 = n2747 ^ n2716 ;
  assign n2743 = n2713 ^ n2712 ;
  assign n2744 = n2715 & ~n2743 ;
  assign n2745 = n2744 ^ n2714 ;
  assign n2749 = n2748 ^ n2745 ;
  assign n2740 = n2707 ^ n2706 ;
  assign n2741 = n2709 & ~n2740 ;
  assign n2742 = n2741 ^ n2708 ;
  assign n2750 = n2749 ^ n2742 ;
  assign n2778 = n2753 ^ n2750 ;
  assign n2779 = n2765 & ~n2778 ;
  assign n2780 = n2779 ^ n2764 ;
  assign n2775 = n2759 ^ n2756 ;
  assign n2776 = n2763 & ~n2775 ;
  assign n2777 = n2776 ^ n2762 ;
  assign n2781 = n2780 ^ n2777 ;
  assign n2772 = n2745 ^ n2742 ;
  assign n2773 = n2749 & ~n2772 ;
  assign n2774 = n2773 ^ n2748 ;
  assign n2788 = n2777 ^ n2774 ;
  assign n2789 = n2781 & ~n2788 ;
  assign n2790 = n2789 ^ n2780 ;
  assign n2782 = n2781 ^ n2774 ;
  assign n2766 = n2765 ^ n2750 ;
  assign n2734 = n2733 ^ n2718 ;
  assign n2705 = x513 ^ x97 ;
  assign n2735 = n2734 ^ n2705 ;
  assign n2662 = x517 ^ x101 ;
  assign n2661 = x516 ^ x100 ;
  assign n2663 = n2662 ^ n2661 ;
  assign n2660 = x518 ^ x102 ;
  assign n2664 = n2663 ^ n2660 ;
  assign n2656 = x520 ^ x104 ;
  assign n2655 = x519 ^ x103 ;
  assign n2657 = n2656 ^ n2655 ;
  assign n2654 = x521 ^ x105 ;
  assign n2658 = n2657 ^ n2654 ;
  assign n2653 = x515 ^ x99 ;
  assign n2659 = n2658 ^ n2653 ;
  assign n2665 = n2664 ^ n2659 ;
  assign n2648 = x524 ^ x108 ;
  assign n2647 = x523 ^ x107 ;
  assign n2649 = n2648 ^ n2647 ;
  assign n2646 = x525 ^ x109 ;
  assign n2650 = n2649 ^ n2646 ;
  assign n2642 = x527 ^ x111 ;
  assign n2641 = x526 ^ x110 ;
  assign n2643 = n2642 ^ n2641 ;
  assign n2640 = x528 ^ x112 ;
  assign n2644 = n2643 ^ n2640 ;
  assign n2639 = x522 ^ x106 ;
  assign n2645 = n2644 ^ n2639 ;
  assign n2651 = n2650 ^ n2645 ;
  assign n2638 = x514 ^ x98 ;
  assign n2652 = n2651 ^ n2638 ;
  assign n2736 = n2665 ^ n2652 ;
  assign n2737 = n2736 ^ n2705 ;
  assign n2738 = n2735 & ~n2737 ;
  assign n2739 = n2738 ^ n2734 ;
  assign n2767 = n2766 ^ n2739 ;
  assign n2687 = n2655 ^ n2654 ;
  assign n2688 = n2657 & ~n2687 ;
  assign n2689 = n2688 ^ n2656 ;
  assign n2684 = n2664 ^ n2658 ;
  assign n2685 = ~n2659 & n2684 ;
  assign n2686 = n2685 ^ n2664 ;
  assign n2690 = n2689 ^ n2686 ;
  assign n2681 = n2661 ^ n2660 ;
  assign n2682 = n2663 & ~n2681 ;
  assign n2683 = n2682 ^ n2662 ;
  assign n2691 = n2690 ^ n2683 ;
  assign n2675 = n2650 ^ n2644 ;
  assign n2676 = ~n2645 & n2675 ;
  assign n2677 = n2676 ^ n2650 ;
  assign n2672 = n2641 ^ n2640 ;
  assign n2673 = n2643 & ~n2672 ;
  assign n2674 = n2673 ^ n2642 ;
  assign n2678 = n2677 ^ n2674 ;
  assign n2669 = n2647 ^ n2646 ;
  assign n2670 = n2649 & ~n2669 ;
  assign n2671 = n2670 ^ n2648 ;
  assign n2679 = n2678 ^ n2671 ;
  assign n2666 = n2665 ^ n2638 ;
  assign n2667 = n2652 & ~n2666 ;
  assign n2668 = n2667 ^ n2651 ;
  assign n2680 = n2679 ^ n2668 ;
  assign n2768 = n2691 ^ n2680 ;
  assign n2769 = n2768 ^ n2766 ;
  assign n2770 = n2767 & ~n2769 ;
  assign n2771 = n2770 ^ n2739 ;
  assign n2783 = n2782 ^ n2771 ;
  assign n2699 = n2686 ^ n2683 ;
  assign n2700 = n2690 & ~n2699 ;
  assign n2701 = n2700 ^ n2689 ;
  assign n2695 = n2674 ^ n2671 ;
  assign n2696 = n2678 & ~n2695 ;
  assign n2697 = n2696 ^ n2677 ;
  assign n2692 = n2691 ^ n2668 ;
  assign n2693 = n2680 & ~n2692 ;
  assign n2694 = n2693 ^ n2679 ;
  assign n2698 = n2697 ^ n2694 ;
  assign n2784 = n2701 ^ n2698 ;
  assign n2785 = n2784 ^ n2771 ;
  assign n2786 = n2783 & ~n2785 ;
  assign n2787 = n2786 ^ n2782 ;
  assign n2791 = n2790 ^ n2787 ;
  assign n2702 = n2701 ^ n2697 ;
  assign n2703 = ~n2698 & n2702 ;
  assign n2704 = n2703 ^ n2701 ;
  assign n2792 = n2791 ^ n2704 ;
  assign n2793 = n2768 ^ n2767 ;
  assign n2794 = n2736 ^ n2735 ;
  assign n2795 = x512 ^ x96 ;
  assign n2796 = n2794 & n2795 ;
  assign n2797 = n2793 & n2796 ;
  assign n2798 = n2784 ^ n2783 ;
  assign n2799 = n2797 & n2798 ;
  assign n2800 = n2792 & n2799 ;
  assign n2801 = n2787 ^ n2704 ;
  assign n2802 = n2791 & ~n2801 ;
  assign n2803 = n2802 ^ n2790 ;
  assign n2804 = n2800 & n2803 ;
  assign n2805 = ~n2637 & ~n2804 ;
  assign n2806 = n2805 ^ n2637 ;
  assign n2807 = n2635 ^ n2633 ;
  assign n2808 = n2807 ^ n2632 ;
  assign n2809 = ~n2806 & n2808 ;
  assign n2810 = ~n2635 & n2809 ;
  assign n2811 = n2810 ^ n2809 ;
  assign n2812 = n2811 ^ n2635 ;
  assign n2813 = n2812 ^ n2809 ;
  assign n2814 = n2808 ^ n2806 ;
  assign n2815 = n2814 ^ n2809 ;
  assign n2906 = x543 ^ x95 ;
  assign n2904 = x542 ^ x94 ;
  assign n2903 = x541 ^ x93 ;
  assign n2905 = n2904 ^ n2903 ;
  assign n2907 = n2906 ^ n2905 ;
  assign n2902 = x537 ^ x89 ;
  assign n2908 = n2907 ^ n2902 ;
  assign n2900 = x540 ^ x92 ;
  assign n2898 = x539 ^ x91 ;
  assign n2897 = x538 ^ x90 ;
  assign n2899 = n2898 ^ n2897 ;
  assign n2901 = n2900 ^ n2899 ;
  assign n2938 = n2902 ^ n2901 ;
  assign n2939 = n2908 & ~n2938 ;
  assign n2940 = n2939 ^ n2907 ;
  assign n2935 = n2906 ^ n2904 ;
  assign n2936 = ~n2905 & n2935 ;
  assign n2937 = n2936 ^ n2906 ;
  assign n2941 = n2940 ^ n2937 ;
  assign n2932 = n2900 ^ n2898 ;
  assign n2933 = ~n2899 & n2932 ;
  assign n2934 = n2933 ^ n2900 ;
  assign n2942 = n2941 ^ n2934 ;
  assign n2910 = x529 ^ x81 ;
  assign n2909 = n2908 ^ n2901 ;
  assign n2911 = n2910 ^ n2909 ;
  assign n2892 = x535 ^ x87 ;
  assign n2891 = x534 ^ x86 ;
  assign n2893 = n2892 ^ n2891 ;
  assign n2890 = x536 ^ x88 ;
  assign n2894 = n2893 ^ n2890 ;
  assign n2889 = x530 ^ x82 ;
  assign n2895 = n2894 ^ n2889 ;
  assign n2886 = x532 ^ x84 ;
  assign n2885 = x531 ^ x83 ;
  assign n2887 = n2886 ^ n2885 ;
  assign n2884 = x533 ^ x85 ;
  assign n2888 = n2887 ^ n2884 ;
  assign n2896 = n2895 ^ n2888 ;
  assign n2929 = n2909 ^ n2896 ;
  assign n2930 = n2911 & ~n2929 ;
  assign n2931 = n2930 ^ n2910 ;
  assign n2943 = n2942 ^ n2931 ;
  assign n2924 = n2889 ^ n2888 ;
  assign n2925 = n2895 & ~n2924 ;
  assign n2926 = n2925 ^ n2894 ;
  assign n2921 = n2891 ^ n2890 ;
  assign n2922 = n2893 & ~n2921 ;
  assign n2923 = n2922 ^ n2892 ;
  assign n2927 = n2926 ^ n2923 ;
  assign n2918 = n2885 ^ n2884 ;
  assign n2919 = n2887 & ~n2918 ;
  assign n2920 = n2919 ^ n2886 ;
  assign n2928 = n2927 ^ n2920 ;
  assign n2956 = n2931 ^ n2928 ;
  assign n2957 = n2943 & ~n2956 ;
  assign n2958 = n2957 ^ n2942 ;
  assign n2953 = n2937 ^ n2934 ;
  assign n2954 = n2941 & ~n2953 ;
  assign n2955 = n2954 ^ n2940 ;
  assign n2959 = n2958 ^ n2955 ;
  assign n2950 = n2923 ^ n2920 ;
  assign n2951 = n2927 & ~n2950 ;
  assign n2952 = n2951 ^ n2926 ;
  assign n2966 = n2955 ^ n2952 ;
  assign n2967 = n2959 & ~n2966 ;
  assign n2968 = n2967 ^ n2958 ;
  assign n2960 = n2959 ^ n2952 ;
  assign n2944 = n2943 ^ n2928 ;
  assign n2912 = n2911 ^ n2896 ;
  assign n2883 = x513 ^ x65 ;
  assign n2913 = n2912 ^ n2883 ;
  assign n2840 = x517 ^ x69 ;
  assign n2839 = x516 ^ x68 ;
  assign n2841 = n2840 ^ n2839 ;
  assign n2838 = x518 ^ x70 ;
  assign n2842 = n2841 ^ n2838 ;
  assign n2834 = x520 ^ x72 ;
  assign n2833 = x519 ^ x71 ;
  assign n2835 = n2834 ^ n2833 ;
  assign n2832 = x521 ^ x73 ;
  assign n2836 = n2835 ^ n2832 ;
  assign n2831 = x515 ^ x67 ;
  assign n2837 = n2836 ^ n2831 ;
  assign n2843 = n2842 ^ n2837 ;
  assign n2826 = x524 ^ x76 ;
  assign n2825 = x523 ^ x75 ;
  assign n2827 = n2826 ^ n2825 ;
  assign n2824 = x525 ^ x77 ;
  assign n2828 = n2827 ^ n2824 ;
  assign n2820 = x527 ^ x79 ;
  assign n2819 = x526 ^ x78 ;
  assign n2821 = n2820 ^ n2819 ;
  assign n2818 = x528 ^ x80 ;
  assign n2822 = n2821 ^ n2818 ;
  assign n2817 = x522 ^ x74 ;
  assign n2823 = n2822 ^ n2817 ;
  assign n2829 = n2828 ^ n2823 ;
  assign n2816 = x514 ^ x66 ;
  assign n2830 = n2829 ^ n2816 ;
  assign n2914 = n2843 ^ n2830 ;
  assign n2915 = n2914 ^ n2883 ;
  assign n2916 = n2913 & ~n2915 ;
  assign n2917 = n2916 ^ n2912 ;
  assign n2945 = n2944 ^ n2917 ;
  assign n2865 = n2833 ^ n2832 ;
  assign n2866 = n2835 & ~n2865 ;
  assign n2867 = n2866 ^ n2834 ;
  assign n2862 = n2842 ^ n2836 ;
  assign n2863 = ~n2837 & n2862 ;
  assign n2864 = n2863 ^ n2842 ;
  assign n2868 = n2867 ^ n2864 ;
  assign n2859 = n2839 ^ n2838 ;
  assign n2860 = n2841 & ~n2859 ;
  assign n2861 = n2860 ^ n2840 ;
  assign n2869 = n2868 ^ n2861 ;
  assign n2853 = n2828 ^ n2822 ;
  assign n2854 = ~n2823 & n2853 ;
  assign n2855 = n2854 ^ n2828 ;
  assign n2850 = n2819 ^ n2818 ;
  assign n2851 = n2821 & ~n2850 ;
  assign n2852 = n2851 ^ n2820 ;
  assign n2856 = n2855 ^ n2852 ;
  assign n2847 = n2825 ^ n2824 ;
  assign n2848 = n2827 & ~n2847 ;
  assign n2849 = n2848 ^ n2826 ;
  assign n2857 = n2856 ^ n2849 ;
  assign n2844 = n2843 ^ n2816 ;
  assign n2845 = n2830 & ~n2844 ;
  assign n2846 = n2845 ^ n2829 ;
  assign n2858 = n2857 ^ n2846 ;
  assign n2946 = n2869 ^ n2858 ;
  assign n2947 = n2946 ^ n2944 ;
  assign n2948 = n2945 & ~n2947 ;
  assign n2949 = n2948 ^ n2917 ;
  assign n2961 = n2960 ^ n2949 ;
  assign n2877 = n2864 ^ n2861 ;
  assign n2878 = n2868 & ~n2877 ;
  assign n2879 = n2878 ^ n2867 ;
  assign n2873 = n2852 ^ n2849 ;
  assign n2874 = n2856 & ~n2873 ;
  assign n2875 = n2874 ^ n2855 ;
  assign n2870 = n2869 ^ n2846 ;
  assign n2871 = n2858 & ~n2870 ;
  assign n2872 = n2871 ^ n2857 ;
  assign n2876 = n2875 ^ n2872 ;
  assign n2962 = n2879 ^ n2876 ;
  assign n2963 = n2962 ^ n2949 ;
  assign n2964 = n2961 & ~n2963 ;
  assign n2965 = n2964 ^ n2960 ;
  assign n2969 = n2968 ^ n2965 ;
  assign n2880 = n2879 ^ n2875 ;
  assign n2881 = ~n2876 & n2880 ;
  assign n2882 = n2881 ^ n2879 ;
  assign n2970 = n2969 ^ n2882 ;
  assign n2971 = n2946 ^ n2945 ;
  assign n2972 = n2914 ^ n2913 ;
  assign n2973 = x512 ^ x64 ;
  assign n2974 = n2972 & n2973 ;
  assign n2975 = n2971 & n2974 ;
  assign n2976 = n2962 ^ n2961 ;
  assign n2977 = n2975 & n2976 ;
  assign n2978 = n2970 & n2977 ;
  assign n2979 = n2965 ^ n2882 ;
  assign n2980 = n2969 & ~n2979 ;
  assign n2981 = n2980 ^ n2968 ;
  assign n2982 = n2978 & n2981 ;
  assign n2983 = ~n2815 & ~n2982 ;
  assign n2984 = n2983 ^ n2815 ;
  assign n2985 = ~n2813 & n2984 ;
  assign n3080 = x543 ^ x63 ;
  assign n3078 = x542 ^ x62 ;
  assign n3077 = x541 ^ x61 ;
  assign n3079 = n3078 ^ n3077 ;
  assign n3081 = n3080 ^ n3079 ;
  assign n3076 = x537 ^ x57 ;
  assign n3082 = n3081 ^ n3076 ;
  assign n3074 = x540 ^ x60 ;
  assign n3072 = x539 ^ x59 ;
  assign n3071 = x538 ^ x58 ;
  assign n3073 = n3072 ^ n3071 ;
  assign n3075 = n3074 ^ n3073 ;
  assign n3112 = n3076 ^ n3075 ;
  assign n3113 = n3082 & ~n3112 ;
  assign n3114 = n3113 ^ n3081 ;
  assign n3109 = n3080 ^ n3078 ;
  assign n3110 = ~n3079 & n3109 ;
  assign n3111 = n3110 ^ n3080 ;
  assign n3115 = n3114 ^ n3111 ;
  assign n3106 = n3074 ^ n3072 ;
  assign n3107 = ~n3073 & n3106 ;
  assign n3108 = n3107 ^ n3074 ;
  assign n3116 = n3115 ^ n3108 ;
  assign n3084 = x529 ^ x49 ;
  assign n3083 = n3082 ^ n3075 ;
  assign n3085 = n3084 ^ n3083 ;
  assign n3066 = x535 ^ x55 ;
  assign n3065 = x534 ^ x54 ;
  assign n3067 = n3066 ^ n3065 ;
  assign n3064 = x536 ^ x56 ;
  assign n3068 = n3067 ^ n3064 ;
  assign n3063 = x530 ^ x50 ;
  assign n3069 = n3068 ^ n3063 ;
  assign n3060 = x532 ^ x52 ;
  assign n3059 = x531 ^ x51 ;
  assign n3061 = n3060 ^ n3059 ;
  assign n3058 = x533 ^ x53 ;
  assign n3062 = n3061 ^ n3058 ;
  assign n3070 = n3069 ^ n3062 ;
  assign n3103 = n3083 ^ n3070 ;
  assign n3104 = n3085 & ~n3103 ;
  assign n3105 = n3104 ^ n3084 ;
  assign n3117 = n3116 ^ n3105 ;
  assign n3098 = n3063 ^ n3062 ;
  assign n3099 = n3069 & ~n3098 ;
  assign n3100 = n3099 ^ n3068 ;
  assign n3095 = n3065 ^ n3064 ;
  assign n3096 = n3067 & ~n3095 ;
  assign n3097 = n3096 ^ n3066 ;
  assign n3101 = n3100 ^ n3097 ;
  assign n3092 = n3059 ^ n3058 ;
  assign n3093 = n3061 & ~n3092 ;
  assign n3094 = n3093 ^ n3060 ;
  assign n3102 = n3101 ^ n3094 ;
  assign n3130 = n3105 ^ n3102 ;
  assign n3131 = n3117 & ~n3130 ;
  assign n3132 = n3131 ^ n3116 ;
  assign n3127 = n3111 ^ n3108 ;
  assign n3128 = n3115 & ~n3127 ;
  assign n3129 = n3128 ^ n3114 ;
  assign n3133 = n3132 ^ n3129 ;
  assign n3124 = n3097 ^ n3094 ;
  assign n3125 = n3101 & ~n3124 ;
  assign n3126 = n3125 ^ n3100 ;
  assign n3140 = n3129 ^ n3126 ;
  assign n3141 = n3133 & ~n3140 ;
  assign n3142 = n3141 ^ n3132 ;
  assign n3134 = n3133 ^ n3126 ;
  assign n3118 = n3117 ^ n3102 ;
  assign n3086 = n3085 ^ n3070 ;
  assign n3057 = x513 ^ x33 ;
  assign n3087 = n3086 ^ n3057 ;
  assign n3014 = x517 ^ x37 ;
  assign n3013 = x516 ^ x36 ;
  assign n3015 = n3014 ^ n3013 ;
  assign n3012 = x518 ^ x38 ;
  assign n3016 = n3015 ^ n3012 ;
  assign n3008 = x520 ^ x40 ;
  assign n3007 = x519 ^ x39 ;
  assign n3009 = n3008 ^ n3007 ;
  assign n3006 = x521 ^ x41 ;
  assign n3010 = n3009 ^ n3006 ;
  assign n3005 = x515 ^ x35 ;
  assign n3011 = n3010 ^ n3005 ;
  assign n3017 = n3016 ^ n3011 ;
  assign n3000 = x524 ^ x44 ;
  assign n2999 = x523 ^ x43 ;
  assign n3001 = n3000 ^ n2999 ;
  assign n2998 = x525 ^ x45 ;
  assign n3002 = n3001 ^ n2998 ;
  assign n2994 = x527 ^ x47 ;
  assign n2993 = x526 ^ x46 ;
  assign n2995 = n2994 ^ n2993 ;
  assign n2992 = x528 ^ x48 ;
  assign n2996 = n2995 ^ n2992 ;
  assign n2991 = x522 ^ x42 ;
  assign n2997 = n2996 ^ n2991 ;
  assign n3003 = n3002 ^ n2997 ;
  assign n2990 = x514 ^ x34 ;
  assign n3004 = n3003 ^ n2990 ;
  assign n3088 = n3017 ^ n3004 ;
  assign n3089 = n3088 ^ n3057 ;
  assign n3090 = n3087 & ~n3089 ;
  assign n3091 = n3090 ^ n3086 ;
  assign n3119 = n3118 ^ n3091 ;
  assign n3039 = n3007 ^ n3006 ;
  assign n3040 = n3009 & ~n3039 ;
  assign n3041 = n3040 ^ n3008 ;
  assign n3036 = n3016 ^ n3010 ;
  assign n3037 = ~n3011 & n3036 ;
  assign n3038 = n3037 ^ n3016 ;
  assign n3042 = n3041 ^ n3038 ;
  assign n3033 = n3013 ^ n3012 ;
  assign n3034 = n3015 & ~n3033 ;
  assign n3035 = n3034 ^ n3014 ;
  assign n3043 = n3042 ^ n3035 ;
  assign n3027 = n3002 ^ n2996 ;
  assign n3028 = ~n2997 & n3027 ;
  assign n3029 = n3028 ^ n3002 ;
  assign n3024 = n2993 ^ n2992 ;
  assign n3025 = n2995 & ~n3024 ;
  assign n3026 = n3025 ^ n2994 ;
  assign n3030 = n3029 ^ n3026 ;
  assign n3021 = n2999 ^ n2998 ;
  assign n3022 = n3001 & ~n3021 ;
  assign n3023 = n3022 ^ n3000 ;
  assign n3031 = n3030 ^ n3023 ;
  assign n3018 = n3017 ^ n2990 ;
  assign n3019 = n3004 & ~n3018 ;
  assign n3020 = n3019 ^ n3003 ;
  assign n3032 = n3031 ^ n3020 ;
  assign n3120 = n3043 ^ n3032 ;
  assign n3121 = n3120 ^ n3118 ;
  assign n3122 = n3119 & ~n3121 ;
  assign n3123 = n3122 ^ n3091 ;
  assign n3135 = n3134 ^ n3123 ;
  assign n3051 = n3038 ^ n3035 ;
  assign n3052 = n3042 & ~n3051 ;
  assign n3053 = n3052 ^ n3041 ;
  assign n3047 = n3026 ^ n3023 ;
  assign n3048 = n3030 & ~n3047 ;
  assign n3049 = n3048 ^ n3029 ;
  assign n3044 = n3043 ^ n3020 ;
  assign n3045 = n3032 & ~n3044 ;
  assign n3046 = n3045 ^ n3031 ;
  assign n3050 = n3049 ^ n3046 ;
  assign n3136 = n3053 ^ n3050 ;
  assign n3137 = n3136 ^ n3123 ;
  assign n3138 = n3135 & ~n3137 ;
  assign n3139 = n3138 ^ n3134 ;
  assign n3143 = n3142 ^ n3139 ;
  assign n3054 = n3053 ^ n3049 ;
  assign n3055 = ~n3050 & n3054 ;
  assign n3056 = n3055 ^ n3053 ;
  assign n3144 = n3143 ^ n3056 ;
  assign n3145 = n3120 ^ n3119 ;
  assign n3146 = n3088 ^ n3087 ;
  assign n3147 = x512 ^ x32 ;
  assign n3148 = n3146 & n3147 ;
  assign n3149 = n3145 & n3148 ;
  assign n3150 = n3136 ^ n3135 ;
  assign n3151 = n3149 & n3150 ;
  assign n3152 = n3144 & n3151 ;
  assign n3153 = n3139 ^ n3056 ;
  assign n3154 = n3143 & ~n3153 ;
  assign n3155 = n3154 ^ n3142 ;
  assign n3156 = n3152 & n3155 ;
  assign n3157 = ~n2985 & ~n3156 ;
  assign n3158 = n3157 ^ n2985 ;
  assign n2986 = n2984 ^ n2813 ;
  assign n2987 = n2986 ^ n2985 ;
  assign n2988 = n2811 & ~n2987 ;
  assign n3159 = n2988 ^ n2987 ;
  assign n3160 = ~n3158 & n3159 ;
  assign n2989 = n2988 ^ n2811 ;
  assign n3162 = n3160 ^ n2989 ;
  assign n3161 = ~n2989 & n3160 ;
  assign n3163 = n3162 ^ n3161 ;
  assign n3337 = n3163 ^ n2989 ;
  assign n3164 = n3163 ^ n3160 ;
  assign n3165 = n3159 ^ n3158 ;
  assign n3166 = n3165 ^ n3160 ;
  assign n3256 = x541 ^ x29 ;
  assign n3255 = x542 ^ x30 ;
  assign n3257 = n3256 ^ n3255 ;
  assign n3254 = x543 ^ x31 ;
  assign n3289 = n3255 ^ n3254 ;
  assign n3290 = n3257 & ~n3289 ;
  assign n3291 = n3290 ^ n3256 ;
  assign n3259 = x537 ^ x25 ;
  assign n3258 = n3257 ^ n3254 ;
  assign n3260 = n3259 ^ n3258 ;
  assign n3251 = x539 ^ x27 ;
  assign n3250 = x538 ^ x26 ;
  assign n3252 = n3251 ^ n3250 ;
  assign n3249 = x540 ^ x28 ;
  assign n3253 = n3252 ^ n3249 ;
  assign n3286 = n3258 ^ n3253 ;
  assign n3287 = n3260 & ~n3286 ;
  assign n3288 = n3287 ^ n3259 ;
  assign n3292 = n3291 ^ n3288 ;
  assign n3283 = n3250 ^ n3249 ;
  assign n3284 = n3252 & ~n3283 ;
  assign n3285 = n3284 ^ n3251 ;
  assign n3307 = n3288 ^ n3285 ;
  assign n3308 = n3292 & ~n3307 ;
  assign n3309 = n3308 ^ n3291 ;
  assign n3293 = n3292 ^ n3285 ;
  assign n3261 = n3260 ^ n3253 ;
  assign n3248 = x529 ^ x17 ;
  assign n3262 = n3261 ^ n3248 ;
  assign n3243 = x535 ^ x23 ;
  assign n3242 = x534 ^ x22 ;
  assign n3244 = n3243 ^ n3242 ;
  assign n3241 = x536 ^ x24 ;
  assign n3245 = n3244 ^ n3241 ;
  assign n3240 = x530 ^ x18 ;
  assign n3246 = n3245 ^ n3240 ;
  assign n3237 = x532 ^ x20 ;
  assign n3236 = x531 ^ x19 ;
  assign n3238 = n3237 ^ n3236 ;
  assign n3235 = x533 ^ x21 ;
  assign n3239 = n3238 ^ n3235 ;
  assign n3247 = n3246 ^ n3239 ;
  assign n3280 = n3248 ^ n3247 ;
  assign n3281 = n3262 & ~n3280 ;
  assign n3282 = n3281 ^ n3261 ;
  assign n3294 = n3293 ^ n3282 ;
  assign n3275 = n3240 ^ n3239 ;
  assign n3276 = n3246 & ~n3275 ;
  assign n3277 = n3276 ^ n3245 ;
  assign n3272 = n3242 ^ n3241 ;
  assign n3273 = n3244 & ~n3272 ;
  assign n3274 = n3273 ^ n3243 ;
  assign n3278 = n3277 ^ n3274 ;
  assign n3269 = n3236 ^ n3235 ;
  assign n3270 = n3238 & ~n3269 ;
  assign n3271 = n3270 ^ n3237 ;
  assign n3279 = n3278 ^ n3271 ;
  assign n3304 = n3293 ^ n3279 ;
  assign n3305 = n3294 & ~n3304 ;
  assign n3306 = n3305 ^ n3282 ;
  assign n3310 = n3309 ^ n3306 ;
  assign n3301 = n3274 ^ n3271 ;
  assign n3302 = n3278 & ~n3301 ;
  assign n3303 = n3302 ^ n3277 ;
  assign n3317 = n3306 ^ n3303 ;
  assign n3318 = n3310 & ~n3317 ;
  assign n3319 = n3318 ^ n3309 ;
  assign n3311 = n3310 ^ n3303 ;
  assign n3295 = n3294 ^ n3279 ;
  assign n3263 = n3262 ^ n3247 ;
  assign n3234 = x513 ^ x1 ;
  assign n3264 = n3263 ^ n3234 ;
  assign n3204 = x517 ^ x5 ;
  assign n3203 = x516 ^ x4 ;
  assign n3205 = n3204 ^ n3203 ;
  assign n3202 = x518 ^ x6 ;
  assign n3206 = n3205 ^ n3202 ;
  assign n3198 = x520 ^ x8 ;
  assign n3197 = x519 ^ x7 ;
  assign n3199 = n3198 ^ n3197 ;
  assign n3196 = x521 ^ x9 ;
  assign n3200 = n3199 ^ n3196 ;
  assign n3195 = x515 ^ x3 ;
  assign n3201 = n3200 ^ n3195 ;
  assign n3207 = n3206 ^ n3201 ;
  assign n3193 = x514 ^ x2 ;
  assign n3179 = x524 ^ x12 ;
  assign n3178 = x523 ^ x11 ;
  assign n3180 = n3179 ^ n3178 ;
  assign n3177 = x525 ^ x13 ;
  assign n3181 = n3180 ^ n3177 ;
  assign n3170 = x528 ^ x16 ;
  assign n3168 = x527 ^ x15 ;
  assign n3167 = x526 ^ x14 ;
  assign n3169 = n3168 ^ n3167 ;
  assign n3175 = n3170 ^ n3169 ;
  assign n3174 = x522 ^ x10 ;
  assign n3176 = n3175 ^ n3174 ;
  assign n3192 = n3181 ^ n3176 ;
  assign n3194 = n3193 ^ n3192 ;
  assign n3265 = n3207 ^ n3194 ;
  assign n3266 = n3265 ^ n3234 ;
  assign n3267 = n3264 & ~n3266 ;
  assign n3268 = n3267 ^ n3263 ;
  assign n3296 = n3295 ^ n3268 ;
  assign n3219 = n3197 ^ n3196 ;
  assign n3220 = n3199 & ~n3219 ;
  assign n3221 = n3220 ^ n3198 ;
  assign n3216 = n3206 ^ n3200 ;
  assign n3217 = ~n3201 & n3216 ;
  assign n3218 = n3217 ^ n3206 ;
  assign n3222 = n3221 ^ n3218 ;
  assign n3213 = n3203 ^ n3202 ;
  assign n3214 = n3205 & ~n3213 ;
  assign n3215 = n3214 ^ n3204 ;
  assign n3223 = n3222 ^ n3215 ;
  assign n3186 = n3178 ^ n3177 ;
  assign n3187 = n3180 & ~n3186 ;
  assign n3188 = n3187 ^ n3179 ;
  assign n3182 = n3181 ^ n3174 ;
  assign n3183 = n3176 & ~n3182 ;
  assign n3184 = n3183 ^ n3175 ;
  assign n3171 = n3170 ^ n3167 ;
  assign n3172 = n3169 & ~n3171 ;
  assign n3173 = n3172 ^ n3168 ;
  assign n3185 = n3184 ^ n3173 ;
  assign n3211 = n3188 ^ n3185 ;
  assign n3208 = n3207 ^ n3192 ;
  assign n3209 = n3194 & ~n3208 ;
  assign n3210 = n3209 ^ n3193 ;
  assign n3212 = n3211 ^ n3210 ;
  assign n3297 = n3223 ^ n3212 ;
  assign n3298 = n3297 ^ n3295 ;
  assign n3299 = n3296 & ~n3298 ;
  assign n3300 = n3299 ^ n3268 ;
  assign n3312 = n3311 ^ n3300 ;
  assign n3228 = n3218 ^ n3215 ;
  assign n3229 = n3222 & ~n3228 ;
  assign n3230 = n3229 ^ n3221 ;
  assign n3224 = n3223 ^ n3211 ;
  assign n3225 = n3212 & ~n3224 ;
  assign n3226 = n3225 ^ n3210 ;
  assign n3189 = n3188 ^ n3173 ;
  assign n3190 = n3185 & ~n3189 ;
  assign n3191 = n3190 ^ n3184 ;
  assign n3227 = n3226 ^ n3191 ;
  assign n3313 = n3230 ^ n3227 ;
  assign n3314 = n3313 ^ n3300 ;
  assign n3315 = n3312 & ~n3314 ;
  assign n3316 = n3315 ^ n3311 ;
  assign n3320 = n3319 ^ n3316 ;
  assign n3231 = n3230 ^ n3191 ;
  assign n3232 = n3227 & ~n3231 ;
  assign n3233 = n3232 ^ n3226 ;
  assign n3321 = n3320 ^ n3233 ;
  assign n3322 = n3297 ^ n3296 ;
  assign n3323 = n3265 ^ n3264 ;
  assign n3324 = x512 ^ x0 ;
  assign n3325 = n3323 & n3324 ;
  assign n3326 = n3322 & n3325 ;
  assign n3327 = n3313 ^ n3312 ;
  assign n3328 = n3326 & n3327 ;
  assign n3329 = n3321 & n3328 ;
  assign n3330 = n3319 ^ n3233 ;
  assign n3331 = ~n3320 & n3330 ;
  assign n3332 = n3331 ^ n3233 ;
  assign n3333 = n3329 & n3332 ;
  assign n3334 = ~n3166 & ~n3333 ;
  assign n3335 = n3334 ^ n3166 ;
  assign n3336 = n3164 & ~n3335 ;
  assign n3338 = n3337 ^ n3336 ;
  assign n3343 = n710 ^ n707 ;
  assign n3344 = n3343 ^ n878 ;
  assign n3345 = n878 & ~n3343 ;
  assign n3346 = n3345 ^ n881 ;
  assign n3347 = n3345 ^ n3344 ;
  assign n3349 = n706 ^ n695 ;
  assign n3348 = n876 ^ n875 ;
  assign n3350 = n3349 ^ n3348 ;
  assign n3352 = n874 ^ n869 ;
  assign n3351 = n694 ^ n689 ;
  assign n3353 = n3352 ^ n3351 ;
  assign n3357 = n693 ^ n690 ;
  assign n3354 = n692 ^ n691 ;
  assign n3355 = n872 ^ n871 ;
  assign n3356 = ~n3354 & n3355 ;
  assign n3358 = n3357 ^ n3356 ;
  assign n3359 = n873 ^ n870 ;
  assign n3360 = n3359 ^ n3356 ;
  assign n3361 = ~n3358 & ~n3360 ;
  assign n3362 = n3361 ^ n3357 ;
  assign n3363 = n3362 ^ n3352 ;
  assign n3364 = ~n3353 & n3363 ;
  assign n3365 = n3364 ^ n3351 ;
  assign n3366 = n3365 ^ n3349 ;
  assign n3367 = ~n3350 & n3366 ;
  assign n3368 = n3367 ^ n3349 ;
  assign n3369 = ~n3347 & ~n3368 ;
  assign n3370 = ~n3346 & ~n3369 ;
  assign n3371 = n1051 & ~n3370 ;
  assign n3372 = n3344 & ~n3371 ;
  assign n3415 = n3372 ^ n3343 ;
  assign n3375 = n1048 ^ n1045 ;
  assign n3342 = n878 ^ n711 ;
  assign n3373 = n3372 ^ n3342 ;
  assign n3374 = n3373 ^ n711 ;
  assign n3376 = n3375 ^ n3374 ;
  assign n3379 = n1044 ^ n1037 ;
  assign n3377 = n3350 & ~n3371 ;
  assign n3378 = n3377 ^ n3348 ;
  assign n3380 = n3379 ^ n3378 ;
  assign n3382 = n3353 & ~n3371 ;
  assign n3383 = n3382 ^ n3353 ;
  assign n3384 = n3383 ^ n3351 ;
  assign n3381 = n1043 ^ n1042 ;
  assign n3385 = n3384 ^ n3381 ;
  assign n3387 = n3359 ^ n3357 ;
  assign n3388 = n3371 & n3387 ;
  assign n3389 = n3388 ^ n3387 ;
  assign n3390 = n3389 ^ n3359 ;
  assign n3386 = n1041 ^ n1038 ;
  assign n3391 = n3390 ^ n3386 ;
  assign n3392 = n1040 ^ n1039 ;
  assign n3393 = n3355 ^ n3354 ;
  assign n3394 = ~n3371 & n3393 ;
  assign n3395 = n3394 ^ n3393 ;
  assign n3396 = n3395 ^ n3354 ;
  assign n3397 = n3392 & ~n3396 ;
  assign n3398 = n3397 ^ n3390 ;
  assign n3399 = ~n3391 & ~n3398 ;
  assign n3400 = n3399 ^ n3390 ;
  assign n3401 = n3400 ^ n3384 ;
  assign n3402 = ~n3385 & n3401 ;
  assign n3403 = n3402 ^ n3384 ;
  assign n3404 = n3403 ^ n3379 ;
  assign n3405 = ~n3380 & ~n3404 ;
  assign n3406 = n3405 ^ n3379 ;
  assign n3407 = n3406 ^ n3374 ;
  assign n3408 = ~n3376 & n3407 ;
  assign n3409 = n3408 ^ n3375 ;
  assign n3410 = n3409 ^ n1049 ;
  assign n3411 = ~n1057 & ~n3410 ;
  assign n3412 = n3411 ^ n882 ;
  assign n3413 = n3376 & n3412 ;
  assign n3414 = n3413 ^ n3374 ;
  assign n3416 = n3415 ^ n3414 ;
  assign n3417 = n3414 & ~n3415 ;
  assign n3418 = n3417 ^ n1053 ;
  assign n3419 = n3417 ^ n3416 ;
  assign n3421 = n3380 & n3412 ;
  assign n3422 = n3421 ^ n3378 ;
  assign n3420 = n3377 ^ n3349 ;
  assign n3423 = n3422 ^ n3420 ;
  assign n3425 = n3385 & n3412 ;
  assign n3426 = n3425 ^ n3385 ;
  assign n3427 = n3426 ^ n3381 ;
  assign n3424 = n3382 ^ n3351 ;
  assign n3428 = n3427 ^ n3424 ;
  assign n3430 = n3391 & n3412 ;
  assign n3431 = n3430 ^ n3391 ;
  assign n3432 = n3431 ^ n3386 ;
  assign n3429 = n3388 ^ n3359 ;
  assign n3433 = n3432 ^ n3429 ;
  assign n3434 = n3394 ^ n3354 ;
  assign n3435 = n3396 ^ n3392 ;
  assign n3436 = n3412 & n3435 ;
  assign n3437 = n3436 ^ n3435 ;
  assign n3438 = n3437 ^ n3392 ;
  assign n3439 = ~n3434 & n3438 ;
  assign n3440 = n3439 ^ n3432 ;
  assign n3441 = ~n3433 & n3440 ;
  assign n3442 = n3441 ^ n3432 ;
  assign n3443 = n3442 ^ n3424 ;
  assign n3444 = ~n3428 & ~n3443 ;
  assign n3445 = n3444 ^ n3424 ;
  assign n3446 = n3445 ^ n3422 ;
  assign n3447 = ~n3423 & ~n3446 ;
  assign n3448 = n3447 ^ n3422 ;
  assign n3449 = ~n3419 & n3448 ;
  assign n3450 = ~n3418 & ~n3449 ;
  assign n3451 = n1055 & ~n3450 ;
  assign n3452 = n3416 & ~n3451 ;
  assign n3532 = n3452 ^ n3415 ;
  assign n3455 = n1224 ^ n1221 ;
  assign n3454 = n3413 ^ n3375 ;
  assign n3456 = n3455 ^ n3454 ;
  assign n3457 = n3454 & ~n3455 ;
  assign n3458 = ~n1226 & ~n3457 ;
  assign n3460 = n1220 ^ n1213 ;
  assign n3459 = n3421 ^ n3379 ;
  assign n3461 = n3460 ^ n3459 ;
  assign n3463 = n1219 ^ n1218 ;
  assign n3462 = n3425 ^ n3381 ;
  assign n3464 = n3463 ^ n3462 ;
  assign n3466 = n3430 ^ n3386 ;
  assign n3465 = n1217 ^ n1214 ;
  assign n3467 = n3466 ^ n3465 ;
  assign n3468 = n1216 ^ n1215 ;
  assign n3469 = n3436 ^ n3392 ;
  assign n3470 = n3468 & ~n3469 ;
  assign n3471 = n3470 ^ n3466 ;
  assign n3472 = ~n3467 & ~n3471 ;
  assign n3473 = n3472 ^ n3466 ;
  assign n3474 = n3473 ^ n3462 ;
  assign n3475 = ~n3464 & ~n3474 ;
  assign n3476 = n3475 ^ n3463 ;
  assign n3477 = n3476 ^ n3460 ;
  assign n3478 = ~n3461 & n3477 ;
  assign n3479 = n3478 ^ n3460 ;
  assign n3480 = n3458 & n3479 ;
  assign n3481 = n3456 ^ n1225 ;
  assign n3482 = n3481 ^ n3457 ;
  assign n3483 = ~n1058 & n3482 ;
  assign n3484 = ~n3480 & ~n3483 ;
  assign n3485 = n3456 & ~n3484 ;
  assign n3486 = n3485 ^ n3455 ;
  assign n3453 = n3452 ^ n3414 ;
  assign n3487 = n3486 ^ n3453 ;
  assign n3490 = n3461 & n3484 ;
  assign n3491 = n3490 ^ n3459 ;
  assign n3488 = n3423 & ~n3451 ;
  assign n3489 = n3488 ^ n3422 ;
  assign n3492 = n3491 ^ n3489 ;
  assign n3495 = n3428 & ~n3451 ;
  assign n3496 = n3495 ^ n3428 ;
  assign n3497 = n3496 ^ n3424 ;
  assign n3493 = n3464 & ~n3484 ;
  assign n3494 = n3493 ^ n3463 ;
  assign n3498 = n3497 ^ n3494 ;
  assign n3502 = n3467 & ~n3484 ;
  assign n3503 = n3502 ^ n3465 ;
  assign n3499 = n3433 & ~n3451 ;
  assign n3500 = n3499 ^ n3433 ;
  assign n3501 = n3500 ^ n3429 ;
  assign n3504 = n3503 ^ n3501 ;
  assign n3505 = n3469 ^ n3468 ;
  assign n3506 = ~n3484 & n3505 ;
  assign n3507 = n3506 ^ n3468 ;
  assign n3508 = n3438 ^ n3434 ;
  assign n3509 = ~n3451 & n3508 ;
  assign n3510 = n3509 ^ n3508 ;
  assign n3511 = n3510 ^ n3434 ;
  assign n3512 = n3507 & ~n3511 ;
  assign n3513 = n3512 ^ n3503 ;
  assign n3514 = ~n3504 & n3513 ;
  assign n3515 = n3514 ^ n3503 ;
  assign n3516 = n3515 ^ n3497 ;
  assign n3517 = ~n3498 & ~n3516 ;
  assign n3518 = n3517 ^ n3497 ;
  assign n3519 = n3518 ^ n3491 ;
  assign n3520 = ~n3492 & n3519 ;
  assign n3521 = n3520 ^ n3489 ;
  assign n3522 = n3521 ^ n3486 ;
  assign n3523 = ~n3487 & n3522 ;
  assign n3524 = n3523 ^ n3453 ;
  assign n3525 = n3524 ^ n1227 ;
  assign n3526 = n1229 & n3525 ;
  assign n3527 = n3526 ^ n1056 ;
  assign n3528 = n3487 & n3527 ;
  assign n3529 = n3528 ^ n3453 ;
  assign n3530 = n3529 ^ n3486 ;
  assign n3531 = n3530 ^ n3453 ;
  assign n3533 = n3532 ^ n3531 ;
  assign n3534 = n1228 ^ n1054 ;
  assign n3536 = n3492 & n3527 ;
  assign n3537 = n3536 ^ n3492 ;
  assign n3538 = n3537 ^ n3489 ;
  assign n3535 = n3488 ^ n3420 ;
  assign n3539 = n3538 ^ n3535 ;
  assign n3543 = n3495 ^ n3424 ;
  assign n3540 = n3498 & ~n3527 ;
  assign n3541 = n3540 ^ n3498 ;
  assign n3542 = n3541 ^ n3494 ;
  assign n3544 = n3543 ^ n3542 ;
  assign n3546 = n3504 & n3527 ;
  assign n3547 = n3546 ^ n3504 ;
  assign n3548 = n3547 ^ n3501 ;
  assign n3545 = n3499 ^ n3429 ;
  assign n3549 = n3548 ^ n3545 ;
  assign n3550 = n3511 ^ n3507 ;
  assign n3551 = ~n3527 & n3550 ;
  assign n3552 = n3551 ^ n3550 ;
  assign n3553 = n3552 ^ n3507 ;
  assign n3554 = n3509 ^ n3434 ;
  assign n3555 = n3553 & ~n3554 ;
  assign n3556 = n3555 ^ n3548 ;
  assign n3557 = ~n3549 & n3556 ;
  assign n3558 = n3557 ^ n3548 ;
  assign n3559 = n3558 ^ n3542 ;
  assign n3560 = ~n3544 & n3559 ;
  assign n3561 = n3560 ^ n3542 ;
  assign n3562 = n3561 ^ n3538 ;
  assign n3563 = ~n3539 & n3562 ;
  assign n3564 = n3563 ^ n3538 ;
  assign n3565 = n3564 ^ n3532 ;
  assign n3566 = ~n3533 & ~n3565 ;
  assign n3567 = n3566 ^ n3532 ;
  assign n3568 = n3567 ^ n1228 ;
  assign n3569 = ~n3534 & n3568 ;
  assign n3570 = n3569 ^ n1054 ;
  assign n3571 = n3533 & n3570 ;
  assign n3572 = n3571 ^ n3532 ;
  assign n3605 = n3571 ^ n3531 ;
  assign n3573 = n1396 ^ n1393 ;
  assign n3574 = n3573 ^ n3529 ;
  assign n3575 = n3529 & ~n3573 ;
  assign n3576 = ~n1398 & ~n3575 ;
  assign n3578 = n3536 ^ n3489 ;
  assign n3577 = n1392 ^ n1385 ;
  assign n3579 = n3578 ^ n3577 ;
  assign n3581 = n1391 ^ n1390 ;
  assign n3580 = n3540 ^ n3494 ;
  assign n3582 = n3581 ^ n3580 ;
  assign n3584 = n1389 ^ n1386 ;
  assign n3583 = n3546 ^ n3501 ;
  assign n3585 = n3584 ^ n3583 ;
  assign n3586 = n1388 ^ n1387 ;
  assign n3587 = n3551 ^ n3507 ;
  assign n3588 = n3586 & ~n3587 ;
  assign n3589 = n3588 ^ n3584 ;
  assign n3590 = ~n3585 & n3589 ;
  assign n3591 = n3590 ^ n3584 ;
  assign n3592 = n3591 ^ n3580 ;
  assign n3593 = ~n3582 & n3592 ;
  assign n3594 = n3593 ^ n3581 ;
  assign n3595 = n3594 ^ n3578 ;
  assign n3596 = ~n3579 & ~n3595 ;
  assign n3597 = n3596 ^ n3578 ;
  assign n3598 = n3576 & ~n3597 ;
  assign n3599 = n3574 ^ n1397 ;
  assign n3600 = n3599 ^ n3575 ;
  assign n3601 = n1230 & n3600 ;
  assign n3602 = ~n3598 & ~n3601 ;
  assign n3603 = n3574 & n3602 ;
  assign n3604 = n3603 ^ n3529 ;
  assign n3606 = n3605 ^ n3604 ;
  assign n3609 = n3539 & n3570 ;
  assign n3610 = n3609 ^ n3538 ;
  assign n3607 = n3579 & ~n3602 ;
  assign n3608 = n3607 ^ n3577 ;
  assign n3611 = n3610 ^ n3608 ;
  assign n3615 = n3582 & ~n3602 ;
  assign n3616 = n3615 ^ n3581 ;
  assign n3612 = n3544 & ~n3570 ;
  assign n3613 = n3612 ^ n3544 ;
  assign n3614 = n3613 ^ n3542 ;
  assign n3617 = n3616 ^ n3614 ;
  assign n3620 = n3549 & n3570 ;
  assign n3621 = n3620 ^ n3549 ;
  assign n3622 = n3621 ^ n3545 ;
  assign n3618 = n3585 & n3602 ;
  assign n3619 = n3618 ^ n3583 ;
  assign n3623 = n3622 ^ n3619 ;
  assign n3624 = n3587 ^ n3586 ;
  assign n3625 = ~n3602 & n3624 ;
  assign n3626 = n3625 ^ n3586 ;
  assign n3627 = n3554 ^ n3553 ;
  assign n3628 = ~n3570 & n3627 ;
  assign n3629 = n3628 ^ n3627 ;
  assign n3630 = n3629 ^ n3553 ;
  assign n3631 = n3626 & ~n3630 ;
  assign n3632 = n3631 ^ n3622 ;
  assign n3633 = ~n3623 & ~n3632 ;
  assign n3634 = n3633 ^ n3622 ;
  assign n3635 = n3634 ^ n3616 ;
  assign n3636 = ~n3617 & ~n3635 ;
  assign n3637 = n3636 ^ n3616 ;
  assign n3638 = n3637 ^ n3608 ;
  assign n3639 = ~n3611 & ~n3638 ;
  assign n3640 = n3639 ^ n3610 ;
  assign n3641 = n3640 ^ n3604 ;
  assign n3642 = ~n3606 & n3641 ;
  assign n3643 = n3642 ^ n3605 ;
  assign n3644 = n3643 ^ n1399 ;
  assign n3645 = n1405 & ~n3644 ;
  assign n3646 = n3645 ^ n1403 ;
  assign n3647 = n3606 & ~n3646 ;
  assign n3648 = n3647 ^ n3605 ;
  assign n3649 = n3648 ^ n3604 ;
  assign n3650 = n3649 ^ n3605 ;
  assign n3692 = ~n3572 & n3650 ;
  assign n3693 = n1576 & n3692 ;
  assign n3651 = n3650 ^ n3572 ;
  assign n3652 = n1404 ^ n1401 ;
  assign n3656 = n3609 ^ n3535 ;
  assign n3653 = n3611 & ~n3646 ;
  assign n3654 = n3653 ^ n3611 ;
  assign n3655 = n3654 ^ n3610 ;
  assign n3657 = n3656 ^ n3655 ;
  assign n3659 = n3617 & ~n3646 ;
  assign n3660 = n3659 ^ n3617 ;
  assign n3661 = n3660 ^ n3614 ;
  assign n3658 = n3612 ^ n3542 ;
  assign n3662 = n3661 ^ n3658 ;
  assign n3666 = n3620 ^ n3545 ;
  assign n3663 = n3623 & n3646 ;
  assign n3664 = n3663 ^ n3623 ;
  assign n3665 = n3664 ^ n3619 ;
  assign n3667 = n3666 ^ n3665 ;
  assign n3668 = n3628 ^ n3553 ;
  assign n3669 = n3630 ^ n3626 ;
  assign n3670 = n3646 & n3669 ;
  assign n3671 = n3670 ^ n3669 ;
  assign n3672 = n3671 ^ n3626 ;
  assign n3673 = ~n3668 & n3672 ;
  assign n3674 = n3673 ^ n3665 ;
  assign n3675 = ~n3667 & n3674 ;
  assign n3676 = n3675 ^ n3665 ;
  assign n3677 = n3676 ^ n3661 ;
  assign n3678 = ~n3662 & n3677 ;
  assign n3679 = n3678 ^ n3661 ;
  assign n3680 = n3679 ^ n3656 ;
  assign n3681 = ~n3657 & ~n3680 ;
  assign n3682 = n3681 ^ n3656 ;
  assign n3683 = n3682 ^ n3650 ;
  assign n3684 = ~n3651 & n3683 ;
  assign n3685 = n3684 ^ n3572 ;
  assign n3686 = n3685 ^ n1401 ;
  assign n3687 = ~n3652 & ~n3686 ;
  assign n3688 = n3687 ^ n1404 ;
  assign n3689 = n3651 & ~n3688 ;
  assign n3690 = n3572 & ~n3689 ;
  assign n3808 = n3693 ^ n3690 ;
  assign n3695 = n1572 ^ n1569 ;
  assign n3696 = n3695 ^ n3648 ;
  assign n3698 = n3696 ^ n1573 ;
  assign n3697 = n3648 & ~n3695 ;
  assign n3699 = n3698 ^ n3697 ;
  assign n3700 = n1406 & n3699 ;
  assign n3701 = ~n1574 & ~n3697 ;
  assign n3703 = n1568 ^ n1561 ;
  assign n3702 = n3653 ^ n3610 ;
  assign n3704 = n3703 ^ n3702 ;
  assign n3706 = n3659 ^ n3614 ;
  assign n3705 = n1567 ^ n1566 ;
  assign n3707 = n3706 ^ n3705 ;
  assign n3709 = n1565 ^ n1562 ;
  assign n3708 = n3663 ^ n3619 ;
  assign n3710 = n3709 ^ n3708 ;
  assign n3711 = n1564 ^ n1563 ;
  assign n3712 = n3670 ^ n3626 ;
  assign n3713 = n3711 & ~n3712 ;
  assign n3714 = n3713 ^ n3709 ;
  assign n3715 = ~n3710 & n3714 ;
  assign n3716 = n3715 ^ n3709 ;
  assign n3717 = n3716 ^ n3705 ;
  assign n3718 = ~n3707 & n3717 ;
  assign n3719 = n3718 ^ n3705 ;
  assign n3720 = n3719 ^ n3703 ;
  assign n3721 = ~n3704 & n3720 ;
  assign n3722 = n3721 ^ n3703 ;
  assign n3723 = n3701 & n3722 ;
  assign n3724 = ~n3700 & ~n3723 ;
  assign n3725 = n3696 & ~n3724 ;
  assign n3726 = n3725 ^ n3695 ;
  assign n3691 = n3690 ^ n3651 ;
  assign n3694 = n3693 ^ n3691 ;
  assign n3727 = n3726 ^ n3694 ;
  assign n3730 = n3657 & ~n3688 ;
  assign n3731 = n3730 ^ n3655 ;
  assign n3728 = n3704 & ~n3724 ;
  assign n3729 = n3728 ^ n3703 ;
  assign n3732 = n3731 ^ n3729 ;
  assign n3736 = n3707 & ~n3724 ;
  assign n3737 = n3736 ^ n3705 ;
  assign n3733 = n3662 & ~n3688 ;
  assign n3734 = n3733 ^ n3662 ;
  assign n3735 = n3734 ^ n3658 ;
  assign n3738 = n3737 ^ n3735 ;
  assign n3741 = n3667 & n3688 ;
  assign n3742 = n3741 ^ n3667 ;
  assign n3743 = n3742 ^ n3665 ;
  assign n3739 = n3710 & n3724 ;
  assign n3740 = n3739 ^ n3708 ;
  assign n3744 = n3743 ^ n3740 ;
  assign n3745 = n3712 ^ n3711 ;
  assign n3746 = ~n3724 & n3745 ;
  assign n3747 = n3746 ^ n3711 ;
  assign n3748 = n3672 ^ n3668 ;
  assign n3749 = ~n3688 & n3748 ;
  assign n3750 = n3749 ^ n3748 ;
  assign n3751 = n3750 ^ n3668 ;
  assign n3752 = n3747 & ~n3751 ;
  assign n3753 = n3752 ^ n3743 ;
  assign n3754 = ~n3744 & ~n3753 ;
  assign n3755 = n3754 ^ n3743 ;
  assign n3756 = n3755 ^ n3737 ;
  assign n3757 = ~n3738 & ~n3756 ;
  assign n3758 = n3757 ^ n3737 ;
  assign n3759 = n3758 ^ n3731 ;
  assign n3760 = ~n3732 & n3759 ;
  assign n3761 = n3760 ^ n3729 ;
  assign n3762 = n3761 ^ n3726 ;
  assign n3763 = ~n3727 & ~n3762 ;
  assign n3764 = n3763 ^ n3694 ;
  assign n3765 = n3764 ^ n1577 ;
  assign n3766 = n1584 & ~n3765 ;
  assign n3767 = n3766 ^ n1575 ;
  assign n3768 = n3727 & ~n3767 ;
  assign n3769 = n3768 ^ n3694 ;
  assign n3806 = n3769 ^ n3726 ;
  assign n3807 = n3806 ^ n3694 ;
  assign n3809 = n3808 ^ n3807 ;
  assign n3810 = n1579 ^ n1578 ;
  assign n3776 = n3732 & ~n3767 ;
  assign n3812 = n3776 ^ n3732 ;
  assign n3813 = n3812 ^ n3731 ;
  assign n3811 = n3730 ^ n3656 ;
  assign n3814 = n3813 ^ n3811 ;
  assign n3781 = n3738 & ~n3767 ;
  assign n3816 = n3781 ^ n3738 ;
  assign n3817 = n3816 ^ n3735 ;
  assign n3815 = n3733 ^ n3658 ;
  assign n3818 = n3817 ^ n3815 ;
  assign n3821 = n3741 ^ n3665 ;
  assign n3784 = n3744 & n3767 ;
  assign n3819 = n3784 ^ n3744 ;
  assign n3820 = n3819 ^ n3740 ;
  assign n3822 = n3821 ^ n3820 ;
  assign n3789 = n3751 ^ n3747 ;
  assign n3790 = n3767 & n3789 ;
  assign n3823 = n3790 ^ n3789 ;
  assign n3824 = n3823 ^ n3747 ;
  assign n3825 = n3749 ^ n3668 ;
  assign n3826 = n3824 & ~n3825 ;
  assign n3827 = n3826 ^ n3820 ;
  assign n3828 = ~n3822 & n3827 ;
  assign n3829 = n3828 ^ n3820 ;
  assign n3830 = n3829 ^ n3817 ;
  assign n3831 = ~n3818 & n3830 ;
  assign n3832 = n3831 ^ n3817 ;
  assign n3833 = n3832 ^ n3813 ;
  assign n3834 = ~n3814 & n3833 ;
  assign n3835 = n3834 ^ n3813 ;
  assign n3836 = n3835 ^ n3808 ;
  assign n3837 = ~n3809 & ~n3836 ;
  assign n3838 = n3837 ^ n3808 ;
  assign n3839 = n3838 ^ n1579 ;
  assign n3840 = ~n3810 & ~n3839 ;
  assign n3841 = n3840 ^ n1578 ;
  assign n3842 = n3809 & ~n3841 ;
  assign n3889 = n3842 ^ n3808 ;
  assign n3843 = n3842 ^ n3807 ;
  assign n3341 = n1751 ^ n1748 ;
  assign n3770 = n3769 ^ n3341 ;
  assign n3772 = n3770 ^ n1752 ;
  assign n3771 = ~n3341 & n3769 ;
  assign n3773 = n3772 ^ n3771 ;
  assign n3774 = n1585 & n3773 ;
  assign n3775 = ~n1753 & ~n3771 ;
  assign n3778 = n1747 ^ n1740 ;
  assign n3777 = n3776 ^ n3731 ;
  assign n3779 = n3778 ^ n3777 ;
  assign n3782 = n3781 ^ n3735 ;
  assign n3780 = n1746 ^ n1745 ;
  assign n3783 = n3782 ^ n3780 ;
  assign n3786 = n1744 ^ n1741 ;
  assign n3785 = n3784 ^ n3740 ;
  assign n3787 = n3786 ^ n3785 ;
  assign n3788 = n1743 ^ n1742 ;
  assign n3791 = n3790 ^ n3747 ;
  assign n3792 = n3788 & ~n3791 ;
  assign n3793 = n3792 ^ n3786 ;
  assign n3794 = ~n3787 & n3793 ;
  assign n3795 = n3794 ^ n3786 ;
  assign n3796 = n3795 ^ n3780 ;
  assign n3797 = ~n3783 & n3796 ;
  assign n3798 = n3797 ^ n3780 ;
  assign n3799 = n3798 ^ n3778 ;
  assign n3800 = ~n3779 & n3799 ;
  assign n3801 = n3800 ^ n3778 ;
  assign n3802 = n3775 & n3801 ;
  assign n3803 = ~n3774 & ~n3802 ;
  assign n3804 = n3770 & ~n3803 ;
  assign n3805 = n3804 ^ n3341 ;
  assign n3844 = n3843 ^ n3805 ;
  assign n3847 = n3779 & ~n3803 ;
  assign n3848 = n3847 ^ n3778 ;
  assign n3845 = n3814 & ~n3841 ;
  assign n3846 = n3845 ^ n3813 ;
  assign n3849 = n3848 ^ n3846 ;
  assign n3853 = n3783 & ~n3803 ;
  assign n3854 = n3853 ^ n3780 ;
  assign n3850 = n3818 & ~n3841 ;
  assign n3851 = n3850 ^ n3818 ;
  assign n3852 = n3851 ^ n3815 ;
  assign n3855 = n3854 ^ n3852 ;
  assign n3858 = n3822 & n3841 ;
  assign n3859 = n3858 ^ n3822 ;
  assign n3860 = n3859 ^ n3820 ;
  assign n3856 = n3787 & n3803 ;
  assign n3857 = n3856 ^ n3785 ;
  assign n3861 = n3860 ^ n3857 ;
  assign n3862 = n3791 ^ n3788 ;
  assign n3863 = ~n3803 & n3862 ;
  assign n3864 = n3863 ^ n3788 ;
  assign n3865 = n3825 ^ n3824 ;
  assign n3866 = n3841 & n3865 ;
  assign n3867 = n3866 ^ n3865 ;
  assign n3868 = n3867 ^ n3824 ;
  assign n3869 = n3864 & ~n3868 ;
  assign n3870 = n3869 ^ n3860 ;
  assign n3871 = ~n3861 & ~n3870 ;
  assign n3872 = n3871 ^ n3860 ;
  assign n3873 = n3872 ^ n3854 ;
  assign n3874 = ~n3855 & ~n3873 ;
  assign n3875 = n3874 ^ n3854 ;
  assign n3876 = n3875 ^ n3846 ;
  assign n3877 = ~n3849 & n3876 ;
  assign n3878 = n3877 ^ n3848 ;
  assign n3879 = n3878 ^ n3805 ;
  assign n3880 = ~n3844 & ~n3879 ;
  assign n3881 = n3880 ^ n3843 ;
  assign n3882 = n3881 ^ n1754 ;
  assign n3883 = n1760 & ~n3882 ;
  assign n3884 = n3883 ^ n1583 ;
  assign n3885 = n3844 & ~n3884 ;
  assign n3886 = n3885 ^ n3843 ;
  assign n3887 = n3886 ^ n3805 ;
  assign n3888 = n3887 ^ n3843 ;
  assign n3890 = n3889 ^ n3888 ;
  assign n3891 = n1755 ^ n1581 ;
  assign n3893 = n3849 & ~n3884 ;
  assign n3894 = n3893 ^ n3849 ;
  assign n3895 = n3894 ^ n3846 ;
  assign n3892 = n3845 ^ n3811 ;
  assign n3896 = n3895 ^ n3892 ;
  assign n3898 = n3855 & ~n3884 ;
  assign n3899 = n3898 ^ n3855 ;
  assign n3900 = n3899 ^ n3852 ;
  assign n3897 = n3850 ^ n3815 ;
  assign n3901 = n3900 ^ n3897 ;
  assign n3908 = n3861 & n3884 ;
  assign n3909 = n3908 ^ n3861 ;
  assign n3910 = n3909 ^ n3857 ;
  assign n3902 = n3868 ^ n3864 ;
  assign n3903 = n3884 & n3902 ;
  assign n3904 = n3903 ^ n3902 ;
  assign n3905 = n3904 ^ n3864 ;
  assign n3906 = n3866 ^ n3824 ;
  assign n3907 = n3905 & ~n3906 ;
  assign n3911 = n3910 ^ n3907 ;
  assign n3912 = n3858 ^ n3820 ;
  assign n3913 = n3912 ^ n3907 ;
  assign n3914 = n3911 & ~n3913 ;
  assign n3915 = n3914 ^ n3907 ;
  assign n3916 = n3915 ^ n3900 ;
  assign n3917 = ~n3901 & n3916 ;
  assign n3918 = n3917 ^ n3900 ;
  assign n3919 = n3918 ^ n3895 ;
  assign n3920 = ~n3896 & n3919 ;
  assign n3921 = n3920 ^ n3895 ;
  assign n3922 = n3921 ^ n3889 ;
  assign n3923 = ~n3890 & ~n3922 ;
  assign n3924 = n3923 ^ n3889 ;
  assign n3925 = n3924 ^ n1755 ;
  assign n3926 = ~n3891 & n3925 ;
  assign n3927 = n3926 ^ n1581 ;
  assign n3928 = n3890 & n3927 ;
  assign n3929 = n3928 ^ n3889 ;
  assign n3962 = n3928 ^ n3888 ;
  assign n3930 = n1927 ^ n1924 ;
  assign n3931 = n3930 ^ n3886 ;
  assign n3933 = n3931 ^ n1928 ;
  assign n3932 = n3886 & ~n3930 ;
  assign n3934 = n3933 ^ n3932 ;
  assign n3935 = n1761 & n3934 ;
  assign n3936 = ~n1929 & ~n3932 ;
  assign n3938 = n1923 ^ n1916 ;
  assign n3937 = n3893 ^ n3846 ;
  assign n3939 = n3938 ^ n3937 ;
  assign n3941 = n3898 ^ n3852 ;
  assign n3940 = n1922 ^ n1921 ;
  assign n3942 = n3941 ^ n3940 ;
  assign n3944 = n3908 ^ n3857 ;
  assign n3943 = n1920 ^ n1917 ;
  assign n3945 = n3944 ^ n3943 ;
  assign n3946 = n1919 ^ n1918 ;
  assign n3947 = n3903 ^ n3864 ;
  assign n3948 = n3946 & ~n3947 ;
  assign n3949 = n3948 ^ n3944 ;
  assign n3950 = ~n3945 & ~n3949 ;
  assign n3951 = n3950 ^ n3944 ;
  assign n3952 = n3951 ^ n3940 ;
  assign n3953 = ~n3942 & ~n3952 ;
  assign n3954 = n3953 ^ n3940 ;
  assign n3955 = n3954 ^ n3938 ;
  assign n3956 = ~n3939 & n3955 ;
  assign n3957 = n3956 ^ n3938 ;
  assign n3958 = n3936 & n3957 ;
  assign n3959 = ~n3935 & ~n3958 ;
  assign n3960 = n3931 & ~n3959 ;
  assign n3961 = n3960 ^ n3930 ;
  assign n3963 = n3962 ^ n3961 ;
  assign n3966 = n3939 & ~n3959 ;
  assign n3967 = n3966 ^ n3938 ;
  assign n3964 = n3896 & n3927 ;
  assign n3965 = n3964 ^ n3895 ;
  assign n3968 = n3967 ^ n3965 ;
  assign n3972 = n3942 & ~n3959 ;
  assign n3973 = n3972 ^ n3940 ;
  assign n3969 = n3901 & n3927 ;
  assign n3970 = n3969 ^ n3901 ;
  assign n3971 = n3970 ^ n3897 ;
  assign n3974 = n3973 ^ n3971 ;
  assign n3977 = n3912 ^ n3910 ;
  assign n3978 = ~n3927 & n3977 ;
  assign n3979 = n3978 ^ n3977 ;
  assign n3980 = n3979 ^ n3910 ;
  assign n3975 = n3945 & ~n3959 ;
  assign n3976 = n3975 ^ n3943 ;
  assign n3981 = n3980 ^ n3976 ;
  assign n3982 = n3906 ^ n3905 ;
  assign n3983 = ~n3927 & n3982 ;
  assign n3984 = n3983 ^ n3982 ;
  assign n3985 = n3984 ^ n3905 ;
  assign n3986 = n3947 ^ n3946 ;
  assign n3987 = ~n3959 & n3986 ;
  assign n3988 = n3987 ^ n3946 ;
  assign n3989 = ~n3985 & n3988 ;
  assign n3990 = n3989 ^ n3980 ;
  assign n3991 = ~n3981 & ~n3990 ;
  assign n3992 = n3991 ^ n3980 ;
  assign n3993 = n3992 ^ n3973 ;
  assign n3994 = ~n3974 & ~n3993 ;
  assign n3995 = n3994 ^ n3973 ;
  assign n3996 = n3995 ^ n3967 ;
  assign n3997 = ~n3968 & ~n3996 ;
  assign n3998 = n3997 ^ n3965 ;
  assign n3999 = n3998 ^ n3961 ;
  assign n4000 = ~n3963 & n3999 ;
  assign n4001 = n4000 ^ n3962 ;
  assign n4002 = n4001 ^ n1930 ;
  assign n4003 = n1934 & ~n4002 ;
  assign n4004 = n4003 ^ n1759 ;
  assign n4005 = n3963 & ~n4004 ;
  assign n4006 = n4005 ^ n3962 ;
  assign n4007 = n4006 ^ n3961 ;
  assign n4008 = n4007 ^ n3962 ;
  assign n4050 = n3929 & ~n4008 ;
  assign n4009 = n4008 ^ n3929 ;
  assign n4051 = n4050 ^ n4009 ;
  assign n4052 = n1932 & n4051 ;
  assign n4010 = n1931 ^ n1757 ;
  assign n4012 = n3968 & ~n4004 ;
  assign n4013 = n4012 ^ n3968 ;
  assign n4014 = n4013 ^ n3965 ;
  assign n4011 = n3964 ^ n3892 ;
  assign n4015 = n4014 ^ n4011 ;
  assign n4017 = n3974 & ~n4004 ;
  assign n4018 = n4017 ^ n3974 ;
  assign n4019 = n4018 ^ n3971 ;
  assign n4016 = n3969 ^ n3897 ;
  assign n4020 = n4019 ^ n4016 ;
  assign n4027 = n3981 & n4004 ;
  assign n4028 = n4027 ^ n3981 ;
  assign n4029 = n4028 ^ n3976 ;
  assign n4021 = n3988 ^ n3985 ;
  assign n4022 = ~n4004 & n4021 ;
  assign n4023 = n4022 ^ n4021 ;
  assign n4024 = n4023 ^ n3985 ;
  assign n4025 = n3983 ^ n3905 ;
  assign n4026 = n4024 & ~n4025 ;
  assign n4030 = n4029 ^ n4026 ;
  assign n4031 = n3978 ^ n3910 ;
  assign n4032 = n4031 ^ n4026 ;
  assign n4033 = n4030 & ~n4032 ;
  assign n4034 = n4033 ^ n4026 ;
  assign n4035 = n4034 ^ n4019 ;
  assign n4036 = ~n4020 & n4035 ;
  assign n4037 = n4036 ^ n4019 ;
  assign n4038 = n4037 ^ n4011 ;
  assign n4039 = ~n4015 & ~n4038 ;
  assign n4040 = n4039 ^ n4011 ;
  assign n4041 = n4040 ^ n4008 ;
  assign n4042 = ~n4009 & n4041 ;
  assign n4043 = n4042 ^ n3929 ;
  assign n4044 = n4043 ^ n1757 ;
  assign n4045 = ~n4010 & ~n4044 ;
  assign n4046 = n4045 ^ n1931 ;
  assign n4047 = n4009 & ~n4046 ;
  assign n4048 = n3929 & ~n4047 ;
  assign n4168 = n4052 ^ n4048 ;
  assign n4054 = n2101 ^ n2098 ;
  assign n4055 = n4054 ^ n4006 ;
  assign n4057 = n4055 ^ n2102 ;
  assign n4056 = n4006 & ~n4054 ;
  assign n4058 = n4057 ^ n4056 ;
  assign n4059 = n1935 & n4058 ;
  assign n4060 = ~n2103 & ~n4056 ;
  assign n4062 = n2097 ^ n2090 ;
  assign n4061 = n4012 ^ n3965 ;
  assign n4063 = n4062 ^ n4061 ;
  assign n4065 = n4017 ^ n3971 ;
  assign n4064 = n2096 ^ n2095 ;
  assign n4066 = n4065 ^ n4064 ;
  assign n4068 = n4027 ^ n3976 ;
  assign n4067 = n2094 ^ n2091 ;
  assign n4069 = n4068 ^ n4067 ;
  assign n4070 = n2093 ^ n2092 ;
  assign n4071 = n4022 ^ n3985 ;
  assign n4072 = n4070 & ~n4071 ;
  assign n4073 = n4072 ^ n4068 ;
  assign n4074 = ~n4069 & ~n4073 ;
  assign n4075 = n4074 ^ n4068 ;
  assign n4076 = n4075 ^ n4064 ;
  assign n4077 = ~n4066 & ~n4076 ;
  assign n4078 = n4077 ^ n4064 ;
  assign n4079 = n4078 ^ n4062 ;
  assign n4080 = ~n4063 & n4079 ;
  assign n4081 = n4080 ^ n4062 ;
  assign n4082 = n4060 & n4081 ;
  assign n4083 = ~n4059 & ~n4082 ;
  assign n4084 = n4055 & ~n4083 ;
  assign n4085 = n4084 ^ n4054 ;
  assign n4049 = n4048 ^ n4009 ;
  assign n4053 = n4052 ^ n4049 ;
  assign n4086 = n4085 ^ n4053 ;
  assign n4089 = n4015 & ~n4046 ;
  assign n4090 = n4089 ^ n4014 ;
  assign n4087 = n4063 & ~n4083 ;
  assign n4088 = n4087 ^ n4062 ;
  assign n4091 = n4090 ^ n4088 ;
  assign n4095 = n4066 & ~n4083 ;
  assign n4096 = n4095 ^ n4064 ;
  assign n4092 = n4020 & ~n4046 ;
  assign n4093 = n4092 ^ n4020 ;
  assign n4094 = n4093 ^ n4016 ;
  assign n4097 = n4096 ^ n4094 ;
  assign n4102 = n4069 & ~n4083 ;
  assign n4103 = n4102 ^ n4067 ;
  assign n4098 = n4031 ^ n4029 ;
  assign n4099 = ~n4046 & n4098 ;
  assign n4100 = n4099 ^ n4098 ;
  assign n4101 = n4100 ^ n4031 ;
  assign n4104 = n4103 ^ n4101 ;
  assign n4105 = n4025 ^ n4024 ;
  assign n4106 = n4046 & n4105 ;
  assign n4107 = n4106 ^ n4105 ;
  assign n4108 = n4107 ^ n4024 ;
  assign n4109 = n4071 ^ n4070 ;
  assign n4110 = ~n4083 & n4109 ;
  assign n4111 = n4110 ^ n4070 ;
  assign n4112 = ~n4108 & n4111 ;
  assign n4113 = n4112 ^ n4103 ;
  assign n4114 = ~n4104 & n4113 ;
  assign n4115 = n4114 ^ n4103 ;
  assign n4116 = n4115 ^ n4096 ;
  assign n4117 = ~n4097 & n4116 ;
  assign n4118 = n4117 ^ n4096 ;
  assign n4119 = n4118 ^ n4088 ;
  assign n4120 = ~n4091 & ~n4119 ;
  assign n4121 = n4120 ^ n4090 ;
  assign n4122 = n4121 ^ n4085 ;
  assign n4123 = ~n4086 & n4122 ;
  assign n4124 = n4123 ^ n4053 ;
  assign n4125 = n4124 ^ n1933 ;
  assign n4126 = n2109 & ~n4125 ;
  assign n4127 = n4126 ^ n2104 ;
  assign n4128 = n4086 & ~n4127 ;
  assign n4129 = n4128 ^ n4053 ;
  assign n4166 = n4129 ^ n4085 ;
  assign n4167 = n4166 ^ n4053 ;
  assign n4169 = n4168 ^ n4167 ;
  assign n4170 = n2106 ^ n2105 ;
  assign n4136 = n4091 & ~n4127 ;
  assign n4172 = n4136 ^ n4091 ;
  assign n4173 = n4172 ^ n4090 ;
  assign n4171 = n4089 ^ n4011 ;
  assign n4174 = n4173 ^ n4171 ;
  assign n4141 = n4097 & ~n4127 ;
  assign n4176 = n4141 ^ n4097 ;
  assign n4177 = n4176 ^ n4094 ;
  assign n4175 = n4092 ^ n4016 ;
  assign n4178 = n4177 ^ n4175 ;
  assign n4145 = n4104 & ~n4127 ;
  assign n4183 = n4145 ^ n4104 ;
  assign n4184 = n4183 ^ n4101 ;
  assign n4179 = n4106 ^ n4024 ;
  assign n4149 = n4111 ^ n4108 ;
  assign n4150 = ~n4127 & n4149 ;
  assign n4180 = n4150 ^ n4149 ;
  assign n4181 = n4180 ^ n4108 ;
  assign n4182 = ~n4179 & n4181 ;
  assign n4185 = n4184 ^ n4182 ;
  assign n4186 = n4099 ^ n4031 ;
  assign n4187 = n4186 ^ n4182 ;
  assign n4188 = n4185 & ~n4187 ;
  assign n4189 = n4188 ^ n4182 ;
  assign n4190 = n4189 ^ n4177 ;
  assign n4191 = ~n4178 & n4190 ;
  assign n4192 = n4191 ^ n4177 ;
  assign n4193 = n4192 ^ n4173 ;
  assign n4194 = ~n4174 & n4193 ;
  assign n4195 = n4194 ^ n4173 ;
  assign n4196 = n4195 ^ n4168 ;
  assign n4197 = ~n4169 & ~n4196 ;
  assign n4198 = n4197 ^ n4168 ;
  assign n4199 = n4198 ^ n2106 ;
  assign n4200 = ~n4170 & ~n4199 ;
  assign n4201 = n4200 ^ n2105 ;
  assign n4202 = n4169 & ~n4201 ;
  assign n4250 = n4202 ^ n4168 ;
  assign n4203 = n4202 ^ n4167 ;
  assign n3340 = n2276 ^ n2273 ;
  assign n4130 = n4129 ^ n3340 ;
  assign n4132 = n4130 ^ n2277 ;
  assign n4131 = ~n3340 & n4129 ;
  assign n4133 = n4132 ^ n4131 ;
  assign n4134 = n2110 & n4133 ;
  assign n4135 = ~n2278 & ~n4131 ;
  assign n4138 = n2272 ^ n2265 ;
  assign n4137 = n4136 ^ n4090 ;
  assign n4139 = n4138 ^ n4137 ;
  assign n4142 = n4141 ^ n4094 ;
  assign n4140 = n2271 ^ n2270 ;
  assign n4143 = n4142 ^ n4140 ;
  assign n4146 = n4145 ^ n4101 ;
  assign n4144 = n2269 ^ n2266 ;
  assign n4147 = n4146 ^ n4144 ;
  assign n4148 = n2268 ^ n2267 ;
  assign n4151 = n4150 ^ n4108 ;
  assign n4152 = n4148 & ~n4151 ;
  assign n4153 = n4152 ^ n4146 ;
  assign n4154 = ~n4147 & ~n4153 ;
  assign n4155 = n4154 ^ n4146 ;
  assign n4156 = n4155 ^ n4140 ;
  assign n4157 = ~n4143 & ~n4156 ;
  assign n4158 = n4157 ^ n4140 ;
  assign n4159 = n4158 ^ n4138 ;
  assign n4160 = ~n4139 & n4159 ;
  assign n4161 = n4160 ^ n4138 ;
  assign n4162 = n4135 & n4161 ;
  assign n4163 = ~n4134 & ~n4162 ;
  assign n4164 = n4130 & ~n4163 ;
  assign n4165 = n4164 ^ n3340 ;
  assign n4204 = n4203 ^ n4165 ;
  assign n4207 = n4174 & ~n4201 ;
  assign n4208 = n4207 ^ n4173 ;
  assign n4205 = n4139 & ~n4163 ;
  assign n4206 = n4205 ^ n4138 ;
  assign n4209 = n4208 ^ n4206 ;
  assign n4213 = n4143 & ~n4163 ;
  assign n4214 = n4213 ^ n4140 ;
  assign n4210 = n4178 & ~n4201 ;
  assign n4211 = n4210 ^ n4178 ;
  assign n4212 = n4211 ^ n4175 ;
  assign n4215 = n4214 ^ n4212 ;
  assign n4218 = n4186 ^ n4184 ;
  assign n4219 = ~n4201 & n4218 ;
  assign n4220 = n4219 ^ n4218 ;
  assign n4221 = n4220 ^ n4186 ;
  assign n4216 = n4147 & ~n4163 ;
  assign n4217 = n4216 ^ n4144 ;
  assign n4222 = n4221 ^ n4217 ;
  assign n4223 = n4181 ^ n4179 ;
  assign n4224 = ~n4201 & n4223 ;
  assign n4225 = n4224 ^ n4223 ;
  assign n4226 = n4225 ^ n4179 ;
  assign n4227 = n4151 ^ n4148 ;
  assign n4228 = ~n4163 & n4227 ;
  assign n4229 = n4228 ^ n4148 ;
  assign n4230 = ~n4226 & n4229 ;
  assign n4231 = n4230 ^ n4221 ;
  assign n4232 = ~n4222 & ~n4231 ;
  assign n4233 = n4232 ^ n4221 ;
  assign n4234 = n4233 ^ n4214 ;
  assign n4235 = ~n4215 & ~n4234 ;
  assign n4236 = n4235 ^ n4214 ;
  assign n4237 = n4236 ^ n4208 ;
  assign n4238 = ~n4209 & n4237 ;
  assign n4239 = n4238 ^ n4206 ;
  assign n4240 = n4239 ^ n4165 ;
  assign n4241 = ~n4204 & ~n4240 ;
  assign n4242 = n4241 ^ n4203 ;
  assign n4243 = n4242 ^ n2279 ;
  assign n4244 = n2285 & ~n4243 ;
  assign n4245 = n4244 ^ n2281 ;
  assign n4246 = n4204 & ~n4245 ;
  assign n4247 = n4246 ^ n4203 ;
  assign n4248 = n4247 ^ n4165 ;
  assign n4249 = n4248 ^ n4203 ;
  assign n4251 = n4250 ^ n4249 ;
  assign n4252 = n2282 ^ n2108 ;
  assign n4254 = n4209 & ~n4245 ;
  assign n4255 = n4254 ^ n4209 ;
  assign n4256 = n4255 ^ n4208 ;
  assign n4253 = n4207 ^ n4171 ;
  assign n4257 = n4256 ^ n4253 ;
  assign n4259 = n4215 & ~n4245 ;
  assign n4260 = n4259 ^ n4215 ;
  assign n4261 = n4260 ^ n4212 ;
  assign n4258 = n4210 ^ n4175 ;
  assign n4262 = n4261 ^ n4258 ;
  assign n4269 = n4222 & n4245 ;
  assign n4270 = n4269 ^ n4222 ;
  assign n4271 = n4270 ^ n4217 ;
  assign n4263 = n4229 ^ n4226 ;
  assign n4264 = ~n4245 & n4263 ;
  assign n4265 = n4264 ^ n4263 ;
  assign n4266 = n4265 ^ n4226 ;
  assign n4267 = n4224 ^ n4179 ;
  assign n4268 = n4266 & ~n4267 ;
  assign n4272 = n4271 ^ n4268 ;
  assign n4273 = n4219 ^ n4186 ;
  assign n4274 = n4273 ^ n4268 ;
  assign n4275 = n4272 & ~n4274 ;
  assign n4276 = n4275 ^ n4268 ;
  assign n4277 = n4276 ^ n4261 ;
  assign n4278 = ~n4262 & n4277 ;
  assign n4279 = n4278 ^ n4261 ;
  assign n4280 = n4279 ^ n4256 ;
  assign n4281 = ~n4257 & n4280 ;
  assign n4282 = n4281 ^ n4256 ;
  assign n4283 = n4282 ^ n4250 ;
  assign n4284 = ~n4251 & ~n4283 ;
  assign n4285 = n4284 ^ n4250 ;
  assign n4286 = n4285 ^ n2282 ;
  assign n4287 = ~n4252 & n4286 ;
  assign n4288 = n4287 ^ n2108 ;
  assign n4289 = n4251 & n4288 ;
  assign n4290 = n4289 ^ n4250 ;
  assign n4323 = n4289 ^ n4249 ;
  assign n4291 = n2452 ^ n2449 ;
  assign n4292 = n4291 ^ n4247 ;
  assign n4294 = n4292 ^ n2453 ;
  assign n4293 = n4247 & ~n4291 ;
  assign n4295 = n4294 ^ n4293 ;
  assign n4296 = n2286 & n4295 ;
  assign n4297 = ~n2454 & ~n4293 ;
  assign n4299 = n2448 ^ n2441 ;
  assign n4298 = n4254 ^ n4208 ;
  assign n4300 = n4299 ^ n4298 ;
  assign n4302 = n4259 ^ n4212 ;
  assign n4301 = n2447 ^ n2446 ;
  assign n4303 = n4302 ^ n4301 ;
  assign n4305 = n4269 ^ n4217 ;
  assign n4304 = n2445 ^ n2442 ;
  assign n4306 = n4305 ^ n4304 ;
  assign n4307 = n2444 ^ n2443 ;
  assign n4308 = n4264 ^ n4226 ;
  assign n4309 = n4307 & ~n4308 ;
  assign n4310 = n4309 ^ n4305 ;
  assign n4311 = ~n4306 & ~n4310 ;
  assign n4312 = n4311 ^ n4305 ;
  assign n4313 = n4312 ^ n4301 ;
  assign n4314 = ~n4303 & ~n4313 ;
  assign n4315 = n4314 ^ n4301 ;
  assign n4316 = n4315 ^ n4299 ;
  assign n4317 = ~n4300 & n4316 ;
  assign n4318 = n4317 ^ n4299 ;
  assign n4319 = n4297 & n4318 ;
  assign n4320 = ~n4296 & ~n4319 ;
  assign n4321 = n4292 & ~n4320 ;
  assign n4322 = n4321 ^ n4291 ;
  assign n4324 = n4323 ^ n4322 ;
  assign n4327 = n4300 & ~n4320 ;
  assign n4328 = n4327 ^ n4299 ;
  assign n4325 = n4257 & n4288 ;
  assign n4326 = n4325 ^ n4256 ;
  assign n4329 = n4328 ^ n4326 ;
  assign n4333 = n4303 & ~n4320 ;
  assign n4334 = n4333 ^ n4301 ;
  assign n4330 = n4262 & n4288 ;
  assign n4331 = n4330 ^ n4262 ;
  assign n4332 = n4331 ^ n4258 ;
  assign n4335 = n4334 ^ n4332 ;
  assign n4340 = n4306 & ~n4320 ;
  assign n4341 = n4340 ^ n4304 ;
  assign n4336 = n4273 ^ n4271 ;
  assign n4337 = n4288 & n4336 ;
  assign n4338 = n4337 ^ n4336 ;
  assign n4339 = n4338 ^ n4273 ;
  assign n4342 = n4341 ^ n4339 ;
  assign n4343 = n4267 ^ n4266 ;
  assign n4344 = ~n4288 & n4343 ;
  assign n4345 = n4344 ^ n4343 ;
  assign n4346 = n4345 ^ n4266 ;
  assign n4347 = n4308 ^ n4307 ;
  assign n4348 = ~n4320 & n4347 ;
  assign n4349 = n4348 ^ n4307 ;
  assign n4350 = ~n4346 & n4349 ;
  assign n4351 = n4350 ^ n4341 ;
  assign n4352 = ~n4342 & n4351 ;
  assign n4353 = n4352 ^ n4341 ;
  assign n4354 = n4353 ^ n4334 ;
  assign n4355 = ~n4335 & n4354 ;
  assign n4356 = n4355 ^ n4334 ;
  assign n4357 = n4356 ^ n4326 ;
  assign n4358 = ~n4329 & n4357 ;
  assign n4359 = n4358 ^ n4328 ;
  assign n4360 = n4359 ^ n4322 ;
  assign n4361 = ~n4324 & ~n4360 ;
  assign n4362 = n4361 ^ n4323 ;
  assign n4363 = n4362 ^ n2455 ;
  assign n4364 = n2461 & ~n4363 ;
  assign n4365 = n4364 ^ n2457 ;
  assign n4366 = n4324 & ~n4365 ;
  assign n4367 = n4366 ^ n4323 ;
  assign n4368 = n4367 ^ n4322 ;
  assign n4369 = n4368 ^ n4323 ;
  assign n4411 = n4290 & ~n4369 ;
  assign n4370 = n4369 ^ n4290 ;
  assign n4412 = n4411 ^ n4370 ;
  assign n4413 = n2459 & n4412 ;
  assign n4371 = n2458 ^ n2284 ;
  assign n4373 = n4329 & ~n4365 ;
  assign n4374 = n4373 ^ n4329 ;
  assign n4375 = n4374 ^ n4326 ;
  assign n4372 = n4325 ^ n4253 ;
  assign n4376 = n4375 ^ n4372 ;
  assign n4378 = n4335 & ~n4365 ;
  assign n4379 = n4378 ^ n4335 ;
  assign n4380 = n4379 ^ n4332 ;
  assign n4377 = n4330 ^ n4258 ;
  assign n4381 = n4380 ^ n4377 ;
  assign n4388 = n4342 & ~n4365 ;
  assign n4389 = n4388 ^ n4342 ;
  assign n4390 = n4389 ^ n4339 ;
  assign n4382 = n4344 ^ n4266 ;
  assign n4383 = n4349 ^ n4346 ;
  assign n4384 = ~n4365 & n4383 ;
  assign n4385 = n4384 ^ n4383 ;
  assign n4386 = n4385 ^ n4346 ;
  assign n4387 = ~n4382 & n4386 ;
  assign n4391 = n4390 ^ n4387 ;
  assign n4392 = n4337 ^ n4273 ;
  assign n4393 = n4392 ^ n4387 ;
  assign n4394 = n4391 & ~n4393 ;
  assign n4395 = n4394 ^ n4387 ;
  assign n4396 = n4395 ^ n4380 ;
  assign n4397 = ~n4381 & n4396 ;
  assign n4398 = n4397 ^ n4380 ;
  assign n4399 = n4398 ^ n4372 ;
  assign n4400 = ~n4376 & ~n4399 ;
  assign n4401 = n4400 ^ n4372 ;
  assign n4402 = n4401 ^ n4369 ;
  assign n4403 = ~n4370 & n4402 ;
  assign n4404 = n4403 ^ n4290 ;
  assign n4405 = n4404 ^ n2284 ;
  assign n4406 = ~n4371 & ~n4405 ;
  assign n4407 = n4406 ^ n2458 ;
  assign n4408 = n4370 & ~n4407 ;
  assign n4409 = n4290 & ~n4408 ;
  assign n4529 = n4413 ^ n4409 ;
  assign n4415 = n2628 ^ n2625 ;
  assign n4416 = n4415 ^ n4367 ;
  assign n4418 = n4416 ^ n2629 ;
  assign n4417 = n4367 & ~n4415 ;
  assign n4419 = n4418 ^ n4417 ;
  assign n4420 = n2462 & n4419 ;
  assign n4421 = ~n2630 & ~n4417 ;
  assign n4423 = n2624 ^ n2617 ;
  assign n4422 = n4373 ^ n4326 ;
  assign n4424 = n4423 ^ n4422 ;
  assign n4426 = n4378 ^ n4332 ;
  assign n4425 = n2623 ^ n2622 ;
  assign n4427 = n4426 ^ n4425 ;
  assign n4429 = n4388 ^ n4339 ;
  assign n4428 = n2621 ^ n2618 ;
  assign n4430 = n4429 ^ n4428 ;
  assign n4431 = n2620 ^ n2619 ;
  assign n4432 = n4384 ^ n4346 ;
  assign n4433 = n4431 & ~n4432 ;
  assign n4434 = n4433 ^ n4429 ;
  assign n4435 = ~n4430 & ~n4434 ;
  assign n4436 = n4435 ^ n4429 ;
  assign n4437 = n4436 ^ n4425 ;
  assign n4438 = ~n4427 & ~n4437 ;
  assign n4439 = n4438 ^ n4425 ;
  assign n4440 = n4439 ^ n4423 ;
  assign n4441 = ~n4424 & n4440 ;
  assign n4442 = n4441 ^ n4423 ;
  assign n4443 = n4421 & n4442 ;
  assign n4444 = ~n4420 & ~n4443 ;
  assign n4445 = n4416 & ~n4444 ;
  assign n4446 = n4445 ^ n4415 ;
  assign n4410 = n4409 ^ n4370 ;
  assign n4414 = n4413 ^ n4410 ;
  assign n4447 = n4446 ^ n4414 ;
  assign n4450 = n4424 & ~n4444 ;
  assign n4451 = n4450 ^ n4423 ;
  assign n4448 = n4376 & ~n4407 ;
  assign n4449 = n4448 ^ n4375 ;
  assign n4452 = n4451 ^ n4449 ;
  assign n4456 = n4427 & ~n4444 ;
  assign n4457 = n4456 ^ n4425 ;
  assign n4453 = n4381 & ~n4407 ;
  assign n4454 = n4453 ^ n4381 ;
  assign n4455 = n4454 ^ n4377 ;
  assign n4458 = n4457 ^ n4455 ;
  assign n4461 = n4392 ^ n4390 ;
  assign n4462 = ~n4407 & n4461 ;
  assign n4463 = n4462 ^ n4461 ;
  assign n4464 = n4463 ^ n4392 ;
  assign n4459 = n4430 & ~n4444 ;
  assign n4460 = n4459 ^ n4428 ;
  assign n4465 = n4464 ^ n4460 ;
  assign n4466 = n4386 ^ n4382 ;
  assign n4467 = ~n4407 & n4466 ;
  assign n4468 = n4467 ^ n4466 ;
  assign n4469 = n4468 ^ n4382 ;
  assign n4470 = n4432 ^ n4431 ;
  assign n4471 = ~n4444 & n4470 ;
  assign n4472 = n4471 ^ n4431 ;
  assign n4473 = ~n4469 & n4472 ;
  assign n4474 = n4473 ^ n4464 ;
  assign n4475 = ~n4465 & ~n4474 ;
  assign n4476 = n4475 ^ n4464 ;
  assign n4477 = n4476 ^ n4457 ;
  assign n4478 = ~n4458 & ~n4477 ;
  assign n4479 = n4478 ^ n4457 ;
  assign n4480 = n4479 ^ n4451 ;
  assign n4481 = ~n4452 & ~n4480 ;
  assign n4482 = n4481 ^ n4449 ;
  assign n4483 = n4482 ^ n4446 ;
  assign n4484 = ~n4447 & n4483 ;
  assign n4485 = n4484 ^ n4414 ;
  assign n4486 = n4485 ^ n2460 ;
  assign n4487 = n2636 & ~n4486 ;
  assign n4488 = n4487 ^ n2631 ;
  assign n4489 = n4447 & ~n4488 ;
  assign n4490 = n4489 ^ n4414 ;
  assign n4527 = n4490 ^ n4446 ;
  assign n4528 = n4527 ^ n4414 ;
  assign n4530 = n4529 ^ n4528 ;
  assign n4531 = n2633 ^ n2632 ;
  assign n4497 = n4452 & ~n4488 ;
  assign n4533 = n4497 ^ n4452 ;
  assign n4534 = n4533 ^ n4449 ;
  assign n4532 = n4448 ^ n4372 ;
  assign n4535 = n4534 ^ n4532 ;
  assign n4502 = n4458 & ~n4488 ;
  assign n4537 = n4502 ^ n4458 ;
  assign n4538 = n4537 ^ n4455 ;
  assign n4536 = n4453 ^ n4377 ;
  assign n4539 = n4538 ^ n4536 ;
  assign n4506 = n4465 & n4488 ;
  assign n4544 = n4506 ^ n4465 ;
  assign n4545 = n4544 ^ n4460 ;
  assign n4510 = n4472 ^ n4469 ;
  assign n4511 = ~n4488 & n4510 ;
  assign n4540 = n4511 ^ n4510 ;
  assign n4541 = n4540 ^ n4469 ;
  assign n4542 = n4467 ^ n4382 ;
  assign n4543 = n4541 & ~n4542 ;
  assign n4546 = n4545 ^ n4543 ;
  assign n4547 = n4462 ^ n4392 ;
  assign n4548 = n4547 ^ n4543 ;
  assign n4549 = n4546 & ~n4548 ;
  assign n4550 = n4549 ^ n4543 ;
  assign n4551 = n4550 ^ n4538 ;
  assign n4552 = ~n4539 & n4551 ;
  assign n4553 = n4552 ^ n4538 ;
  assign n4554 = n4553 ^ n4534 ;
  assign n4555 = ~n4535 & n4554 ;
  assign n4556 = n4555 ^ n4534 ;
  assign n4557 = n4556 ^ n4529 ;
  assign n4558 = ~n4530 & ~n4557 ;
  assign n4559 = n4558 ^ n4529 ;
  assign n4560 = n4559 ^ n2633 ;
  assign n4561 = ~n4531 & ~n4560 ;
  assign n4562 = n4561 ^ n2632 ;
  assign n4563 = n4530 & ~n4562 ;
  assign n4611 = n4563 ^ n4529 ;
  assign n4564 = n4563 ^ n4528 ;
  assign n3339 = n2803 ^ n2800 ;
  assign n4491 = n4490 ^ n3339 ;
  assign n4493 = n4491 ^ n2804 ;
  assign n4492 = ~n3339 & n4490 ;
  assign n4494 = n4493 ^ n4492 ;
  assign n4495 = n2637 & n4494 ;
  assign n4496 = ~n2805 & ~n4492 ;
  assign n4499 = n2799 ^ n2792 ;
  assign n4498 = n4497 ^ n4449 ;
  assign n4500 = n4499 ^ n4498 ;
  assign n4503 = n4502 ^ n4455 ;
  assign n4501 = n2798 ^ n2797 ;
  assign n4504 = n4503 ^ n4501 ;
  assign n4507 = n4506 ^ n4460 ;
  assign n4505 = n2796 ^ n2793 ;
  assign n4508 = n4507 ^ n4505 ;
  assign n4509 = n2795 ^ n2794 ;
  assign n4512 = n4511 ^ n4469 ;
  assign n4513 = n4509 & ~n4512 ;
  assign n4514 = n4513 ^ n4507 ;
  assign n4515 = ~n4508 & ~n4514 ;
  assign n4516 = n4515 ^ n4507 ;
  assign n4517 = n4516 ^ n4501 ;
  assign n4518 = ~n4504 & ~n4517 ;
  assign n4519 = n4518 ^ n4501 ;
  assign n4520 = n4519 ^ n4499 ;
  assign n4521 = ~n4500 & n4520 ;
  assign n4522 = n4521 ^ n4499 ;
  assign n4523 = n4496 & n4522 ;
  assign n4524 = ~n4495 & ~n4523 ;
  assign n4525 = n4491 & ~n4524 ;
  assign n4526 = n4525 ^ n3339 ;
  assign n4565 = n4564 ^ n4526 ;
  assign n4568 = n4535 & ~n4562 ;
  assign n4569 = n4568 ^ n4534 ;
  assign n4566 = n4500 & ~n4524 ;
  assign n4567 = n4566 ^ n4499 ;
  assign n4570 = n4569 ^ n4567 ;
  assign n4574 = n4504 & ~n4524 ;
  assign n4575 = n4574 ^ n4501 ;
  assign n4571 = n4539 & ~n4562 ;
  assign n4572 = n4571 ^ n4539 ;
  assign n4573 = n4572 ^ n4536 ;
  assign n4576 = n4575 ^ n4573 ;
  assign n4581 = n4508 & ~n4524 ;
  assign n4582 = n4581 ^ n4505 ;
  assign n4577 = n4547 ^ n4545 ;
  assign n4578 = ~n4562 & n4577 ;
  assign n4579 = n4578 ^ n4577 ;
  assign n4580 = n4579 ^ n4547 ;
  assign n4583 = n4582 ^ n4580 ;
  assign n4584 = n4542 ^ n4541 ;
  assign n4585 = n4562 & n4584 ;
  assign n4586 = n4585 ^ n4584 ;
  assign n4587 = n4586 ^ n4541 ;
  assign n4588 = n4512 ^ n4509 ;
  assign n4589 = ~n4524 & n4588 ;
  assign n4590 = n4589 ^ n4509 ;
  assign n4591 = ~n4587 & n4590 ;
  assign n4592 = n4591 ^ n4582 ;
  assign n4593 = ~n4583 & n4592 ;
  assign n4594 = n4593 ^ n4582 ;
  assign n4595 = n4594 ^ n4575 ;
  assign n4596 = ~n4576 & n4595 ;
  assign n4597 = n4596 ^ n4575 ;
  assign n4598 = n4597 ^ n4567 ;
  assign n4599 = ~n4570 & ~n4598 ;
  assign n4600 = n4599 ^ n4569 ;
  assign n4601 = n4600 ^ n4526 ;
  assign n4602 = ~n4565 & n4601 ;
  assign n4603 = n4602 ^ n4564 ;
  assign n4604 = n4603 ^ n2806 ;
  assign n4605 = n2814 & ~n4604 ;
  assign n4606 = n4605 ^ n2808 ;
  assign n4607 = n4565 & ~n4606 ;
  assign n4608 = n4607 ^ n4564 ;
  assign n4609 = n4608 ^ n4526 ;
  assign n4610 = n4609 ^ n4564 ;
  assign n4612 = n4611 ^ n4610 ;
  assign n4613 = n2809 ^ n2635 ;
  assign n4615 = n4570 & ~n4606 ;
  assign n4616 = n4615 ^ n4570 ;
  assign n4617 = n4616 ^ n4569 ;
  assign n4614 = n4568 ^ n4532 ;
  assign n4618 = n4617 ^ n4614 ;
  assign n4620 = n4576 & ~n4606 ;
  assign n4621 = n4620 ^ n4576 ;
  assign n4622 = n4621 ^ n4573 ;
  assign n4619 = n4571 ^ n4536 ;
  assign n4623 = n4622 ^ n4619 ;
  assign n4630 = n4583 & ~n4606 ;
  assign n4631 = n4630 ^ n4583 ;
  assign n4632 = n4631 ^ n4580 ;
  assign n4624 = n4585 ^ n4541 ;
  assign n4625 = n4590 ^ n4587 ;
  assign n4626 = ~n4606 & n4625 ;
  assign n4627 = n4626 ^ n4625 ;
  assign n4628 = n4627 ^ n4587 ;
  assign n4629 = ~n4624 & n4628 ;
  assign n4633 = n4632 ^ n4629 ;
  assign n4634 = n4578 ^ n4547 ;
  assign n4635 = n4634 ^ n4629 ;
  assign n4636 = n4633 & ~n4635 ;
  assign n4637 = n4636 ^ n4629 ;
  assign n4638 = n4637 ^ n4622 ;
  assign n4639 = ~n4623 & n4638 ;
  assign n4640 = n4639 ^ n4622 ;
  assign n4641 = n4640 ^ n4617 ;
  assign n4642 = ~n4618 & n4641 ;
  assign n4643 = n4642 ^ n4617 ;
  assign n4644 = n4643 ^ n4611 ;
  assign n4645 = ~n4612 & ~n4644 ;
  assign n4646 = n4645 ^ n4611 ;
  assign n4647 = n4646 ^ n2809 ;
  assign n4648 = ~n4613 & n4647 ;
  assign n4649 = n4648 ^ n2635 ;
  assign n4650 = n4612 & n4649 ;
  assign n4684 = n4650 ^ n4610 ;
  assign n4652 = n2981 ^ n2978 ;
  assign n4653 = n4652 ^ n4608 ;
  assign n4655 = n4653 ^ n2982 ;
  assign n4654 = n4608 & ~n4652 ;
  assign n4656 = n4655 ^ n4654 ;
  assign n4657 = n2815 & n4656 ;
  assign n4658 = ~n2983 & ~n4654 ;
  assign n4660 = n2977 ^ n2970 ;
  assign n4659 = n4615 ^ n4569 ;
  assign n4661 = n4660 ^ n4659 ;
  assign n4663 = n4620 ^ n4573 ;
  assign n4662 = n2976 ^ n2975 ;
  assign n4664 = n4663 ^ n4662 ;
  assign n4666 = n4630 ^ n4580 ;
  assign n4665 = n2974 ^ n2971 ;
  assign n4667 = n4666 ^ n4665 ;
  assign n4668 = n2973 ^ n2972 ;
  assign n4669 = n4626 ^ n4587 ;
  assign n4670 = n4668 & ~n4669 ;
  assign n4671 = n4670 ^ n4666 ;
  assign n4672 = ~n4667 & ~n4671 ;
  assign n4673 = n4672 ^ n4666 ;
  assign n4674 = n4673 ^ n4662 ;
  assign n4675 = ~n4664 & ~n4674 ;
  assign n4676 = n4675 ^ n4662 ;
  assign n4677 = n4676 ^ n4660 ;
  assign n4678 = ~n4661 & n4677 ;
  assign n4679 = n4678 ^ n4660 ;
  assign n4680 = n4658 & n4679 ;
  assign n4681 = ~n4657 & ~n4680 ;
  assign n4682 = n4653 & ~n4681 ;
  assign n4683 = n4682 ^ n4652 ;
  assign n4685 = n4684 ^ n4683 ;
  assign n4688 = n4618 & n4649 ;
  assign n4689 = n4688 ^ n4617 ;
  assign n4686 = n4661 & ~n4681 ;
  assign n4687 = n4686 ^ n4660 ;
  assign n4690 = n4689 ^ n4687 ;
  assign n4694 = n4664 & ~n4681 ;
  assign n4695 = n4694 ^ n4662 ;
  assign n4691 = n4623 & n4649 ;
  assign n4692 = n4691 ^ n4623 ;
  assign n4693 = n4692 ^ n4619 ;
  assign n4696 = n4695 ^ n4693 ;
  assign n4699 = n4634 ^ n4632 ;
  assign n4700 = n4649 & n4699 ;
  assign n4701 = n4700 ^ n4699 ;
  assign n4702 = n4701 ^ n4634 ;
  assign n4697 = n4667 & ~n4681 ;
  assign n4698 = n4697 ^ n4665 ;
  assign n4703 = n4702 ^ n4698 ;
  assign n4704 = n4628 ^ n4624 ;
  assign n4705 = n4649 & n4704 ;
  assign n4706 = n4705 ^ n4704 ;
  assign n4707 = n4706 ^ n4624 ;
  assign n4708 = n4669 ^ n4668 ;
  assign n4709 = ~n4681 & n4708 ;
  assign n4710 = n4709 ^ n4668 ;
  assign n4711 = ~n4707 & n4710 ;
  assign n4712 = n4711 ^ n4702 ;
  assign n4713 = ~n4703 & ~n4712 ;
  assign n4714 = n4713 ^ n4702 ;
  assign n4715 = n4714 ^ n4695 ;
  assign n4716 = ~n4696 & ~n4715 ;
  assign n4717 = n4716 ^ n4695 ;
  assign n4718 = n4717 ^ n4689 ;
  assign n4719 = ~n4690 & n4718 ;
  assign n4720 = n4719 ^ n4687 ;
  assign n4721 = n4720 ^ n4683 ;
  assign n4722 = ~n4685 & ~n4721 ;
  assign n4723 = n4722 ^ n4684 ;
  assign n4724 = n4723 ^ n2984 ;
  assign n4725 = n2986 & ~n4724 ;
  assign n4726 = n4725 ^ n2813 ;
  assign n4727 = n4685 & ~n4726 ;
  assign n4728 = n4727 ^ n4684 ;
  assign n4729 = n4728 ^ n4683 ;
  assign n4730 = n4729 ^ n4684 ;
  assign n4651 = n4650 ^ n4611 ;
  assign n4734 = n4730 ^ n4651 ;
  assign n4731 = ~n4651 & n4730 ;
  assign n4735 = n4734 ^ n4731 ;
  assign n4736 = n2987 ^ n2811 ;
  assign n4738 = n4690 & ~n4726 ;
  assign n4739 = n4738 ^ n4690 ;
  assign n4740 = n4739 ^ n4689 ;
  assign n4737 = n4688 ^ n4614 ;
  assign n4741 = n4740 ^ n4737 ;
  assign n4743 = n4696 & ~n4726 ;
  assign n4744 = n4743 ^ n4696 ;
  assign n4745 = n4744 ^ n4693 ;
  assign n4742 = n4691 ^ n4619 ;
  assign n4746 = n4745 ^ n4742 ;
  assign n4753 = n4703 & n4726 ;
  assign n4754 = n4753 ^ n4703 ;
  assign n4755 = n4754 ^ n4698 ;
  assign n4747 = n4710 ^ n4707 ;
  assign n4748 = ~n4726 & n4747 ;
  assign n4749 = n4748 ^ n4747 ;
  assign n4750 = n4749 ^ n4707 ;
  assign n4751 = n4705 ^ n4624 ;
  assign n4752 = n4750 & ~n4751 ;
  assign n4756 = n4755 ^ n4752 ;
  assign n4757 = n4700 ^ n4634 ;
  assign n4758 = n4757 ^ n4752 ;
  assign n4759 = n4756 & ~n4758 ;
  assign n4760 = n4759 ^ n4752 ;
  assign n4761 = n4760 ^ n4745 ;
  assign n4762 = ~n4746 & n4761 ;
  assign n4763 = n4762 ^ n4745 ;
  assign n4764 = n4763 ^ n4737 ;
  assign n4765 = ~n4741 & ~n4764 ;
  assign n4766 = n4765 ^ n4737 ;
  assign n4767 = n4766 ^ n4730 ;
  assign n4768 = ~n4734 & n4767 ;
  assign n4769 = n4768 ^ n4651 ;
  assign n4770 = n4769 ^ n2811 ;
  assign n4771 = ~n4736 & ~n4770 ;
  assign n4772 = n4771 ^ n2987 ;
  assign n4773 = n4735 & ~n4772 ;
  assign n4732 = n2988 & n4731 ;
  assign n4733 = n4732 ^ n4651 ;
  assign n4774 = n4773 ^ n4733 ;
  assign n4777 = n3155 ^ n3152 ;
  assign n4778 = n4777 ^ n4728 ;
  assign n4780 = n4778 ^ n3156 ;
  assign n4779 = n4728 & ~n4777 ;
  assign n4781 = n4780 ^ n4779 ;
  assign n4782 = n2985 & n4781 ;
  assign n4783 = ~n3157 & ~n4779 ;
  assign n4785 = n3151 ^ n3144 ;
  assign n4784 = n4738 ^ n4689 ;
  assign n4786 = n4785 ^ n4784 ;
  assign n4788 = n4743 ^ n4693 ;
  assign n4787 = n3150 ^ n3149 ;
  assign n4789 = n4788 ^ n4787 ;
  assign n4791 = n4753 ^ n4698 ;
  assign n4790 = n3148 ^ n3145 ;
  assign n4792 = n4791 ^ n4790 ;
  assign n4793 = n3147 ^ n3146 ;
  assign n4794 = n4748 ^ n4707 ;
  assign n4795 = n4793 & ~n4794 ;
  assign n4796 = n4795 ^ n4791 ;
  assign n4797 = ~n4792 & ~n4796 ;
  assign n4798 = n4797 ^ n4791 ;
  assign n4799 = n4798 ^ n4787 ;
  assign n4800 = ~n4789 & ~n4799 ;
  assign n4801 = n4800 ^ n4787 ;
  assign n4802 = n4801 ^ n4785 ;
  assign n4803 = ~n4786 & n4802 ;
  assign n4804 = n4803 ^ n4785 ;
  assign n4805 = n4783 & n4804 ;
  assign n4806 = ~n4782 & ~n4805 ;
  assign n4807 = n4778 & ~n4806 ;
  assign n4808 = n4807 ^ n4777 ;
  assign n4775 = n4773 ^ n4730 ;
  assign n4776 = n4775 ^ n4732 ;
  assign n4809 = n4808 ^ n4776 ;
  assign n4812 = n4786 & ~n4806 ;
  assign n4813 = n4812 ^ n4785 ;
  assign n4810 = n4741 & ~n4772 ;
  assign n4811 = n4810 ^ n4740 ;
  assign n4814 = n4813 ^ n4811 ;
  assign n4818 = n4789 & ~n4806 ;
  assign n4819 = n4818 ^ n4787 ;
  assign n4815 = n4746 & ~n4772 ;
  assign n4816 = n4815 ^ n4746 ;
  assign n4817 = n4816 ^ n4742 ;
  assign n4820 = n4819 ^ n4817 ;
  assign n4825 = n4792 & ~n4806 ;
  assign n4826 = n4825 ^ n4790 ;
  assign n4821 = n4757 ^ n4755 ;
  assign n4822 = ~n4772 & n4821 ;
  assign n4823 = n4822 ^ n4821 ;
  assign n4824 = n4823 ^ n4757 ;
  assign n4827 = n4826 ^ n4824 ;
  assign n4828 = n4751 ^ n4750 ;
  assign n4829 = n4772 & n4828 ;
  assign n4830 = n4829 ^ n4828 ;
  assign n4831 = n4830 ^ n4750 ;
  assign n4832 = n4794 ^ n4793 ;
  assign n4833 = ~n4806 & n4832 ;
  assign n4834 = n4833 ^ n4793 ;
  assign n4835 = ~n4831 & n4834 ;
  assign n4836 = n4835 ^ n4826 ;
  assign n4837 = ~n4827 & n4836 ;
  assign n4838 = n4837 ^ n4826 ;
  assign n4839 = n4838 ^ n4819 ;
  assign n4840 = ~n4820 & n4839 ;
  assign n4841 = n4840 ^ n4819 ;
  assign n4842 = n4841 ^ n4811 ;
  assign n4843 = ~n4814 & n4842 ;
  assign n4844 = n4843 ^ n4813 ;
  assign n4845 = n4844 ^ n4808 ;
  assign n4846 = ~n4809 & ~n4845 ;
  assign n4847 = n4846 ^ n4776 ;
  assign n4848 = n4847 ^ n3159 ;
  assign n4849 = n3165 & ~n4848 ;
  assign n4850 = n4849 ^ n3158 ;
  assign n4851 = n4809 & ~n4850 ;
  assign n4852 = n4851 ^ n4776 ;
  assign n4853 = n4852 ^ n4808 ;
  assign n4854 = n4853 ^ n4776 ;
  assign n4856 = ~n4774 & n4854 ;
  assign n4896 = n3163 & n4856 ;
  assign n4975 = n4896 ^ n4774 ;
  assign n4855 = n4854 ^ n4774 ;
  assign n4857 = n4856 ^ n4855 ;
  assign n4859 = n4814 & ~n4850 ;
  assign n4860 = n4859 ^ n4814 ;
  assign n4861 = n4860 ^ n4811 ;
  assign n4858 = n4810 ^ n4737 ;
  assign n4862 = n4861 ^ n4858 ;
  assign n4864 = n4820 & ~n4850 ;
  assign n4865 = n4864 ^ n4820 ;
  assign n4866 = n4865 ^ n4817 ;
  assign n4863 = n4815 ^ n4742 ;
  assign n4867 = n4866 ^ n4863 ;
  assign n4874 = n4827 & ~n4850 ;
  assign n4875 = n4874 ^ n4827 ;
  assign n4876 = n4875 ^ n4824 ;
  assign n4868 = n4829 ^ n4750 ;
  assign n4869 = n4834 ^ n4831 ;
  assign n4870 = ~n4850 & n4869 ;
  assign n4871 = n4870 ^ n4869 ;
  assign n4872 = n4871 ^ n4831 ;
  assign n4873 = ~n4868 & n4872 ;
  assign n4877 = n4876 ^ n4873 ;
  assign n4878 = n4822 ^ n4757 ;
  assign n4879 = n4878 ^ n4873 ;
  assign n4880 = n4877 & ~n4879 ;
  assign n4881 = n4880 ^ n4873 ;
  assign n4882 = n4881 ^ n4866 ;
  assign n4883 = ~n4867 & n4882 ;
  assign n4884 = n4883 ^ n4866 ;
  assign n4885 = n4884 ^ n4858 ;
  assign n4886 = ~n4862 & ~n4885 ;
  assign n4887 = n4886 ^ n4858 ;
  assign n4888 = n4887 ^ n4774 ;
  assign n4889 = ~n4855 & ~n4888 ;
  assign n4890 = n4889 ^ n4854 ;
  assign n4891 = n4890 ^ n3160 ;
  assign n4892 = ~n3162 & ~n4891 ;
  assign n4893 = n4892 ^ n2989 ;
  assign n4894 = n4857 & n4893 ;
  assign n4976 = n4975 ^ n4894 ;
  assign n4898 = n3332 ^ n3329 ;
  assign n4899 = n4898 ^ n4852 ;
  assign n4901 = n4899 ^ n3333 ;
  assign n4900 = n4852 & ~n4898 ;
  assign n4902 = n4901 ^ n4900 ;
  assign n4903 = n3166 & n4902 ;
  assign n4904 = ~n3334 & ~n4900 ;
  assign n4906 = n3328 ^ n3321 ;
  assign n4905 = n4859 ^ n4811 ;
  assign n4907 = n4906 ^ n4905 ;
  assign n4909 = n4864 ^ n4817 ;
  assign n4908 = n3327 ^ n3326 ;
  assign n4910 = n4909 ^ n4908 ;
  assign n4912 = n3325 ^ n3322 ;
  assign n4911 = n4874 ^ n4824 ;
  assign n4913 = n4912 ^ n4911 ;
  assign n4914 = n3324 ^ n3323 ;
  assign n4915 = n4870 ^ n4831 ;
  assign n4916 = n4914 & ~n4915 ;
  assign n4917 = n4916 ^ n4912 ;
  assign n4918 = ~n4913 & n4917 ;
  assign n4919 = n4918 ^ n4912 ;
  assign n4920 = n4919 ^ n4908 ;
  assign n4921 = ~n4910 & n4920 ;
  assign n4922 = n4921 ^ n4908 ;
  assign n4923 = n4922 ^ n4906 ;
  assign n4924 = ~n4907 & n4923 ;
  assign n4925 = n4924 ^ n4906 ;
  assign n4926 = n4904 & n4925 ;
  assign n4927 = ~n4903 & ~n4926 ;
  assign n4928 = n4899 & ~n4927 ;
  assign n4929 = n4928 ^ n4898 ;
  assign n4895 = n4894 ^ n4854 ;
  assign n4897 = n4896 ^ n4895 ;
  assign n4930 = n4929 ^ n4897 ;
  assign n4931 = n3335 ^ n3164 ;
  assign n4934 = n4907 & ~n4927 ;
  assign n4935 = n4934 ^ n4906 ;
  assign n4932 = n4862 & n4893 ;
  assign n4933 = n4932 ^ n4861 ;
  assign n4936 = n4935 ^ n4933 ;
  assign n4940 = n4910 & ~n4927 ;
  assign n4941 = n4940 ^ n4908 ;
  assign n4937 = n4867 & n4893 ;
  assign n4938 = n4937 ^ n4867 ;
  assign n4939 = n4938 ^ n4863 ;
  assign n4942 = n4941 ^ n4939 ;
  assign n4945 = n4878 ^ n4876 ;
  assign n4946 = n4893 & n4945 ;
  assign n4947 = n4946 ^ n4945 ;
  assign n4948 = n4947 ^ n4878 ;
  assign n4943 = n4913 & n4927 ;
  assign n4944 = n4943 ^ n4911 ;
  assign n4949 = n4948 ^ n4944 ;
  assign n4950 = n4915 ^ n4914 ;
  assign n4951 = ~n4927 & n4950 ;
  assign n4952 = n4951 ^ n4914 ;
  assign n4953 = n4872 ^ n4868 ;
  assign n4954 = n4893 & n4953 ;
  assign n4955 = n4954 ^ n4953 ;
  assign n4956 = n4955 ^ n4868 ;
  assign n4957 = n4952 & ~n4956 ;
  assign n4958 = n4957 ^ n4948 ;
  assign n4959 = ~n4949 & ~n4958 ;
  assign n4960 = n4959 ^ n4948 ;
  assign n4961 = n4960 ^ n4941 ;
  assign n4962 = ~n4942 & ~n4961 ;
  assign n4963 = n4962 ^ n4941 ;
  assign n4964 = n4963 ^ n4935 ;
  assign n4965 = ~n4936 & ~n4964 ;
  assign n4966 = n4965 ^ n4933 ;
  assign n4967 = n4966 ^ n4929 ;
  assign n4968 = ~n4930 & n4967 ;
  assign n4969 = n4968 ^ n4897 ;
  assign n4970 = n4969 ^ n3335 ;
  assign n4971 = n4931 & ~n4970 ;
  assign n4972 = n4971 ^ n3164 ;
  assign n4973 = n4930 & n4972 ;
  assign n4974 = n4973 ^ n4897 ;
  assign n4977 = n4976 ^ n4974 ;
  assign n4980 = n4932 ^ n4858 ;
  assign n4978 = n4936 & n4972 ;
  assign n4979 = n4978 ^ n4933 ;
  assign n4981 = n4980 ^ n4979 ;
  assign n4983 = n4942 & n4972 ;
  assign n4984 = n4983 ^ n4939 ;
  assign n4982 = n4937 ^ n4863 ;
  assign n4985 = n4984 ^ n4982 ;
  assign n4987 = n4949 & ~n4972 ;
  assign n4988 = n4987 ^ n4944 ;
  assign n4986 = n4946 ^ n4878 ;
  assign n4989 = n4988 ^ n4986 ;
  assign n4990 = n4954 ^ n4868 ;
  assign n4991 = n4956 ^ n4952 ;
  assign n4992 = n4972 & n4991 ;
  assign n4993 = n4992 ^ n4956 ;
  assign n4994 = ~n4990 & n4993 ;
  assign n4995 = n4994 ^ n4988 ;
  assign n4996 = ~n4989 & n4995 ;
  assign n4997 = n4996 ^ n4988 ;
  assign n4998 = n4997 ^ n4984 ;
  assign n4999 = ~n4985 & n4998 ;
  assign n5000 = n4999 ^ n4984 ;
  assign n5001 = n5000 ^ n4979 ;
  assign n5002 = ~n4981 & n5001 ;
  assign n5003 = n5002 ^ n4979 ;
  assign n5004 = n5003 ^ n4974 ;
  assign n5005 = ~n4977 & ~n5004 ;
  assign n5006 = n5005 ^ n4976 ;
  assign n5007 = n5006 ^ n3336 ;
  assign n5008 = ~n3338 & n5007 ;
  assign n5009 = n5008 ^ n3337 ;
  assign n5010 = x480 ^ x448 ;
  assign n5011 = n3371 & n5010 ;
  assign n5018 = n5011 ^ x448 ;
  assign n5012 = n5011 ^ n5010 ;
  assign n5013 = n5012 ^ x448 ;
  assign n5014 = n5013 ^ x416 ;
  assign n5015 = n3412 & n5014 ;
  assign n5016 = n5015 ^ n5014 ;
  assign n5017 = n5016 ^ x416 ;
  assign n5019 = n5018 ^ n5017 ;
  assign n5020 = n3451 & n5019 ;
  assign n5035 = n5020 ^ n5017 ;
  assign n5023 = n5015 ^ x416 ;
  assign n5024 = n5023 ^ x384 ;
  assign n5025 = ~n3484 & n5024 ;
  assign n5026 = n5025 ^ x384 ;
  assign n5021 = n5020 ^ n5019 ;
  assign n5022 = n5021 ^ n5017 ;
  assign n5027 = n5026 ^ n5022 ;
  assign n5028 = ~n3527 & n5027 ;
  assign n5034 = n5028 ^ n5022 ;
  assign n5036 = n5035 ^ n5034 ;
  assign n5037 = ~n3570 & n5036 ;
  assign n5038 = n5037 ^ n5036 ;
  assign n5039 = n5038 ^ n5034 ;
  assign n5029 = n5028 ^ n5027 ;
  assign n5030 = n5029 ^ n5022 ;
  assign n5031 = n5030 ^ x352 ;
  assign n5032 = ~n3602 & n5031 ;
  assign n5033 = n5032 ^ x352 ;
  assign n5040 = n5039 ^ n5033 ;
  assign n5041 = ~n3646 & n5040 ;
  assign n5048 = n5041 ^ n5033 ;
  assign n5047 = n5037 ^ n5034 ;
  assign n5049 = n5048 ^ n5047 ;
  assign n5050 = ~n3688 & n5049 ;
  assign n5057 = n5050 ^ n5047 ;
  assign n5051 = n5050 ^ n5049 ;
  assign n5052 = n5051 ^ n5047 ;
  assign n5042 = n5041 ^ n5040 ;
  assign n5043 = n5042 ^ n5033 ;
  assign n5044 = n5043 ^ x320 ;
  assign n5045 = ~n3724 & n5044 ;
  assign n5046 = n5045 ^ x320 ;
  assign n5053 = n5052 ^ n5046 ;
  assign n5054 = n3767 & n5053 ;
  assign n5055 = n5054 ^ n5053 ;
  assign n5056 = n5055 ^ n5046 ;
  assign n5058 = n5057 ^ n5056 ;
  assign n5059 = n3841 & n5058 ;
  assign n5070 = n5059 ^ n5056 ;
  assign n5062 = n5054 ^ n5046 ;
  assign n5063 = n5062 ^ x288 ;
  assign n5064 = ~n3803 & n5063 ;
  assign n5065 = n5064 ^ x288 ;
  assign n5060 = n5059 ^ n5058 ;
  assign n5061 = n5060 ^ n5056 ;
  assign n5066 = n5065 ^ n5061 ;
  assign n5067 = ~n3884 & n5066 ;
  assign n5068 = n5067 ^ n5066 ;
  assign n5069 = n5068 ^ n5061 ;
  assign n5071 = n5070 ^ n5069 ;
  assign n5072 = ~n3927 & n5071 ;
  assign n5087 = n5072 ^ n5069 ;
  assign n5075 = n5067 ^ n5061 ;
  assign n5076 = n5075 ^ x256 ;
  assign n5077 = ~n3959 & n5076 ;
  assign n5078 = n5077 ^ x256 ;
  assign n5073 = n5072 ^ n5071 ;
  assign n5074 = n5073 ^ n5069 ;
  assign n5079 = n5078 ^ n5074 ;
  assign n5080 = n4004 & n5079 ;
  assign n5086 = n5080 ^ n5074 ;
  assign n5088 = n5087 ^ n5086 ;
  assign n5089 = n4046 & n5088 ;
  assign n5096 = n5089 ^ n5086 ;
  assign n5090 = n5089 ^ n5088 ;
  assign n5091 = n5090 ^ n5086 ;
  assign n5081 = n5080 ^ n5079 ;
  assign n5082 = n5081 ^ n5074 ;
  assign n5083 = n5082 ^ x224 ;
  assign n5084 = ~n4083 & n5083 ;
  assign n5085 = n5084 ^ x224 ;
  assign n5092 = n5091 ^ n5085 ;
  assign n5093 = n4127 & n5092 ;
  assign n5094 = n5093 ^ n5092 ;
  assign n5095 = n5094 ^ n5085 ;
  assign n5097 = n5096 ^ n5095 ;
  assign n5098 = n4201 & n5097 ;
  assign n5109 = n5098 ^ n5095 ;
  assign n5101 = n5093 ^ n5085 ;
  assign n5102 = n5101 ^ x192 ;
  assign n5103 = ~n4163 & n5102 ;
  assign n5104 = n5103 ^ x192 ;
  assign n5099 = n5098 ^ n5097 ;
  assign n5100 = n5099 ^ n5095 ;
  assign n5105 = n5104 ^ n5100 ;
  assign n5106 = ~n4245 & n5105 ;
  assign n5107 = n5106 ^ n5105 ;
  assign n5108 = n5107 ^ n5100 ;
  assign n5110 = n5109 ^ n5108 ;
  assign n5111 = ~n4288 & n5110 ;
  assign n5126 = n5111 ^ n5108 ;
  assign n5114 = n5106 ^ n5100 ;
  assign n5115 = n5114 ^ x160 ;
  assign n5116 = ~n4320 & n5115 ;
  assign n5117 = n5116 ^ x160 ;
  assign n5112 = n5111 ^ n5110 ;
  assign n5113 = n5112 ^ n5108 ;
  assign n5118 = n5117 ^ n5113 ;
  assign n5119 = n4365 & n5118 ;
  assign n5125 = n5119 ^ n5113 ;
  assign n5127 = n5126 ^ n5125 ;
  assign n5128 = n4407 & n5127 ;
  assign n5135 = n5128 ^ n5125 ;
  assign n5129 = n5128 ^ n5127 ;
  assign n5130 = n5129 ^ n5125 ;
  assign n5120 = n5119 ^ n5118 ;
  assign n5121 = n5120 ^ n5113 ;
  assign n5122 = n5121 ^ x128 ;
  assign n5123 = ~n4444 & n5122 ;
  assign n5124 = n5123 ^ x128 ;
  assign n5131 = n5130 ^ n5124 ;
  assign n5132 = n4488 & n5131 ;
  assign n5133 = n5132 ^ n5131 ;
  assign n5134 = n5133 ^ n5124 ;
  assign n5136 = n5135 ^ n5134 ;
  assign n5137 = n4562 & n5136 ;
  assign n5148 = n5137 ^ n5134 ;
  assign n5140 = n5132 ^ n5124 ;
  assign n5141 = n5140 ^ x96 ;
  assign n5142 = ~n4524 & n5141 ;
  assign n5143 = n5142 ^ x96 ;
  assign n5138 = n5137 ^ n5136 ;
  assign n5139 = n5138 ^ n5134 ;
  assign n5144 = n5143 ^ n5139 ;
  assign n5145 = ~n4606 & n5144 ;
  assign n5146 = n5145 ^ n5144 ;
  assign n5147 = n5146 ^ n5139 ;
  assign n5149 = n5148 ^ n5147 ;
  assign n5150 = ~n4649 & n5149 ;
  assign n5161 = n5150 ^ n5147 ;
  assign n5153 = n5145 ^ n5139 ;
  assign n5154 = n5153 ^ x64 ;
  assign n5155 = ~n4681 & n5154 ;
  assign n5156 = n5155 ^ x64 ;
  assign n5151 = n5150 ^ n5149 ;
  assign n5152 = n5151 ^ n5147 ;
  assign n5157 = n5156 ^ n5152 ;
  assign n5158 = ~n4726 & n5157 ;
  assign n5159 = n5158 ^ n5157 ;
  assign n5160 = n5159 ^ n5152 ;
  assign n5162 = n5161 ^ n5160 ;
  assign n5163 = n4772 & n5162 ;
  assign n5178 = n5163 ^ n5160 ;
  assign n5166 = n5158 ^ n5152 ;
  assign n5167 = n5166 ^ x32 ;
  assign n5168 = ~n4806 & n5167 ;
  assign n5169 = n5168 ^ x32 ;
  assign n5164 = n5163 ^ n5162 ;
  assign n5165 = n5164 ^ n5160 ;
  assign n5170 = n5169 ^ n5165 ;
  assign n5171 = n4850 & n5170 ;
  assign n5177 = n5171 ^ n5165 ;
  assign n5179 = n5178 ^ n5177 ;
  assign n5180 = ~n4893 & n5179 ;
  assign n5187 = n5180 ^ n5177 ;
  assign n5181 = n5180 ^ n5179 ;
  assign n5182 = n5181 ^ n5177 ;
  assign n5172 = n5171 ^ n5170 ;
  assign n5173 = n5172 ^ n5165 ;
  assign n5174 = n5173 ^ x0 ;
  assign n5175 = ~n4927 & n5174 ;
  assign n5176 = n5175 ^ x0 ;
  assign n5183 = n5182 ^ n5176 ;
  assign n5184 = n4972 & n5183 ;
  assign n5185 = n5184 ^ n5183 ;
  assign n5186 = n5185 ^ n5176 ;
  assign n5188 = n5187 ^ n5186 ;
  assign n5189 = n5009 & n5188 ;
  assign n5190 = n5189 ^ n5188 ;
  assign n5191 = n5190 ^ n5186 ;
  assign n5192 = x481 ^ x449 ;
  assign n5193 = n3371 & n5192 ;
  assign n5200 = n5193 ^ x449 ;
  assign n5194 = n5193 ^ n5192 ;
  assign n5195 = n5194 ^ x449 ;
  assign n5196 = n5195 ^ x417 ;
  assign n5197 = n3412 & n5196 ;
  assign n5198 = n5197 ^ n5196 ;
  assign n5199 = n5198 ^ x417 ;
  assign n5201 = n5200 ^ n5199 ;
  assign n5202 = n3451 & n5201 ;
  assign n5217 = n5202 ^ n5199 ;
  assign n5205 = n5197 ^ x417 ;
  assign n5206 = n5205 ^ x385 ;
  assign n5207 = ~n3484 & n5206 ;
  assign n5208 = n5207 ^ x385 ;
  assign n5203 = n5202 ^ n5201 ;
  assign n5204 = n5203 ^ n5199 ;
  assign n5209 = n5208 ^ n5204 ;
  assign n5210 = ~n3527 & n5209 ;
  assign n5216 = n5210 ^ n5204 ;
  assign n5218 = n5217 ^ n5216 ;
  assign n5219 = ~n3570 & n5218 ;
  assign n5220 = n5219 ^ n5218 ;
  assign n5221 = n5220 ^ n5216 ;
  assign n5211 = n5210 ^ n5209 ;
  assign n5212 = n5211 ^ n5204 ;
  assign n5213 = n5212 ^ x353 ;
  assign n5214 = ~n3602 & n5213 ;
  assign n5215 = n5214 ^ x353 ;
  assign n5222 = n5221 ^ n5215 ;
  assign n5223 = ~n3646 & n5222 ;
  assign n5230 = n5223 ^ n5215 ;
  assign n5229 = n5219 ^ n5216 ;
  assign n5231 = n5230 ^ n5229 ;
  assign n5232 = ~n3688 & n5231 ;
  assign n5239 = n5232 ^ n5229 ;
  assign n5233 = n5232 ^ n5231 ;
  assign n5234 = n5233 ^ n5229 ;
  assign n5224 = n5223 ^ n5222 ;
  assign n5225 = n5224 ^ n5215 ;
  assign n5226 = n5225 ^ x321 ;
  assign n5227 = ~n3724 & n5226 ;
  assign n5228 = n5227 ^ x321 ;
  assign n5235 = n5234 ^ n5228 ;
  assign n5236 = n3767 & n5235 ;
  assign n5237 = n5236 ^ n5235 ;
  assign n5238 = n5237 ^ n5228 ;
  assign n5240 = n5239 ^ n5238 ;
  assign n5241 = n3841 & n5240 ;
  assign n5252 = n5241 ^ n5238 ;
  assign n5244 = n5236 ^ n5228 ;
  assign n5245 = n5244 ^ x289 ;
  assign n5246 = ~n3803 & n5245 ;
  assign n5247 = n5246 ^ x289 ;
  assign n5242 = n5241 ^ n5240 ;
  assign n5243 = n5242 ^ n5238 ;
  assign n5248 = n5247 ^ n5243 ;
  assign n5249 = ~n3884 & n5248 ;
  assign n5250 = n5249 ^ n5248 ;
  assign n5251 = n5250 ^ n5243 ;
  assign n5253 = n5252 ^ n5251 ;
  assign n5254 = ~n3927 & n5253 ;
  assign n5269 = n5254 ^ n5251 ;
  assign n5257 = n5249 ^ n5243 ;
  assign n5258 = n5257 ^ x257 ;
  assign n5259 = ~n3959 & n5258 ;
  assign n5260 = n5259 ^ x257 ;
  assign n5255 = n5254 ^ n5253 ;
  assign n5256 = n5255 ^ n5251 ;
  assign n5261 = n5260 ^ n5256 ;
  assign n5262 = n4004 & n5261 ;
  assign n5268 = n5262 ^ n5256 ;
  assign n5270 = n5269 ^ n5268 ;
  assign n5271 = n4046 & n5270 ;
  assign n5278 = n5271 ^ n5268 ;
  assign n5272 = n5271 ^ n5270 ;
  assign n5273 = n5272 ^ n5268 ;
  assign n5263 = n5262 ^ n5261 ;
  assign n5264 = n5263 ^ n5256 ;
  assign n5265 = n5264 ^ x225 ;
  assign n5266 = ~n4083 & n5265 ;
  assign n5267 = n5266 ^ x225 ;
  assign n5274 = n5273 ^ n5267 ;
  assign n5275 = n4127 & n5274 ;
  assign n5276 = n5275 ^ n5274 ;
  assign n5277 = n5276 ^ n5267 ;
  assign n5279 = n5278 ^ n5277 ;
  assign n5280 = n4201 & n5279 ;
  assign n5291 = n5280 ^ n5277 ;
  assign n5283 = n5275 ^ n5267 ;
  assign n5284 = n5283 ^ x193 ;
  assign n5285 = ~n4163 & n5284 ;
  assign n5286 = n5285 ^ x193 ;
  assign n5281 = n5280 ^ n5279 ;
  assign n5282 = n5281 ^ n5277 ;
  assign n5287 = n5286 ^ n5282 ;
  assign n5288 = ~n4245 & n5287 ;
  assign n5289 = n5288 ^ n5287 ;
  assign n5290 = n5289 ^ n5282 ;
  assign n5292 = n5291 ^ n5290 ;
  assign n5293 = ~n4288 & n5292 ;
  assign n5308 = n5293 ^ n5290 ;
  assign n5296 = n5288 ^ n5282 ;
  assign n5297 = n5296 ^ x161 ;
  assign n5298 = ~n4320 & n5297 ;
  assign n5299 = n5298 ^ x161 ;
  assign n5294 = n5293 ^ n5292 ;
  assign n5295 = n5294 ^ n5290 ;
  assign n5300 = n5299 ^ n5295 ;
  assign n5301 = n4365 & n5300 ;
  assign n5307 = n5301 ^ n5295 ;
  assign n5309 = n5308 ^ n5307 ;
  assign n5310 = n4407 & n5309 ;
  assign n5317 = n5310 ^ n5307 ;
  assign n5311 = n5310 ^ n5309 ;
  assign n5312 = n5311 ^ n5307 ;
  assign n5302 = n5301 ^ n5300 ;
  assign n5303 = n5302 ^ n5295 ;
  assign n5304 = n5303 ^ x129 ;
  assign n5305 = ~n4444 & n5304 ;
  assign n5306 = n5305 ^ x129 ;
  assign n5313 = n5312 ^ n5306 ;
  assign n5314 = n4488 & n5313 ;
  assign n5315 = n5314 ^ n5313 ;
  assign n5316 = n5315 ^ n5306 ;
  assign n5318 = n5317 ^ n5316 ;
  assign n5319 = n4562 & n5318 ;
  assign n5330 = n5319 ^ n5316 ;
  assign n5322 = n5314 ^ n5306 ;
  assign n5323 = n5322 ^ x97 ;
  assign n5324 = ~n4524 & n5323 ;
  assign n5325 = n5324 ^ x97 ;
  assign n5320 = n5319 ^ n5318 ;
  assign n5321 = n5320 ^ n5316 ;
  assign n5326 = n5325 ^ n5321 ;
  assign n5327 = ~n4606 & n5326 ;
  assign n5328 = n5327 ^ n5326 ;
  assign n5329 = n5328 ^ n5321 ;
  assign n5331 = n5330 ^ n5329 ;
  assign n5332 = ~n4649 & n5331 ;
  assign n5347 = n5332 ^ n5329 ;
  assign n5335 = n5327 ^ n5321 ;
  assign n5336 = n5335 ^ x65 ;
  assign n5337 = ~n4681 & n5336 ;
  assign n5338 = n5337 ^ x65 ;
  assign n5333 = n5332 ^ n5331 ;
  assign n5334 = n5333 ^ n5329 ;
  assign n5339 = n5338 ^ n5334 ;
  assign n5340 = n4726 & n5339 ;
  assign n5346 = n5340 ^ n5334 ;
  assign n5348 = n5347 ^ n5346 ;
  assign n5349 = n4772 & n5348 ;
  assign n5356 = n5349 ^ n5346 ;
  assign n5350 = n5349 ^ n5348 ;
  assign n5351 = n5350 ^ n5346 ;
  assign n5341 = n5340 ^ n5339 ;
  assign n5342 = n5341 ^ n5334 ;
  assign n5343 = n5342 ^ x33 ;
  assign n5344 = ~n4806 & n5343 ;
  assign n5345 = n5344 ^ x33 ;
  assign n5352 = n5351 ^ n5345 ;
  assign n5353 = n4850 & n5352 ;
  assign n5354 = n5353 ^ n5352 ;
  assign n5355 = n5354 ^ n5345 ;
  assign n5357 = n5356 ^ n5355 ;
  assign n5358 = ~n4893 & n5357 ;
  assign n5369 = n5358 ^ n5355 ;
  assign n5361 = n5353 ^ n5345 ;
  assign n5362 = n5361 ^ x1 ;
  assign n5363 = ~n4927 & n5362 ;
  assign n5364 = n5363 ^ x1 ;
  assign n5359 = n5358 ^ n5357 ;
  assign n5360 = n5359 ^ n5355 ;
  assign n5365 = n5364 ^ n5360 ;
  assign n5366 = ~n4972 & n5365 ;
  assign n5367 = n5366 ^ n5365 ;
  assign n5368 = n5367 ^ n5360 ;
  assign n5370 = n5369 ^ n5368 ;
  assign n5371 = n5009 & n5370 ;
  assign n5372 = n5371 ^ n5370 ;
  assign n5373 = n5372 ^ n5368 ;
  assign n5374 = x482 ^ x450 ;
  assign n5375 = n3371 & n5374 ;
  assign n5382 = n5375 ^ x450 ;
  assign n5376 = n5375 ^ n5374 ;
  assign n5377 = n5376 ^ x450 ;
  assign n5378 = n5377 ^ x418 ;
  assign n5379 = n3412 & n5378 ;
  assign n5380 = n5379 ^ n5378 ;
  assign n5381 = n5380 ^ x418 ;
  assign n5383 = n5382 ^ n5381 ;
  assign n5384 = n3451 & n5383 ;
  assign n5399 = n5384 ^ n5381 ;
  assign n5387 = n5379 ^ x418 ;
  assign n5388 = n5387 ^ x386 ;
  assign n5389 = ~n3484 & n5388 ;
  assign n5390 = n5389 ^ x386 ;
  assign n5385 = n5384 ^ n5383 ;
  assign n5386 = n5385 ^ n5381 ;
  assign n5391 = n5390 ^ n5386 ;
  assign n5392 = ~n3527 & n5391 ;
  assign n5398 = n5392 ^ n5386 ;
  assign n5400 = n5399 ^ n5398 ;
  assign n5401 = ~n3570 & n5400 ;
  assign n5402 = n5401 ^ n5400 ;
  assign n5403 = n5402 ^ n5398 ;
  assign n5393 = n5392 ^ n5391 ;
  assign n5394 = n5393 ^ n5386 ;
  assign n5395 = n5394 ^ x354 ;
  assign n5396 = ~n3602 & n5395 ;
  assign n5397 = n5396 ^ x354 ;
  assign n5404 = n5403 ^ n5397 ;
  assign n5405 = ~n3646 & n5404 ;
  assign n5412 = n5405 ^ n5397 ;
  assign n5411 = n5401 ^ n5398 ;
  assign n5413 = n5412 ^ n5411 ;
  assign n5414 = ~n3688 & n5413 ;
  assign n5421 = n5414 ^ n5411 ;
  assign n5415 = n5414 ^ n5413 ;
  assign n5416 = n5415 ^ n5411 ;
  assign n5406 = n5405 ^ n5404 ;
  assign n5407 = n5406 ^ n5397 ;
  assign n5408 = n5407 ^ x322 ;
  assign n5409 = ~n3724 & n5408 ;
  assign n5410 = n5409 ^ x322 ;
  assign n5417 = n5416 ^ n5410 ;
  assign n5418 = n3767 & n5417 ;
  assign n5419 = n5418 ^ n5417 ;
  assign n5420 = n5419 ^ n5410 ;
  assign n5422 = n5421 ^ n5420 ;
  assign n5423 = n3841 & n5422 ;
  assign n5434 = n5423 ^ n5420 ;
  assign n5426 = n5418 ^ n5410 ;
  assign n5427 = n5426 ^ x290 ;
  assign n5428 = ~n3803 & n5427 ;
  assign n5429 = n5428 ^ x290 ;
  assign n5424 = n5423 ^ n5422 ;
  assign n5425 = n5424 ^ n5420 ;
  assign n5430 = n5429 ^ n5425 ;
  assign n5431 = ~n3884 & n5430 ;
  assign n5432 = n5431 ^ n5430 ;
  assign n5433 = n5432 ^ n5425 ;
  assign n5435 = n5434 ^ n5433 ;
  assign n5436 = ~n3927 & n5435 ;
  assign n5451 = n5436 ^ n5433 ;
  assign n5439 = n5431 ^ n5425 ;
  assign n5440 = n5439 ^ x258 ;
  assign n5441 = ~n3959 & n5440 ;
  assign n5442 = n5441 ^ x258 ;
  assign n5437 = n5436 ^ n5435 ;
  assign n5438 = n5437 ^ n5433 ;
  assign n5443 = n5442 ^ n5438 ;
  assign n5444 = n4004 & n5443 ;
  assign n5450 = n5444 ^ n5438 ;
  assign n5452 = n5451 ^ n5450 ;
  assign n5453 = n4046 & n5452 ;
  assign n5460 = n5453 ^ n5450 ;
  assign n5454 = n5453 ^ n5452 ;
  assign n5455 = n5454 ^ n5450 ;
  assign n5445 = n5444 ^ n5443 ;
  assign n5446 = n5445 ^ n5438 ;
  assign n5447 = n5446 ^ x226 ;
  assign n5448 = ~n4083 & n5447 ;
  assign n5449 = n5448 ^ x226 ;
  assign n5456 = n5455 ^ n5449 ;
  assign n5457 = n4127 & n5456 ;
  assign n5458 = n5457 ^ n5456 ;
  assign n5459 = n5458 ^ n5449 ;
  assign n5461 = n5460 ^ n5459 ;
  assign n5462 = n4201 & n5461 ;
  assign n5473 = n5462 ^ n5459 ;
  assign n5465 = n5457 ^ n5449 ;
  assign n5466 = n5465 ^ x194 ;
  assign n5467 = ~n4163 & n5466 ;
  assign n5468 = n5467 ^ x194 ;
  assign n5463 = n5462 ^ n5461 ;
  assign n5464 = n5463 ^ n5459 ;
  assign n5469 = n5468 ^ n5464 ;
  assign n5470 = ~n4245 & n5469 ;
  assign n5471 = n5470 ^ n5469 ;
  assign n5472 = n5471 ^ n5464 ;
  assign n5474 = n5473 ^ n5472 ;
  assign n5475 = ~n4288 & n5474 ;
  assign n5490 = n5475 ^ n5472 ;
  assign n5478 = n5470 ^ n5464 ;
  assign n5479 = n5478 ^ x162 ;
  assign n5480 = ~n4320 & n5479 ;
  assign n5481 = n5480 ^ x162 ;
  assign n5476 = n5475 ^ n5474 ;
  assign n5477 = n5476 ^ n5472 ;
  assign n5482 = n5481 ^ n5477 ;
  assign n5483 = n4365 & n5482 ;
  assign n5489 = n5483 ^ n5477 ;
  assign n5491 = n5490 ^ n5489 ;
  assign n5492 = n4407 & n5491 ;
  assign n5499 = n5492 ^ n5489 ;
  assign n5493 = n5492 ^ n5491 ;
  assign n5494 = n5493 ^ n5489 ;
  assign n5484 = n5483 ^ n5482 ;
  assign n5485 = n5484 ^ n5477 ;
  assign n5486 = n5485 ^ x130 ;
  assign n5487 = ~n4444 & n5486 ;
  assign n5488 = n5487 ^ x130 ;
  assign n5495 = n5494 ^ n5488 ;
  assign n5496 = n4488 & n5495 ;
  assign n5497 = n5496 ^ n5495 ;
  assign n5498 = n5497 ^ n5488 ;
  assign n5500 = n5499 ^ n5498 ;
  assign n5501 = n4562 & n5500 ;
  assign n5512 = n5501 ^ n5498 ;
  assign n5504 = n5496 ^ n5488 ;
  assign n5505 = n5504 ^ x98 ;
  assign n5506 = ~n4524 & n5505 ;
  assign n5507 = n5506 ^ x98 ;
  assign n5502 = n5501 ^ n5500 ;
  assign n5503 = n5502 ^ n5498 ;
  assign n5508 = n5507 ^ n5503 ;
  assign n5509 = ~n4606 & n5508 ;
  assign n5510 = n5509 ^ n5508 ;
  assign n5511 = n5510 ^ n5503 ;
  assign n5513 = n5512 ^ n5511 ;
  assign n5514 = ~n4649 & n5513 ;
  assign n5529 = n5514 ^ n5511 ;
  assign n5517 = n5509 ^ n5503 ;
  assign n5518 = n5517 ^ x66 ;
  assign n5519 = ~n4681 & n5518 ;
  assign n5520 = n5519 ^ x66 ;
  assign n5515 = n5514 ^ n5513 ;
  assign n5516 = n5515 ^ n5511 ;
  assign n5521 = n5520 ^ n5516 ;
  assign n5522 = n4726 & n5521 ;
  assign n5528 = n5522 ^ n5516 ;
  assign n5530 = n5529 ^ n5528 ;
  assign n5531 = n4772 & n5530 ;
  assign n5538 = n5531 ^ n5528 ;
  assign n5532 = n5531 ^ n5530 ;
  assign n5533 = n5532 ^ n5528 ;
  assign n5523 = n5522 ^ n5521 ;
  assign n5524 = n5523 ^ n5516 ;
  assign n5525 = n5524 ^ x34 ;
  assign n5526 = ~n4806 & n5525 ;
  assign n5527 = n5526 ^ x34 ;
  assign n5534 = n5533 ^ n5527 ;
  assign n5535 = n4850 & n5534 ;
  assign n5536 = n5535 ^ n5534 ;
  assign n5537 = n5536 ^ n5527 ;
  assign n5539 = n5538 ^ n5537 ;
  assign n5540 = ~n4893 & n5539 ;
  assign n5551 = n5540 ^ n5537 ;
  assign n5543 = n5535 ^ n5527 ;
  assign n5544 = n5543 ^ x2 ;
  assign n5545 = ~n4927 & n5544 ;
  assign n5546 = n5545 ^ x2 ;
  assign n5541 = n5540 ^ n5539 ;
  assign n5542 = n5541 ^ n5537 ;
  assign n5547 = n5546 ^ n5542 ;
  assign n5548 = ~n4972 & n5547 ;
  assign n5549 = n5548 ^ n5547 ;
  assign n5550 = n5549 ^ n5542 ;
  assign n5552 = n5551 ^ n5550 ;
  assign n5553 = n5009 & n5552 ;
  assign n5554 = n5553 ^ n5552 ;
  assign n5555 = n5554 ^ n5550 ;
  assign n5556 = x483 ^ x451 ;
  assign n5557 = n3371 & n5556 ;
  assign n5564 = n5557 ^ x451 ;
  assign n5558 = n5557 ^ n5556 ;
  assign n5559 = n5558 ^ x451 ;
  assign n5560 = n5559 ^ x419 ;
  assign n5561 = n3412 & n5560 ;
  assign n5562 = n5561 ^ n5560 ;
  assign n5563 = n5562 ^ x419 ;
  assign n5565 = n5564 ^ n5563 ;
  assign n5566 = n3451 & n5565 ;
  assign n5581 = n5566 ^ n5563 ;
  assign n5569 = n5561 ^ x419 ;
  assign n5570 = n5569 ^ x387 ;
  assign n5571 = ~n3484 & n5570 ;
  assign n5572 = n5571 ^ x387 ;
  assign n5567 = n5566 ^ n5565 ;
  assign n5568 = n5567 ^ n5563 ;
  assign n5573 = n5572 ^ n5568 ;
  assign n5574 = ~n3527 & n5573 ;
  assign n5580 = n5574 ^ n5568 ;
  assign n5582 = n5581 ^ n5580 ;
  assign n5583 = ~n3570 & n5582 ;
  assign n5584 = n5583 ^ n5582 ;
  assign n5585 = n5584 ^ n5580 ;
  assign n5575 = n5574 ^ n5573 ;
  assign n5576 = n5575 ^ n5568 ;
  assign n5577 = n5576 ^ x355 ;
  assign n5578 = ~n3602 & n5577 ;
  assign n5579 = n5578 ^ x355 ;
  assign n5586 = n5585 ^ n5579 ;
  assign n5587 = ~n3646 & n5586 ;
  assign n5594 = n5587 ^ n5579 ;
  assign n5593 = n5583 ^ n5580 ;
  assign n5595 = n5594 ^ n5593 ;
  assign n5596 = ~n3688 & n5595 ;
  assign n5603 = n5596 ^ n5593 ;
  assign n5597 = n5596 ^ n5595 ;
  assign n5598 = n5597 ^ n5593 ;
  assign n5588 = n5587 ^ n5586 ;
  assign n5589 = n5588 ^ n5579 ;
  assign n5590 = n5589 ^ x323 ;
  assign n5591 = ~n3724 & n5590 ;
  assign n5592 = n5591 ^ x323 ;
  assign n5599 = n5598 ^ n5592 ;
  assign n5600 = n3767 & n5599 ;
  assign n5601 = n5600 ^ n5599 ;
  assign n5602 = n5601 ^ n5592 ;
  assign n5604 = n5603 ^ n5602 ;
  assign n5605 = n3841 & n5604 ;
  assign n5616 = n5605 ^ n5602 ;
  assign n5608 = n5600 ^ n5592 ;
  assign n5609 = n5608 ^ x291 ;
  assign n5610 = ~n3803 & n5609 ;
  assign n5611 = n5610 ^ x291 ;
  assign n5606 = n5605 ^ n5604 ;
  assign n5607 = n5606 ^ n5602 ;
  assign n5612 = n5611 ^ n5607 ;
  assign n5613 = ~n3884 & n5612 ;
  assign n5614 = n5613 ^ n5612 ;
  assign n5615 = n5614 ^ n5607 ;
  assign n5617 = n5616 ^ n5615 ;
  assign n5618 = ~n3927 & n5617 ;
  assign n5633 = n5618 ^ n5615 ;
  assign n5621 = n5613 ^ n5607 ;
  assign n5622 = n5621 ^ x259 ;
  assign n5623 = ~n3959 & n5622 ;
  assign n5624 = n5623 ^ x259 ;
  assign n5619 = n5618 ^ n5617 ;
  assign n5620 = n5619 ^ n5615 ;
  assign n5625 = n5624 ^ n5620 ;
  assign n5626 = n4004 & n5625 ;
  assign n5632 = n5626 ^ n5620 ;
  assign n5634 = n5633 ^ n5632 ;
  assign n5635 = n4046 & n5634 ;
  assign n5642 = n5635 ^ n5632 ;
  assign n5636 = n5635 ^ n5634 ;
  assign n5637 = n5636 ^ n5632 ;
  assign n5627 = n5626 ^ n5625 ;
  assign n5628 = n5627 ^ n5620 ;
  assign n5629 = n5628 ^ x227 ;
  assign n5630 = ~n4083 & n5629 ;
  assign n5631 = n5630 ^ x227 ;
  assign n5638 = n5637 ^ n5631 ;
  assign n5639 = n4127 & n5638 ;
  assign n5640 = n5639 ^ n5638 ;
  assign n5641 = n5640 ^ n5631 ;
  assign n5643 = n5642 ^ n5641 ;
  assign n5644 = n4201 & n5643 ;
  assign n5655 = n5644 ^ n5641 ;
  assign n5647 = n5639 ^ n5631 ;
  assign n5648 = n5647 ^ x195 ;
  assign n5649 = ~n4163 & n5648 ;
  assign n5650 = n5649 ^ x195 ;
  assign n5645 = n5644 ^ n5643 ;
  assign n5646 = n5645 ^ n5641 ;
  assign n5651 = n5650 ^ n5646 ;
  assign n5652 = ~n4245 & n5651 ;
  assign n5653 = n5652 ^ n5651 ;
  assign n5654 = n5653 ^ n5646 ;
  assign n5656 = n5655 ^ n5654 ;
  assign n5657 = ~n4288 & n5656 ;
  assign n5672 = n5657 ^ n5654 ;
  assign n5660 = n5652 ^ n5646 ;
  assign n5661 = n5660 ^ x163 ;
  assign n5662 = ~n4320 & n5661 ;
  assign n5663 = n5662 ^ x163 ;
  assign n5658 = n5657 ^ n5656 ;
  assign n5659 = n5658 ^ n5654 ;
  assign n5664 = n5663 ^ n5659 ;
  assign n5665 = n4365 & n5664 ;
  assign n5671 = n5665 ^ n5659 ;
  assign n5673 = n5672 ^ n5671 ;
  assign n5674 = n4407 & n5673 ;
  assign n5681 = n5674 ^ n5671 ;
  assign n5675 = n5674 ^ n5673 ;
  assign n5676 = n5675 ^ n5671 ;
  assign n5666 = n5665 ^ n5664 ;
  assign n5667 = n5666 ^ n5659 ;
  assign n5668 = n5667 ^ x131 ;
  assign n5669 = ~n4444 & n5668 ;
  assign n5670 = n5669 ^ x131 ;
  assign n5677 = n5676 ^ n5670 ;
  assign n5678 = n4488 & n5677 ;
  assign n5679 = n5678 ^ n5677 ;
  assign n5680 = n5679 ^ n5670 ;
  assign n5682 = n5681 ^ n5680 ;
  assign n5683 = n4562 & n5682 ;
  assign n5694 = n5683 ^ n5680 ;
  assign n5686 = n5678 ^ n5670 ;
  assign n5687 = n5686 ^ x99 ;
  assign n5688 = ~n4524 & n5687 ;
  assign n5689 = n5688 ^ x99 ;
  assign n5684 = n5683 ^ n5682 ;
  assign n5685 = n5684 ^ n5680 ;
  assign n5690 = n5689 ^ n5685 ;
  assign n5691 = ~n4606 & n5690 ;
  assign n5692 = n5691 ^ n5690 ;
  assign n5693 = n5692 ^ n5685 ;
  assign n5695 = n5694 ^ n5693 ;
  assign n5696 = ~n4649 & n5695 ;
  assign n5711 = n5696 ^ n5693 ;
  assign n5699 = n5691 ^ n5685 ;
  assign n5700 = n5699 ^ x67 ;
  assign n5701 = ~n4681 & n5700 ;
  assign n5702 = n5701 ^ x67 ;
  assign n5697 = n5696 ^ n5695 ;
  assign n5698 = n5697 ^ n5693 ;
  assign n5703 = n5702 ^ n5698 ;
  assign n5704 = n4726 & n5703 ;
  assign n5710 = n5704 ^ n5698 ;
  assign n5712 = n5711 ^ n5710 ;
  assign n5713 = n4772 & n5712 ;
  assign n5720 = n5713 ^ n5710 ;
  assign n5714 = n5713 ^ n5712 ;
  assign n5715 = n5714 ^ n5710 ;
  assign n5705 = n5704 ^ n5703 ;
  assign n5706 = n5705 ^ n5698 ;
  assign n5707 = n5706 ^ x35 ;
  assign n5708 = ~n4806 & n5707 ;
  assign n5709 = n5708 ^ x35 ;
  assign n5716 = n5715 ^ n5709 ;
  assign n5717 = n4850 & n5716 ;
  assign n5718 = n5717 ^ n5716 ;
  assign n5719 = n5718 ^ n5709 ;
  assign n5721 = n5720 ^ n5719 ;
  assign n5722 = ~n4893 & n5721 ;
  assign n5733 = n5722 ^ n5719 ;
  assign n5725 = n5717 ^ n5709 ;
  assign n5726 = n5725 ^ x3 ;
  assign n5727 = ~n4927 & n5726 ;
  assign n5728 = n5727 ^ x3 ;
  assign n5723 = n5722 ^ n5721 ;
  assign n5724 = n5723 ^ n5719 ;
  assign n5729 = n5728 ^ n5724 ;
  assign n5730 = ~n4972 & n5729 ;
  assign n5731 = n5730 ^ n5729 ;
  assign n5732 = n5731 ^ n5724 ;
  assign n5734 = n5733 ^ n5732 ;
  assign n5735 = n5009 & n5734 ;
  assign n5736 = n5735 ^ n5734 ;
  assign n5737 = n5736 ^ n5732 ;
  assign n5738 = x484 ^ x452 ;
  assign n5739 = n3371 & n5738 ;
  assign n5746 = n5739 ^ x452 ;
  assign n5740 = n5739 ^ n5738 ;
  assign n5741 = n5740 ^ x452 ;
  assign n5742 = n5741 ^ x420 ;
  assign n5743 = n3412 & n5742 ;
  assign n5744 = n5743 ^ n5742 ;
  assign n5745 = n5744 ^ x420 ;
  assign n5747 = n5746 ^ n5745 ;
  assign n5748 = n3451 & n5747 ;
  assign n5763 = n5748 ^ n5745 ;
  assign n5751 = n5743 ^ x420 ;
  assign n5752 = n5751 ^ x388 ;
  assign n5753 = ~n3484 & n5752 ;
  assign n5754 = n5753 ^ x388 ;
  assign n5749 = n5748 ^ n5747 ;
  assign n5750 = n5749 ^ n5745 ;
  assign n5755 = n5754 ^ n5750 ;
  assign n5756 = ~n3527 & n5755 ;
  assign n5762 = n5756 ^ n5750 ;
  assign n5764 = n5763 ^ n5762 ;
  assign n5765 = ~n3570 & n5764 ;
  assign n5766 = n5765 ^ n5764 ;
  assign n5767 = n5766 ^ n5762 ;
  assign n5757 = n5756 ^ n5755 ;
  assign n5758 = n5757 ^ n5750 ;
  assign n5759 = n5758 ^ x356 ;
  assign n5760 = ~n3602 & n5759 ;
  assign n5761 = n5760 ^ x356 ;
  assign n5768 = n5767 ^ n5761 ;
  assign n5769 = ~n3646 & n5768 ;
  assign n5776 = n5769 ^ n5761 ;
  assign n5775 = n5765 ^ n5762 ;
  assign n5777 = n5776 ^ n5775 ;
  assign n5778 = ~n3688 & n5777 ;
  assign n5785 = n5778 ^ n5775 ;
  assign n5779 = n5778 ^ n5777 ;
  assign n5780 = n5779 ^ n5775 ;
  assign n5770 = n5769 ^ n5768 ;
  assign n5771 = n5770 ^ n5761 ;
  assign n5772 = n5771 ^ x324 ;
  assign n5773 = ~n3724 & n5772 ;
  assign n5774 = n5773 ^ x324 ;
  assign n5781 = n5780 ^ n5774 ;
  assign n5782 = n3767 & n5781 ;
  assign n5783 = n5782 ^ n5781 ;
  assign n5784 = n5783 ^ n5774 ;
  assign n5786 = n5785 ^ n5784 ;
  assign n5787 = n3841 & n5786 ;
  assign n5798 = n5787 ^ n5784 ;
  assign n5790 = n5782 ^ n5774 ;
  assign n5791 = n5790 ^ x292 ;
  assign n5792 = ~n3803 & n5791 ;
  assign n5793 = n5792 ^ x292 ;
  assign n5788 = n5787 ^ n5786 ;
  assign n5789 = n5788 ^ n5784 ;
  assign n5794 = n5793 ^ n5789 ;
  assign n5795 = ~n3884 & n5794 ;
  assign n5796 = n5795 ^ n5794 ;
  assign n5797 = n5796 ^ n5789 ;
  assign n5799 = n5798 ^ n5797 ;
  assign n5800 = ~n3927 & n5799 ;
  assign n5815 = n5800 ^ n5797 ;
  assign n5803 = n5795 ^ n5789 ;
  assign n5804 = n5803 ^ x260 ;
  assign n5805 = ~n3959 & n5804 ;
  assign n5806 = n5805 ^ x260 ;
  assign n5801 = n5800 ^ n5799 ;
  assign n5802 = n5801 ^ n5797 ;
  assign n5807 = n5806 ^ n5802 ;
  assign n5808 = n4004 & n5807 ;
  assign n5814 = n5808 ^ n5802 ;
  assign n5816 = n5815 ^ n5814 ;
  assign n5817 = n4046 & n5816 ;
  assign n5824 = n5817 ^ n5814 ;
  assign n5818 = n5817 ^ n5816 ;
  assign n5819 = n5818 ^ n5814 ;
  assign n5809 = n5808 ^ n5807 ;
  assign n5810 = n5809 ^ n5802 ;
  assign n5811 = n5810 ^ x228 ;
  assign n5812 = ~n4083 & n5811 ;
  assign n5813 = n5812 ^ x228 ;
  assign n5820 = n5819 ^ n5813 ;
  assign n5821 = n4127 & n5820 ;
  assign n5822 = n5821 ^ n5820 ;
  assign n5823 = n5822 ^ n5813 ;
  assign n5825 = n5824 ^ n5823 ;
  assign n5826 = n4201 & n5825 ;
  assign n5837 = n5826 ^ n5823 ;
  assign n5829 = n5821 ^ n5813 ;
  assign n5830 = n5829 ^ x196 ;
  assign n5831 = ~n4163 & n5830 ;
  assign n5832 = n5831 ^ x196 ;
  assign n5827 = n5826 ^ n5825 ;
  assign n5828 = n5827 ^ n5823 ;
  assign n5833 = n5832 ^ n5828 ;
  assign n5834 = ~n4245 & n5833 ;
  assign n5835 = n5834 ^ n5833 ;
  assign n5836 = n5835 ^ n5828 ;
  assign n5838 = n5837 ^ n5836 ;
  assign n5839 = ~n4288 & n5838 ;
  assign n5854 = n5839 ^ n5836 ;
  assign n5842 = n5834 ^ n5828 ;
  assign n5843 = n5842 ^ x164 ;
  assign n5844 = ~n4320 & n5843 ;
  assign n5845 = n5844 ^ x164 ;
  assign n5840 = n5839 ^ n5838 ;
  assign n5841 = n5840 ^ n5836 ;
  assign n5846 = n5845 ^ n5841 ;
  assign n5847 = n4365 & n5846 ;
  assign n5853 = n5847 ^ n5841 ;
  assign n5855 = n5854 ^ n5853 ;
  assign n5856 = n4407 & n5855 ;
  assign n5863 = n5856 ^ n5853 ;
  assign n5857 = n5856 ^ n5855 ;
  assign n5858 = n5857 ^ n5853 ;
  assign n5848 = n5847 ^ n5846 ;
  assign n5849 = n5848 ^ n5841 ;
  assign n5850 = n5849 ^ x132 ;
  assign n5851 = ~n4444 & n5850 ;
  assign n5852 = n5851 ^ x132 ;
  assign n5859 = n5858 ^ n5852 ;
  assign n5860 = n4488 & n5859 ;
  assign n5861 = n5860 ^ n5859 ;
  assign n5862 = n5861 ^ n5852 ;
  assign n5864 = n5863 ^ n5862 ;
  assign n5865 = n4562 & n5864 ;
  assign n5876 = n5865 ^ n5862 ;
  assign n5868 = n5860 ^ n5852 ;
  assign n5869 = n5868 ^ x100 ;
  assign n5870 = ~n4524 & n5869 ;
  assign n5871 = n5870 ^ x100 ;
  assign n5866 = n5865 ^ n5864 ;
  assign n5867 = n5866 ^ n5862 ;
  assign n5872 = n5871 ^ n5867 ;
  assign n5873 = ~n4606 & n5872 ;
  assign n5874 = n5873 ^ n5872 ;
  assign n5875 = n5874 ^ n5867 ;
  assign n5877 = n5876 ^ n5875 ;
  assign n5878 = ~n4649 & n5877 ;
  assign n5893 = n5878 ^ n5875 ;
  assign n5881 = n5873 ^ n5867 ;
  assign n5882 = n5881 ^ x68 ;
  assign n5883 = ~n4681 & n5882 ;
  assign n5884 = n5883 ^ x68 ;
  assign n5879 = n5878 ^ n5877 ;
  assign n5880 = n5879 ^ n5875 ;
  assign n5885 = n5884 ^ n5880 ;
  assign n5886 = n4726 & n5885 ;
  assign n5892 = n5886 ^ n5880 ;
  assign n5894 = n5893 ^ n5892 ;
  assign n5895 = n4772 & n5894 ;
  assign n5902 = n5895 ^ n5892 ;
  assign n5896 = n5895 ^ n5894 ;
  assign n5897 = n5896 ^ n5892 ;
  assign n5887 = n5886 ^ n5885 ;
  assign n5888 = n5887 ^ n5880 ;
  assign n5889 = n5888 ^ x36 ;
  assign n5890 = ~n4806 & n5889 ;
  assign n5891 = n5890 ^ x36 ;
  assign n5898 = n5897 ^ n5891 ;
  assign n5899 = n4850 & n5898 ;
  assign n5900 = n5899 ^ n5898 ;
  assign n5901 = n5900 ^ n5891 ;
  assign n5903 = n5902 ^ n5901 ;
  assign n5904 = ~n4893 & n5903 ;
  assign n5915 = n5904 ^ n5901 ;
  assign n5907 = n5899 ^ n5891 ;
  assign n5908 = n5907 ^ x4 ;
  assign n5909 = ~n4927 & n5908 ;
  assign n5910 = n5909 ^ x4 ;
  assign n5905 = n5904 ^ n5903 ;
  assign n5906 = n5905 ^ n5901 ;
  assign n5911 = n5910 ^ n5906 ;
  assign n5912 = ~n4972 & n5911 ;
  assign n5913 = n5912 ^ n5911 ;
  assign n5914 = n5913 ^ n5906 ;
  assign n5916 = n5915 ^ n5914 ;
  assign n5917 = n5009 & n5916 ;
  assign n5918 = n5917 ^ n5916 ;
  assign n5919 = n5918 ^ n5914 ;
  assign n5920 = x485 ^ x453 ;
  assign n5921 = n3371 & n5920 ;
  assign n5928 = n5921 ^ x453 ;
  assign n5922 = n5921 ^ n5920 ;
  assign n5923 = n5922 ^ x453 ;
  assign n5924 = n5923 ^ x421 ;
  assign n5925 = n3412 & n5924 ;
  assign n5926 = n5925 ^ n5924 ;
  assign n5927 = n5926 ^ x421 ;
  assign n5929 = n5928 ^ n5927 ;
  assign n5930 = n3451 & n5929 ;
  assign n5945 = n5930 ^ n5927 ;
  assign n5933 = n5925 ^ x421 ;
  assign n5934 = n5933 ^ x389 ;
  assign n5935 = ~n3484 & n5934 ;
  assign n5936 = n5935 ^ x389 ;
  assign n5931 = n5930 ^ n5929 ;
  assign n5932 = n5931 ^ n5927 ;
  assign n5937 = n5936 ^ n5932 ;
  assign n5938 = ~n3527 & n5937 ;
  assign n5944 = n5938 ^ n5932 ;
  assign n5946 = n5945 ^ n5944 ;
  assign n5947 = ~n3570 & n5946 ;
  assign n5948 = n5947 ^ n5946 ;
  assign n5949 = n5948 ^ n5944 ;
  assign n5939 = n5938 ^ n5937 ;
  assign n5940 = n5939 ^ n5932 ;
  assign n5941 = n5940 ^ x357 ;
  assign n5942 = ~n3602 & n5941 ;
  assign n5943 = n5942 ^ x357 ;
  assign n5950 = n5949 ^ n5943 ;
  assign n5951 = ~n3646 & n5950 ;
  assign n5958 = n5951 ^ n5943 ;
  assign n5957 = n5947 ^ n5944 ;
  assign n5959 = n5958 ^ n5957 ;
  assign n5960 = ~n3688 & n5959 ;
  assign n5967 = n5960 ^ n5957 ;
  assign n5961 = n5960 ^ n5959 ;
  assign n5962 = n5961 ^ n5957 ;
  assign n5952 = n5951 ^ n5950 ;
  assign n5953 = n5952 ^ n5943 ;
  assign n5954 = n5953 ^ x325 ;
  assign n5955 = ~n3724 & n5954 ;
  assign n5956 = n5955 ^ x325 ;
  assign n5963 = n5962 ^ n5956 ;
  assign n5964 = n3767 & n5963 ;
  assign n5965 = n5964 ^ n5963 ;
  assign n5966 = n5965 ^ n5956 ;
  assign n5968 = n5967 ^ n5966 ;
  assign n5969 = n3841 & n5968 ;
  assign n5980 = n5969 ^ n5966 ;
  assign n5972 = n5964 ^ n5956 ;
  assign n5973 = n5972 ^ x293 ;
  assign n5974 = ~n3803 & n5973 ;
  assign n5975 = n5974 ^ x293 ;
  assign n5970 = n5969 ^ n5968 ;
  assign n5971 = n5970 ^ n5966 ;
  assign n5976 = n5975 ^ n5971 ;
  assign n5977 = ~n3884 & n5976 ;
  assign n5978 = n5977 ^ n5976 ;
  assign n5979 = n5978 ^ n5971 ;
  assign n5981 = n5980 ^ n5979 ;
  assign n5982 = ~n3927 & n5981 ;
  assign n5997 = n5982 ^ n5979 ;
  assign n5985 = n5977 ^ n5971 ;
  assign n5986 = n5985 ^ x261 ;
  assign n5987 = ~n3959 & n5986 ;
  assign n5988 = n5987 ^ x261 ;
  assign n5983 = n5982 ^ n5981 ;
  assign n5984 = n5983 ^ n5979 ;
  assign n5989 = n5988 ^ n5984 ;
  assign n5990 = n4004 & n5989 ;
  assign n5996 = n5990 ^ n5984 ;
  assign n5998 = n5997 ^ n5996 ;
  assign n5999 = n4046 & n5998 ;
  assign n6006 = n5999 ^ n5996 ;
  assign n6000 = n5999 ^ n5998 ;
  assign n6001 = n6000 ^ n5996 ;
  assign n5991 = n5990 ^ n5989 ;
  assign n5992 = n5991 ^ n5984 ;
  assign n5993 = n5992 ^ x229 ;
  assign n5994 = ~n4083 & n5993 ;
  assign n5995 = n5994 ^ x229 ;
  assign n6002 = n6001 ^ n5995 ;
  assign n6003 = n4127 & n6002 ;
  assign n6004 = n6003 ^ n6002 ;
  assign n6005 = n6004 ^ n5995 ;
  assign n6007 = n6006 ^ n6005 ;
  assign n6008 = n4201 & n6007 ;
  assign n6019 = n6008 ^ n6005 ;
  assign n6011 = n6003 ^ n5995 ;
  assign n6012 = n6011 ^ x197 ;
  assign n6013 = ~n4163 & n6012 ;
  assign n6014 = n6013 ^ x197 ;
  assign n6009 = n6008 ^ n6007 ;
  assign n6010 = n6009 ^ n6005 ;
  assign n6015 = n6014 ^ n6010 ;
  assign n6016 = ~n4245 & n6015 ;
  assign n6017 = n6016 ^ n6015 ;
  assign n6018 = n6017 ^ n6010 ;
  assign n6020 = n6019 ^ n6018 ;
  assign n6021 = ~n4288 & n6020 ;
  assign n6036 = n6021 ^ n6018 ;
  assign n6024 = n6016 ^ n6010 ;
  assign n6025 = n6024 ^ x165 ;
  assign n6026 = ~n4320 & n6025 ;
  assign n6027 = n6026 ^ x165 ;
  assign n6022 = n6021 ^ n6020 ;
  assign n6023 = n6022 ^ n6018 ;
  assign n6028 = n6027 ^ n6023 ;
  assign n6029 = n4365 & n6028 ;
  assign n6035 = n6029 ^ n6023 ;
  assign n6037 = n6036 ^ n6035 ;
  assign n6038 = n4407 & n6037 ;
  assign n6045 = n6038 ^ n6035 ;
  assign n6039 = n6038 ^ n6037 ;
  assign n6040 = n6039 ^ n6035 ;
  assign n6030 = n6029 ^ n6028 ;
  assign n6031 = n6030 ^ n6023 ;
  assign n6032 = n6031 ^ x133 ;
  assign n6033 = ~n4444 & n6032 ;
  assign n6034 = n6033 ^ x133 ;
  assign n6041 = n6040 ^ n6034 ;
  assign n6042 = n4488 & n6041 ;
  assign n6043 = n6042 ^ n6041 ;
  assign n6044 = n6043 ^ n6034 ;
  assign n6046 = n6045 ^ n6044 ;
  assign n6047 = n4562 & n6046 ;
  assign n6058 = n6047 ^ n6044 ;
  assign n6050 = n6042 ^ n6034 ;
  assign n6051 = n6050 ^ x101 ;
  assign n6052 = ~n4524 & n6051 ;
  assign n6053 = n6052 ^ x101 ;
  assign n6048 = n6047 ^ n6046 ;
  assign n6049 = n6048 ^ n6044 ;
  assign n6054 = n6053 ^ n6049 ;
  assign n6055 = ~n4606 & n6054 ;
  assign n6056 = n6055 ^ n6054 ;
  assign n6057 = n6056 ^ n6049 ;
  assign n6059 = n6058 ^ n6057 ;
  assign n6060 = ~n4649 & n6059 ;
  assign n6075 = n6060 ^ n6057 ;
  assign n6063 = n6055 ^ n6049 ;
  assign n6064 = n6063 ^ x69 ;
  assign n6065 = ~n4681 & n6064 ;
  assign n6066 = n6065 ^ x69 ;
  assign n6061 = n6060 ^ n6059 ;
  assign n6062 = n6061 ^ n6057 ;
  assign n6067 = n6066 ^ n6062 ;
  assign n6068 = n4726 & n6067 ;
  assign n6074 = n6068 ^ n6062 ;
  assign n6076 = n6075 ^ n6074 ;
  assign n6077 = n4772 & n6076 ;
  assign n6084 = n6077 ^ n6074 ;
  assign n6078 = n6077 ^ n6076 ;
  assign n6079 = n6078 ^ n6074 ;
  assign n6069 = n6068 ^ n6067 ;
  assign n6070 = n6069 ^ n6062 ;
  assign n6071 = n6070 ^ x37 ;
  assign n6072 = ~n4806 & n6071 ;
  assign n6073 = n6072 ^ x37 ;
  assign n6080 = n6079 ^ n6073 ;
  assign n6081 = n4850 & n6080 ;
  assign n6082 = n6081 ^ n6080 ;
  assign n6083 = n6082 ^ n6073 ;
  assign n6085 = n6084 ^ n6083 ;
  assign n6086 = ~n4893 & n6085 ;
  assign n6097 = n6086 ^ n6083 ;
  assign n6089 = n6081 ^ n6073 ;
  assign n6090 = n6089 ^ x5 ;
  assign n6091 = ~n4927 & n6090 ;
  assign n6092 = n6091 ^ x5 ;
  assign n6087 = n6086 ^ n6085 ;
  assign n6088 = n6087 ^ n6083 ;
  assign n6093 = n6092 ^ n6088 ;
  assign n6094 = ~n4972 & n6093 ;
  assign n6095 = n6094 ^ n6093 ;
  assign n6096 = n6095 ^ n6088 ;
  assign n6098 = n6097 ^ n6096 ;
  assign n6099 = n5009 & n6098 ;
  assign n6100 = n6099 ^ n6098 ;
  assign n6101 = n6100 ^ n6096 ;
  assign n6102 = x486 ^ x454 ;
  assign n6103 = n3371 & n6102 ;
  assign n6110 = n6103 ^ x454 ;
  assign n6104 = n6103 ^ n6102 ;
  assign n6105 = n6104 ^ x454 ;
  assign n6106 = n6105 ^ x422 ;
  assign n6107 = n3412 & n6106 ;
  assign n6108 = n6107 ^ n6106 ;
  assign n6109 = n6108 ^ x422 ;
  assign n6111 = n6110 ^ n6109 ;
  assign n6112 = n3451 & n6111 ;
  assign n6127 = n6112 ^ n6109 ;
  assign n6115 = n6107 ^ x422 ;
  assign n6116 = n6115 ^ x390 ;
  assign n6117 = ~n3484 & n6116 ;
  assign n6118 = n6117 ^ x390 ;
  assign n6113 = n6112 ^ n6111 ;
  assign n6114 = n6113 ^ n6109 ;
  assign n6119 = n6118 ^ n6114 ;
  assign n6120 = ~n3527 & n6119 ;
  assign n6126 = n6120 ^ n6114 ;
  assign n6128 = n6127 ^ n6126 ;
  assign n6129 = ~n3570 & n6128 ;
  assign n6130 = n6129 ^ n6128 ;
  assign n6131 = n6130 ^ n6126 ;
  assign n6121 = n6120 ^ n6119 ;
  assign n6122 = n6121 ^ n6114 ;
  assign n6123 = n6122 ^ x358 ;
  assign n6124 = ~n3602 & n6123 ;
  assign n6125 = n6124 ^ x358 ;
  assign n6132 = n6131 ^ n6125 ;
  assign n6133 = ~n3646 & n6132 ;
  assign n6140 = n6133 ^ n6125 ;
  assign n6139 = n6129 ^ n6126 ;
  assign n6141 = n6140 ^ n6139 ;
  assign n6142 = ~n3688 & n6141 ;
  assign n6149 = n6142 ^ n6139 ;
  assign n6143 = n6142 ^ n6141 ;
  assign n6144 = n6143 ^ n6139 ;
  assign n6134 = n6133 ^ n6132 ;
  assign n6135 = n6134 ^ n6125 ;
  assign n6136 = n6135 ^ x326 ;
  assign n6137 = ~n3724 & n6136 ;
  assign n6138 = n6137 ^ x326 ;
  assign n6145 = n6144 ^ n6138 ;
  assign n6146 = n3767 & n6145 ;
  assign n6147 = n6146 ^ n6145 ;
  assign n6148 = n6147 ^ n6138 ;
  assign n6150 = n6149 ^ n6148 ;
  assign n6151 = n3841 & n6150 ;
  assign n6162 = n6151 ^ n6148 ;
  assign n6154 = n6146 ^ n6138 ;
  assign n6155 = n6154 ^ x294 ;
  assign n6156 = ~n3803 & n6155 ;
  assign n6157 = n6156 ^ x294 ;
  assign n6152 = n6151 ^ n6150 ;
  assign n6153 = n6152 ^ n6148 ;
  assign n6158 = n6157 ^ n6153 ;
  assign n6159 = ~n3884 & n6158 ;
  assign n6160 = n6159 ^ n6158 ;
  assign n6161 = n6160 ^ n6153 ;
  assign n6163 = n6162 ^ n6161 ;
  assign n6164 = ~n3927 & n6163 ;
  assign n6179 = n6164 ^ n6161 ;
  assign n6167 = n6159 ^ n6153 ;
  assign n6168 = n6167 ^ x262 ;
  assign n6169 = ~n3959 & n6168 ;
  assign n6170 = n6169 ^ x262 ;
  assign n6165 = n6164 ^ n6163 ;
  assign n6166 = n6165 ^ n6161 ;
  assign n6171 = n6170 ^ n6166 ;
  assign n6172 = n4004 & n6171 ;
  assign n6178 = n6172 ^ n6166 ;
  assign n6180 = n6179 ^ n6178 ;
  assign n6181 = n4046 & n6180 ;
  assign n6188 = n6181 ^ n6178 ;
  assign n6182 = n6181 ^ n6180 ;
  assign n6183 = n6182 ^ n6178 ;
  assign n6173 = n6172 ^ n6171 ;
  assign n6174 = n6173 ^ n6166 ;
  assign n6175 = n6174 ^ x230 ;
  assign n6176 = ~n4083 & n6175 ;
  assign n6177 = n6176 ^ x230 ;
  assign n6184 = n6183 ^ n6177 ;
  assign n6185 = n4127 & n6184 ;
  assign n6186 = n6185 ^ n6184 ;
  assign n6187 = n6186 ^ n6177 ;
  assign n6189 = n6188 ^ n6187 ;
  assign n6190 = n4201 & n6189 ;
  assign n6201 = n6190 ^ n6187 ;
  assign n6193 = n6185 ^ n6177 ;
  assign n6194 = n6193 ^ x198 ;
  assign n6195 = ~n4163 & n6194 ;
  assign n6196 = n6195 ^ x198 ;
  assign n6191 = n6190 ^ n6189 ;
  assign n6192 = n6191 ^ n6187 ;
  assign n6197 = n6196 ^ n6192 ;
  assign n6198 = ~n4245 & n6197 ;
  assign n6199 = n6198 ^ n6197 ;
  assign n6200 = n6199 ^ n6192 ;
  assign n6202 = n6201 ^ n6200 ;
  assign n6203 = ~n4288 & n6202 ;
  assign n6218 = n6203 ^ n6200 ;
  assign n6206 = n6198 ^ n6192 ;
  assign n6207 = n6206 ^ x166 ;
  assign n6208 = ~n4320 & n6207 ;
  assign n6209 = n6208 ^ x166 ;
  assign n6204 = n6203 ^ n6202 ;
  assign n6205 = n6204 ^ n6200 ;
  assign n6210 = n6209 ^ n6205 ;
  assign n6211 = n4365 & n6210 ;
  assign n6217 = n6211 ^ n6205 ;
  assign n6219 = n6218 ^ n6217 ;
  assign n6220 = n4407 & n6219 ;
  assign n6227 = n6220 ^ n6217 ;
  assign n6221 = n6220 ^ n6219 ;
  assign n6222 = n6221 ^ n6217 ;
  assign n6212 = n6211 ^ n6210 ;
  assign n6213 = n6212 ^ n6205 ;
  assign n6214 = n6213 ^ x134 ;
  assign n6215 = ~n4444 & n6214 ;
  assign n6216 = n6215 ^ x134 ;
  assign n6223 = n6222 ^ n6216 ;
  assign n6224 = n4488 & n6223 ;
  assign n6225 = n6224 ^ n6223 ;
  assign n6226 = n6225 ^ n6216 ;
  assign n6228 = n6227 ^ n6226 ;
  assign n6229 = n4562 & n6228 ;
  assign n6240 = n6229 ^ n6226 ;
  assign n6232 = n6224 ^ n6216 ;
  assign n6233 = n6232 ^ x102 ;
  assign n6234 = ~n4524 & n6233 ;
  assign n6235 = n6234 ^ x102 ;
  assign n6230 = n6229 ^ n6228 ;
  assign n6231 = n6230 ^ n6226 ;
  assign n6236 = n6235 ^ n6231 ;
  assign n6237 = ~n4606 & n6236 ;
  assign n6238 = n6237 ^ n6236 ;
  assign n6239 = n6238 ^ n6231 ;
  assign n6241 = n6240 ^ n6239 ;
  assign n6242 = ~n4649 & n6241 ;
  assign n6257 = n6242 ^ n6239 ;
  assign n6245 = n6237 ^ n6231 ;
  assign n6246 = n6245 ^ x70 ;
  assign n6247 = ~n4681 & n6246 ;
  assign n6248 = n6247 ^ x70 ;
  assign n6243 = n6242 ^ n6241 ;
  assign n6244 = n6243 ^ n6239 ;
  assign n6249 = n6248 ^ n6244 ;
  assign n6250 = n4726 & n6249 ;
  assign n6256 = n6250 ^ n6244 ;
  assign n6258 = n6257 ^ n6256 ;
  assign n6259 = n4772 & n6258 ;
  assign n6266 = n6259 ^ n6256 ;
  assign n6260 = n6259 ^ n6258 ;
  assign n6261 = n6260 ^ n6256 ;
  assign n6251 = n6250 ^ n6249 ;
  assign n6252 = n6251 ^ n6244 ;
  assign n6253 = n6252 ^ x38 ;
  assign n6254 = ~n4806 & n6253 ;
  assign n6255 = n6254 ^ x38 ;
  assign n6262 = n6261 ^ n6255 ;
  assign n6263 = n4850 & n6262 ;
  assign n6264 = n6263 ^ n6262 ;
  assign n6265 = n6264 ^ n6255 ;
  assign n6267 = n6266 ^ n6265 ;
  assign n6268 = ~n4893 & n6267 ;
  assign n6279 = n6268 ^ n6265 ;
  assign n6271 = n6263 ^ n6255 ;
  assign n6272 = n6271 ^ x6 ;
  assign n6273 = ~n4927 & n6272 ;
  assign n6274 = n6273 ^ x6 ;
  assign n6269 = n6268 ^ n6267 ;
  assign n6270 = n6269 ^ n6265 ;
  assign n6275 = n6274 ^ n6270 ;
  assign n6276 = ~n4972 & n6275 ;
  assign n6277 = n6276 ^ n6275 ;
  assign n6278 = n6277 ^ n6270 ;
  assign n6280 = n6279 ^ n6278 ;
  assign n6281 = n5009 & n6280 ;
  assign n6282 = n6281 ^ n6280 ;
  assign n6283 = n6282 ^ n6278 ;
  assign n6284 = x487 ^ x455 ;
  assign n6285 = n3371 & n6284 ;
  assign n6292 = n6285 ^ x455 ;
  assign n6286 = n6285 ^ n6284 ;
  assign n6287 = n6286 ^ x455 ;
  assign n6288 = n6287 ^ x423 ;
  assign n6289 = n3412 & n6288 ;
  assign n6290 = n6289 ^ n6288 ;
  assign n6291 = n6290 ^ x423 ;
  assign n6293 = n6292 ^ n6291 ;
  assign n6294 = n3451 & n6293 ;
  assign n6309 = n6294 ^ n6291 ;
  assign n6297 = n6289 ^ x423 ;
  assign n6298 = n6297 ^ x391 ;
  assign n6299 = ~n3484 & n6298 ;
  assign n6300 = n6299 ^ x391 ;
  assign n6295 = n6294 ^ n6293 ;
  assign n6296 = n6295 ^ n6291 ;
  assign n6301 = n6300 ^ n6296 ;
  assign n6302 = ~n3527 & n6301 ;
  assign n6308 = n6302 ^ n6296 ;
  assign n6310 = n6309 ^ n6308 ;
  assign n6311 = ~n3570 & n6310 ;
  assign n6312 = n6311 ^ n6310 ;
  assign n6313 = n6312 ^ n6308 ;
  assign n6303 = n6302 ^ n6301 ;
  assign n6304 = n6303 ^ n6296 ;
  assign n6305 = n6304 ^ x359 ;
  assign n6306 = ~n3602 & n6305 ;
  assign n6307 = n6306 ^ x359 ;
  assign n6314 = n6313 ^ n6307 ;
  assign n6315 = ~n3646 & n6314 ;
  assign n6322 = n6315 ^ n6307 ;
  assign n6321 = n6311 ^ n6308 ;
  assign n6323 = n6322 ^ n6321 ;
  assign n6324 = ~n3688 & n6323 ;
  assign n6331 = n6324 ^ n6321 ;
  assign n6325 = n6324 ^ n6323 ;
  assign n6326 = n6325 ^ n6321 ;
  assign n6316 = n6315 ^ n6314 ;
  assign n6317 = n6316 ^ n6307 ;
  assign n6318 = n6317 ^ x327 ;
  assign n6319 = ~n3724 & n6318 ;
  assign n6320 = n6319 ^ x327 ;
  assign n6327 = n6326 ^ n6320 ;
  assign n6328 = n3767 & n6327 ;
  assign n6329 = n6328 ^ n6327 ;
  assign n6330 = n6329 ^ n6320 ;
  assign n6332 = n6331 ^ n6330 ;
  assign n6333 = n3841 & n6332 ;
  assign n6344 = n6333 ^ n6330 ;
  assign n6336 = n6328 ^ n6320 ;
  assign n6337 = n6336 ^ x295 ;
  assign n6338 = ~n3803 & n6337 ;
  assign n6339 = n6338 ^ x295 ;
  assign n6334 = n6333 ^ n6332 ;
  assign n6335 = n6334 ^ n6330 ;
  assign n6340 = n6339 ^ n6335 ;
  assign n6341 = ~n3884 & n6340 ;
  assign n6342 = n6341 ^ n6340 ;
  assign n6343 = n6342 ^ n6335 ;
  assign n6345 = n6344 ^ n6343 ;
  assign n6346 = ~n3927 & n6345 ;
  assign n6361 = n6346 ^ n6343 ;
  assign n6349 = n6341 ^ n6335 ;
  assign n6350 = n6349 ^ x263 ;
  assign n6351 = ~n3959 & n6350 ;
  assign n6352 = n6351 ^ x263 ;
  assign n6347 = n6346 ^ n6345 ;
  assign n6348 = n6347 ^ n6343 ;
  assign n6353 = n6352 ^ n6348 ;
  assign n6354 = n4004 & n6353 ;
  assign n6360 = n6354 ^ n6348 ;
  assign n6362 = n6361 ^ n6360 ;
  assign n6363 = n4046 & n6362 ;
  assign n6370 = n6363 ^ n6360 ;
  assign n6364 = n6363 ^ n6362 ;
  assign n6365 = n6364 ^ n6360 ;
  assign n6355 = n6354 ^ n6353 ;
  assign n6356 = n6355 ^ n6348 ;
  assign n6357 = n6356 ^ x231 ;
  assign n6358 = ~n4083 & n6357 ;
  assign n6359 = n6358 ^ x231 ;
  assign n6366 = n6365 ^ n6359 ;
  assign n6367 = n4127 & n6366 ;
  assign n6368 = n6367 ^ n6366 ;
  assign n6369 = n6368 ^ n6359 ;
  assign n6371 = n6370 ^ n6369 ;
  assign n6372 = n4201 & n6371 ;
  assign n6383 = n6372 ^ n6369 ;
  assign n6375 = n6367 ^ n6359 ;
  assign n6376 = n6375 ^ x199 ;
  assign n6377 = ~n4163 & n6376 ;
  assign n6378 = n6377 ^ x199 ;
  assign n6373 = n6372 ^ n6371 ;
  assign n6374 = n6373 ^ n6369 ;
  assign n6379 = n6378 ^ n6374 ;
  assign n6380 = ~n4245 & n6379 ;
  assign n6381 = n6380 ^ n6379 ;
  assign n6382 = n6381 ^ n6374 ;
  assign n6384 = n6383 ^ n6382 ;
  assign n6385 = ~n4288 & n6384 ;
  assign n6400 = n6385 ^ n6382 ;
  assign n6388 = n6380 ^ n6374 ;
  assign n6389 = n6388 ^ x167 ;
  assign n6390 = ~n4320 & n6389 ;
  assign n6391 = n6390 ^ x167 ;
  assign n6386 = n6385 ^ n6384 ;
  assign n6387 = n6386 ^ n6382 ;
  assign n6392 = n6391 ^ n6387 ;
  assign n6393 = n4365 & n6392 ;
  assign n6399 = n6393 ^ n6387 ;
  assign n6401 = n6400 ^ n6399 ;
  assign n6402 = n4407 & n6401 ;
  assign n6409 = n6402 ^ n6399 ;
  assign n6403 = n6402 ^ n6401 ;
  assign n6404 = n6403 ^ n6399 ;
  assign n6394 = n6393 ^ n6392 ;
  assign n6395 = n6394 ^ n6387 ;
  assign n6396 = n6395 ^ x135 ;
  assign n6397 = ~n4444 & n6396 ;
  assign n6398 = n6397 ^ x135 ;
  assign n6405 = n6404 ^ n6398 ;
  assign n6406 = n4488 & n6405 ;
  assign n6407 = n6406 ^ n6405 ;
  assign n6408 = n6407 ^ n6398 ;
  assign n6410 = n6409 ^ n6408 ;
  assign n6411 = n4562 & n6410 ;
  assign n6422 = n6411 ^ n6408 ;
  assign n6414 = n6406 ^ n6398 ;
  assign n6415 = n6414 ^ x103 ;
  assign n6416 = ~n4524 & n6415 ;
  assign n6417 = n6416 ^ x103 ;
  assign n6412 = n6411 ^ n6410 ;
  assign n6413 = n6412 ^ n6408 ;
  assign n6418 = n6417 ^ n6413 ;
  assign n6419 = ~n4606 & n6418 ;
  assign n6420 = n6419 ^ n6418 ;
  assign n6421 = n6420 ^ n6413 ;
  assign n6423 = n6422 ^ n6421 ;
  assign n6424 = ~n4649 & n6423 ;
  assign n6439 = n6424 ^ n6421 ;
  assign n6427 = n6419 ^ n6413 ;
  assign n6428 = n6427 ^ x71 ;
  assign n6429 = ~n4681 & n6428 ;
  assign n6430 = n6429 ^ x71 ;
  assign n6425 = n6424 ^ n6423 ;
  assign n6426 = n6425 ^ n6421 ;
  assign n6431 = n6430 ^ n6426 ;
  assign n6432 = n4726 & n6431 ;
  assign n6438 = n6432 ^ n6426 ;
  assign n6440 = n6439 ^ n6438 ;
  assign n6441 = n4772 & n6440 ;
  assign n6448 = n6441 ^ n6438 ;
  assign n6442 = n6441 ^ n6440 ;
  assign n6443 = n6442 ^ n6438 ;
  assign n6433 = n6432 ^ n6431 ;
  assign n6434 = n6433 ^ n6426 ;
  assign n6435 = n6434 ^ x39 ;
  assign n6436 = ~n4806 & n6435 ;
  assign n6437 = n6436 ^ x39 ;
  assign n6444 = n6443 ^ n6437 ;
  assign n6445 = n4850 & n6444 ;
  assign n6446 = n6445 ^ n6444 ;
  assign n6447 = n6446 ^ n6437 ;
  assign n6449 = n6448 ^ n6447 ;
  assign n6450 = ~n4893 & n6449 ;
  assign n6461 = n6450 ^ n6447 ;
  assign n6453 = n6445 ^ n6437 ;
  assign n6454 = n6453 ^ x7 ;
  assign n6455 = ~n4927 & n6454 ;
  assign n6456 = n6455 ^ x7 ;
  assign n6451 = n6450 ^ n6449 ;
  assign n6452 = n6451 ^ n6447 ;
  assign n6457 = n6456 ^ n6452 ;
  assign n6458 = ~n4972 & n6457 ;
  assign n6459 = n6458 ^ n6457 ;
  assign n6460 = n6459 ^ n6452 ;
  assign n6462 = n6461 ^ n6460 ;
  assign n6463 = n5009 & n6462 ;
  assign n6464 = n6463 ^ n6462 ;
  assign n6465 = n6464 ^ n6460 ;
  assign n6466 = x488 ^ x456 ;
  assign n6467 = n3371 & n6466 ;
  assign n6474 = n6467 ^ x456 ;
  assign n6468 = n6467 ^ n6466 ;
  assign n6469 = n6468 ^ x456 ;
  assign n6470 = n6469 ^ x424 ;
  assign n6471 = n3412 & n6470 ;
  assign n6472 = n6471 ^ n6470 ;
  assign n6473 = n6472 ^ x424 ;
  assign n6475 = n6474 ^ n6473 ;
  assign n6476 = n3451 & n6475 ;
  assign n6491 = n6476 ^ n6473 ;
  assign n6479 = n6471 ^ x424 ;
  assign n6480 = n6479 ^ x392 ;
  assign n6481 = ~n3484 & n6480 ;
  assign n6482 = n6481 ^ x392 ;
  assign n6477 = n6476 ^ n6475 ;
  assign n6478 = n6477 ^ n6473 ;
  assign n6483 = n6482 ^ n6478 ;
  assign n6484 = ~n3527 & n6483 ;
  assign n6490 = n6484 ^ n6478 ;
  assign n6492 = n6491 ^ n6490 ;
  assign n6493 = ~n3570 & n6492 ;
  assign n6494 = n6493 ^ n6492 ;
  assign n6495 = n6494 ^ n6490 ;
  assign n6485 = n6484 ^ n6483 ;
  assign n6486 = n6485 ^ n6478 ;
  assign n6487 = n6486 ^ x360 ;
  assign n6488 = ~n3602 & n6487 ;
  assign n6489 = n6488 ^ x360 ;
  assign n6496 = n6495 ^ n6489 ;
  assign n6497 = ~n3646 & n6496 ;
  assign n6504 = n6497 ^ n6489 ;
  assign n6503 = n6493 ^ n6490 ;
  assign n6505 = n6504 ^ n6503 ;
  assign n6506 = ~n3688 & n6505 ;
  assign n6513 = n6506 ^ n6503 ;
  assign n6507 = n6506 ^ n6505 ;
  assign n6508 = n6507 ^ n6503 ;
  assign n6498 = n6497 ^ n6496 ;
  assign n6499 = n6498 ^ n6489 ;
  assign n6500 = n6499 ^ x328 ;
  assign n6501 = ~n3724 & n6500 ;
  assign n6502 = n6501 ^ x328 ;
  assign n6509 = n6508 ^ n6502 ;
  assign n6510 = n3767 & n6509 ;
  assign n6511 = n6510 ^ n6509 ;
  assign n6512 = n6511 ^ n6502 ;
  assign n6514 = n6513 ^ n6512 ;
  assign n6515 = n3841 & n6514 ;
  assign n6526 = n6515 ^ n6512 ;
  assign n6518 = n6510 ^ n6502 ;
  assign n6519 = n6518 ^ x296 ;
  assign n6520 = ~n3803 & n6519 ;
  assign n6521 = n6520 ^ x296 ;
  assign n6516 = n6515 ^ n6514 ;
  assign n6517 = n6516 ^ n6512 ;
  assign n6522 = n6521 ^ n6517 ;
  assign n6523 = ~n3884 & n6522 ;
  assign n6524 = n6523 ^ n6522 ;
  assign n6525 = n6524 ^ n6517 ;
  assign n6527 = n6526 ^ n6525 ;
  assign n6528 = ~n3927 & n6527 ;
  assign n6543 = n6528 ^ n6525 ;
  assign n6531 = n6523 ^ n6517 ;
  assign n6532 = n6531 ^ x264 ;
  assign n6533 = ~n3959 & n6532 ;
  assign n6534 = n6533 ^ x264 ;
  assign n6529 = n6528 ^ n6527 ;
  assign n6530 = n6529 ^ n6525 ;
  assign n6535 = n6534 ^ n6530 ;
  assign n6536 = n4004 & n6535 ;
  assign n6542 = n6536 ^ n6530 ;
  assign n6544 = n6543 ^ n6542 ;
  assign n6545 = n4046 & n6544 ;
  assign n6552 = n6545 ^ n6542 ;
  assign n6546 = n6545 ^ n6544 ;
  assign n6547 = n6546 ^ n6542 ;
  assign n6537 = n6536 ^ n6535 ;
  assign n6538 = n6537 ^ n6530 ;
  assign n6539 = n6538 ^ x232 ;
  assign n6540 = ~n4083 & n6539 ;
  assign n6541 = n6540 ^ x232 ;
  assign n6548 = n6547 ^ n6541 ;
  assign n6549 = n4127 & n6548 ;
  assign n6550 = n6549 ^ n6548 ;
  assign n6551 = n6550 ^ n6541 ;
  assign n6553 = n6552 ^ n6551 ;
  assign n6554 = n4201 & n6553 ;
  assign n6565 = n6554 ^ n6551 ;
  assign n6557 = n6549 ^ n6541 ;
  assign n6558 = n6557 ^ x200 ;
  assign n6559 = ~n4163 & n6558 ;
  assign n6560 = n6559 ^ x200 ;
  assign n6555 = n6554 ^ n6553 ;
  assign n6556 = n6555 ^ n6551 ;
  assign n6561 = n6560 ^ n6556 ;
  assign n6562 = ~n4245 & n6561 ;
  assign n6563 = n6562 ^ n6561 ;
  assign n6564 = n6563 ^ n6556 ;
  assign n6566 = n6565 ^ n6564 ;
  assign n6567 = ~n4288 & n6566 ;
  assign n6582 = n6567 ^ n6564 ;
  assign n6570 = n6562 ^ n6556 ;
  assign n6571 = n6570 ^ x168 ;
  assign n6572 = ~n4320 & n6571 ;
  assign n6573 = n6572 ^ x168 ;
  assign n6568 = n6567 ^ n6566 ;
  assign n6569 = n6568 ^ n6564 ;
  assign n6574 = n6573 ^ n6569 ;
  assign n6575 = n4365 & n6574 ;
  assign n6581 = n6575 ^ n6569 ;
  assign n6583 = n6582 ^ n6581 ;
  assign n6584 = n4407 & n6583 ;
  assign n6591 = n6584 ^ n6581 ;
  assign n6585 = n6584 ^ n6583 ;
  assign n6586 = n6585 ^ n6581 ;
  assign n6576 = n6575 ^ n6574 ;
  assign n6577 = n6576 ^ n6569 ;
  assign n6578 = n6577 ^ x136 ;
  assign n6579 = ~n4444 & n6578 ;
  assign n6580 = n6579 ^ x136 ;
  assign n6587 = n6586 ^ n6580 ;
  assign n6588 = n4488 & n6587 ;
  assign n6589 = n6588 ^ n6587 ;
  assign n6590 = n6589 ^ n6580 ;
  assign n6592 = n6591 ^ n6590 ;
  assign n6593 = n4562 & n6592 ;
  assign n6604 = n6593 ^ n6590 ;
  assign n6596 = n6588 ^ n6580 ;
  assign n6597 = n6596 ^ x104 ;
  assign n6598 = ~n4524 & n6597 ;
  assign n6599 = n6598 ^ x104 ;
  assign n6594 = n6593 ^ n6592 ;
  assign n6595 = n6594 ^ n6590 ;
  assign n6600 = n6599 ^ n6595 ;
  assign n6601 = ~n4606 & n6600 ;
  assign n6602 = n6601 ^ n6600 ;
  assign n6603 = n6602 ^ n6595 ;
  assign n6605 = n6604 ^ n6603 ;
  assign n6606 = ~n4649 & n6605 ;
  assign n6621 = n6606 ^ n6603 ;
  assign n6609 = n6601 ^ n6595 ;
  assign n6610 = n6609 ^ x72 ;
  assign n6611 = ~n4681 & n6610 ;
  assign n6612 = n6611 ^ x72 ;
  assign n6607 = n6606 ^ n6605 ;
  assign n6608 = n6607 ^ n6603 ;
  assign n6613 = n6612 ^ n6608 ;
  assign n6614 = n4726 & n6613 ;
  assign n6620 = n6614 ^ n6608 ;
  assign n6622 = n6621 ^ n6620 ;
  assign n6623 = n4772 & n6622 ;
  assign n6630 = n6623 ^ n6620 ;
  assign n6624 = n6623 ^ n6622 ;
  assign n6625 = n6624 ^ n6620 ;
  assign n6615 = n6614 ^ n6613 ;
  assign n6616 = n6615 ^ n6608 ;
  assign n6617 = n6616 ^ x40 ;
  assign n6618 = ~n4806 & n6617 ;
  assign n6619 = n6618 ^ x40 ;
  assign n6626 = n6625 ^ n6619 ;
  assign n6627 = n4850 & n6626 ;
  assign n6628 = n6627 ^ n6626 ;
  assign n6629 = n6628 ^ n6619 ;
  assign n6631 = n6630 ^ n6629 ;
  assign n6632 = ~n4893 & n6631 ;
  assign n6643 = n6632 ^ n6629 ;
  assign n6635 = n6627 ^ n6619 ;
  assign n6636 = n6635 ^ x8 ;
  assign n6637 = ~n4927 & n6636 ;
  assign n6638 = n6637 ^ x8 ;
  assign n6633 = n6632 ^ n6631 ;
  assign n6634 = n6633 ^ n6629 ;
  assign n6639 = n6638 ^ n6634 ;
  assign n6640 = ~n4972 & n6639 ;
  assign n6641 = n6640 ^ n6639 ;
  assign n6642 = n6641 ^ n6634 ;
  assign n6644 = n6643 ^ n6642 ;
  assign n6645 = n5009 & n6644 ;
  assign n6646 = n6645 ^ n6644 ;
  assign n6647 = n6646 ^ n6642 ;
  assign n6648 = x489 ^ x457 ;
  assign n6649 = n3371 & n6648 ;
  assign n6656 = n6649 ^ x457 ;
  assign n6650 = n6649 ^ n6648 ;
  assign n6651 = n6650 ^ x457 ;
  assign n6652 = n6651 ^ x425 ;
  assign n6653 = n3412 & n6652 ;
  assign n6654 = n6653 ^ n6652 ;
  assign n6655 = n6654 ^ x425 ;
  assign n6657 = n6656 ^ n6655 ;
  assign n6658 = n3451 & n6657 ;
  assign n6673 = n6658 ^ n6655 ;
  assign n6661 = n6653 ^ x425 ;
  assign n6662 = n6661 ^ x393 ;
  assign n6663 = ~n3484 & n6662 ;
  assign n6664 = n6663 ^ x393 ;
  assign n6659 = n6658 ^ n6657 ;
  assign n6660 = n6659 ^ n6655 ;
  assign n6665 = n6664 ^ n6660 ;
  assign n6666 = ~n3527 & n6665 ;
  assign n6672 = n6666 ^ n6660 ;
  assign n6674 = n6673 ^ n6672 ;
  assign n6675 = ~n3570 & n6674 ;
  assign n6676 = n6675 ^ n6674 ;
  assign n6677 = n6676 ^ n6672 ;
  assign n6667 = n6666 ^ n6665 ;
  assign n6668 = n6667 ^ n6660 ;
  assign n6669 = n6668 ^ x361 ;
  assign n6670 = ~n3602 & n6669 ;
  assign n6671 = n6670 ^ x361 ;
  assign n6678 = n6677 ^ n6671 ;
  assign n6679 = ~n3646 & n6678 ;
  assign n6686 = n6679 ^ n6671 ;
  assign n6685 = n6675 ^ n6672 ;
  assign n6687 = n6686 ^ n6685 ;
  assign n6688 = ~n3688 & n6687 ;
  assign n6695 = n6688 ^ n6685 ;
  assign n6689 = n6688 ^ n6687 ;
  assign n6690 = n6689 ^ n6685 ;
  assign n6680 = n6679 ^ n6678 ;
  assign n6681 = n6680 ^ n6671 ;
  assign n6682 = n6681 ^ x329 ;
  assign n6683 = ~n3724 & n6682 ;
  assign n6684 = n6683 ^ x329 ;
  assign n6691 = n6690 ^ n6684 ;
  assign n6692 = n3767 & n6691 ;
  assign n6693 = n6692 ^ n6691 ;
  assign n6694 = n6693 ^ n6684 ;
  assign n6696 = n6695 ^ n6694 ;
  assign n6697 = n3841 & n6696 ;
  assign n6708 = n6697 ^ n6694 ;
  assign n6700 = n6692 ^ n6684 ;
  assign n6701 = n6700 ^ x297 ;
  assign n6702 = ~n3803 & n6701 ;
  assign n6703 = n6702 ^ x297 ;
  assign n6698 = n6697 ^ n6696 ;
  assign n6699 = n6698 ^ n6694 ;
  assign n6704 = n6703 ^ n6699 ;
  assign n6705 = ~n3884 & n6704 ;
  assign n6706 = n6705 ^ n6704 ;
  assign n6707 = n6706 ^ n6699 ;
  assign n6709 = n6708 ^ n6707 ;
  assign n6710 = ~n3927 & n6709 ;
  assign n6725 = n6710 ^ n6707 ;
  assign n6713 = n6705 ^ n6699 ;
  assign n6714 = n6713 ^ x265 ;
  assign n6715 = ~n3959 & n6714 ;
  assign n6716 = n6715 ^ x265 ;
  assign n6711 = n6710 ^ n6709 ;
  assign n6712 = n6711 ^ n6707 ;
  assign n6717 = n6716 ^ n6712 ;
  assign n6718 = n4004 & n6717 ;
  assign n6724 = n6718 ^ n6712 ;
  assign n6726 = n6725 ^ n6724 ;
  assign n6727 = n4046 & n6726 ;
  assign n6734 = n6727 ^ n6724 ;
  assign n6728 = n6727 ^ n6726 ;
  assign n6729 = n6728 ^ n6724 ;
  assign n6719 = n6718 ^ n6717 ;
  assign n6720 = n6719 ^ n6712 ;
  assign n6721 = n6720 ^ x233 ;
  assign n6722 = ~n4083 & n6721 ;
  assign n6723 = n6722 ^ x233 ;
  assign n6730 = n6729 ^ n6723 ;
  assign n6731 = n4127 & n6730 ;
  assign n6732 = n6731 ^ n6730 ;
  assign n6733 = n6732 ^ n6723 ;
  assign n6735 = n6734 ^ n6733 ;
  assign n6736 = n4201 & n6735 ;
  assign n6747 = n6736 ^ n6733 ;
  assign n6739 = n6731 ^ n6723 ;
  assign n6740 = n6739 ^ x201 ;
  assign n6741 = ~n4163 & n6740 ;
  assign n6742 = n6741 ^ x201 ;
  assign n6737 = n6736 ^ n6735 ;
  assign n6738 = n6737 ^ n6733 ;
  assign n6743 = n6742 ^ n6738 ;
  assign n6744 = ~n4245 & n6743 ;
  assign n6745 = n6744 ^ n6743 ;
  assign n6746 = n6745 ^ n6738 ;
  assign n6748 = n6747 ^ n6746 ;
  assign n6749 = ~n4288 & n6748 ;
  assign n6764 = n6749 ^ n6746 ;
  assign n6752 = n6744 ^ n6738 ;
  assign n6753 = n6752 ^ x169 ;
  assign n6754 = ~n4320 & n6753 ;
  assign n6755 = n6754 ^ x169 ;
  assign n6750 = n6749 ^ n6748 ;
  assign n6751 = n6750 ^ n6746 ;
  assign n6756 = n6755 ^ n6751 ;
  assign n6757 = n4365 & n6756 ;
  assign n6763 = n6757 ^ n6751 ;
  assign n6765 = n6764 ^ n6763 ;
  assign n6766 = n4407 & n6765 ;
  assign n6773 = n6766 ^ n6763 ;
  assign n6767 = n6766 ^ n6765 ;
  assign n6768 = n6767 ^ n6763 ;
  assign n6758 = n6757 ^ n6756 ;
  assign n6759 = n6758 ^ n6751 ;
  assign n6760 = n6759 ^ x137 ;
  assign n6761 = ~n4444 & n6760 ;
  assign n6762 = n6761 ^ x137 ;
  assign n6769 = n6768 ^ n6762 ;
  assign n6770 = n4488 & n6769 ;
  assign n6771 = n6770 ^ n6769 ;
  assign n6772 = n6771 ^ n6762 ;
  assign n6774 = n6773 ^ n6772 ;
  assign n6775 = n4562 & n6774 ;
  assign n6786 = n6775 ^ n6772 ;
  assign n6778 = n6770 ^ n6762 ;
  assign n6779 = n6778 ^ x105 ;
  assign n6780 = ~n4524 & n6779 ;
  assign n6781 = n6780 ^ x105 ;
  assign n6776 = n6775 ^ n6774 ;
  assign n6777 = n6776 ^ n6772 ;
  assign n6782 = n6781 ^ n6777 ;
  assign n6783 = ~n4606 & n6782 ;
  assign n6784 = n6783 ^ n6782 ;
  assign n6785 = n6784 ^ n6777 ;
  assign n6787 = n6786 ^ n6785 ;
  assign n6788 = ~n4649 & n6787 ;
  assign n6803 = n6788 ^ n6785 ;
  assign n6791 = n6783 ^ n6777 ;
  assign n6792 = n6791 ^ x73 ;
  assign n6793 = ~n4681 & n6792 ;
  assign n6794 = n6793 ^ x73 ;
  assign n6789 = n6788 ^ n6787 ;
  assign n6790 = n6789 ^ n6785 ;
  assign n6795 = n6794 ^ n6790 ;
  assign n6796 = n4726 & n6795 ;
  assign n6802 = n6796 ^ n6790 ;
  assign n6804 = n6803 ^ n6802 ;
  assign n6805 = n4772 & n6804 ;
  assign n6812 = n6805 ^ n6802 ;
  assign n6806 = n6805 ^ n6804 ;
  assign n6807 = n6806 ^ n6802 ;
  assign n6797 = n6796 ^ n6795 ;
  assign n6798 = n6797 ^ n6790 ;
  assign n6799 = n6798 ^ x41 ;
  assign n6800 = ~n4806 & n6799 ;
  assign n6801 = n6800 ^ x41 ;
  assign n6808 = n6807 ^ n6801 ;
  assign n6809 = n4850 & n6808 ;
  assign n6810 = n6809 ^ n6808 ;
  assign n6811 = n6810 ^ n6801 ;
  assign n6813 = n6812 ^ n6811 ;
  assign n6814 = ~n4893 & n6813 ;
  assign n6825 = n6814 ^ n6811 ;
  assign n6817 = n6809 ^ n6801 ;
  assign n6818 = n6817 ^ x9 ;
  assign n6819 = ~n4927 & n6818 ;
  assign n6820 = n6819 ^ x9 ;
  assign n6815 = n6814 ^ n6813 ;
  assign n6816 = n6815 ^ n6811 ;
  assign n6821 = n6820 ^ n6816 ;
  assign n6822 = ~n4972 & n6821 ;
  assign n6823 = n6822 ^ n6821 ;
  assign n6824 = n6823 ^ n6816 ;
  assign n6826 = n6825 ^ n6824 ;
  assign n6827 = n5009 & n6826 ;
  assign n6828 = n6827 ^ n6826 ;
  assign n6829 = n6828 ^ n6824 ;
  assign n6830 = x490 ^ x458 ;
  assign n6831 = n3371 & n6830 ;
  assign n6838 = n6831 ^ x458 ;
  assign n6832 = n6831 ^ n6830 ;
  assign n6833 = n6832 ^ x458 ;
  assign n6834 = n6833 ^ x426 ;
  assign n6835 = n3412 & n6834 ;
  assign n6836 = n6835 ^ n6834 ;
  assign n6837 = n6836 ^ x426 ;
  assign n6839 = n6838 ^ n6837 ;
  assign n6840 = n3451 & n6839 ;
  assign n6855 = n6840 ^ n6837 ;
  assign n6843 = n6835 ^ x426 ;
  assign n6844 = n6843 ^ x394 ;
  assign n6845 = ~n3484 & n6844 ;
  assign n6846 = n6845 ^ x394 ;
  assign n6841 = n6840 ^ n6839 ;
  assign n6842 = n6841 ^ n6837 ;
  assign n6847 = n6846 ^ n6842 ;
  assign n6848 = ~n3527 & n6847 ;
  assign n6854 = n6848 ^ n6842 ;
  assign n6856 = n6855 ^ n6854 ;
  assign n6857 = ~n3570 & n6856 ;
  assign n6858 = n6857 ^ n6856 ;
  assign n6859 = n6858 ^ n6854 ;
  assign n6849 = n6848 ^ n6847 ;
  assign n6850 = n6849 ^ n6842 ;
  assign n6851 = n6850 ^ x362 ;
  assign n6852 = ~n3602 & n6851 ;
  assign n6853 = n6852 ^ x362 ;
  assign n6860 = n6859 ^ n6853 ;
  assign n6861 = ~n3646 & n6860 ;
  assign n6868 = n6861 ^ n6853 ;
  assign n6867 = n6857 ^ n6854 ;
  assign n6869 = n6868 ^ n6867 ;
  assign n6870 = ~n3688 & n6869 ;
  assign n6877 = n6870 ^ n6867 ;
  assign n6871 = n6870 ^ n6869 ;
  assign n6872 = n6871 ^ n6867 ;
  assign n6862 = n6861 ^ n6860 ;
  assign n6863 = n6862 ^ n6853 ;
  assign n6864 = n6863 ^ x330 ;
  assign n6865 = ~n3724 & n6864 ;
  assign n6866 = n6865 ^ x330 ;
  assign n6873 = n6872 ^ n6866 ;
  assign n6874 = n3767 & n6873 ;
  assign n6875 = n6874 ^ n6873 ;
  assign n6876 = n6875 ^ n6866 ;
  assign n6878 = n6877 ^ n6876 ;
  assign n6879 = n3841 & n6878 ;
  assign n6890 = n6879 ^ n6876 ;
  assign n6882 = n6874 ^ n6866 ;
  assign n6883 = n6882 ^ x298 ;
  assign n6884 = ~n3803 & n6883 ;
  assign n6885 = n6884 ^ x298 ;
  assign n6880 = n6879 ^ n6878 ;
  assign n6881 = n6880 ^ n6876 ;
  assign n6886 = n6885 ^ n6881 ;
  assign n6887 = ~n3884 & n6886 ;
  assign n6888 = n6887 ^ n6886 ;
  assign n6889 = n6888 ^ n6881 ;
  assign n6891 = n6890 ^ n6889 ;
  assign n6892 = ~n3927 & n6891 ;
  assign n6907 = n6892 ^ n6889 ;
  assign n6895 = n6887 ^ n6881 ;
  assign n6896 = n6895 ^ x266 ;
  assign n6897 = ~n3959 & n6896 ;
  assign n6898 = n6897 ^ x266 ;
  assign n6893 = n6892 ^ n6891 ;
  assign n6894 = n6893 ^ n6889 ;
  assign n6899 = n6898 ^ n6894 ;
  assign n6900 = n4004 & n6899 ;
  assign n6906 = n6900 ^ n6894 ;
  assign n6908 = n6907 ^ n6906 ;
  assign n6909 = n4046 & n6908 ;
  assign n6916 = n6909 ^ n6906 ;
  assign n6910 = n6909 ^ n6908 ;
  assign n6911 = n6910 ^ n6906 ;
  assign n6901 = n6900 ^ n6899 ;
  assign n6902 = n6901 ^ n6894 ;
  assign n6903 = n6902 ^ x234 ;
  assign n6904 = ~n4083 & n6903 ;
  assign n6905 = n6904 ^ x234 ;
  assign n6912 = n6911 ^ n6905 ;
  assign n6913 = n4127 & n6912 ;
  assign n6914 = n6913 ^ n6912 ;
  assign n6915 = n6914 ^ n6905 ;
  assign n6917 = n6916 ^ n6915 ;
  assign n6918 = n4201 & n6917 ;
  assign n6929 = n6918 ^ n6915 ;
  assign n6921 = n6913 ^ n6905 ;
  assign n6922 = n6921 ^ x202 ;
  assign n6923 = ~n4163 & n6922 ;
  assign n6924 = n6923 ^ x202 ;
  assign n6919 = n6918 ^ n6917 ;
  assign n6920 = n6919 ^ n6915 ;
  assign n6925 = n6924 ^ n6920 ;
  assign n6926 = ~n4245 & n6925 ;
  assign n6927 = n6926 ^ n6925 ;
  assign n6928 = n6927 ^ n6920 ;
  assign n6930 = n6929 ^ n6928 ;
  assign n6931 = ~n4288 & n6930 ;
  assign n6946 = n6931 ^ n6928 ;
  assign n6934 = n6926 ^ n6920 ;
  assign n6935 = n6934 ^ x170 ;
  assign n6936 = ~n4320 & n6935 ;
  assign n6937 = n6936 ^ x170 ;
  assign n6932 = n6931 ^ n6930 ;
  assign n6933 = n6932 ^ n6928 ;
  assign n6938 = n6937 ^ n6933 ;
  assign n6939 = n4365 & n6938 ;
  assign n6945 = n6939 ^ n6933 ;
  assign n6947 = n6946 ^ n6945 ;
  assign n6948 = n4407 & n6947 ;
  assign n6955 = n6948 ^ n6945 ;
  assign n6949 = n6948 ^ n6947 ;
  assign n6950 = n6949 ^ n6945 ;
  assign n6940 = n6939 ^ n6938 ;
  assign n6941 = n6940 ^ n6933 ;
  assign n6942 = n6941 ^ x138 ;
  assign n6943 = ~n4444 & n6942 ;
  assign n6944 = n6943 ^ x138 ;
  assign n6951 = n6950 ^ n6944 ;
  assign n6952 = n4488 & n6951 ;
  assign n6953 = n6952 ^ n6951 ;
  assign n6954 = n6953 ^ n6944 ;
  assign n6956 = n6955 ^ n6954 ;
  assign n6957 = n4562 & n6956 ;
  assign n6968 = n6957 ^ n6954 ;
  assign n6960 = n6952 ^ n6944 ;
  assign n6961 = n6960 ^ x106 ;
  assign n6962 = ~n4524 & n6961 ;
  assign n6963 = n6962 ^ x106 ;
  assign n6958 = n6957 ^ n6956 ;
  assign n6959 = n6958 ^ n6954 ;
  assign n6964 = n6963 ^ n6959 ;
  assign n6965 = ~n4606 & n6964 ;
  assign n6966 = n6965 ^ n6964 ;
  assign n6967 = n6966 ^ n6959 ;
  assign n6969 = n6968 ^ n6967 ;
  assign n6970 = ~n4649 & n6969 ;
  assign n6985 = n6970 ^ n6967 ;
  assign n6973 = n6965 ^ n6959 ;
  assign n6974 = n6973 ^ x74 ;
  assign n6975 = ~n4681 & n6974 ;
  assign n6976 = n6975 ^ x74 ;
  assign n6971 = n6970 ^ n6969 ;
  assign n6972 = n6971 ^ n6967 ;
  assign n6977 = n6976 ^ n6972 ;
  assign n6978 = n4726 & n6977 ;
  assign n6984 = n6978 ^ n6972 ;
  assign n6986 = n6985 ^ n6984 ;
  assign n6987 = n4772 & n6986 ;
  assign n6994 = n6987 ^ n6984 ;
  assign n6988 = n6987 ^ n6986 ;
  assign n6989 = n6988 ^ n6984 ;
  assign n6979 = n6978 ^ n6977 ;
  assign n6980 = n6979 ^ n6972 ;
  assign n6981 = n6980 ^ x42 ;
  assign n6982 = ~n4806 & n6981 ;
  assign n6983 = n6982 ^ x42 ;
  assign n6990 = n6989 ^ n6983 ;
  assign n6991 = n4850 & n6990 ;
  assign n6992 = n6991 ^ n6990 ;
  assign n6993 = n6992 ^ n6983 ;
  assign n6995 = n6994 ^ n6993 ;
  assign n6996 = ~n4893 & n6995 ;
  assign n7007 = n6996 ^ n6993 ;
  assign n6999 = n6991 ^ n6983 ;
  assign n7000 = n6999 ^ x10 ;
  assign n7001 = ~n4927 & n7000 ;
  assign n7002 = n7001 ^ x10 ;
  assign n6997 = n6996 ^ n6995 ;
  assign n6998 = n6997 ^ n6993 ;
  assign n7003 = n7002 ^ n6998 ;
  assign n7004 = ~n4972 & n7003 ;
  assign n7005 = n7004 ^ n7003 ;
  assign n7006 = n7005 ^ n6998 ;
  assign n7008 = n7007 ^ n7006 ;
  assign n7009 = n5009 & n7008 ;
  assign n7010 = n7009 ^ n7008 ;
  assign n7011 = n7010 ^ n7006 ;
  assign n7012 = x491 ^ x459 ;
  assign n7013 = n3371 & n7012 ;
  assign n7020 = n7013 ^ x459 ;
  assign n7014 = n7013 ^ n7012 ;
  assign n7015 = n7014 ^ x459 ;
  assign n7016 = n7015 ^ x427 ;
  assign n7017 = n3412 & n7016 ;
  assign n7018 = n7017 ^ n7016 ;
  assign n7019 = n7018 ^ x427 ;
  assign n7021 = n7020 ^ n7019 ;
  assign n7022 = n3451 & n7021 ;
  assign n7037 = n7022 ^ n7019 ;
  assign n7025 = n7017 ^ x427 ;
  assign n7026 = n7025 ^ x395 ;
  assign n7027 = ~n3484 & n7026 ;
  assign n7028 = n7027 ^ x395 ;
  assign n7023 = n7022 ^ n7021 ;
  assign n7024 = n7023 ^ n7019 ;
  assign n7029 = n7028 ^ n7024 ;
  assign n7030 = ~n3527 & n7029 ;
  assign n7036 = n7030 ^ n7024 ;
  assign n7038 = n7037 ^ n7036 ;
  assign n7039 = ~n3570 & n7038 ;
  assign n7040 = n7039 ^ n7038 ;
  assign n7041 = n7040 ^ n7036 ;
  assign n7031 = n7030 ^ n7029 ;
  assign n7032 = n7031 ^ n7024 ;
  assign n7033 = n7032 ^ x363 ;
  assign n7034 = ~n3602 & n7033 ;
  assign n7035 = n7034 ^ x363 ;
  assign n7042 = n7041 ^ n7035 ;
  assign n7043 = ~n3646 & n7042 ;
  assign n7050 = n7043 ^ n7035 ;
  assign n7049 = n7039 ^ n7036 ;
  assign n7051 = n7050 ^ n7049 ;
  assign n7052 = ~n3688 & n7051 ;
  assign n7059 = n7052 ^ n7049 ;
  assign n7053 = n7052 ^ n7051 ;
  assign n7054 = n7053 ^ n7049 ;
  assign n7044 = n7043 ^ n7042 ;
  assign n7045 = n7044 ^ n7035 ;
  assign n7046 = n7045 ^ x331 ;
  assign n7047 = ~n3724 & n7046 ;
  assign n7048 = n7047 ^ x331 ;
  assign n7055 = n7054 ^ n7048 ;
  assign n7056 = n3767 & n7055 ;
  assign n7057 = n7056 ^ n7055 ;
  assign n7058 = n7057 ^ n7048 ;
  assign n7060 = n7059 ^ n7058 ;
  assign n7061 = n3841 & n7060 ;
  assign n7072 = n7061 ^ n7058 ;
  assign n7064 = n7056 ^ n7048 ;
  assign n7065 = n7064 ^ x299 ;
  assign n7066 = ~n3803 & n7065 ;
  assign n7067 = n7066 ^ x299 ;
  assign n7062 = n7061 ^ n7060 ;
  assign n7063 = n7062 ^ n7058 ;
  assign n7068 = n7067 ^ n7063 ;
  assign n7069 = ~n3884 & n7068 ;
  assign n7070 = n7069 ^ n7068 ;
  assign n7071 = n7070 ^ n7063 ;
  assign n7073 = n7072 ^ n7071 ;
  assign n7074 = ~n3927 & n7073 ;
  assign n7089 = n7074 ^ n7071 ;
  assign n7077 = n7069 ^ n7063 ;
  assign n7078 = n7077 ^ x267 ;
  assign n7079 = ~n3959 & n7078 ;
  assign n7080 = n7079 ^ x267 ;
  assign n7075 = n7074 ^ n7073 ;
  assign n7076 = n7075 ^ n7071 ;
  assign n7081 = n7080 ^ n7076 ;
  assign n7082 = n4004 & n7081 ;
  assign n7088 = n7082 ^ n7076 ;
  assign n7090 = n7089 ^ n7088 ;
  assign n7091 = n4046 & n7090 ;
  assign n7098 = n7091 ^ n7088 ;
  assign n7092 = n7091 ^ n7090 ;
  assign n7093 = n7092 ^ n7088 ;
  assign n7083 = n7082 ^ n7081 ;
  assign n7084 = n7083 ^ n7076 ;
  assign n7085 = n7084 ^ x235 ;
  assign n7086 = ~n4083 & n7085 ;
  assign n7087 = n7086 ^ x235 ;
  assign n7094 = n7093 ^ n7087 ;
  assign n7095 = n4127 & n7094 ;
  assign n7096 = n7095 ^ n7094 ;
  assign n7097 = n7096 ^ n7087 ;
  assign n7099 = n7098 ^ n7097 ;
  assign n7100 = n4201 & n7099 ;
  assign n7111 = n7100 ^ n7097 ;
  assign n7103 = n7095 ^ n7087 ;
  assign n7104 = n7103 ^ x203 ;
  assign n7105 = ~n4163 & n7104 ;
  assign n7106 = n7105 ^ x203 ;
  assign n7101 = n7100 ^ n7099 ;
  assign n7102 = n7101 ^ n7097 ;
  assign n7107 = n7106 ^ n7102 ;
  assign n7108 = ~n4245 & n7107 ;
  assign n7109 = n7108 ^ n7107 ;
  assign n7110 = n7109 ^ n7102 ;
  assign n7112 = n7111 ^ n7110 ;
  assign n7113 = ~n4288 & n7112 ;
  assign n7128 = n7113 ^ n7110 ;
  assign n7116 = n7108 ^ n7102 ;
  assign n7117 = n7116 ^ x171 ;
  assign n7118 = ~n4320 & n7117 ;
  assign n7119 = n7118 ^ x171 ;
  assign n7114 = n7113 ^ n7112 ;
  assign n7115 = n7114 ^ n7110 ;
  assign n7120 = n7119 ^ n7115 ;
  assign n7121 = n4365 & n7120 ;
  assign n7127 = n7121 ^ n7115 ;
  assign n7129 = n7128 ^ n7127 ;
  assign n7130 = n4407 & n7129 ;
  assign n7137 = n7130 ^ n7127 ;
  assign n7131 = n7130 ^ n7129 ;
  assign n7132 = n7131 ^ n7127 ;
  assign n7122 = n7121 ^ n7120 ;
  assign n7123 = n7122 ^ n7115 ;
  assign n7124 = n7123 ^ x139 ;
  assign n7125 = ~n4444 & n7124 ;
  assign n7126 = n7125 ^ x139 ;
  assign n7133 = n7132 ^ n7126 ;
  assign n7134 = n4488 & n7133 ;
  assign n7135 = n7134 ^ n7133 ;
  assign n7136 = n7135 ^ n7126 ;
  assign n7138 = n7137 ^ n7136 ;
  assign n7139 = n4562 & n7138 ;
  assign n7150 = n7139 ^ n7136 ;
  assign n7142 = n7134 ^ n7126 ;
  assign n7143 = n7142 ^ x107 ;
  assign n7144 = ~n4524 & n7143 ;
  assign n7145 = n7144 ^ x107 ;
  assign n7140 = n7139 ^ n7138 ;
  assign n7141 = n7140 ^ n7136 ;
  assign n7146 = n7145 ^ n7141 ;
  assign n7147 = ~n4606 & n7146 ;
  assign n7148 = n7147 ^ n7146 ;
  assign n7149 = n7148 ^ n7141 ;
  assign n7151 = n7150 ^ n7149 ;
  assign n7152 = ~n4649 & n7151 ;
  assign n7167 = n7152 ^ n7149 ;
  assign n7155 = n7147 ^ n7141 ;
  assign n7156 = n7155 ^ x75 ;
  assign n7157 = ~n4681 & n7156 ;
  assign n7158 = n7157 ^ x75 ;
  assign n7153 = n7152 ^ n7151 ;
  assign n7154 = n7153 ^ n7149 ;
  assign n7159 = n7158 ^ n7154 ;
  assign n7160 = n4726 & n7159 ;
  assign n7166 = n7160 ^ n7154 ;
  assign n7168 = n7167 ^ n7166 ;
  assign n7169 = n4772 & n7168 ;
  assign n7176 = n7169 ^ n7166 ;
  assign n7170 = n7169 ^ n7168 ;
  assign n7171 = n7170 ^ n7166 ;
  assign n7161 = n7160 ^ n7159 ;
  assign n7162 = n7161 ^ n7154 ;
  assign n7163 = n7162 ^ x43 ;
  assign n7164 = ~n4806 & n7163 ;
  assign n7165 = n7164 ^ x43 ;
  assign n7172 = n7171 ^ n7165 ;
  assign n7173 = n4850 & n7172 ;
  assign n7174 = n7173 ^ n7172 ;
  assign n7175 = n7174 ^ n7165 ;
  assign n7177 = n7176 ^ n7175 ;
  assign n7178 = ~n4893 & n7177 ;
  assign n7189 = n7178 ^ n7175 ;
  assign n7181 = n7173 ^ n7165 ;
  assign n7182 = n7181 ^ x11 ;
  assign n7183 = ~n4927 & n7182 ;
  assign n7184 = n7183 ^ x11 ;
  assign n7179 = n7178 ^ n7177 ;
  assign n7180 = n7179 ^ n7175 ;
  assign n7185 = n7184 ^ n7180 ;
  assign n7186 = ~n4972 & n7185 ;
  assign n7187 = n7186 ^ n7185 ;
  assign n7188 = n7187 ^ n7180 ;
  assign n7190 = n7189 ^ n7188 ;
  assign n7191 = n5009 & n7190 ;
  assign n7192 = n7191 ^ n7190 ;
  assign n7193 = n7192 ^ n7188 ;
  assign n7194 = x492 ^ x460 ;
  assign n7195 = n3371 & n7194 ;
  assign n7202 = n7195 ^ x460 ;
  assign n7196 = n7195 ^ n7194 ;
  assign n7197 = n7196 ^ x460 ;
  assign n7198 = n7197 ^ x428 ;
  assign n7199 = n3412 & n7198 ;
  assign n7200 = n7199 ^ n7198 ;
  assign n7201 = n7200 ^ x428 ;
  assign n7203 = n7202 ^ n7201 ;
  assign n7204 = n3451 & n7203 ;
  assign n7219 = n7204 ^ n7201 ;
  assign n7207 = n7199 ^ x428 ;
  assign n7208 = n7207 ^ x396 ;
  assign n7209 = ~n3484 & n7208 ;
  assign n7210 = n7209 ^ x396 ;
  assign n7205 = n7204 ^ n7203 ;
  assign n7206 = n7205 ^ n7201 ;
  assign n7211 = n7210 ^ n7206 ;
  assign n7212 = ~n3527 & n7211 ;
  assign n7218 = n7212 ^ n7206 ;
  assign n7220 = n7219 ^ n7218 ;
  assign n7221 = ~n3570 & n7220 ;
  assign n7222 = n7221 ^ n7220 ;
  assign n7223 = n7222 ^ n7218 ;
  assign n7213 = n7212 ^ n7211 ;
  assign n7214 = n7213 ^ n7206 ;
  assign n7215 = n7214 ^ x364 ;
  assign n7216 = ~n3602 & n7215 ;
  assign n7217 = n7216 ^ x364 ;
  assign n7224 = n7223 ^ n7217 ;
  assign n7225 = ~n3646 & n7224 ;
  assign n7232 = n7225 ^ n7217 ;
  assign n7231 = n7221 ^ n7218 ;
  assign n7233 = n7232 ^ n7231 ;
  assign n7234 = ~n3688 & n7233 ;
  assign n7241 = n7234 ^ n7231 ;
  assign n7235 = n7234 ^ n7233 ;
  assign n7236 = n7235 ^ n7231 ;
  assign n7226 = n7225 ^ n7224 ;
  assign n7227 = n7226 ^ n7217 ;
  assign n7228 = n7227 ^ x332 ;
  assign n7229 = ~n3724 & n7228 ;
  assign n7230 = n7229 ^ x332 ;
  assign n7237 = n7236 ^ n7230 ;
  assign n7238 = n3767 & n7237 ;
  assign n7239 = n7238 ^ n7237 ;
  assign n7240 = n7239 ^ n7230 ;
  assign n7242 = n7241 ^ n7240 ;
  assign n7243 = n3841 & n7242 ;
  assign n7254 = n7243 ^ n7240 ;
  assign n7246 = n7238 ^ n7230 ;
  assign n7247 = n7246 ^ x300 ;
  assign n7248 = ~n3803 & n7247 ;
  assign n7249 = n7248 ^ x300 ;
  assign n7244 = n7243 ^ n7242 ;
  assign n7245 = n7244 ^ n7240 ;
  assign n7250 = n7249 ^ n7245 ;
  assign n7251 = ~n3884 & n7250 ;
  assign n7252 = n7251 ^ n7250 ;
  assign n7253 = n7252 ^ n7245 ;
  assign n7255 = n7254 ^ n7253 ;
  assign n7256 = ~n3927 & n7255 ;
  assign n7271 = n7256 ^ n7253 ;
  assign n7259 = n7251 ^ n7245 ;
  assign n7260 = n7259 ^ x268 ;
  assign n7261 = ~n3959 & n7260 ;
  assign n7262 = n7261 ^ x268 ;
  assign n7257 = n7256 ^ n7255 ;
  assign n7258 = n7257 ^ n7253 ;
  assign n7263 = n7262 ^ n7258 ;
  assign n7264 = n4004 & n7263 ;
  assign n7270 = n7264 ^ n7258 ;
  assign n7272 = n7271 ^ n7270 ;
  assign n7273 = n4046 & n7272 ;
  assign n7280 = n7273 ^ n7270 ;
  assign n7274 = n7273 ^ n7272 ;
  assign n7275 = n7274 ^ n7270 ;
  assign n7265 = n7264 ^ n7263 ;
  assign n7266 = n7265 ^ n7258 ;
  assign n7267 = n7266 ^ x236 ;
  assign n7268 = ~n4083 & n7267 ;
  assign n7269 = n7268 ^ x236 ;
  assign n7276 = n7275 ^ n7269 ;
  assign n7277 = n4127 & n7276 ;
  assign n7278 = n7277 ^ n7276 ;
  assign n7279 = n7278 ^ n7269 ;
  assign n7281 = n7280 ^ n7279 ;
  assign n7282 = n4201 & n7281 ;
  assign n7293 = n7282 ^ n7279 ;
  assign n7285 = n7277 ^ n7269 ;
  assign n7286 = n7285 ^ x204 ;
  assign n7287 = ~n4163 & n7286 ;
  assign n7288 = n7287 ^ x204 ;
  assign n7283 = n7282 ^ n7281 ;
  assign n7284 = n7283 ^ n7279 ;
  assign n7289 = n7288 ^ n7284 ;
  assign n7290 = ~n4245 & n7289 ;
  assign n7291 = n7290 ^ n7289 ;
  assign n7292 = n7291 ^ n7284 ;
  assign n7294 = n7293 ^ n7292 ;
  assign n7295 = ~n4288 & n7294 ;
  assign n7310 = n7295 ^ n7292 ;
  assign n7298 = n7290 ^ n7284 ;
  assign n7299 = n7298 ^ x172 ;
  assign n7300 = ~n4320 & n7299 ;
  assign n7301 = n7300 ^ x172 ;
  assign n7296 = n7295 ^ n7294 ;
  assign n7297 = n7296 ^ n7292 ;
  assign n7302 = n7301 ^ n7297 ;
  assign n7303 = n4365 & n7302 ;
  assign n7309 = n7303 ^ n7297 ;
  assign n7311 = n7310 ^ n7309 ;
  assign n7312 = n4407 & n7311 ;
  assign n7319 = n7312 ^ n7309 ;
  assign n7313 = n7312 ^ n7311 ;
  assign n7314 = n7313 ^ n7309 ;
  assign n7304 = n7303 ^ n7302 ;
  assign n7305 = n7304 ^ n7297 ;
  assign n7306 = n7305 ^ x140 ;
  assign n7307 = ~n4444 & n7306 ;
  assign n7308 = n7307 ^ x140 ;
  assign n7315 = n7314 ^ n7308 ;
  assign n7316 = n4488 & n7315 ;
  assign n7317 = n7316 ^ n7315 ;
  assign n7318 = n7317 ^ n7308 ;
  assign n7320 = n7319 ^ n7318 ;
  assign n7321 = n4562 & n7320 ;
  assign n7332 = n7321 ^ n7318 ;
  assign n7324 = n7316 ^ n7308 ;
  assign n7325 = n7324 ^ x108 ;
  assign n7326 = ~n4524 & n7325 ;
  assign n7327 = n7326 ^ x108 ;
  assign n7322 = n7321 ^ n7320 ;
  assign n7323 = n7322 ^ n7318 ;
  assign n7328 = n7327 ^ n7323 ;
  assign n7329 = ~n4606 & n7328 ;
  assign n7330 = n7329 ^ n7328 ;
  assign n7331 = n7330 ^ n7323 ;
  assign n7333 = n7332 ^ n7331 ;
  assign n7334 = ~n4649 & n7333 ;
  assign n7349 = n7334 ^ n7331 ;
  assign n7337 = n7329 ^ n7323 ;
  assign n7338 = n7337 ^ x76 ;
  assign n7339 = ~n4681 & n7338 ;
  assign n7340 = n7339 ^ x76 ;
  assign n7335 = n7334 ^ n7333 ;
  assign n7336 = n7335 ^ n7331 ;
  assign n7341 = n7340 ^ n7336 ;
  assign n7342 = n4726 & n7341 ;
  assign n7348 = n7342 ^ n7336 ;
  assign n7350 = n7349 ^ n7348 ;
  assign n7351 = n4772 & n7350 ;
  assign n7358 = n7351 ^ n7348 ;
  assign n7352 = n7351 ^ n7350 ;
  assign n7353 = n7352 ^ n7348 ;
  assign n7343 = n7342 ^ n7341 ;
  assign n7344 = n7343 ^ n7336 ;
  assign n7345 = n7344 ^ x44 ;
  assign n7346 = ~n4806 & n7345 ;
  assign n7347 = n7346 ^ x44 ;
  assign n7354 = n7353 ^ n7347 ;
  assign n7355 = n4850 & n7354 ;
  assign n7356 = n7355 ^ n7354 ;
  assign n7357 = n7356 ^ n7347 ;
  assign n7359 = n7358 ^ n7357 ;
  assign n7360 = ~n4893 & n7359 ;
  assign n7371 = n7360 ^ n7357 ;
  assign n7363 = n7355 ^ n7347 ;
  assign n7364 = n7363 ^ x12 ;
  assign n7365 = ~n4927 & n7364 ;
  assign n7366 = n7365 ^ x12 ;
  assign n7361 = n7360 ^ n7359 ;
  assign n7362 = n7361 ^ n7357 ;
  assign n7367 = n7366 ^ n7362 ;
  assign n7368 = ~n4972 & n7367 ;
  assign n7369 = n7368 ^ n7367 ;
  assign n7370 = n7369 ^ n7362 ;
  assign n7372 = n7371 ^ n7370 ;
  assign n7373 = n5009 & n7372 ;
  assign n7374 = n7373 ^ n7372 ;
  assign n7375 = n7374 ^ n7370 ;
  assign n7376 = x493 ^ x461 ;
  assign n7377 = n3371 & n7376 ;
  assign n7384 = n7377 ^ x461 ;
  assign n7378 = n7377 ^ n7376 ;
  assign n7379 = n7378 ^ x461 ;
  assign n7380 = n7379 ^ x429 ;
  assign n7381 = n3412 & n7380 ;
  assign n7382 = n7381 ^ n7380 ;
  assign n7383 = n7382 ^ x429 ;
  assign n7385 = n7384 ^ n7383 ;
  assign n7386 = n3451 & n7385 ;
  assign n7401 = n7386 ^ n7383 ;
  assign n7389 = n7381 ^ x429 ;
  assign n7390 = n7389 ^ x397 ;
  assign n7391 = ~n3484 & n7390 ;
  assign n7392 = n7391 ^ x397 ;
  assign n7387 = n7386 ^ n7385 ;
  assign n7388 = n7387 ^ n7383 ;
  assign n7393 = n7392 ^ n7388 ;
  assign n7394 = ~n3527 & n7393 ;
  assign n7400 = n7394 ^ n7388 ;
  assign n7402 = n7401 ^ n7400 ;
  assign n7403 = ~n3570 & n7402 ;
  assign n7404 = n7403 ^ n7402 ;
  assign n7405 = n7404 ^ n7400 ;
  assign n7395 = n7394 ^ n7393 ;
  assign n7396 = n7395 ^ n7388 ;
  assign n7397 = n7396 ^ x365 ;
  assign n7398 = ~n3602 & n7397 ;
  assign n7399 = n7398 ^ x365 ;
  assign n7406 = n7405 ^ n7399 ;
  assign n7407 = ~n3646 & n7406 ;
  assign n7414 = n7407 ^ n7399 ;
  assign n7413 = n7403 ^ n7400 ;
  assign n7415 = n7414 ^ n7413 ;
  assign n7416 = ~n3688 & n7415 ;
  assign n7423 = n7416 ^ n7413 ;
  assign n7417 = n7416 ^ n7415 ;
  assign n7418 = n7417 ^ n7413 ;
  assign n7408 = n7407 ^ n7406 ;
  assign n7409 = n7408 ^ n7399 ;
  assign n7410 = n7409 ^ x333 ;
  assign n7411 = ~n3724 & n7410 ;
  assign n7412 = n7411 ^ x333 ;
  assign n7419 = n7418 ^ n7412 ;
  assign n7420 = n3767 & n7419 ;
  assign n7421 = n7420 ^ n7419 ;
  assign n7422 = n7421 ^ n7412 ;
  assign n7424 = n7423 ^ n7422 ;
  assign n7425 = n3841 & n7424 ;
  assign n7436 = n7425 ^ n7422 ;
  assign n7428 = n7420 ^ n7412 ;
  assign n7429 = n7428 ^ x301 ;
  assign n7430 = ~n3803 & n7429 ;
  assign n7431 = n7430 ^ x301 ;
  assign n7426 = n7425 ^ n7424 ;
  assign n7427 = n7426 ^ n7422 ;
  assign n7432 = n7431 ^ n7427 ;
  assign n7433 = ~n3884 & n7432 ;
  assign n7434 = n7433 ^ n7432 ;
  assign n7435 = n7434 ^ n7427 ;
  assign n7437 = n7436 ^ n7435 ;
  assign n7438 = ~n3927 & n7437 ;
  assign n7453 = n7438 ^ n7435 ;
  assign n7441 = n7433 ^ n7427 ;
  assign n7442 = n7441 ^ x269 ;
  assign n7443 = ~n3959 & n7442 ;
  assign n7444 = n7443 ^ x269 ;
  assign n7439 = n7438 ^ n7437 ;
  assign n7440 = n7439 ^ n7435 ;
  assign n7445 = n7444 ^ n7440 ;
  assign n7446 = n4004 & n7445 ;
  assign n7452 = n7446 ^ n7440 ;
  assign n7454 = n7453 ^ n7452 ;
  assign n7455 = n4046 & n7454 ;
  assign n7462 = n7455 ^ n7452 ;
  assign n7456 = n7455 ^ n7454 ;
  assign n7457 = n7456 ^ n7452 ;
  assign n7447 = n7446 ^ n7445 ;
  assign n7448 = n7447 ^ n7440 ;
  assign n7449 = n7448 ^ x237 ;
  assign n7450 = ~n4083 & n7449 ;
  assign n7451 = n7450 ^ x237 ;
  assign n7458 = n7457 ^ n7451 ;
  assign n7459 = n4127 & n7458 ;
  assign n7460 = n7459 ^ n7458 ;
  assign n7461 = n7460 ^ n7451 ;
  assign n7463 = n7462 ^ n7461 ;
  assign n7464 = n4201 & n7463 ;
  assign n7475 = n7464 ^ n7461 ;
  assign n7467 = n7459 ^ n7451 ;
  assign n7468 = n7467 ^ x205 ;
  assign n7469 = ~n4163 & n7468 ;
  assign n7470 = n7469 ^ x205 ;
  assign n7465 = n7464 ^ n7463 ;
  assign n7466 = n7465 ^ n7461 ;
  assign n7471 = n7470 ^ n7466 ;
  assign n7472 = ~n4245 & n7471 ;
  assign n7473 = n7472 ^ n7471 ;
  assign n7474 = n7473 ^ n7466 ;
  assign n7476 = n7475 ^ n7474 ;
  assign n7477 = ~n4288 & n7476 ;
  assign n7492 = n7477 ^ n7474 ;
  assign n7480 = n7472 ^ n7466 ;
  assign n7481 = n7480 ^ x173 ;
  assign n7482 = ~n4320 & n7481 ;
  assign n7483 = n7482 ^ x173 ;
  assign n7478 = n7477 ^ n7476 ;
  assign n7479 = n7478 ^ n7474 ;
  assign n7484 = n7483 ^ n7479 ;
  assign n7485 = n4365 & n7484 ;
  assign n7491 = n7485 ^ n7479 ;
  assign n7493 = n7492 ^ n7491 ;
  assign n7494 = n4407 & n7493 ;
  assign n7501 = n7494 ^ n7491 ;
  assign n7495 = n7494 ^ n7493 ;
  assign n7496 = n7495 ^ n7491 ;
  assign n7486 = n7485 ^ n7484 ;
  assign n7487 = n7486 ^ n7479 ;
  assign n7488 = n7487 ^ x141 ;
  assign n7489 = ~n4444 & n7488 ;
  assign n7490 = n7489 ^ x141 ;
  assign n7497 = n7496 ^ n7490 ;
  assign n7498 = n4488 & n7497 ;
  assign n7499 = n7498 ^ n7497 ;
  assign n7500 = n7499 ^ n7490 ;
  assign n7502 = n7501 ^ n7500 ;
  assign n7503 = n4562 & n7502 ;
  assign n7514 = n7503 ^ n7500 ;
  assign n7506 = n7498 ^ n7490 ;
  assign n7507 = n7506 ^ x109 ;
  assign n7508 = ~n4524 & n7507 ;
  assign n7509 = n7508 ^ x109 ;
  assign n7504 = n7503 ^ n7502 ;
  assign n7505 = n7504 ^ n7500 ;
  assign n7510 = n7509 ^ n7505 ;
  assign n7511 = ~n4606 & n7510 ;
  assign n7512 = n7511 ^ n7510 ;
  assign n7513 = n7512 ^ n7505 ;
  assign n7515 = n7514 ^ n7513 ;
  assign n7516 = ~n4649 & n7515 ;
  assign n7531 = n7516 ^ n7513 ;
  assign n7519 = n7511 ^ n7505 ;
  assign n7520 = n7519 ^ x77 ;
  assign n7521 = ~n4681 & n7520 ;
  assign n7522 = n7521 ^ x77 ;
  assign n7517 = n7516 ^ n7515 ;
  assign n7518 = n7517 ^ n7513 ;
  assign n7523 = n7522 ^ n7518 ;
  assign n7524 = n4726 & n7523 ;
  assign n7530 = n7524 ^ n7518 ;
  assign n7532 = n7531 ^ n7530 ;
  assign n7533 = n4772 & n7532 ;
  assign n7540 = n7533 ^ n7530 ;
  assign n7534 = n7533 ^ n7532 ;
  assign n7535 = n7534 ^ n7530 ;
  assign n7525 = n7524 ^ n7523 ;
  assign n7526 = n7525 ^ n7518 ;
  assign n7527 = n7526 ^ x45 ;
  assign n7528 = ~n4806 & n7527 ;
  assign n7529 = n7528 ^ x45 ;
  assign n7536 = n7535 ^ n7529 ;
  assign n7537 = n4850 & n7536 ;
  assign n7538 = n7537 ^ n7536 ;
  assign n7539 = n7538 ^ n7529 ;
  assign n7541 = n7540 ^ n7539 ;
  assign n7542 = ~n4893 & n7541 ;
  assign n7553 = n7542 ^ n7539 ;
  assign n7545 = n7537 ^ n7529 ;
  assign n7546 = n7545 ^ x13 ;
  assign n7547 = ~n4927 & n7546 ;
  assign n7548 = n7547 ^ x13 ;
  assign n7543 = n7542 ^ n7541 ;
  assign n7544 = n7543 ^ n7539 ;
  assign n7549 = n7548 ^ n7544 ;
  assign n7550 = ~n4972 & n7549 ;
  assign n7551 = n7550 ^ n7549 ;
  assign n7552 = n7551 ^ n7544 ;
  assign n7554 = n7553 ^ n7552 ;
  assign n7555 = n5009 & n7554 ;
  assign n7556 = n7555 ^ n7554 ;
  assign n7557 = n7556 ^ n7552 ;
  assign n7558 = x494 ^ x462 ;
  assign n7559 = n3371 & n7558 ;
  assign n7566 = n7559 ^ x462 ;
  assign n7560 = n7559 ^ n7558 ;
  assign n7561 = n7560 ^ x462 ;
  assign n7562 = n7561 ^ x430 ;
  assign n7563 = n3412 & n7562 ;
  assign n7564 = n7563 ^ n7562 ;
  assign n7565 = n7564 ^ x430 ;
  assign n7567 = n7566 ^ n7565 ;
  assign n7568 = n3451 & n7567 ;
  assign n7583 = n7568 ^ n7565 ;
  assign n7571 = n7563 ^ x430 ;
  assign n7572 = n7571 ^ x398 ;
  assign n7573 = ~n3484 & n7572 ;
  assign n7574 = n7573 ^ x398 ;
  assign n7569 = n7568 ^ n7567 ;
  assign n7570 = n7569 ^ n7565 ;
  assign n7575 = n7574 ^ n7570 ;
  assign n7576 = ~n3527 & n7575 ;
  assign n7582 = n7576 ^ n7570 ;
  assign n7584 = n7583 ^ n7582 ;
  assign n7585 = ~n3570 & n7584 ;
  assign n7586 = n7585 ^ n7584 ;
  assign n7587 = n7586 ^ n7582 ;
  assign n7577 = n7576 ^ n7575 ;
  assign n7578 = n7577 ^ n7570 ;
  assign n7579 = n7578 ^ x366 ;
  assign n7580 = ~n3602 & n7579 ;
  assign n7581 = n7580 ^ x366 ;
  assign n7588 = n7587 ^ n7581 ;
  assign n7589 = ~n3646 & n7588 ;
  assign n7596 = n7589 ^ n7581 ;
  assign n7595 = n7585 ^ n7582 ;
  assign n7597 = n7596 ^ n7595 ;
  assign n7598 = ~n3688 & n7597 ;
  assign n7605 = n7598 ^ n7595 ;
  assign n7599 = n7598 ^ n7597 ;
  assign n7600 = n7599 ^ n7595 ;
  assign n7590 = n7589 ^ n7588 ;
  assign n7591 = n7590 ^ n7581 ;
  assign n7592 = n7591 ^ x334 ;
  assign n7593 = ~n3724 & n7592 ;
  assign n7594 = n7593 ^ x334 ;
  assign n7601 = n7600 ^ n7594 ;
  assign n7602 = n3767 & n7601 ;
  assign n7603 = n7602 ^ n7601 ;
  assign n7604 = n7603 ^ n7594 ;
  assign n7606 = n7605 ^ n7604 ;
  assign n7607 = n3841 & n7606 ;
  assign n7618 = n7607 ^ n7604 ;
  assign n7610 = n7602 ^ n7594 ;
  assign n7611 = n7610 ^ x302 ;
  assign n7612 = ~n3803 & n7611 ;
  assign n7613 = n7612 ^ x302 ;
  assign n7608 = n7607 ^ n7606 ;
  assign n7609 = n7608 ^ n7604 ;
  assign n7614 = n7613 ^ n7609 ;
  assign n7615 = ~n3884 & n7614 ;
  assign n7616 = n7615 ^ n7614 ;
  assign n7617 = n7616 ^ n7609 ;
  assign n7619 = n7618 ^ n7617 ;
  assign n7620 = ~n3927 & n7619 ;
  assign n7635 = n7620 ^ n7617 ;
  assign n7623 = n7615 ^ n7609 ;
  assign n7624 = n7623 ^ x270 ;
  assign n7625 = ~n3959 & n7624 ;
  assign n7626 = n7625 ^ x270 ;
  assign n7621 = n7620 ^ n7619 ;
  assign n7622 = n7621 ^ n7617 ;
  assign n7627 = n7626 ^ n7622 ;
  assign n7628 = n4004 & n7627 ;
  assign n7634 = n7628 ^ n7622 ;
  assign n7636 = n7635 ^ n7634 ;
  assign n7637 = n4046 & n7636 ;
  assign n7644 = n7637 ^ n7634 ;
  assign n7638 = n7637 ^ n7636 ;
  assign n7639 = n7638 ^ n7634 ;
  assign n7629 = n7628 ^ n7627 ;
  assign n7630 = n7629 ^ n7622 ;
  assign n7631 = n7630 ^ x238 ;
  assign n7632 = ~n4083 & n7631 ;
  assign n7633 = n7632 ^ x238 ;
  assign n7640 = n7639 ^ n7633 ;
  assign n7641 = n4127 & n7640 ;
  assign n7642 = n7641 ^ n7640 ;
  assign n7643 = n7642 ^ n7633 ;
  assign n7645 = n7644 ^ n7643 ;
  assign n7646 = n4201 & n7645 ;
  assign n7657 = n7646 ^ n7643 ;
  assign n7649 = n7641 ^ n7633 ;
  assign n7650 = n7649 ^ x206 ;
  assign n7651 = ~n4163 & n7650 ;
  assign n7652 = n7651 ^ x206 ;
  assign n7647 = n7646 ^ n7645 ;
  assign n7648 = n7647 ^ n7643 ;
  assign n7653 = n7652 ^ n7648 ;
  assign n7654 = ~n4245 & n7653 ;
  assign n7655 = n7654 ^ n7653 ;
  assign n7656 = n7655 ^ n7648 ;
  assign n7658 = n7657 ^ n7656 ;
  assign n7659 = ~n4288 & n7658 ;
  assign n7674 = n7659 ^ n7656 ;
  assign n7662 = n7654 ^ n7648 ;
  assign n7663 = n7662 ^ x174 ;
  assign n7664 = ~n4320 & n7663 ;
  assign n7665 = n7664 ^ x174 ;
  assign n7660 = n7659 ^ n7658 ;
  assign n7661 = n7660 ^ n7656 ;
  assign n7666 = n7665 ^ n7661 ;
  assign n7667 = n4365 & n7666 ;
  assign n7673 = n7667 ^ n7661 ;
  assign n7675 = n7674 ^ n7673 ;
  assign n7676 = n4407 & n7675 ;
  assign n7683 = n7676 ^ n7673 ;
  assign n7677 = n7676 ^ n7675 ;
  assign n7678 = n7677 ^ n7673 ;
  assign n7668 = n7667 ^ n7666 ;
  assign n7669 = n7668 ^ n7661 ;
  assign n7670 = n7669 ^ x142 ;
  assign n7671 = ~n4444 & n7670 ;
  assign n7672 = n7671 ^ x142 ;
  assign n7679 = n7678 ^ n7672 ;
  assign n7680 = n4488 & n7679 ;
  assign n7681 = n7680 ^ n7679 ;
  assign n7682 = n7681 ^ n7672 ;
  assign n7684 = n7683 ^ n7682 ;
  assign n7685 = n4562 & n7684 ;
  assign n7696 = n7685 ^ n7682 ;
  assign n7688 = n7680 ^ n7672 ;
  assign n7689 = n7688 ^ x110 ;
  assign n7690 = ~n4524 & n7689 ;
  assign n7691 = n7690 ^ x110 ;
  assign n7686 = n7685 ^ n7684 ;
  assign n7687 = n7686 ^ n7682 ;
  assign n7692 = n7691 ^ n7687 ;
  assign n7693 = ~n4606 & n7692 ;
  assign n7694 = n7693 ^ n7692 ;
  assign n7695 = n7694 ^ n7687 ;
  assign n7697 = n7696 ^ n7695 ;
  assign n7698 = ~n4649 & n7697 ;
  assign n7713 = n7698 ^ n7695 ;
  assign n7701 = n7693 ^ n7687 ;
  assign n7702 = n7701 ^ x78 ;
  assign n7703 = ~n4681 & n7702 ;
  assign n7704 = n7703 ^ x78 ;
  assign n7699 = n7698 ^ n7697 ;
  assign n7700 = n7699 ^ n7695 ;
  assign n7705 = n7704 ^ n7700 ;
  assign n7706 = n4726 & n7705 ;
  assign n7712 = n7706 ^ n7700 ;
  assign n7714 = n7713 ^ n7712 ;
  assign n7715 = n4772 & n7714 ;
  assign n7722 = n7715 ^ n7712 ;
  assign n7716 = n7715 ^ n7714 ;
  assign n7717 = n7716 ^ n7712 ;
  assign n7707 = n7706 ^ n7705 ;
  assign n7708 = n7707 ^ n7700 ;
  assign n7709 = n7708 ^ x46 ;
  assign n7710 = ~n4806 & n7709 ;
  assign n7711 = n7710 ^ x46 ;
  assign n7718 = n7717 ^ n7711 ;
  assign n7719 = n4850 & n7718 ;
  assign n7720 = n7719 ^ n7718 ;
  assign n7721 = n7720 ^ n7711 ;
  assign n7723 = n7722 ^ n7721 ;
  assign n7724 = ~n4893 & n7723 ;
  assign n7735 = n7724 ^ n7721 ;
  assign n7727 = n7719 ^ n7711 ;
  assign n7728 = n7727 ^ x14 ;
  assign n7729 = ~n4927 & n7728 ;
  assign n7730 = n7729 ^ x14 ;
  assign n7725 = n7724 ^ n7723 ;
  assign n7726 = n7725 ^ n7721 ;
  assign n7731 = n7730 ^ n7726 ;
  assign n7732 = ~n4972 & n7731 ;
  assign n7733 = n7732 ^ n7731 ;
  assign n7734 = n7733 ^ n7726 ;
  assign n7736 = n7735 ^ n7734 ;
  assign n7737 = n5009 & n7736 ;
  assign n7738 = n7737 ^ n7736 ;
  assign n7739 = n7738 ^ n7734 ;
  assign n7740 = x495 ^ x463 ;
  assign n7741 = n3371 & n7740 ;
  assign n7748 = n7741 ^ x463 ;
  assign n7742 = n7741 ^ n7740 ;
  assign n7743 = n7742 ^ x463 ;
  assign n7744 = n7743 ^ x431 ;
  assign n7745 = n3412 & n7744 ;
  assign n7746 = n7745 ^ n7744 ;
  assign n7747 = n7746 ^ x431 ;
  assign n7749 = n7748 ^ n7747 ;
  assign n7750 = n3451 & n7749 ;
  assign n7765 = n7750 ^ n7747 ;
  assign n7753 = n7745 ^ x431 ;
  assign n7754 = n7753 ^ x399 ;
  assign n7755 = ~n3484 & n7754 ;
  assign n7756 = n7755 ^ x399 ;
  assign n7751 = n7750 ^ n7749 ;
  assign n7752 = n7751 ^ n7747 ;
  assign n7757 = n7756 ^ n7752 ;
  assign n7758 = ~n3527 & n7757 ;
  assign n7764 = n7758 ^ n7752 ;
  assign n7766 = n7765 ^ n7764 ;
  assign n7767 = ~n3570 & n7766 ;
  assign n7768 = n7767 ^ n7766 ;
  assign n7769 = n7768 ^ n7764 ;
  assign n7759 = n7758 ^ n7757 ;
  assign n7760 = n7759 ^ n7752 ;
  assign n7761 = n7760 ^ x367 ;
  assign n7762 = ~n3602 & n7761 ;
  assign n7763 = n7762 ^ x367 ;
  assign n7770 = n7769 ^ n7763 ;
  assign n7771 = ~n3646 & n7770 ;
  assign n7778 = n7771 ^ n7763 ;
  assign n7777 = n7767 ^ n7764 ;
  assign n7779 = n7778 ^ n7777 ;
  assign n7780 = ~n3688 & n7779 ;
  assign n7787 = n7780 ^ n7777 ;
  assign n7781 = n7780 ^ n7779 ;
  assign n7782 = n7781 ^ n7777 ;
  assign n7772 = n7771 ^ n7770 ;
  assign n7773 = n7772 ^ n7763 ;
  assign n7774 = n7773 ^ x335 ;
  assign n7775 = ~n3724 & n7774 ;
  assign n7776 = n7775 ^ x335 ;
  assign n7783 = n7782 ^ n7776 ;
  assign n7784 = n3767 & n7783 ;
  assign n7785 = n7784 ^ n7783 ;
  assign n7786 = n7785 ^ n7776 ;
  assign n7788 = n7787 ^ n7786 ;
  assign n7789 = n3841 & n7788 ;
  assign n7800 = n7789 ^ n7786 ;
  assign n7792 = n7784 ^ n7776 ;
  assign n7793 = n7792 ^ x303 ;
  assign n7794 = ~n3803 & n7793 ;
  assign n7795 = n7794 ^ x303 ;
  assign n7790 = n7789 ^ n7788 ;
  assign n7791 = n7790 ^ n7786 ;
  assign n7796 = n7795 ^ n7791 ;
  assign n7797 = ~n3884 & n7796 ;
  assign n7798 = n7797 ^ n7796 ;
  assign n7799 = n7798 ^ n7791 ;
  assign n7801 = n7800 ^ n7799 ;
  assign n7802 = ~n3927 & n7801 ;
  assign n7817 = n7802 ^ n7799 ;
  assign n7805 = n7797 ^ n7791 ;
  assign n7806 = n7805 ^ x271 ;
  assign n7807 = ~n3959 & n7806 ;
  assign n7808 = n7807 ^ x271 ;
  assign n7803 = n7802 ^ n7801 ;
  assign n7804 = n7803 ^ n7799 ;
  assign n7809 = n7808 ^ n7804 ;
  assign n7810 = n4004 & n7809 ;
  assign n7816 = n7810 ^ n7804 ;
  assign n7818 = n7817 ^ n7816 ;
  assign n7819 = n4046 & n7818 ;
  assign n7826 = n7819 ^ n7816 ;
  assign n7820 = n7819 ^ n7818 ;
  assign n7821 = n7820 ^ n7816 ;
  assign n7811 = n7810 ^ n7809 ;
  assign n7812 = n7811 ^ n7804 ;
  assign n7813 = n7812 ^ x239 ;
  assign n7814 = ~n4083 & n7813 ;
  assign n7815 = n7814 ^ x239 ;
  assign n7822 = n7821 ^ n7815 ;
  assign n7823 = n4127 & n7822 ;
  assign n7824 = n7823 ^ n7822 ;
  assign n7825 = n7824 ^ n7815 ;
  assign n7827 = n7826 ^ n7825 ;
  assign n7828 = n4201 & n7827 ;
  assign n7839 = n7828 ^ n7825 ;
  assign n7831 = n7823 ^ n7815 ;
  assign n7832 = n7831 ^ x207 ;
  assign n7833 = ~n4163 & n7832 ;
  assign n7834 = n7833 ^ x207 ;
  assign n7829 = n7828 ^ n7827 ;
  assign n7830 = n7829 ^ n7825 ;
  assign n7835 = n7834 ^ n7830 ;
  assign n7836 = ~n4245 & n7835 ;
  assign n7837 = n7836 ^ n7835 ;
  assign n7838 = n7837 ^ n7830 ;
  assign n7840 = n7839 ^ n7838 ;
  assign n7841 = ~n4288 & n7840 ;
  assign n7856 = n7841 ^ n7838 ;
  assign n7844 = n7836 ^ n7830 ;
  assign n7845 = n7844 ^ x175 ;
  assign n7846 = ~n4320 & n7845 ;
  assign n7847 = n7846 ^ x175 ;
  assign n7842 = n7841 ^ n7840 ;
  assign n7843 = n7842 ^ n7838 ;
  assign n7848 = n7847 ^ n7843 ;
  assign n7849 = n4365 & n7848 ;
  assign n7855 = n7849 ^ n7843 ;
  assign n7857 = n7856 ^ n7855 ;
  assign n7858 = n4407 & n7857 ;
  assign n7865 = n7858 ^ n7855 ;
  assign n7859 = n7858 ^ n7857 ;
  assign n7860 = n7859 ^ n7855 ;
  assign n7850 = n7849 ^ n7848 ;
  assign n7851 = n7850 ^ n7843 ;
  assign n7852 = n7851 ^ x143 ;
  assign n7853 = ~n4444 & n7852 ;
  assign n7854 = n7853 ^ x143 ;
  assign n7861 = n7860 ^ n7854 ;
  assign n7862 = n4488 & n7861 ;
  assign n7863 = n7862 ^ n7861 ;
  assign n7864 = n7863 ^ n7854 ;
  assign n7866 = n7865 ^ n7864 ;
  assign n7867 = n4562 & n7866 ;
  assign n7878 = n7867 ^ n7864 ;
  assign n7870 = n7862 ^ n7854 ;
  assign n7871 = n7870 ^ x111 ;
  assign n7872 = ~n4524 & n7871 ;
  assign n7873 = n7872 ^ x111 ;
  assign n7868 = n7867 ^ n7866 ;
  assign n7869 = n7868 ^ n7864 ;
  assign n7874 = n7873 ^ n7869 ;
  assign n7875 = ~n4606 & n7874 ;
  assign n7876 = n7875 ^ n7874 ;
  assign n7877 = n7876 ^ n7869 ;
  assign n7879 = n7878 ^ n7877 ;
  assign n7880 = ~n4649 & n7879 ;
  assign n7895 = n7880 ^ n7877 ;
  assign n7883 = n7875 ^ n7869 ;
  assign n7884 = n7883 ^ x79 ;
  assign n7885 = ~n4681 & n7884 ;
  assign n7886 = n7885 ^ x79 ;
  assign n7881 = n7880 ^ n7879 ;
  assign n7882 = n7881 ^ n7877 ;
  assign n7887 = n7886 ^ n7882 ;
  assign n7888 = n4726 & n7887 ;
  assign n7894 = n7888 ^ n7882 ;
  assign n7896 = n7895 ^ n7894 ;
  assign n7897 = n4772 & n7896 ;
  assign n7904 = n7897 ^ n7894 ;
  assign n7898 = n7897 ^ n7896 ;
  assign n7899 = n7898 ^ n7894 ;
  assign n7889 = n7888 ^ n7887 ;
  assign n7890 = n7889 ^ n7882 ;
  assign n7891 = n7890 ^ x47 ;
  assign n7892 = ~n4806 & n7891 ;
  assign n7893 = n7892 ^ x47 ;
  assign n7900 = n7899 ^ n7893 ;
  assign n7901 = n4850 & n7900 ;
  assign n7902 = n7901 ^ n7900 ;
  assign n7903 = n7902 ^ n7893 ;
  assign n7905 = n7904 ^ n7903 ;
  assign n7906 = ~n4893 & n7905 ;
  assign n7917 = n7906 ^ n7903 ;
  assign n7909 = n7901 ^ n7893 ;
  assign n7910 = n7909 ^ x15 ;
  assign n7911 = ~n4927 & n7910 ;
  assign n7912 = n7911 ^ x15 ;
  assign n7907 = n7906 ^ n7905 ;
  assign n7908 = n7907 ^ n7903 ;
  assign n7913 = n7912 ^ n7908 ;
  assign n7914 = ~n4972 & n7913 ;
  assign n7915 = n7914 ^ n7913 ;
  assign n7916 = n7915 ^ n7908 ;
  assign n7918 = n7917 ^ n7916 ;
  assign n7919 = n5009 & n7918 ;
  assign n7920 = n7919 ^ n7918 ;
  assign n7921 = n7920 ^ n7916 ;
  assign n7922 = x496 ^ x464 ;
  assign n7923 = n3371 & n7922 ;
  assign n7930 = n7923 ^ x464 ;
  assign n7924 = n7923 ^ n7922 ;
  assign n7925 = n7924 ^ x464 ;
  assign n7926 = n7925 ^ x432 ;
  assign n7927 = n3412 & n7926 ;
  assign n7928 = n7927 ^ n7926 ;
  assign n7929 = n7928 ^ x432 ;
  assign n7931 = n7930 ^ n7929 ;
  assign n7932 = n3451 & n7931 ;
  assign n7947 = n7932 ^ n7929 ;
  assign n7935 = n7927 ^ x432 ;
  assign n7936 = n7935 ^ x400 ;
  assign n7937 = ~n3484 & n7936 ;
  assign n7938 = n7937 ^ x400 ;
  assign n7933 = n7932 ^ n7931 ;
  assign n7934 = n7933 ^ n7929 ;
  assign n7939 = n7938 ^ n7934 ;
  assign n7940 = ~n3527 & n7939 ;
  assign n7946 = n7940 ^ n7934 ;
  assign n7948 = n7947 ^ n7946 ;
  assign n7949 = ~n3570 & n7948 ;
  assign n7950 = n7949 ^ n7948 ;
  assign n7951 = n7950 ^ n7946 ;
  assign n7941 = n7940 ^ n7939 ;
  assign n7942 = n7941 ^ n7934 ;
  assign n7943 = n7942 ^ x368 ;
  assign n7944 = ~n3602 & n7943 ;
  assign n7945 = n7944 ^ x368 ;
  assign n7952 = n7951 ^ n7945 ;
  assign n7953 = ~n3646 & n7952 ;
  assign n7960 = n7953 ^ n7945 ;
  assign n7959 = n7949 ^ n7946 ;
  assign n7961 = n7960 ^ n7959 ;
  assign n7962 = ~n3688 & n7961 ;
  assign n7969 = n7962 ^ n7959 ;
  assign n7963 = n7962 ^ n7961 ;
  assign n7964 = n7963 ^ n7959 ;
  assign n7954 = n7953 ^ n7952 ;
  assign n7955 = n7954 ^ n7945 ;
  assign n7956 = n7955 ^ x336 ;
  assign n7957 = ~n3724 & n7956 ;
  assign n7958 = n7957 ^ x336 ;
  assign n7965 = n7964 ^ n7958 ;
  assign n7966 = n3767 & n7965 ;
  assign n7967 = n7966 ^ n7965 ;
  assign n7968 = n7967 ^ n7958 ;
  assign n7970 = n7969 ^ n7968 ;
  assign n7971 = n3841 & n7970 ;
  assign n7982 = n7971 ^ n7968 ;
  assign n7974 = n7966 ^ n7958 ;
  assign n7975 = n7974 ^ x304 ;
  assign n7976 = ~n3803 & n7975 ;
  assign n7977 = n7976 ^ x304 ;
  assign n7972 = n7971 ^ n7970 ;
  assign n7973 = n7972 ^ n7968 ;
  assign n7978 = n7977 ^ n7973 ;
  assign n7979 = ~n3884 & n7978 ;
  assign n7980 = n7979 ^ n7978 ;
  assign n7981 = n7980 ^ n7973 ;
  assign n7983 = n7982 ^ n7981 ;
  assign n7984 = ~n3927 & n7983 ;
  assign n7999 = n7984 ^ n7981 ;
  assign n7987 = n7979 ^ n7973 ;
  assign n7988 = n7987 ^ x272 ;
  assign n7989 = ~n3959 & n7988 ;
  assign n7990 = n7989 ^ x272 ;
  assign n7985 = n7984 ^ n7983 ;
  assign n7986 = n7985 ^ n7981 ;
  assign n7991 = n7990 ^ n7986 ;
  assign n7992 = n4004 & n7991 ;
  assign n7998 = n7992 ^ n7986 ;
  assign n8000 = n7999 ^ n7998 ;
  assign n8001 = n4046 & n8000 ;
  assign n8008 = n8001 ^ n7998 ;
  assign n8002 = n8001 ^ n8000 ;
  assign n8003 = n8002 ^ n7998 ;
  assign n7993 = n7992 ^ n7991 ;
  assign n7994 = n7993 ^ n7986 ;
  assign n7995 = n7994 ^ x240 ;
  assign n7996 = ~n4083 & n7995 ;
  assign n7997 = n7996 ^ x240 ;
  assign n8004 = n8003 ^ n7997 ;
  assign n8005 = n4127 & n8004 ;
  assign n8006 = n8005 ^ n8004 ;
  assign n8007 = n8006 ^ n7997 ;
  assign n8009 = n8008 ^ n8007 ;
  assign n8010 = n4201 & n8009 ;
  assign n8021 = n8010 ^ n8007 ;
  assign n8013 = n8005 ^ n7997 ;
  assign n8014 = n8013 ^ x208 ;
  assign n8015 = ~n4163 & n8014 ;
  assign n8016 = n8015 ^ x208 ;
  assign n8011 = n8010 ^ n8009 ;
  assign n8012 = n8011 ^ n8007 ;
  assign n8017 = n8016 ^ n8012 ;
  assign n8018 = ~n4245 & n8017 ;
  assign n8019 = n8018 ^ n8017 ;
  assign n8020 = n8019 ^ n8012 ;
  assign n8022 = n8021 ^ n8020 ;
  assign n8023 = ~n4288 & n8022 ;
  assign n8038 = n8023 ^ n8020 ;
  assign n8026 = n8018 ^ n8012 ;
  assign n8027 = n8026 ^ x176 ;
  assign n8028 = ~n4320 & n8027 ;
  assign n8029 = n8028 ^ x176 ;
  assign n8024 = n8023 ^ n8022 ;
  assign n8025 = n8024 ^ n8020 ;
  assign n8030 = n8029 ^ n8025 ;
  assign n8031 = n4365 & n8030 ;
  assign n8037 = n8031 ^ n8025 ;
  assign n8039 = n8038 ^ n8037 ;
  assign n8040 = n4407 & n8039 ;
  assign n8047 = n8040 ^ n8037 ;
  assign n8041 = n8040 ^ n8039 ;
  assign n8042 = n8041 ^ n8037 ;
  assign n8032 = n8031 ^ n8030 ;
  assign n8033 = n8032 ^ n8025 ;
  assign n8034 = n8033 ^ x144 ;
  assign n8035 = ~n4444 & n8034 ;
  assign n8036 = n8035 ^ x144 ;
  assign n8043 = n8042 ^ n8036 ;
  assign n8044 = n4488 & n8043 ;
  assign n8045 = n8044 ^ n8043 ;
  assign n8046 = n8045 ^ n8036 ;
  assign n8048 = n8047 ^ n8046 ;
  assign n8049 = n4562 & n8048 ;
  assign n8060 = n8049 ^ n8046 ;
  assign n8052 = n8044 ^ n8036 ;
  assign n8053 = n8052 ^ x112 ;
  assign n8054 = ~n4524 & n8053 ;
  assign n8055 = n8054 ^ x112 ;
  assign n8050 = n8049 ^ n8048 ;
  assign n8051 = n8050 ^ n8046 ;
  assign n8056 = n8055 ^ n8051 ;
  assign n8057 = ~n4606 & n8056 ;
  assign n8058 = n8057 ^ n8056 ;
  assign n8059 = n8058 ^ n8051 ;
  assign n8061 = n8060 ^ n8059 ;
  assign n8062 = ~n4649 & n8061 ;
  assign n8077 = n8062 ^ n8059 ;
  assign n8065 = n8057 ^ n8051 ;
  assign n8066 = n8065 ^ x80 ;
  assign n8067 = ~n4681 & n8066 ;
  assign n8068 = n8067 ^ x80 ;
  assign n8063 = n8062 ^ n8061 ;
  assign n8064 = n8063 ^ n8059 ;
  assign n8069 = n8068 ^ n8064 ;
  assign n8070 = n4726 & n8069 ;
  assign n8076 = n8070 ^ n8064 ;
  assign n8078 = n8077 ^ n8076 ;
  assign n8079 = n4772 & n8078 ;
  assign n8086 = n8079 ^ n8076 ;
  assign n8080 = n8079 ^ n8078 ;
  assign n8081 = n8080 ^ n8076 ;
  assign n8071 = n8070 ^ n8069 ;
  assign n8072 = n8071 ^ n8064 ;
  assign n8073 = n8072 ^ x48 ;
  assign n8074 = ~n4806 & n8073 ;
  assign n8075 = n8074 ^ x48 ;
  assign n8082 = n8081 ^ n8075 ;
  assign n8083 = n4850 & n8082 ;
  assign n8084 = n8083 ^ n8082 ;
  assign n8085 = n8084 ^ n8075 ;
  assign n8087 = n8086 ^ n8085 ;
  assign n8088 = ~n4893 & n8087 ;
  assign n8099 = n8088 ^ n8085 ;
  assign n8091 = n8083 ^ n8075 ;
  assign n8092 = n8091 ^ x16 ;
  assign n8093 = ~n4927 & n8092 ;
  assign n8094 = n8093 ^ x16 ;
  assign n8089 = n8088 ^ n8087 ;
  assign n8090 = n8089 ^ n8085 ;
  assign n8095 = n8094 ^ n8090 ;
  assign n8096 = ~n4972 & n8095 ;
  assign n8097 = n8096 ^ n8095 ;
  assign n8098 = n8097 ^ n8090 ;
  assign n8100 = n8099 ^ n8098 ;
  assign n8101 = n5009 & n8100 ;
  assign n8102 = n8101 ^ n8100 ;
  assign n8103 = n8102 ^ n8098 ;
  assign n8104 = x497 ^ x465 ;
  assign n8105 = n3371 & n8104 ;
  assign n8112 = n8105 ^ x465 ;
  assign n8106 = n8105 ^ n8104 ;
  assign n8107 = n8106 ^ x465 ;
  assign n8108 = n8107 ^ x433 ;
  assign n8109 = n3412 & n8108 ;
  assign n8110 = n8109 ^ n8108 ;
  assign n8111 = n8110 ^ x433 ;
  assign n8113 = n8112 ^ n8111 ;
  assign n8114 = n3451 & n8113 ;
  assign n8129 = n8114 ^ n8111 ;
  assign n8117 = n8109 ^ x433 ;
  assign n8118 = n8117 ^ x401 ;
  assign n8119 = ~n3484 & n8118 ;
  assign n8120 = n8119 ^ x401 ;
  assign n8115 = n8114 ^ n8113 ;
  assign n8116 = n8115 ^ n8111 ;
  assign n8121 = n8120 ^ n8116 ;
  assign n8122 = ~n3527 & n8121 ;
  assign n8128 = n8122 ^ n8116 ;
  assign n8130 = n8129 ^ n8128 ;
  assign n8131 = ~n3570 & n8130 ;
  assign n8132 = n8131 ^ n8130 ;
  assign n8133 = n8132 ^ n8128 ;
  assign n8123 = n8122 ^ n8121 ;
  assign n8124 = n8123 ^ n8116 ;
  assign n8125 = n8124 ^ x369 ;
  assign n8126 = ~n3602 & n8125 ;
  assign n8127 = n8126 ^ x369 ;
  assign n8134 = n8133 ^ n8127 ;
  assign n8135 = ~n3646 & n8134 ;
  assign n8142 = n8135 ^ n8127 ;
  assign n8141 = n8131 ^ n8128 ;
  assign n8143 = n8142 ^ n8141 ;
  assign n8144 = ~n3688 & n8143 ;
  assign n8151 = n8144 ^ n8141 ;
  assign n8145 = n8144 ^ n8143 ;
  assign n8146 = n8145 ^ n8141 ;
  assign n8136 = n8135 ^ n8134 ;
  assign n8137 = n8136 ^ n8127 ;
  assign n8138 = n8137 ^ x337 ;
  assign n8139 = ~n3724 & n8138 ;
  assign n8140 = n8139 ^ x337 ;
  assign n8147 = n8146 ^ n8140 ;
  assign n8148 = n3767 & n8147 ;
  assign n8149 = n8148 ^ n8147 ;
  assign n8150 = n8149 ^ n8140 ;
  assign n8152 = n8151 ^ n8150 ;
  assign n8153 = n3841 & n8152 ;
  assign n8164 = n8153 ^ n8150 ;
  assign n8156 = n8148 ^ n8140 ;
  assign n8157 = n8156 ^ x305 ;
  assign n8158 = ~n3803 & n8157 ;
  assign n8159 = n8158 ^ x305 ;
  assign n8154 = n8153 ^ n8152 ;
  assign n8155 = n8154 ^ n8150 ;
  assign n8160 = n8159 ^ n8155 ;
  assign n8161 = ~n3884 & n8160 ;
  assign n8162 = n8161 ^ n8160 ;
  assign n8163 = n8162 ^ n8155 ;
  assign n8165 = n8164 ^ n8163 ;
  assign n8166 = ~n3927 & n8165 ;
  assign n8181 = n8166 ^ n8163 ;
  assign n8169 = n8161 ^ n8155 ;
  assign n8170 = n8169 ^ x273 ;
  assign n8171 = ~n3959 & n8170 ;
  assign n8172 = n8171 ^ x273 ;
  assign n8167 = n8166 ^ n8165 ;
  assign n8168 = n8167 ^ n8163 ;
  assign n8173 = n8172 ^ n8168 ;
  assign n8174 = n4004 & n8173 ;
  assign n8180 = n8174 ^ n8168 ;
  assign n8182 = n8181 ^ n8180 ;
  assign n8183 = n4046 & n8182 ;
  assign n8190 = n8183 ^ n8180 ;
  assign n8184 = n8183 ^ n8182 ;
  assign n8185 = n8184 ^ n8180 ;
  assign n8175 = n8174 ^ n8173 ;
  assign n8176 = n8175 ^ n8168 ;
  assign n8177 = n8176 ^ x241 ;
  assign n8178 = ~n4083 & n8177 ;
  assign n8179 = n8178 ^ x241 ;
  assign n8186 = n8185 ^ n8179 ;
  assign n8187 = n4127 & n8186 ;
  assign n8188 = n8187 ^ n8186 ;
  assign n8189 = n8188 ^ n8179 ;
  assign n8191 = n8190 ^ n8189 ;
  assign n8192 = n4201 & n8191 ;
  assign n8203 = n8192 ^ n8189 ;
  assign n8195 = n8187 ^ n8179 ;
  assign n8196 = n8195 ^ x209 ;
  assign n8197 = ~n4163 & n8196 ;
  assign n8198 = n8197 ^ x209 ;
  assign n8193 = n8192 ^ n8191 ;
  assign n8194 = n8193 ^ n8189 ;
  assign n8199 = n8198 ^ n8194 ;
  assign n8200 = ~n4245 & n8199 ;
  assign n8201 = n8200 ^ n8199 ;
  assign n8202 = n8201 ^ n8194 ;
  assign n8204 = n8203 ^ n8202 ;
  assign n8205 = ~n4288 & n8204 ;
  assign n8220 = n8205 ^ n8202 ;
  assign n8208 = n8200 ^ n8194 ;
  assign n8209 = n8208 ^ x177 ;
  assign n8210 = ~n4320 & n8209 ;
  assign n8211 = n8210 ^ x177 ;
  assign n8206 = n8205 ^ n8204 ;
  assign n8207 = n8206 ^ n8202 ;
  assign n8212 = n8211 ^ n8207 ;
  assign n8213 = n4365 & n8212 ;
  assign n8219 = n8213 ^ n8207 ;
  assign n8221 = n8220 ^ n8219 ;
  assign n8222 = n4407 & n8221 ;
  assign n8229 = n8222 ^ n8219 ;
  assign n8223 = n8222 ^ n8221 ;
  assign n8224 = n8223 ^ n8219 ;
  assign n8214 = n8213 ^ n8212 ;
  assign n8215 = n8214 ^ n8207 ;
  assign n8216 = n8215 ^ x145 ;
  assign n8217 = ~n4444 & n8216 ;
  assign n8218 = n8217 ^ x145 ;
  assign n8225 = n8224 ^ n8218 ;
  assign n8226 = n4488 & n8225 ;
  assign n8227 = n8226 ^ n8225 ;
  assign n8228 = n8227 ^ n8218 ;
  assign n8230 = n8229 ^ n8228 ;
  assign n8231 = n4562 & n8230 ;
  assign n8242 = n8231 ^ n8228 ;
  assign n8234 = n8226 ^ n8218 ;
  assign n8235 = n8234 ^ x113 ;
  assign n8236 = ~n4524 & n8235 ;
  assign n8237 = n8236 ^ x113 ;
  assign n8232 = n8231 ^ n8230 ;
  assign n8233 = n8232 ^ n8228 ;
  assign n8238 = n8237 ^ n8233 ;
  assign n8239 = ~n4606 & n8238 ;
  assign n8240 = n8239 ^ n8238 ;
  assign n8241 = n8240 ^ n8233 ;
  assign n8243 = n8242 ^ n8241 ;
  assign n8244 = ~n4649 & n8243 ;
  assign n8259 = n8244 ^ n8241 ;
  assign n8247 = n8239 ^ n8233 ;
  assign n8248 = n8247 ^ x81 ;
  assign n8249 = ~n4681 & n8248 ;
  assign n8250 = n8249 ^ x81 ;
  assign n8245 = n8244 ^ n8243 ;
  assign n8246 = n8245 ^ n8241 ;
  assign n8251 = n8250 ^ n8246 ;
  assign n8252 = n4726 & n8251 ;
  assign n8258 = n8252 ^ n8246 ;
  assign n8260 = n8259 ^ n8258 ;
  assign n8261 = n4772 & n8260 ;
  assign n8268 = n8261 ^ n8258 ;
  assign n8262 = n8261 ^ n8260 ;
  assign n8263 = n8262 ^ n8258 ;
  assign n8253 = n8252 ^ n8251 ;
  assign n8254 = n8253 ^ n8246 ;
  assign n8255 = n8254 ^ x49 ;
  assign n8256 = ~n4806 & n8255 ;
  assign n8257 = n8256 ^ x49 ;
  assign n8264 = n8263 ^ n8257 ;
  assign n8265 = n4850 & n8264 ;
  assign n8266 = n8265 ^ n8264 ;
  assign n8267 = n8266 ^ n8257 ;
  assign n8269 = n8268 ^ n8267 ;
  assign n8270 = ~n4893 & n8269 ;
  assign n8281 = n8270 ^ n8267 ;
  assign n8273 = n8265 ^ n8257 ;
  assign n8274 = n8273 ^ x17 ;
  assign n8275 = ~n4927 & n8274 ;
  assign n8276 = n8275 ^ x17 ;
  assign n8271 = n8270 ^ n8269 ;
  assign n8272 = n8271 ^ n8267 ;
  assign n8277 = n8276 ^ n8272 ;
  assign n8278 = ~n4972 & n8277 ;
  assign n8279 = n8278 ^ n8277 ;
  assign n8280 = n8279 ^ n8272 ;
  assign n8282 = n8281 ^ n8280 ;
  assign n8283 = n5009 & n8282 ;
  assign n8284 = n8283 ^ n8282 ;
  assign n8285 = n8284 ^ n8280 ;
  assign n8286 = x498 ^ x466 ;
  assign n8287 = n3371 & n8286 ;
  assign n8294 = n8287 ^ x466 ;
  assign n8288 = n8287 ^ n8286 ;
  assign n8289 = n8288 ^ x466 ;
  assign n8290 = n8289 ^ x434 ;
  assign n8291 = n3412 & n8290 ;
  assign n8292 = n8291 ^ n8290 ;
  assign n8293 = n8292 ^ x434 ;
  assign n8295 = n8294 ^ n8293 ;
  assign n8296 = n3451 & n8295 ;
  assign n8311 = n8296 ^ n8293 ;
  assign n8299 = n8291 ^ x434 ;
  assign n8300 = n8299 ^ x402 ;
  assign n8301 = ~n3484 & n8300 ;
  assign n8302 = n8301 ^ x402 ;
  assign n8297 = n8296 ^ n8295 ;
  assign n8298 = n8297 ^ n8293 ;
  assign n8303 = n8302 ^ n8298 ;
  assign n8304 = ~n3527 & n8303 ;
  assign n8310 = n8304 ^ n8298 ;
  assign n8312 = n8311 ^ n8310 ;
  assign n8313 = ~n3570 & n8312 ;
  assign n8314 = n8313 ^ n8312 ;
  assign n8315 = n8314 ^ n8310 ;
  assign n8305 = n8304 ^ n8303 ;
  assign n8306 = n8305 ^ n8298 ;
  assign n8307 = n8306 ^ x370 ;
  assign n8308 = ~n3602 & n8307 ;
  assign n8309 = n8308 ^ x370 ;
  assign n8316 = n8315 ^ n8309 ;
  assign n8317 = ~n3646 & n8316 ;
  assign n8324 = n8317 ^ n8309 ;
  assign n8323 = n8313 ^ n8310 ;
  assign n8325 = n8324 ^ n8323 ;
  assign n8326 = ~n3688 & n8325 ;
  assign n8333 = n8326 ^ n8323 ;
  assign n8327 = n8326 ^ n8325 ;
  assign n8328 = n8327 ^ n8323 ;
  assign n8318 = n8317 ^ n8316 ;
  assign n8319 = n8318 ^ n8309 ;
  assign n8320 = n8319 ^ x338 ;
  assign n8321 = ~n3724 & n8320 ;
  assign n8322 = n8321 ^ x338 ;
  assign n8329 = n8328 ^ n8322 ;
  assign n8330 = n3767 & n8329 ;
  assign n8331 = n8330 ^ n8329 ;
  assign n8332 = n8331 ^ n8322 ;
  assign n8334 = n8333 ^ n8332 ;
  assign n8335 = n3841 & n8334 ;
  assign n8346 = n8335 ^ n8332 ;
  assign n8338 = n8330 ^ n8322 ;
  assign n8339 = n8338 ^ x306 ;
  assign n8340 = ~n3803 & n8339 ;
  assign n8341 = n8340 ^ x306 ;
  assign n8336 = n8335 ^ n8334 ;
  assign n8337 = n8336 ^ n8332 ;
  assign n8342 = n8341 ^ n8337 ;
  assign n8343 = ~n3884 & n8342 ;
  assign n8344 = n8343 ^ n8342 ;
  assign n8345 = n8344 ^ n8337 ;
  assign n8347 = n8346 ^ n8345 ;
  assign n8348 = ~n3927 & n8347 ;
  assign n8363 = n8348 ^ n8345 ;
  assign n8351 = n8343 ^ n8337 ;
  assign n8352 = n8351 ^ x274 ;
  assign n8353 = ~n3959 & n8352 ;
  assign n8354 = n8353 ^ x274 ;
  assign n8349 = n8348 ^ n8347 ;
  assign n8350 = n8349 ^ n8345 ;
  assign n8355 = n8354 ^ n8350 ;
  assign n8356 = n4004 & n8355 ;
  assign n8362 = n8356 ^ n8350 ;
  assign n8364 = n8363 ^ n8362 ;
  assign n8365 = n4046 & n8364 ;
  assign n8372 = n8365 ^ n8362 ;
  assign n8366 = n8365 ^ n8364 ;
  assign n8367 = n8366 ^ n8362 ;
  assign n8357 = n8356 ^ n8355 ;
  assign n8358 = n8357 ^ n8350 ;
  assign n8359 = n8358 ^ x242 ;
  assign n8360 = ~n4083 & n8359 ;
  assign n8361 = n8360 ^ x242 ;
  assign n8368 = n8367 ^ n8361 ;
  assign n8369 = n4127 & n8368 ;
  assign n8370 = n8369 ^ n8368 ;
  assign n8371 = n8370 ^ n8361 ;
  assign n8373 = n8372 ^ n8371 ;
  assign n8374 = n4201 & n8373 ;
  assign n8385 = n8374 ^ n8371 ;
  assign n8377 = n8369 ^ n8361 ;
  assign n8378 = n8377 ^ x210 ;
  assign n8379 = ~n4163 & n8378 ;
  assign n8380 = n8379 ^ x210 ;
  assign n8375 = n8374 ^ n8373 ;
  assign n8376 = n8375 ^ n8371 ;
  assign n8381 = n8380 ^ n8376 ;
  assign n8382 = ~n4245 & n8381 ;
  assign n8383 = n8382 ^ n8381 ;
  assign n8384 = n8383 ^ n8376 ;
  assign n8386 = n8385 ^ n8384 ;
  assign n8387 = ~n4288 & n8386 ;
  assign n8402 = n8387 ^ n8384 ;
  assign n8390 = n8382 ^ n8376 ;
  assign n8391 = n8390 ^ x178 ;
  assign n8392 = ~n4320 & n8391 ;
  assign n8393 = n8392 ^ x178 ;
  assign n8388 = n8387 ^ n8386 ;
  assign n8389 = n8388 ^ n8384 ;
  assign n8394 = n8393 ^ n8389 ;
  assign n8395 = n4365 & n8394 ;
  assign n8401 = n8395 ^ n8389 ;
  assign n8403 = n8402 ^ n8401 ;
  assign n8404 = n4407 & n8403 ;
  assign n8411 = n8404 ^ n8401 ;
  assign n8405 = n8404 ^ n8403 ;
  assign n8406 = n8405 ^ n8401 ;
  assign n8396 = n8395 ^ n8394 ;
  assign n8397 = n8396 ^ n8389 ;
  assign n8398 = n8397 ^ x146 ;
  assign n8399 = ~n4444 & n8398 ;
  assign n8400 = n8399 ^ x146 ;
  assign n8407 = n8406 ^ n8400 ;
  assign n8408 = n4488 & n8407 ;
  assign n8409 = n8408 ^ n8407 ;
  assign n8410 = n8409 ^ n8400 ;
  assign n8412 = n8411 ^ n8410 ;
  assign n8413 = n4562 & n8412 ;
  assign n8424 = n8413 ^ n8410 ;
  assign n8416 = n8408 ^ n8400 ;
  assign n8417 = n8416 ^ x114 ;
  assign n8418 = ~n4524 & n8417 ;
  assign n8419 = n8418 ^ x114 ;
  assign n8414 = n8413 ^ n8412 ;
  assign n8415 = n8414 ^ n8410 ;
  assign n8420 = n8419 ^ n8415 ;
  assign n8421 = ~n4606 & n8420 ;
  assign n8422 = n8421 ^ n8420 ;
  assign n8423 = n8422 ^ n8415 ;
  assign n8425 = n8424 ^ n8423 ;
  assign n8426 = ~n4649 & n8425 ;
  assign n8441 = n8426 ^ n8423 ;
  assign n8429 = n8421 ^ n8415 ;
  assign n8430 = n8429 ^ x82 ;
  assign n8431 = ~n4681 & n8430 ;
  assign n8432 = n8431 ^ x82 ;
  assign n8427 = n8426 ^ n8425 ;
  assign n8428 = n8427 ^ n8423 ;
  assign n8433 = n8432 ^ n8428 ;
  assign n8434 = n4726 & n8433 ;
  assign n8440 = n8434 ^ n8428 ;
  assign n8442 = n8441 ^ n8440 ;
  assign n8443 = n4772 & n8442 ;
  assign n8450 = n8443 ^ n8440 ;
  assign n8444 = n8443 ^ n8442 ;
  assign n8445 = n8444 ^ n8440 ;
  assign n8435 = n8434 ^ n8433 ;
  assign n8436 = n8435 ^ n8428 ;
  assign n8437 = n8436 ^ x50 ;
  assign n8438 = ~n4806 & n8437 ;
  assign n8439 = n8438 ^ x50 ;
  assign n8446 = n8445 ^ n8439 ;
  assign n8447 = n4850 & n8446 ;
  assign n8448 = n8447 ^ n8446 ;
  assign n8449 = n8448 ^ n8439 ;
  assign n8451 = n8450 ^ n8449 ;
  assign n8452 = ~n4893 & n8451 ;
  assign n8463 = n8452 ^ n8449 ;
  assign n8455 = n8447 ^ n8439 ;
  assign n8456 = n8455 ^ x18 ;
  assign n8457 = ~n4927 & n8456 ;
  assign n8458 = n8457 ^ x18 ;
  assign n8453 = n8452 ^ n8451 ;
  assign n8454 = n8453 ^ n8449 ;
  assign n8459 = n8458 ^ n8454 ;
  assign n8460 = ~n4972 & n8459 ;
  assign n8461 = n8460 ^ n8459 ;
  assign n8462 = n8461 ^ n8454 ;
  assign n8464 = n8463 ^ n8462 ;
  assign n8465 = n5009 & n8464 ;
  assign n8466 = n8465 ^ n8464 ;
  assign n8467 = n8466 ^ n8462 ;
  assign n8468 = x499 ^ x467 ;
  assign n8469 = n3371 & n8468 ;
  assign n8476 = n8469 ^ x467 ;
  assign n8470 = n8469 ^ n8468 ;
  assign n8471 = n8470 ^ x467 ;
  assign n8472 = n8471 ^ x435 ;
  assign n8473 = n3412 & n8472 ;
  assign n8474 = n8473 ^ n8472 ;
  assign n8475 = n8474 ^ x435 ;
  assign n8477 = n8476 ^ n8475 ;
  assign n8478 = n3451 & n8477 ;
  assign n8493 = n8478 ^ n8475 ;
  assign n8481 = n8473 ^ x435 ;
  assign n8482 = n8481 ^ x403 ;
  assign n8483 = ~n3484 & n8482 ;
  assign n8484 = n8483 ^ x403 ;
  assign n8479 = n8478 ^ n8477 ;
  assign n8480 = n8479 ^ n8475 ;
  assign n8485 = n8484 ^ n8480 ;
  assign n8486 = ~n3527 & n8485 ;
  assign n8492 = n8486 ^ n8480 ;
  assign n8494 = n8493 ^ n8492 ;
  assign n8495 = ~n3570 & n8494 ;
  assign n8496 = n8495 ^ n8494 ;
  assign n8497 = n8496 ^ n8492 ;
  assign n8487 = n8486 ^ n8485 ;
  assign n8488 = n8487 ^ n8480 ;
  assign n8489 = n8488 ^ x371 ;
  assign n8490 = ~n3602 & n8489 ;
  assign n8491 = n8490 ^ x371 ;
  assign n8498 = n8497 ^ n8491 ;
  assign n8499 = ~n3646 & n8498 ;
  assign n8506 = n8499 ^ n8491 ;
  assign n8505 = n8495 ^ n8492 ;
  assign n8507 = n8506 ^ n8505 ;
  assign n8508 = ~n3688 & n8507 ;
  assign n8515 = n8508 ^ n8505 ;
  assign n8509 = n8508 ^ n8507 ;
  assign n8510 = n8509 ^ n8505 ;
  assign n8500 = n8499 ^ n8498 ;
  assign n8501 = n8500 ^ n8491 ;
  assign n8502 = n8501 ^ x339 ;
  assign n8503 = ~n3724 & n8502 ;
  assign n8504 = n8503 ^ x339 ;
  assign n8511 = n8510 ^ n8504 ;
  assign n8512 = n3767 & n8511 ;
  assign n8513 = n8512 ^ n8511 ;
  assign n8514 = n8513 ^ n8504 ;
  assign n8516 = n8515 ^ n8514 ;
  assign n8517 = n3841 & n8516 ;
  assign n8528 = n8517 ^ n8514 ;
  assign n8520 = n8512 ^ n8504 ;
  assign n8521 = n8520 ^ x307 ;
  assign n8522 = ~n3803 & n8521 ;
  assign n8523 = n8522 ^ x307 ;
  assign n8518 = n8517 ^ n8516 ;
  assign n8519 = n8518 ^ n8514 ;
  assign n8524 = n8523 ^ n8519 ;
  assign n8525 = ~n3884 & n8524 ;
  assign n8526 = n8525 ^ n8524 ;
  assign n8527 = n8526 ^ n8519 ;
  assign n8529 = n8528 ^ n8527 ;
  assign n8530 = ~n3927 & n8529 ;
  assign n8545 = n8530 ^ n8527 ;
  assign n8533 = n8525 ^ n8519 ;
  assign n8534 = n8533 ^ x275 ;
  assign n8535 = ~n3959 & n8534 ;
  assign n8536 = n8535 ^ x275 ;
  assign n8531 = n8530 ^ n8529 ;
  assign n8532 = n8531 ^ n8527 ;
  assign n8537 = n8536 ^ n8532 ;
  assign n8538 = n4004 & n8537 ;
  assign n8544 = n8538 ^ n8532 ;
  assign n8546 = n8545 ^ n8544 ;
  assign n8547 = n4046 & n8546 ;
  assign n8554 = n8547 ^ n8544 ;
  assign n8548 = n8547 ^ n8546 ;
  assign n8549 = n8548 ^ n8544 ;
  assign n8539 = n8538 ^ n8537 ;
  assign n8540 = n8539 ^ n8532 ;
  assign n8541 = n8540 ^ x243 ;
  assign n8542 = ~n4083 & n8541 ;
  assign n8543 = n8542 ^ x243 ;
  assign n8550 = n8549 ^ n8543 ;
  assign n8551 = n4127 & n8550 ;
  assign n8552 = n8551 ^ n8550 ;
  assign n8553 = n8552 ^ n8543 ;
  assign n8555 = n8554 ^ n8553 ;
  assign n8556 = n4201 & n8555 ;
  assign n8567 = n8556 ^ n8553 ;
  assign n8559 = n8551 ^ n8543 ;
  assign n8560 = n8559 ^ x211 ;
  assign n8561 = ~n4163 & n8560 ;
  assign n8562 = n8561 ^ x211 ;
  assign n8557 = n8556 ^ n8555 ;
  assign n8558 = n8557 ^ n8553 ;
  assign n8563 = n8562 ^ n8558 ;
  assign n8564 = ~n4245 & n8563 ;
  assign n8565 = n8564 ^ n8563 ;
  assign n8566 = n8565 ^ n8558 ;
  assign n8568 = n8567 ^ n8566 ;
  assign n8569 = ~n4288 & n8568 ;
  assign n8584 = n8569 ^ n8566 ;
  assign n8572 = n8564 ^ n8558 ;
  assign n8573 = n8572 ^ x179 ;
  assign n8574 = ~n4320 & n8573 ;
  assign n8575 = n8574 ^ x179 ;
  assign n8570 = n8569 ^ n8568 ;
  assign n8571 = n8570 ^ n8566 ;
  assign n8576 = n8575 ^ n8571 ;
  assign n8577 = n4365 & n8576 ;
  assign n8583 = n8577 ^ n8571 ;
  assign n8585 = n8584 ^ n8583 ;
  assign n8586 = n4407 & n8585 ;
  assign n8593 = n8586 ^ n8583 ;
  assign n8587 = n8586 ^ n8585 ;
  assign n8588 = n8587 ^ n8583 ;
  assign n8578 = n8577 ^ n8576 ;
  assign n8579 = n8578 ^ n8571 ;
  assign n8580 = n8579 ^ x147 ;
  assign n8581 = ~n4444 & n8580 ;
  assign n8582 = n8581 ^ x147 ;
  assign n8589 = n8588 ^ n8582 ;
  assign n8590 = n4488 & n8589 ;
  assign n8591 = n8590 ^ n8589 ;
  assign n8592 = n8591 ^ n8582 ;
  assign n8594 = n8593 ^ n8592 ;
  assign n8595 = n4562 & n8594 ;
  assign n8606 = n8595 ^ n8592 ;
  assign n8598 = n8590 ^ n8582 ;
  assign n8599 = n8598 ^ x115 ;
  assign n8600 = ~n4524 & n8599 ;
  assign n8601 = n8600 ^ x115 ;
  assign n8596 = n8595 ^ n8594 ;
  assign n8597 = n8596 ^ n8592 ;
  assign n8602 = n8601 ^ n8597 ;
  assign n8603 = ~n4606 & n8602 ;
  assign n8604 = n8603 ^ n8602 ;
  assign n8605 = n8604 ^ n8597 ;
  assign n8607 = n8606 ^ n8605 ;
  assign n8608 = ~n4649 & n8607 ;
  assign n8623 = n8608 ^ n8605 ;
  assign n8611 = n8603 ^ n8597 ;
  assign n8612 = n8611 ^ x83 ;
  assign n8613 = ~n4681 & n8612 ;
  assign n8614 = n8613 ^ x83 ;
  assign n8609 = n8608 ^ n8607 ;
  assign n8610 = n8609 ^ n8605 ;
  assign n8615 = n8614 ^ n8610 ;
  assign n8616 = n4726 & n8615 ;
  assign n8622 = n8616 ^ n8610 ;
  assign n8624 = n8623 ^ n8622 ;
  assign n8625 = n4772 & n8624 ;
  assign n8632 = n8625 ^ n8622 ;
  assign n8626 = n8625 ^ n8624 ;
  assign n8627 = n8626 ^ n8622 ;
  assign n8617 = n8616 ^ n8615 ;
  assign n8618 = n8617 ^ n8610 ;
  assign n8619 = n8618 ^ x51 ;
  assign n8620 = ~n4806 & n8619 ;
  assign n8621 = n8620 ^ x51 ;
  assign n8628 = n8627 ^ n8621 ;
  assign n8629 = n4850 & n8628 ;
  assign n8630 = n8629 ^ n8628 ;
  assign n8631 = n8630 ^ n8621 ;
  assign n8633 = n8632 ^ n8631 ;
  assign n8634 = ~n4893 & n8633 ;
  assign n8645 = n8634 ^ n8631 ;
  assign n8637 = n8629 ^ n8621 ;
  assign n8638 = n8637 ^ x19 ;
  assign n8639 = ~n4927 & n8638 ;
  assign n8640 = n8639 ^ x19 ;
  assign n8635 = n8634 ^ n8633 ;
  assign n8636 = n8635 ^ n8631 ;
  assign n8641 = n8640 ^ n8636 ;
  assign n8642 = ~n4972 & n8641 ;
  assign n8643 = n8642 ^ n8641 ;
  assign n8644 = n8643 ^ n8636 ;
  assign n8646 = n8645 ^ n8644 ;
  assign n8647 = n5009 & n8646 ;
  assign n8648 = n8647 ^ n8646 ;
  assign n8649 = n8648 ^ n8644 ;
  assign n8650 = x500 ^ x468 ;
  assign n8651 = n3371 & n8650 ;
  assign n8658 = n8651 ^ x468 ;
  assign n8652 = n8651 ^ n8650 ;
  assign n8653 = n8652 ^ x468 ;
  assign n8654 = n8653 ^ x436 ;
  assign n8655 = n3412 & n8654 ;
  assign n8656 = n8655 ^ n8654 ;
  assign n8657 = n8656 ^ x436 ;
  assign n8659 = n8658 ^ n8657 ;
  assign n8660 = n3451 & n8659 ;
  assign n8675 = n8660 ^ n8657 ;
  assign n8663 = n8655 ^ x436 ;
  assign n8664 = n8663 ^ x404 ;
  assign n8665 = ~n3484 & n8664 ;
  assign n8666 = n8665 ^ x404 ;
  assign n8661 = n8660 ^ n8659 ;
  assign n8662 = n8661 ^ n8657 ;
  assign n8667 = n8666 ^ n8662 ;
  assign n8668 = ~n3527 & n8667 ;
  assign n8674 = n8668 ^ n8662 ;
  assign n8676 = n8675 ^ n8674 ;
  assign n8677 = ~n3570 & n8676 ;
  assign n8678 = n8677 ^ n8676 ;
  assign n8679 = n8678 ^ n8674 ;
  assign n8669 = n8668 ^ n8667 ;
  assign n8670 = n8669 ^ n8662 ;
  assign n8671 = n8670 ^ x372 ;
  assign n8672 = ~n3602 & n8671 ;
  assign n8673 = n8672 ^ x372 ;
  assign n8680 = n8679 ^ n8673 ;
  assign n8681 = ~n3646 & n8680 ;
  assign n8688 = n8681 ^ n8673 ;
  assign n8687 = n8677 ^ n8674 ;
  assign n8689 = n8688 ^ n8687 ;
  assign n8690 = ~n3688 & n8689 ;
  assign n8697 = n8690 ^ n8687 ;
  assign n8691 = n8690 ^ n8689 ;
  assign n8692 = n8691 ^ n8687 ;
  assign n8682 = n8681 ^ n8680 ;
  assign n8683 = n8682 ^ n8673 ;
  assign n8684 = n8683 ^ x340 ;
  assign n8685 = ~n3724 & n8684 ;
  assign n8686 = n8685 ^ x340 ;
  assign n8693 = n8692 ^ n8686 ;
  assign n8694 = n3767 & n8693 ;
  assign n8695 = n8694 ^ n8693 ;
  assign n8696 = n8695 ^ n8686 ;
  assign n8698 = n8697 ^ n8696 ;
  assign n8699 = n3841 & n8698 ;
  assign n8710 = n8699 ^ n8696 ;
  assign n8702 = n8694 ^ n8686 ;
  assign n8703 = n8702 ^ x308 ;
  assign n8704 = ~n3803 & n8703 ;
  assign n8705 = n8704 ^ x308 ;
  assign n8700 = n8699 ^ n8698 ;
  assign n8701 = n8700 ^ n8696 ;
  assign n8706 = n8705 ^ n8701 ;
  assign n8707 = ~n3884 & n8706 ;
  assign n8708 = n8707 ^ n8706 ;
  assign n8709 = n8708 ^ n8701 ;
  assign n8711 = n8710 ^ n8709 ;
  assign n8712 = ~n3927 & n8711 ;
  assign n8727 = n8712 ^ n8709 ;
  assign n8715 = n8707 ^ n8701 ;
  assign n8716 = n8715 ^ x276 ;
  assign n8717 = ~n3959 & n8716 ;
  assign n8718 = n8717 ^ x276 ;
  assign n8713 = n8712 ^ n8711 ;
  assign n8714 = n8713 ^ n8709 ;
  assign n8719 = n8718 ^ n8714 ;
  assign n8720 = n4004 & n8719 ;
  assign n8726 = n8720 ^ n8714 ;
  assign n8728 = n8727 ^ n8726 ;
  assign n8729 = n4046 & n8728 ;
  assign n8736 = n8729 ^ n8726 ;
  assign n8730 = n8729 ^ n8728 ;
  assign n8731 = n8730 ^ n8726 ;
  assign n8721 = n8720 ^ n8719 ;
  assign n8722 = n8721 ^ n8714 ;
  assign n8723 = n8722 ^ x244 ;
  assign n8724 = ~n4083 & n8723 ;
  assign n8725 = n8724 ^ x244 ;
  assign n8732 = n8731 ^ n8725 ;
  assign n8733 = n4127 & n8732 ;
  assign n8734 = n8733 ^ n8732 ;
  assign n8735 = n8734 ^ n8725 ;
  assign n8737 = n8736 ^ n8735 ;
  assign n8738 = n4201 & n8737 ;
  assign n8749 = n8738 ^ n8735 ;
  assign n8741 = n8733 ^ n8725 ;
  assign n8742 = n8741 ^ x212 ;
  assign n8743 = ~n4163 & n8742 ;
  assign n8744 = n8743 ^ x212 ;
  assign n8739 = n8738 ^ n8737 ;
  assign n8740 = n8739 ^ n8735 ;
  assign n8745 = n8744 ^ n8740 ;
  assign n8746 = ~n4245 & n8745 ;
  assign n8747 = n8746 ^ n8745 ;
  assign n8748 = n8747 ^ n8740 ;
  assign n8750 = n8749 ^ n8748 ;
  assign n8751 = ~n4288 & n8750 ;
  assign n8766 = n8751 ^ n8748 ;
  assign n8754 = n8746 ^ n8740 ;
  assign n8755 = n8754 ^ x180 ;
  assign n8756 = ~n4320 & n8755 ;
  assign n8757 = n8756 ^ x180 ;
  assign n8752 = n8751 ^ n8750 ;
  assign n8753 = n8752 ^ n8748 ;
  assign n8758 = n8757 ^ n8753 ;
  assign n8759 = n4365 & n8758 ;
  assign n8765 = n8759 ^ n8753 ;
  assign n8767 = n8766 ^ n8765 ;
  assign n8768 = n4407 & n8767 ;
  assign n8775 = n8768 ^ n8765 ;
  assign n8769 = n8768 ^ n8767 ;
  assign n8770 = n8769 ^ n8765 ;
  assign n8760 = n8759 ^ n8758 ;
  assign n8761 = n8760 ^ n8753 ;
  assign n8762 = n8761 ^ x148 ;
  assign n8763 = ~n4444 & n8762 ;
  assign n8764 = n8763 ^ x148 ;
  assign n8771 = n8770 ^ n8764 ;
  assign n8772 = n4488 & n8771 ;
  assign n8773 = n8772 ^ n8771 ;
  assign n8774 = n8773 ^ n8764 ;
  assign n8776 = n8775 ^ n8774 ;
  assign n8777 = n4562 & n8776 ;
  assign n8788 = n8777 ^ n8774 ;
  assign n8780 = n8772 ^ n8764 ;
  assign n8781 = n8780 ^ x116 ;
  assign n8782 = ~n4524 & n8781 ;
  assign n8783 = n8782 ^ x116 ;
  assign n8778 = n8777 ^ n8776 ;
  assign n8779 = n8778 ^ n8774 ;
  assign n8784 = n8783 ^ n8779 ;
  assign n8785 = ~n4606 & n8784 ;
  assign n8786 = n8785 ^ n8784 ;
  assign n8787 = n8786 ^ n8779 ;
  assign n8789 = n8788 ^ n8787 ;
  assign n8790 = ~n4649 & n8789 ;
  assign n8805 = n8790 ^ n8787 ;
  assign n8793 = n8785 ^ n8779 ;
  assign n8794 = n8793 ^ x84 ;
  assign n8795 = ~n4681 & n8794 ;
  assign n8796 = n8795 ^ x84 ;
  assign n8791 = n8790 ^ n8789 ;
  assign n8792 = n8791 ^ n8787 ;
  assign n8797 = n8796 ^ n8792 ;
  assign n8798 = n4726 & n8797 ;
  assign n8804 = n8798 ^ n8792 ;
  assign n8806 = n8805 ^ n8804 ;
  assign n8807 = n4772 & n8806 ;
  assign n8814 = n8807 ^ n8804 ;
  assign n8808 = n8807 ^ n8806 ;
  assign n8809 = n8808 ^ n8804 ;
  assign n8799 = n8798 ^ n8797 ;
  assign n8800 = n8799 ^ n8792 ;
  assign n8801 = n8800 ^ x52 ;
  assign n8802 = ~n4806 & n8801 ;
  assign n8803 = n8802 ^ x52 ;
  assign n8810 = n8809 ^ n8803 ;
  assign n8811 = n4850 & n8810 ;
  assign n8812 = n8811 ^ n8810 ;
  assign n8813 = n8812 ^ n8803 ;
  assign n8815 = n8814 ^ n8813 ;
  assign n8816 = ~n4893 & n8815 ;
  assign n8827 = n8816 ^ n8813 ;
  assign n8819 = n8811 ^ n8803 ;
  assign n8820 = n8819 ^ x20 ;
  assign n8821 = ~n4927 & n8820 ;
  assign n8822 = n8821 ^ x20 ;
  assign n8817 = n8816 ^ n8815 ;
  assign n8818 = n8817 ^ n8813 ;
  assign n8823 = n8822 ^ n8818 ;
  assign n8824 = ~n4972 & n8823 ;
  assign n8825 = n8824 ^ n8823 ;
  assign n8826 = n8825 ^ n8818 ;
  assign n8828 = n8827 ^ n8826 ;
  assign n8829 = n5009 & n8828 ;
  assign n8830 = n8829 ^ n8828 ;
  assign n8831 = n8830 ^ n8826 ;
  assign n8832 = x501 ^ x469 ;
  assign n8833 = n3371 & n8832 ;
  assign n8840 = n8833 ^ x469 ;
  assign n8834 = n8833 ^ n8832 ;
  assign n8835 = n8834 ^ x469 ;
  assign n8836 = n8835 ^ x437 ;
  assign n8837 = n3412 & n8836 ;
  assign n8838 = n8837 ^ n8836 ;
  assign n8839 = n8838 ^ x437 ;
  assign n8841 = n8840 ^ n8839 ;
  assign n8842 = n3451 & n8841 ;
  assign n8857 = n8842 ^ n8839 ;
  assign n8845 = n8837 ^ x437 ;
  assign n8846 = n8845 ^ x405 ;
  assign n8847 = ~n3484 & n8846 ;
  assign n8848 = n8847 ^ x405 ;
  assign n8843 = n8842 ^ n8841 ;
  assign n8844 = n8843 ^ n8839 ;
  assign n8849 = n8848 ^ n8844 ;
  assign n8850 = ~n3527 & n8849 ;
  assign n8856 = n8850 ^ n8844 ;
  assign n8858 = n8857 ^ n8856 ;
  assign n8859 = ~n3570 & n8858 ;
  assign n8860 = n8859 ^ n8858 ;
  assign n8861 = n8860 ^ n8856 ;
  assign n8851 = n8850 ^ n8849 ;
  assign n8852 = n8851 ^ n8844 ;
  assign n8853 = n8852 ^ x373 ;
  assign n8854 = ~n3602 & n8853 ;
  assign n8855 = n8854 ^ x373 ;
  assign n8862 = n8861 ^ n8855 ;
  assign n8863 = ~n3646 & n8862 ;
  assign n8870 = n8863 ^ n8855 ;
  assign n8869 = n8859 ^ n8856 ;
  assign n8871 = n8870 ^ n8869 ;
  assign n8872 = ~n3688 & n8871 ;
  assign n8879 = n8872 ^ n8869 ;
  assign n8873 = n8872 ^ n8871 ;
  assign n8874 = n8873 ^ n8869 ;
  assign n8864 = n8863 ^ n8862 ;
  assign n8865 = n8864 ^ n8855 ;
  assign n8866 = n8865 ^ x341 ;
  assign n8867 = ~n3724 & n8866 ;
  assign n8868 = n8867 ^ x341 ;
  assign n8875 = n8874 ^ n8868 ;
  assign n8876 = n3767 & n8875 ;
  assign n8877 = n8876 ^ n8875 ;
  assign n8878 = n8877 ^ n8868 ;
  assign n8880 = n8879 ^ n8878 ;
  assign n8881 = n3841 & n8880 ;
  assign n8892 = n8881 ^ n8878 ;
  assign n8884 = n8876 ^ n8868 ;
  assign n8885 = n8884 ^ x309 ;
  assign n8886 = ~n3803 & n8885 ;
  assign n8887 = n8886 ^ x309 ;
  assign n8882 = n8881 ^ n8880 ;
  assign n8883 = n8882 ^ n8878 ;
  assign n8888 = n8887 ^ n8883 ;
  assign n8889 = ~n3884 & n8888 ;
  assign n8890 = n8889 ^ n8888 ;
  assign n8891 = n8890 ^ n8883 ;
  assign n8893 = n8892 ^ n8891 ;
  assign n8894 = ~n3927 & n8893 ;
  assign n8909 = n8894 ^ n8891 ;
  assign n8897 = n8889 ^ n8883 ;
  assign n8898 = n8897 ^ x277 ;
  assign n8899 = ~n3959 & n8898 ;
  assign n8900 = n8899 ^ x277 ;
  assign n8895 = n8894 ^ n8893 ;
  assign n8896 = n8895 ^ n8891 ;
  assign n8901 = n8900 ^ n8896 ;
  assign n8902 = n4004 & n8901 ;
  assign n8908 = n8902 ^ n8896 ;
  assign n8910 = n8909 ^ n8908 ;
  assign n8911 = n4046 & n8910 ;
  assign n8918 = n8911 ^ n8908 ;
  assign n8912 = n8911 ^ n8910 ;
  assign n8913 = n8912 ^ n8908 ;
  assign n8903 = n8902 ^ n8901 ;
  assign n8904 = n8903 ^ n8896 ;
  assign n8905 = n8904 ^ x245 ;
  assign n8906 = ~n4083 & n8905 ;
  assign n8907 = n8906 ^ x245 ;
  assign n8914 = n8913 ^ n8907 ;
  assign n8915 = n4127 & n8914 ;
  assign n8916 = n8915 ^ n8914 ;
  assign n8917 = n8916 ^ n8907 ;
  assign n8919 = n8918 ^ n8917 ;
  assign n8920 = n4201 & n8919 ;
  assign n8931 = n8920 ^ n8917 ;
  assign n8923 = n8915 ^ n8907 ;
  assign n8924 = n8923 ^ x213 ;
  assign n8925 = ~n4163 & n8924 ;
  assign n8926 = n8925 ^ x213 ;
  assign n8921 = n8920 ^ n8919 ;
  assign n8922 = n8921 ^ n8917 ;
  assign n8927 = n8926 ^ n8922 ;
  assign n8928 = ~n4245 & n8927 ;
  assign n8929 = n8928 ^ n8927 ;
  assign n8930 = n8929 ^ n8922 ;
  assign n8932 = n8931 ^ n8930 ;
  assign n8933 = ~n4288 & n8932 ;
  assign n8948 = n8933 ^ n8930 ;
  assign n8936 = n8928 ^ n8922 ;
  assign n8937 = n8936 ^ x181 ;
  assign n8938 = ~n4320 & n8937 ;
  assign n8939 = n8938 ^ x181 ;
  assign n8934 = n8933 ^ n8932 ;
  assign n8935 = n8934 ^ n8930 ;
  assign n8940 = n8939 ^ n8935 ;
  assign n8941 = n4365 & n8940 ;
  assign n8947 = n8941 ^ n8935 ;
  assign n8949 = n8948 ^ n8947 ;
  assign n8950 = n4407 & n8949 ;
  assign n8957 = n8950 ^ n8947 ;
  assign n8951 = n8950 ^ n8949 ;
  assign n8952 = n8951 ^ n8947 ;
  assign n8942 = n8941 ^ n8940 ;
  assign n8943 = n8942 ^ n8935 ;
  assign n8944 = n8943 ^ x149 ;
  assign n8945 = ~n4444 & n8944 ;
  assign n8946 = n8945 ^ x149 ;
  assign n8953 = n8952 ^ n8946 ;
  assign n8954 = n4488 & n8953 ;
  assign n8955 = n8954 ^ n8953 ;
  assign n8956 = n8955 ^ n8946 ;
  assign n8958 = n8957 ^ n8956 ;
  assign n8959 = n4562 & n8958 ;
  assign n8970 = n8959 ^ n8956 ;
  assign n8962 = n8954 ^ n8946 ;
  assign n8963 = n8962 ^ x117 ;
  assign n8964 = ~n4524 & n8963 ;
  assign n8965 = n8964 ^ x117 ;
  assign n8960 = n8959 ^ n8958 ;
  assign n8961 = n8960 ^ n8956 ;
  assign n8966 = n8965 ^ n8961 ;
  assign n8967 = ~n4606 & n8966 ;
  assign n8968 = n8967 ^ n8966 ;
  assign n8969 = n8968 ^ n8961 ;
  assign n8971 = n8970 ^ n8969 ;
  assign n8972 = ~n4649 & n8971 ;
  assign n8987 = n8972 ^ n8969 ;
  assign n8975 = n8967 ^ n8961 ;
  assign n8976 = n8975 ^ x85 ;
  assign n8977 = ~n4681 & n8976 ;
  assign n8978 = n8977 ^ x85 ;
  assign n8973 = n8972 ^ n8971 ;
  assign n8974 = n8973 ^ n8969 ;
  assign n8979 = n8978 ^ n8974 ;
  assign n8980 = n4726 & n8979 ;
  assign n8986 = n8980 ^ n8974 ;
  assign n8988 = n8987 ^ n8986 ;
  assign n8989 = n4772 & n8988 ;
  assign n8996 = n8989 ^ n8986 ;
  assign n8990 = n8989 ^ n8988 ;
  assign n8991 = n8990 ^ n8986 ;
  assign n8981 = n8980 ^ n8979 ;
  assign n8982 = n8981 ^ n8974 ;
  assign n8983 = n8982 ^ x53 ;
  assign n8984 = ~n4806 & n8983 ;
  assign n8985 = n8984 ^ x53 ;
  assign n8992 = n8991 ^ n8985 ;
  assign n8993 = n4850 & n8992 ;
  assign n8994 = n8993 ^ n8992 ;
  assign n8995 = n8994 ^ n8985 ;
  assign n8997 = n8996 ^ n8995 ;
  assign n8998 = ~n4893 & n8997 ;
  assign n9009 = n8998 ^ n8995 ;
  assign n9001 = n8993 ^ n8985 ;
  assign n9002 = n9001 ^ x21 ;
  assign n9003 = ~n4927 & n9002 ;
  assign n9004 = n9003 ^ x21 ;
  assign n8999 = n8998 ^ n8997 ;
  assign n9000 = n8999 ^ n8995 ;
  assign n9005 = n9004 ^ n9000 ;
  assign n9006 = ~n4972 & n9005 ;
  assign n9007 = n9006 ^ n9005 ;
  assign n9008 = n9007 ^ n9000 ;
  assign n9010 = n9009 ^ n9008 ;
  assign n9011 = n5009 & n9010 ;
  assign n9012 = n9011 ^ n9010 ;
  assign n9013 = n9012 ^ n9008 ;
  assign n9014 = x502 ^ x470 ;
  assign n9015 = n3371 & n9014 ;
  assign n9022 = n9015 ^ x470 ;
  assign n9016 = n9015 ^ n9014 ;
  assign n9017 = n9016 ^ x470 ;
  assign n9018 = n9017 ^ x438 ;
  assign n9019 = n3412 & n9018 ;
  assign n9020 = n9019 ^ n9018 ;
  assign n9021 = n9020 ^ x438 ;
  assign n9023 = n9022 ^ n9021 ;
  assign n9024 = n3451 & n9023 ;
  assign n9039 = n9024 ^ n9021 ;
  assign n9027 = n9019 ^ x438 ;
  assign n9028 = n9027 ^ x406 ;
  assign n9029 = ~n3484 & n9028 ;
  assign n9030 = n9029 ^ x406 ;
  assign n9025 = n9024 ^ n9023 ;
  assign n9026 = n9025 ^ n9021 ;
  assign n9031 = n9030 ^ n9026 ;
  assign n9032 = ~n3527 & n9031 ;
  assign n9038 = n9032 ^ n9026 ;
  assign n9040 = n9039 ^ n9038 ;
  assign n9041 = ~n3570 & n9040 ;
  assign n9042 = n9041 ^ n9040 ;
  assign n9043 = n9042 ^ n9038 ;
  assign n9033 = n9032 ^ n9031 ;
  assign n9034 = n9033 ^ n9026 ;
  assign n9035 = n9034 ^ x374 ;
  assign n9036 = ~n3602 & n9035 ;
  assign n9037 = n9036 ^ x374 ;
  assign n9044 = n9043 ^ n9037 ;
  assign n9045 = ~n3646 & n9044 ;
  assign n9052 = n9045 ^ n9037 ;
  assign n9051 = n9041 ^ n9038 ;
  assign n9053 = n9052 ^ n9051 ;
  assign n9054 = ~n3688 & n9053 ;
  assign n9061 = n9054 ^ n9051 ;
  assign n9055 = n9054 ^ n9053 ;
  assign n9056 = n9055 ^ n9051 ;
  assign n9046 = n9045 ^ n9044 ;
  assign n9047 = n9046 ^ n9037 ;
  assign n9048 = n9047 ^ x342 ;
  assign n9049 = ~n3724 & n9048 ;
  assign n9050 = n9049 ^ x342 ;
  assign n9057 = n9056 ^ n9050 ;
  assign n9058 = n3767 & n9057 ;
  assign n9059 = n9058 ^ n9057 ;
  assign n9060 = n9059 ^ n9050 ;
  assign n9062 = n9061 ^ n9060 ;
  assign n9063 = n3841 & n9062 ;
  assign n9074 = n9063 ^ n9060 ;
  assign n9066 = n9058 ^ n9050 ;
  assign n9067 = n9066 ^ x310 ;
  assign n9068 = ~n3803 & n9067 ;
  assign n9069 = n9068 ^ x310 ;
  assign n9064 = n9063 ^ n9062 ;
  assign n9065 = n9064 ^ n9060 ;
  assign n9070 = n9069 ^ n9065 ;
  assign n9071 = ~n3884 & n9070 ;
  assign n9072 = n9071 ^ n9070 ;
  assign n9073 = n9072 ^ n9065 ;
  assign n9075 = n9074 ^ n9073 ;
  assign n9076 = ~n3927 & n9075 ;
  assign n9091 = n9076 ^ n9073 ;
  assign n9079 = n9071 ^ n9065 ;
  assign n9080 = n9079 ^ x278 ;
  assign n9081 = ~n3959 & n9080 ;
  assign n9082 = n9081 ^ x278 ;
  assign n9077 = n9076 ^ n9075 ;
  assign n9078 = n9077 ^ n9073 ;
  assign n9083 = n9082 ^ n9078 ;
  assign n9084 = n4004 & n9083 ;
  assign n9090 = n9084 ^ n9078 ;
  assign n9092 = n9091 ^ n9090 ;
  assign n9093 = n4046 & n9092 ;
  assign n9100 = n9093 ^ n9090 ;
  assign n9094 = n9093 ^ n9092 ;
  assign n9095 = n9094 ^ n9090 ;
  assign n9085 = n9084 ^ n9083 ;
  assign n9086 = n9085 ^ n9078 ;
  assign n9087 = n9086 ^ x246 ;
  assign n9088 = ~n4083 & n9087 ;
  assign n9089 = n9088 ^ x246 ;
  assign n9096 = n9095 ^ n9089 ;
  assign n9097 = n4127 & n9096 ;
  assign n9098 = n9097 ^ n9096 ;
  assign n9099 = n9098 ^ n9089 ;
  assign n9101 = n9100 ^ n9099 ;
  assign n9102 = n4201 & n9101 ;
  assign n9113 = n9102 ^ n9099 ;
  assign n9105 = n9097 ^ n9089 ;
  assign n9106 = n9105 ^ x214 ;
  assign n9107 = ~n4163 & n9106 ;
  assign n9108 = n9107 ^ x214 ;
  assign n9103 = n9102 ^ n9101 ;
  assign n9104 = n9103 ^ n9099 ;
  assign n9109 = n9108 ^ n9104 ;
  assign n9110 = ~n4245 & n9109 ;
  assign n9111 = n9110 ^ n9109 ;
  assign n9112 = n9111 ^ n9104 ;
  assign n9114 = n9113 ^ n9112 ;
  assign n9115 = ~n4288 & n9114 ;
  assign n9130 = n9115 ^ n9112 ;
  assign n9118 = n9110 ^ n9104 ;
  assign n9119 = n9118 ^ x182 ;
  assign n9120 = ~n4320 & n9119 ;
  assign n9121 = n9120 ^ x182 ;
  assign n9116 = n9115 ^ n9114 ;
  assign n9117 = n9116 ^ n9112 ;
  assign n9122 = n9121 ^ n9117 ;
  assign n9123 = n4365 & n9122 ;
  assign n9129 = n9123 ^ n9117 ;
  assign n9131 = n9130 ^ n9129 ;
  assign n9132 = n4407 & n9131 ;
  assign n9139 = n9132 ^ n9129 ;
  assign n9133 = n9132 ^ n9131 ;
  assign n9134 = n9133 ^ n9129 ;
  assign n9124 = n9123 ^ n9122 ;
  assign n9125 = n9124 ^ n9117 ;
  assign n9126 = n9125 ^ x150 ;
  assign n9127 = ~n4444 & n9126 ;
  assign n9128 = n9127 ^ x150 ;
  assign n9135 = n9134 ^ n9128 ;
  assign n9136 = n4488 & n9135 ;
  assign n9137 = n9136 ^ n9135 ;
  assign n9138 = n9137 ^ n9128 ;
  assign n9140 = n9139 ^ n9138 ;
  assign n9141 = n4562 & n9140 ;
  assign n9152 = n9141 ^ n9138 ;
  assign n9144 = n9136 ^ n9128 ;
  assign n9145 = n9144 ^ x118 ;
  assign n9146 = ~n4524 & n9145 ;
  assign n9147 = n9146 ^ x118 ;
  assign n9142 = n9141 ^ n9140 ;
  assign n9143 = n9142 ^ n9138 ;
  assign n9148 = n9147 ^ n9143 ;
  assign n9149 = ~n4606 & n9148 ;
  assign n9150 = n9149 ^ n9148 ;
  assign n9151 = n9150 ^ n9143 ;
  assign n9153 = n9152 ^ n9151 ;
  assign n9154 = ~n4649 & n9153 ;
  assign n9169 = n9154 ^ n9151 ;
  assign n9157 = n9149 ^ n9143 ;
  assign n9158 = n9157 ^ x86 ;
  assign n9159 = ~n4681 & n9158 ;
  assign n9160 = n9159 ^ x86 ;
  assign n9155 = n9154 ^ n9153 ;
  assign n9156 = n9155 ^ n9151 ;
  assign n9161 = n9160 ^ n9156 ;
  assign n9162 = n4726 & n9161 ;
  assign n9168 = n9162 ^ n9156 ;
  assign n9170 = n9169 ^ n9168 ;
  assign n9171 = n4772 & n9170 ;
  assign n9178 = n9171 ^ n9168 ;
  assign n9172 = n9171 ^ n9170 ;
  assign n9173 = n9172 ^ n9168 ;
  assign n9163 = n9162 ^ n9161 ;
  assign n9164 = n9163 ^ n9156 ;
  assign n9165 = n9164 ^ x54 ;
  assign n9166 = ~n4806 & n9165 ;
  assign n9167 = n9166 ^ x54 ;
  assign n9174 = n9173 ^ n9167 ;
  assign n9175 = n4850 & n9174 ;
  assign n9176 = n9175 ^ n9174 ;
  assign n9177 = n9176 ^ n9167 ;
  assign n9179 = n9178 ^ n9177 ;
  assign n9180 = ~n4893 & n9179 ;
  assign n9191 = n9180 ^ n9177 ;
  assign n9183 = n9175 ^ n9167 ;
  assign n9184 = n9183 ^ x22 ;
  assign n9185 = ~n4927 & n9184 ;
  assign n9186 = n9185 ^ x22 ;
  assign n9181 = n9180 ^ n9179 ;
  assign n9182 = n9181 ^ n9177 ;
  assign n9187 = n9186 ^ n9182 ;
  assign n9188 = ~n4972 & n9187 ;
  assign n9189 = n9188 ^ n9187 ;
  assign n9190 = n9189 ^ n9182 ;
  assign n9192 = n9191 ^ n9190 ;
  assign n9193 = n5009 & n9192 ;
  assign n9194 = n9193 ^ n9192 ;
  assign n9195 = n9194 ^ n9190 ;
  assign n9196 = x503 ^ x471 ;
  assign n9197 = n3371 & n9196 ;
  assign n9204 = n9197 ^ x471 ;
  assign n9198 = n9197 ^ n9196 ;
  assign n9199 = n9198 ^ x471 ;
  assign n9200 = n9199 ^ x439 ;
  assign n9201 = n3412 & n9200 ;
  assign n9202 = n9201 ^ n9200 ;
  assign n9203 = n9202 ^ x439 ;
  assign n9205 = n9204 ^ n9203 ;
  assign n9206 = n3451 & n9205 ;
  assign n9221 = n9206 ^ n9203 ;
  assign n9209 = n9201 ^ x439 ;
  assign n9210 = n9209 ^ x407 ;
  assign n9211 = ~n3484 & n9210 ;
  assign n9212 = n9211 ^ x407 ;
  assign n9207 = n9206 ^ n9205 ;
  assign n9208 = n9207 ^ n9203 ;
  assign n9213 = n9212 ^ n9208 ;
  assign n9214 = ~n3527 & n9213 ;
  assign n9220 = n9214 ^ n9208 ;
  assign n9222 = n9221 ^ n9220 ;
  assign n9223 = ~n3570 & n9222 ;
  assign n9224 = n9223 ^ n9222 ;
  assign n9225 = n9224 ^ n9220 ;
  assign n9215 = n9214 ^ n9213 ;
  assign n9216 = n9215 ^ n9208 ;
  assign n9217 = n9216 ^ x375 ;
  assign n9218 = ~n3602 & n9217 ;
  assign n9219 = n9218 ^ x375 ;
  assign n9226 = n9225 ^ n9219 ;
  assign n9227 = ~n3646 & n9226 ;
  assign n9234 = n9227 ^ n9219 ;
  assign n9233 = n9223 ^ n9220 ;
  assign n9235 = n9234 ^ n9233 ;
  assign n9236 = ~n3688 & n9235 ;
  assign n9243 = n9236 ^ n9233 ;
  assign n9237 = n9236 ^ n9235 ;
  assign n9238 = n9237 ^ n9233 ;
  assign n9228 = n9227 ^ n9226 ;
  assign n9229 = n9228 ^ n9219 ;
  assign n9230 = n9229 ^ x343 ;
  assign n9231 = ~n3724 & n9230 ;
  assign n9232 = n9231 ^ x343 ;
  assign n9239 = n9238 ^ n9232 ;
  assign n9240 = n3767 & n9239 ;
  assign n9241 = n9240 ^ n9239 ;
  assign n9242 = n9241 ^ n9232 ;
  assign n9244 = n9243 ^ n9242 ;
  assign n9245 = n3841 & n9244 ;
  assign n9256 = n9245 ^ n9242 ;
  assign n9248 = n9240 ^ n9232 ;
  assign n9249 = n9248 ^ x311 ;
  assign n9250 = ~n3803 & n9249 ;
  assign n9251 = n9250 ^ x311 ;
  assign n9246 = n9245 ^ n9244 ;
  assign n9247 = n9246 ^ n9242 ;
  assign n9252 = n9251 ^ n9247 ;
  assign n9253 = ~n3884 & n9252 ;
  assign n9254 = n9253 ^ n9252 ;
  assign n9255 = n9254 ^ n9247 ;
  assign n9257 = n9256 ^ n9255 ;
  assign n9258 = ~n3927 & n9257 ;
  assign n9273 = n9258 ^ n9255 ;
  assign n9261 = n9253 ^ n9247 ;
  assign n9262 = n9261 ^ x279 ;
  assign n9263 = ~n3959 & n9262 ;
  assign n9264 = n9263 ^ x279 ;
  assign n9259 = n9258 ^ n9257 ;
  assign n9260 = n9259 ^ n9255 ;
  assign n9265 = n9264 ^ n9260 ;
  assign n9266 = n4004 & n9265 ;
  assign n9272 = n9266 ^ n9260 ;
  assign n9274 = n9273 ^ n9272 ;
  assign n9275 = n4046 & n9274 ;
  assign n9282 = n9275 ^ n9272 ;
  assign n9276 = n9275 ^ n9274 ;
  assign n9277 = n9276 ^ n9272 ;
  assign n9267 = n9266 ^ n9265 ;
  assign n9268 = n9267 ^ n9260 ;
  assign n9269 = n9268 ^ x247 ;
  assign n9270 = ~n4083 & n9269 ;
  assign n9271 = n9270 ^ x247 ;
  assign n9278 = n9277 ^ n9271 ;
  assign n9279 = n4127 & n9278 ;
  assign n9280 = n9279 ^ n9278 ;
  assign n9281 = n9280 ^ n9271 ;
  assign n9283 = n9282 ^ n9281 ;
  assign n9284 = n4201 & n9283 ;
  assign n9295 = n9284 ^ n9281 ;
  assign n9287 = n9279 ^ n9271 ;
  assign n9288 = n9287 ^ x215 ;
  assign n9289 = ~n4163 & n9288 ;
  assign n9290 = n9289 ^ x215 ;
  assign n9285 = n9284 ^ n9283 ;
  assign n9286 = n9285 ^ n9281 ;
  assign n9291 = n9290 ^ n9286 ;
  assign n9292 = ~n4245 & n9291 ;
  assign n9293 = n9292 ^ n9291 ;
  assign n9294 = n9293 ^ n9286 ;
  assign n9296 = n9295 ^ n9294 ;
  assign n9297 = ~n4288 & n9296 ;
  assign n9312 = n9297 ^ n9294 ;
  assign n9300 = n9292 ^ n9286 ;
  assign n9301 = n9300 ^ x183 ;
  assign n9302 = ~n4320 & n9301 ;
  assign n9303 = n9302 ^ x183 ;
  assign n9298 = n9297 ^ n9296 ;
  assign n9299 = n9298 ^ n9294 ;
  assign n9304 = n9303 ^ n9299 ;
  assign n9305 = n4365 & n9304 ;
  assign n9311 = n9305 ^ n9299 ;
  assign n9313 = n9312 ^ n9311 ;
  assign n9314 = n4407 & n9313 ;
  assign n9321 = n9314 ^ n9311 ;
  assign n9315 = n9314 ^ n9313 ;
  assign n9316 = n9315 ^ n9311 ;
  assign n9306 = n9305 ^ n9304 ;
  assign n9307 = n9306 ^ n9299 ;
  assign n9308 = n9307 ^ x151 ;
  assign n9309 = ~n4444 & n9308 ;
  assign n9310 = n9309 ^ x151 ;
  assign n9317 = n9316 ^ n9310 ;
  assign n9318 = n4488 & n9317 ;
  assign n9319 = n9318 ^ n9317 ;
  assign n9320 = n9319 ^ n9310 ;
  assign n9322 = n9321 ^ n9320 ;
  assign n9323 = n4562 & n9322 ;
  assign n9334 = n9323 ^ n9320 ;
  assign n9326 = n9318 ^ n9310 ;
  assign n9327 = n9326 ^ x119 ;
  assign n9328 = ~n4524 & n9327 ;
  assign n9329 = n9328 ^ x119 ;
  assign n9324 = n9323 ^ n9322 ;
  assign n9325 = n9324 ^ n9320 ;
  assign n9330 = n9329 ^ n9325 ;
  assign n9331 = ~n4606 & n9330 ;
  assign n9332 = n9331 ^ n9330 ;
  assign n9333 = n9332 ^ n9325 ;
  assign n9335 = n9334 ^ n9333 ;
  assign n9336 = ~n4649 & n9335 ;
  assign n9351 = n9336 ^ n9333 ;
  assign n9339 = n9331 ^ n9325 ;
  assign n9340 = n9339 ^ x87 ;
  assign n9341 = ~n4681 & n9340 ;
  assign n9342 = n9341 ^ x87 ;
  assign n9337 = n9336 ^ n9335 ;
  assign n9338 = n9337 ^ n9333 ;
  assign n9343 = n9342 ^ n9338 ;
  assign n9344 = n4726 & n9343 ;
  assign n9350 = n9344 ^ n9338 ;
  assign n9352 = n9351 ^ n9350 ;
  assign n9353 = n4772 & n9352 ;
  assign n9360 = n9353 ^ n9350 ;
  assign n9354 = n9353 ^ n9352 ;
  assign n9355 = n9354 ^ n9350 ;
  assign n9345 = n9344 ^ n9343 ;
  assign n9346 = n9345 ^ n9338 ;
  assign n9347 = n9346 ^ x55 ;
  assign n9348 = ~n4806 & n9347 ;
  assign n9349 = n9348 ^ x55 ;
  assign n9356 = n9355 ^ n9349 ;
  assign n9357 = n4850 & n9356 ;
  assign n9358 = n9357 ^ n9356 ;
  assign n9359 = n9358 ^ n9349 ;
  assign n9361 = n9360 ^ n9359 ;
  assign n9362 = ~n4893 & n9361 ;
  assign n9373 = n9362 ^ n9359 ;
  assign n9365 = n9357 ^ n9349 ;
  assign n9366 = n9365 ^ x23 ;
  assign n9367 = ~n4927 & n9366 ;
  assign n9368 = n9367 ^ x23 ;
  assign n9363 = n9362 ^ n9361 ;
  assign n9364 = n9363 ^ n9359 ;
  assign n9369 = n9368 ^ n9364 ;
  assign n9370 = ~n4972 & n9369 ;
  assign n9371 = n9370 ^ n9369 ;
  assign n9372 = n9371 ^ n9364 ;
  assign n9374 = n9373 ^ n9372 ;
  assign n9375 = n5009 & n9374 ;
  assign n9376 = n9375 ^ n9374 ;
  assign n9377 = n9376 ^ n9372 ;
  assign n9378 = x504 ^ x472 ;
  assign n9379 = n3371 & n9378 ;
  assign n9386 = n9379 ^ x472 ;
  assign n9380 = n9379 ^ n9378 ;
  assign n9381 = n9380 ^ x472 ;
  assign n9382 = n9381 ^ x440 ;
  assign n9383 = n3412 & n9382 ;
  assign n9384 = n9383 ^ n9382 ;
  assign n9385 = n9384 ^ x440 ;
  assign n9387 = n9386 ^ n9385 ;
  assign n9388 = n3451 & n9387 ;
  assign n9403 = n9388 ^ n9385 ;
  assign n9391 = n9383 ^ x440 ;
  assign n9392 = n9391 ^ x408 ;
  assign n9393 = ~n3484 & n9392 ;
  assign n9394 = n9393 ^ x408 ;
  assign n9389 = n9388 ^ n9387 ;
  assign n9390 = n9389 ^ n9385 ;
  assign n9395 = n9394 ^ n9390 ;
  assign n9396 = ~n3527 & n9395 ;
  assign n9402 = n9396 ^ n9390 ;
  assign n9404 = n9403 ^ n9402 ;
  assign n9405 = ~n3570 & n9404 ;
  assign n9406 = n9405 ^ n9404 ;
  assign n9407 = n9406 ^ n9402 ;
  assign n9397 = n9396 ^ n9395 ;
  assign n9398 = n9397 ^ n9390 ;
  assign n9399 = n9398 ^ x376 ;
  assign n9400 = ~n3602 & n9399 ;
  assign n9401 = n9400 ^ x376 ;
  assign n9408 = n9407 ^ n9401 ;
  assign n9409 = ~n3646 & n9408 ;
  assign n9416 = n9409 ^ n9401 ;
  assign n9415 = n9405 ^ n9402 ;
  assign n9417 = n9416 ^ n9415 ;
  assign n9418 = ~n3688 & n9417 ;
  assign n9425 = n9418 ^ n9415 ;
  assign n9419 = n9418 ^ n9417 ;
  assign n9420 = n9419 ^ n9415 ;
  assign n9410 = n9409 ^ n9408 ;
  assign n9411 = n9410 ^ n9401 ;
  assign n9412 = n9411 ^ x344 ;
  assign n9413 = ~n3724 & n9412 ;
  assign n9414 = n9413 ^ x344 ;
  assign n9421 = n9420 ^ n9414 ;
  assign n9422 = n3767 & n9421 ;
  assign n9423 = n9422 ^ n9421 ;
  assign n9424 = n9423 ^ n9414 ;
  assign n9426 = n9425 ^ n9424 ;
  assign n9427 = n3841 & n9426 ;
  assign n9438 = n9427 ^ n9424 ;
  assign n9430 = n9422 ^ n9414 ;
  assign n9431 = n9430 ^ x312 ;
  assign n9432 = ~n3803 & n9431 ;
  assign n9433 = n9432 ^ x312 ;
  assign n9428 = n9427 ^ n9426 ;
  assign n9429 = n9428 ^ n9424 ;
  assign n9434 = n9433 ^ n9429 ;
  assign n9435 = ~n3884 & n9434 ;
  assign n9436 = n9435 ^ n9434 ;
  assign n9437 = n9436 ^ n9429 ;
  assign n9439 = n9438 ^ n9437 ;
  assign n9440 = ~n3927 & n9439 ;
  assign n9455 = n9440 ^ n9437 ;
  assign n9443 = n9435 ^ n9429 ;
  assign n9444 = n9443 ^ x280 ;
  assign n9445 = ~n3959 & n9444 ;
  assign n9446 = n9445 ^ x280 ;
  assign n9441 = n9440 ^ n9439 ;
  assign n9442 = n9441 ^ n9437 ;
  assign n9447 = n9446 ^ n9442 ;
  assign n9448 = n4004 & n9447 ;
  assign n9454 = n9448 ^ n9442 ;
  assign n9456 = n9455 ^ n9454 ;
  assign n9457 = n4046 & n9456 ;
  assign n9464 = n9457 ^ n9454 ;
  assign n9458 = n9457 ^ n9456 ;
  assign n9459 = n9458 ^ n9454 ;
  assign n9449 = n9448 ^ n9447 ;
  assign n9450 = n9449 ^ n9442 ;
  assign n9451 = n9450 ^ x248 ;
  assign n9452 = ~n4083 & n9451 ;
  assign n9453 = n9452 ^ x248 ;
  assign n9460 = n9459 ^ n9453 ;
  assign n9461 = n4127 & n9460 ;
  assign n9462 = n9461 ^ n9460 ;
  assign n9463 = n9462 ^ n9453 ;
  assign n9465 = n9464 ^ n9463 ;
  assign n9466 = n4201 & n9465 ;
  assign n9477 = n9466 ^ n9463 ;
  assign n9469 = n9461 ^ n9453 ;
  assign n9470 = n9469 ^ x216 ;
  assign n9471 = ~n4163 & n9470 ;
  assign n9472 = n9471 ^ x216 ;
  assign n9467 = n9466 ^ n9465 ;
  assign n9468 = n9467 ^ n9463 ;
  assign n9473 = n9472 ^ n9468 ;
  assign n9474 = ~n4245 & n9473 ;
  assign n9475 = n9474 ^ n9473 ;
  assign n9476 = n9475 ^ n9468 ;
  assign n9478 = n9477 ^ n9476 ;
  assign n9479 = ~n4288 & n9478 ;
  assign n9494 = n9479 ^ n9476 ;
  assign n9482 = n9474 ^ n9468 ;
  assign n9483 = n9482 ^ x184 ;
  assign n9484 = ~n4320 & n9483 ;
  assign n9485 = n9484 ^ x184 ;
  assign n9480 = n9479 ^ n9478 ;
  assign n9481 = n9480 ^ n9476 ;
  assign n9486 = n9485 ^ n9481 ;
  assign n9487 = n4365 & n9486 ;
  assign n9493 = n9487 ^ n9481 ;
  assign n9495 = n9494 ^ n9493 ;
  assign n9496 = n4407 & n9495 ;
  assign n9503 = n9496 ^ n9493 ;
  assign n9497 = n9496 ^ n9495 ;
  assign n9498 = n9497 ^ n9493 ;
  assign n9488 = n9487 ^ n9486 ;
  assign n9489 = n9488 ^ n9481 ;
  assign n9490 = n9489 ^ x152 ;
  assign n9491 = ~n4444 & n9490 ;
  assign n9492 = n9491 ^ x152 ;
  assign n9499 = n9498 ^ n9492 ;
  assign n9500 = n4488 & n9499 ;
  assign n9501 = n9500 ^ n9499 ;
  assign n9502 = n9501 ^ n9492 ;
  assign n9504 = n9503 ^ n9502 ;
  assign n9505 = n4562 & n9504 ;
  assign n9516 = n9505 ^ n9502 ;
  assign n9508 = n9500 ^ n9492 ;
  assign n9509 = n9508 ^ x120 ;
  assign n9510 = ~n4524 & n9509 ;
  assign n9511 = n9510 ^ x120 ;
  assign n9506 = n9505 ^ n9504 ;
  assign n9507 = n9506 ^ n9502 ;
  assign n9512 = n9511 ^ n9507 ;
  assign n9513 = ~n4606 & n9512 ;
  assign n9514 = n9513 ^ n9512 ;
  assign n9515 = n9514 ^ n9507 ;
  assign n9517 = n9516 ^ n9515 ;
  assign n9518 = ~n4649 & n9517 ;
  assign n9533 = n9518 ^ n9515 ;
  assign n9521 = n9513 ^ n9507 ;
  assign n9522 = n9521 ^ x88 ;
  assign n9523 = ~n4681 & n9522 ;
  assign n9524 = n9523 ^ x88 ;
  assign n9519 = n9518 ^ n9517 ;
  assign n9520 = n9519 ^ n9515 ;
  assign n9525 = n9524 ^ n9520 ;
  assign n9526 = n4726 & n9525 ;
  assign n9532 = n9526 ^ n9520 ;
  assign n9534 = n9533 ^ n9532 ;
  assign n9535 = n4772 & n9534 ;
  assign n9542 = n9535 ^ n9532 ;
  assign n9536 = n9535 ^ n9534 ;
  assign n9537 = n9536 ^ n9532 ;
  assign n9527 = n9526 ^ n9525 ;
  assign n9528 = n9527 ^ n9520 ;
  assign n9529 = n9528 ^ x56 ;
  assign n9530 = ~n4806 & n9529 ;
  assign n9531 = n9530 ^ x56 ;
  assign n9538 = n9537 ^ n9531 ;
  assign n9539 = n4850 & n9538 ;
  assign n9540 = n9539 ^ n9538 ;
  assign n9541 = n9540 ^ n9531 ;
  assign n9543 = n9542 ^ n9541 ;
  assign n9544 = ~n4893 & n9543 ;
  assign n9555 = n9544 ^ n9541 ;
  assign n9547 = n9539 ^ n9531 ;
  assign n9548 = n9547 ^ x24 ;
  assign n9549 = ~n4927 & n9548 ;
  assign n9550 = n9549 ^ x24 ;
  assign n9545 = n9544 ^ n9543 ;
  assign n9546 = n9545 ^ n9541 ;
  assign n9551 = n9550 ^ n9546 ;
  assign n9552 = ~n4972 & n9551 ;
  assign n9553 = n9552 ^ n9551 ;
  assign n9554 = n9553 ^ n9546 ;
  assign n9556 = n9555 ^ n9554 ;
  assign n9557 = n5009 & n9556 ;
  assign n9558 = n9557 ^ n9556 ;
  assign n9559 = n9558 ^ n9554 ;
  assign n9560 = x505 ^ x473 ;
  assign n9561 = n3371 & n9560 ;
  assign n9568 = n9561 ^ x473 ;
  assign n9562 = n9561 ^ n9560 ;
  assign n9563 = n9562 ^ x473 ;
  assign n9564 = n9563 ^ x441 ;
  assign n9565 = n3412 & n9564 ;
  assign n9566 = n9565 ^ n9564 ;
  assign n9567 = n9566 ^ x441 ;
  assign n9569 = n9568 ^ n9567 ;
  assign n9570 = n3451 & n9569 ;
  assign n9585 = n9570 ^ n9567 ;
  assign n9573 = n9565 ^ x441 ;
  assign n9574 = n9573 ^ x409 ;
  assign n9575 = ~n3484 & n9574 ;
  assign n9576 = n9575 ^ x409 ;
  assign n9571 = n9570 ^ n9569 ;
  assign n9572 = n9571 ^ n9567 ;
  assign n9577 = n9576 ^ n9572 ;
  assign n9578 = ~n3527 & n9577 ;
  assign n9584 = n9578 ^ n9572 ;
  assign n9586 = n9585 ^ n9584 ;
  assign n9587 = ~n3570 & n9586 ;
  assign n9588 = n9587 ^ n9586 ;
  assign n9589 = n9588 ^ n9584 ;
  assign n9579 = n9578 ^ n9577 ;
  assign n9580 = n9579 ^ n9572 ;
  assign n9581 = n9580 ^ x377 ;
  assign n9582 = ~n3602 & n9581 ;
  assign n9583 = n9582 ^ x377 ;
  assign n9590 = n9589 ^ n9583 ;
  assign n9591 = ~n3646 & n9590 ;
  assign n9598 = n9591 ^ n9583 ;
  assign n9597 = n9587 ^ n9584 ;
  assign n9599 = n9598 ^ n9597 ;
  assign n9600 = ~n3688 & n9599 ;
  assign n9607 = n9600 ^ n9597 ;
  assign n9601 = n9600 ^ n9599 ;
  assign n9602 = n9601 ^ n9597 ;
  assign n9592 = n9591 ^ n9590 ;
  assign n9593 = n9592 ^ n9583 ;
  assign n9594 = n9593 ^ x345 ;
  assign n9595 = ~n3724 & n9594 ;
  assign n9596 = n9595 ^ x345 ;
  assign n9603 = n9602 ^ n9596 ;
  assign n9604 = n3767 & n9603 ;
  assign n9605 = n9604 ^ n9603 ;
  assign n9606 = n9605 ^ n9596 ;
  assign n9608 = n9607 ^ n9606 ;
  assign n9609 = n3841 & n9608 ;
  assign n9620 = n9609 ^ n9606 ;
  assign n9612 = n9604 ^ n9596 ;
  assign n9613 = n9612 ^ x313 ;
  assign n9614 = ~n3803 & n9613 ;
  assign n9615 = n9614 ^ x313 ;
  assign n9610 = n9609 ^ n9608 ;
  assign n9611 = n9610 ^ n9606 ;
  assign n9616 = n9615 ^ n9611 ;
  assign n9617 = ~n3884 & n9616 ;
  assign n9618 = n9617 ^ n9616 ;
  assign n9619 = n9618 ^ n9611 ;
  assign n9621 = n9620 ^ n9619 ;
  assign n9622 = ~n3927 & n9621 ;
  assign n9637 = n9622 ^ n9619 ;
  assign n9625 = n9617 ^ n9611 ;
  assign n9626 = n9625 ^ x281 ;
  assign n9627 = ~n3959 & n9626 ;
  assign n9628 = n9627 ^ x281 ;
  assign n9623 = n9622 ^ n9621 ;
  assign n9624 = n9623 ^ n9619 ;
  assign n9629 = n9628 ^ n9624 ;
  assign n9630 = n4004 & n9629 ;
  assign n9636 = n9630 ^ n9624 ;
  assign n9638 = n9637 ^ n9636 ;
  assign n9639 = n4046 & n9638 ;
  assign n9646 = n9639 ^ n9636 ;
  assign n9640 = n9639 ^ n9638 ;
  assign n9641 = n9640 ^ n9636 ;
  assign n9631 = n9630 ^ n9629 ;
  assign n9632 = n9631 ^ n9624 ;
  assign n9633 = n9632 ^ x249 ;
  assign n9634 = ~n4083 & n9633 ;
  assign n9635 = n9634 ^ x249 ;
  assign n9642 = n9641 ^ n9635 ;
  assign n9643 = n4127 & n9642 ;
  assign n9644 = n9643 ^ n9642 ;
  assign n9645 = n9644 ^ n9635 ;
  assign n9647 = n9646 ^ n9645 ;
  assign n9648 = n4201 & n9647 ;
  assign n9659 = n9648 ^ n9645 ;
  assign n9651 = n9643 ^ n9635 ;
  assign n9652 = n9651 ^ x217 ;
  assign n9653 = ~n4163 & n9652 ;
  assign n9654 = n9653 ^ x217 ;
  assign n9649 = n9648 ^ n9647 ;
  assign n9650 = n9649 ^ n9645 ;
  assign n9655 = n9654 ^ n9650 ;
  assign n9656 = ~n4245 & n9655 ;
  assign n9657 = n9656 ^ n9655 ;
  assign n9658 = n9657 ^ n9650 ;
  assign n9660 = n9659 ^ n9658 ;
  assign n9661 = ~n4288 & n9660 ;
  assign n9676 = n9661 ^ n9658 ;
  assign n9664 = n9656 ^ n9650 ;
  assign n9665 = n9664 ^ x185 ;
  assign n9666 = ~n4320 & n9665 ;
  assign n9667 = n9666 ^ x185 ;
  assign n9662 = n9661 ^ n9660 ;
  assign n9663 = n9662 ^ n9658 ;
  assign n9668 = n9667 ^ n9663 ;
  assign n9669 = n4365 & n9668 ;
  assign n9675 = n9669 ^ n9663 ;
  assign n9677 = n9676 ^ n9675 ;
  assign n9678 = n4407 & n9677 ;
  assign n9685 = n9678 ^ n9675 ;
  assign n9679 = n9678 ^ n9677 ;
  assign n9680 = n9679 ^ n9675 ;
  assign n9670 = n9669 ^ n9668 ;
  assign n9671 = n9670 ^ n9663 ;
  assign n9672 = n9671 ^ x153 ;
  assign n9673 = ~n4444 & n9672 ;
  assign n9674 = n9673 ^ x153 ;
  assign n9681 = n9680 ^ n9674 ;
  assign n9682 = n4488 & n9681 ;
  assign n9683 = n9682 ^ n9681 ;
  assign n9684 = n9683 ^ n9674 ;
  assign n9686 = n9685 ^ n9684 ;
  assign n9687 = n4562 & n9686 ;
  assign n9698 = n9687 ^ n9684 ;
  assign n9690 = n9682 ^ n9674 ;
  assign n9691 = n9690 ^ x121 ;
  assign n9692 = ~n4524 & n9691 ;
  assign n9693 = n9692 ^ x121 ;
  assign n9688 = n9687 ^ n9686 ;
  assign n9689 = n9688 ^ n9684 ;
  assign n9694 = n9693 ^ n9689 ;
  assign n9695 = ~n4606 & n9694 ;
  assign n9696 = n9695 ^ n9694 ;
  assign n9697 = n9696 ^ n9689 ;
  assign n9699 = n9698 ^ n9697 ;
  assign n9700 = ~n4649 & n9699 ;
  assign n9715 = n9700 ^ n9697 ;
  assign n9703 = n9695 ^ n9689 ;
  assign n9704 = n9703 ^ x89 ;
  assign n9705 = ~n4681 & n9704 ;
  assign n9706 = n9705 ^ x89 ;
  assign n9701 = n9700 ^ n9699 ;
  assign n9702 = n9701 ^ n9697 ;
  assign n9707 = n9706 ^ n9702 ;
  assign n9708 = n4726 & n9707 ;
  assign n9714 = n9708 ^ n9702 ;
  assign n9716 = n9715 ^ n9714 ;
  assign n9717 = n4772 & n9716 ;
  assign n9724 = n9717 ^ n9714 ;
  assign n9718 = n9717 ^ n9716 ;
  assign n9719 = n9718 ^ n9714 ;
  assign n9709 = n9708 ^ n9707 ;
  assign n9710 = n9709 ^ n9702 ;
  assign n9711 = n9710 ^ x57 ;
  assign n9712 = ~n4806 & n9711 ;
  assign n9713 = n9712 ^ x57 ;
  assign n9720 = n9719 ^ n9713 ;
  assign n9721 = n4850 & n9720 ;
  assign n9722 = n9721 ^ n9720 ;
  assign n9723 = n9722 ^ n9713 ;
  assign n9725 = n9724 ^ n9723 ;
  assign n9726 = ~n4893 & n9725 ;
  assign n9737 = n9726 ^ n9723 ;
  assign n9729 = n9721 ^ n9713 ;
  assign n9730 = n9729 ^ x25 ;
  assign n9731 = ~n4927 & n9730 ;
  assign n9732 = n9731 ^ x25 ;
  assign n9727 = n9726 ^ n9725 ;
  assign n9728 = n9727 ^ n9723 ;
  assign n9733 = n9732 ^ n9728 ;
  assign n9734 = ~n4972 & n9733 ;
  assign n9735 = n9734 ^ n9733 ;
  assign n9736 = n9735 ^ n9728 ;
  assign n9738 = n9737 ^ n9736 ;
  assign n9739 = n5009 & n9738 ;
  assign n9740 = n9739 ^ n9738 ;
  assign n9741 = n9740 ^ n9736 ;
  assign n9742 = x506 ^ x474 ;
  assign n9743 = n3371 & n9742 ;
  assign n9750 = n9743 ^ x474 ;
  assign n9744 = n9743 ^ n9742 ;
  assign n9745 = n9744 ^ x474 ;
  assign n9746 = n9745 ^ x442 ;
  assign n9747 = n3412 & n9746 ;
  assign n9748 = n9747 ^ n9746 ;
  assign n9749 = n9748 ^ x442 ;
  assign n9751 = n9750 ^ n9749 ;
  assign n9752 = n3451 & n9751 ;
  assign n9767 = n9752 ^ n9749 ;
  assign n9755 = n9747 ^ x442 ;
  assign n9756 = n9755 ^ x410 ;
  assign n9757 = ~n3484 & n9756 ;
  assign n9758 = n9757 ^ x410 ;
  assign n9753 = n9752 ^ n9751 ;
  assign n9754 = n9753 ^ n9749 ;
  assign n9759 = n9758 ^ n9754 ;
  assign n9760 = ~n3527 & n9759 ;
  assign n9766 = n9760 ^ n9754 ;
  assign n9768 = n9767 ^ n9766 ;
  assign n9769 = ~n3570 & n9768 ;
  assign n9770 = n9769 ^ n9768 ;
  assign n9771 = n9770 ^ n9766 ;
  assign n9761 = n9760 ^ n9759 ;
  assign n9762 = n9761 ^ n9754 ;
  assign n9763 = n9762 ^ x378 ;
  assign n9764 = ~n3602 & n9763 ;
  assign n9765 = n9764 ^ x378 ;
  assign n9772 = n9771 ^ n9765 ;
  assign n9773 = ~n3646 & n9772 ;
  assign n9780 = n9773 ^ n9765 ;
  assign n9779 = n9769 ^ n9766 ;
  assign n9781 = n9780 ^ n9779 ;
  assign n9782 = ~n3688 & n9781 ;
  assign n9789 = n9782 ^ n9779 ;
  assign n9783 = n9782 ^ n9781 ;
  assign n9784 = n9783 ^ n9779 ;
  assign n9774 = n9773 ^ n9772 ;
  assign n9775 = n9774 ^ n9765 ;
  assign n9776 = n9775 ^ x346 ;
  assign n9777 = ~n3724 & n9776 ;
  assign n9778 = n9777 ^ x346 ;
  assign n9785 = n9784 ^ n9778 ;
  assign n9786 = n3767 & n9785 ;
  assign n9787 = n9786 ^ n9785 ;
  assign n9788 = n9787 ^ n9778 ;
  assign n9790 = n9789 ^ n9788 ;
  assign n9791 = n3841 & n9790 ;
  assign n9802 = n9791 ^ n9788 ;
  assign n9794 = n9786 ^ n9778 ;
  assign n9795 = n9794 ^ x314 ;
  assign n9796 = ~n3803 & n9795 ;
  assign n9797 = n9796 ^ x314 ;
  assign n9792 = n9791 ^ n9790 ;
  assign n9793 = n9792 ^ n9788 ;
  assign n9798 = n9797 ^ n9793 ;
  assign n9799 = ~n3884 & n9798 ;
  assign n9800 = n9799 ^ n9798 ;
  assign n9801 = n9800 ^ n9793 ;
  assign n9803 = n9802 ^ n9801 ;
  assign n9804 = ~n3927 & n9803 ;
  assign n9819 = n9804 ^ n9801 ;
  assign n9807 = n9799 ^ n9793 ;
  assign n9808 = n9807 ^ x282 ;
  assign n9809 = ~n3959 & n9808 ;
  assign n9810 = n9809 ^ x282 ;
  assign n9805 = n9804 ^ n9803 ;
  assign n9806 = n9805 ^ n9801 ;
  assign n9811 = n9810 ^ n9806 ;
  assign n9812 = n4004 & n9811 ;
  assign n9818 = n9812 ^ n9806 ;
  assign n9820 = n9819 ^ n9818 ;
  assign n9821 = n4046 & n9820 ;
  assign n9828 = n9821 ^ n9818 ;
  assign n9822 = n9821 ^ n9820 ;
  assign n9823 = n9822 ^ n9818 ;
  assign n9813 = n9812 ^ n9811 ;
  assign n9814 = n9813 ^ n9806 ;
  assign n9815 = n9814 ^ x250 ;
  assign n9816 = ~n4083 & n9815 ;
  assign n9817 = n9816 ^ x250 ;
  assign n9824 = n9823 ^ n9817 ;
  assign n9825 = n4127 & n9824 ;
  assign n9826 = n9825 ^ n9824 ;
  assign n9827 = n9826 ^ n9817 ;
  assign n9829 = n9828 ^ n9827 ;
  assign n9830 = n4201 & n9829 ;
  assign n9841 = n9830 ^ n9827 ;
  assign n9833 = n9825 ^ n9817 ;
  assign n9834 = n9833 ^ x218 ;
  assign n9835 = ~n4163 & n9834 ;
  assign n9836 = n9835 ^ x218 ;
  assign n9831 = n9830 ^ n9829 ;
  assign n9832 = n9831 ^ n9827 ;
  assign n9837 = n9836 ^ n9832 ;
  assign n9838 = ~n4245 & n9837 ;
  assign n9839 = n9838 ^ n9837 ;
  assign n9840 = n9839 ^ n9832 ;
  assign n9842 = n9841 ^ n9840 ;
  assign n9843 = ~n4288 & n9842 ;
  assign n9858 = n9843 ^ n9840 ;
  assign n9846 = n9838 ^ n9832 ;
  assign n9847 = n9846 ^ x186 ;
  assign n9848 = ~n4320 & n9847 ;
  assign n9849 = n9848 ^ x186 ;
  assign n9844 = n9843 ^ n9842 ;
  assign n9845 = n9844 ^ n9840 ;
  assign n9850 = n9849 ^ n9845 ;
  assign n9851 = n4365 & n9850 ;
  assign n9857 = n9851 ^ n9845 ;
  assign n9859 = n9858 ^ n9857 ;
  assign n9860 = n4407 & n9859 ;
  assign n9867 = n9860 ^ n9857 ;
  assign n9861 = n9860 ^ n9859 ;
  assign n9862 = n9861 ^ n9857 ;
  assign n9852 = n9851 ^ n9850 ;
  assign n9853 = n9852 ^ n9845 ;
  assign n9854 = n9853 ^ x154 ;
  assign n9855 = ~n4444 & n9854 ;
  assign n9856 = n9855 ^ x154 ;
  assign n9863 = n9862 ^ n9856 ;
  assign n9864 = n4488 & n9863 ;
  assign n9865 = n9864 ^ n9863 ;
  assign n9866 = n9865 ^ n9856 ;
  assign n9868 = n9867 ^ n9866 ;
  assign n9869 = n4562 & n9868 ;
  assign n9880 = n9869 ^ n9866 ;
  assign n9872 = n9864 ^ n9856 ;
  assign n9873 = n9872 ^ x122 ;
  assign n9874 = ~n4524 & n9873 ;
  assign n9875 = n9874 ^ x122 ;
  assign n9870 = n9869 ^ n9868 ;
  assign n9871 = n9870 ^ n9866 ;
  assign n9876 = n9875 ^ n9871 ;
  assign n9877 = ~n4606 & n9876 ;
  assign n9878 = n9877 ^ n9876 ;
  assign n9879 = n9878 ^ n9871 ;
  assign n9881 = n9880 ^ n9879 ;
  assign n9882 = ~n4649 & n9881 ;
  assign n9897 = n9882 ^ n9879 ;
  assign n9885 = n9877 ^ n9871 ;
  assign n9886 = n9885 ^ x90 ;
  assign n9887 = ~n4681 & n9886 ;
  assign n9888 = n9887 ^ x90 ;
  assign n9883 = n9882 ^ n9881 ;
  assign n9884 = n9883 ^ n9879 ;
  assign n9889 = n9888 ^ n9884 ;
  assign n9890 = n4726 & n9889 ;
  assign n9896 = n9890 ^ n9884 ;
  assign n9898 = n9897 ^ n9896 ;
  assign n9899 = n4772 & n9898 ;
  assign n9906 = n9899 ^ n9896 ;
  assign n9900 = n9899 ^ n9898 ;
  assign n9901 = n9900 ^ n9896 ;
  assign n9891 = n9890 ^ n9889 ;
  assign n9892 = n9891 ^ n9884 ;
  assign n9893 = n9892 ^ x58 ;
  assign n9894 = ~n4806 & n9893 ;
  assign n9895 = n9894 ^ x58 ;
  assign n9902 = n9901 ^ n9895 ;
  assign n9903 = n4850 & n9902 ;
  assign n9904 = n9903 ^ n9902 ;
  assign n9905 = n9904 ^ n9895 ;
  assign n9907 = n9906 ^ n9905 ;
  assign n9908 = ~n4893 & n9907 ;
  assign n9919 = n9908 ^ n9905 ;
  assign n9911 = n9903 ^ n9895 ;
  assign n9912 = n9911 ^ x26 ;
  assign n9913 = ~n4927 & n9912 ;
  assign n9914 = n9913 ^ x26 ;
  assign n9909 = n9908 ^ n9907 ;
  assign n9910 = n9909 ^ n9905 ;
  assign n9915 = n9914 ^ n9910 ;
  assign n9916 = ~n4972 & n9915 ;
  assign n9917 = n9916 ^ n9915 ;
  assign n9918 = n9917 ^ n9910 ;
  assign n9920 = n9919 ^ n9918 ;
  assign n9921 = n5009 & n9920 ;
  assign n9922 = n9921 ^ n9920 ;
  assign n9923 = n9922 ^ n9918 ;
  assign n9924 = x507 ^ x475 ;
  assign n9925 = n3371 & n9924 ;
  assign n9932 = n9925 ^ x475 ;
  assign n9926 = n9925 ^ n9924 ;
  assign n9927 = n9926 ^ x475 ;
  assign n9928 = n9927 ^ x443 ;
  assign n9929 = n3412 & n9928 ;
  assign n9930 = n9929 ^ n9928 ;
  assign n9931 = n9930 ^ x443 ;
  assign n9933 = n9932 ^ n9931 ;
  assign n9934 = n3451 & n9933 ;
  assign n9949 = n9934 ^ n9931 ;
  assign n9937 = n9929 ^ x443 ;
  assign n9938 = n9937 ^ x411 ;
  assign n9939 = ~n3484 & n9938 ;
  assign n9940 = n9939 ^ x411 ;
  assign n9935 = n9934 ^ n9933 ;
  assign n9936 = n9935 ^ n9931 ;
  assign n9941 = n9940 ^ n9936 ;
  assign n9942 = ~n3527 & n9941 ;
  assign n9948 = n9942 ^ n9936 ;
  assign n9950 = n9949 ^ n9948 ;
  assign n9951 = ~n3570 & n9950 ;
  assign n9952 = n9951 ^ n9950 ;
  assign n9953 = n9952 ^ n9948 ;
  assign n9943 = n9942 ^ n9941 ;
  assign n9944 = n9943 ^ n9936 ;
  assign n9945 = n9944 ^ x379 ;
  assign n9946 = ~n3602 & n9945 ;
  assign n9947 = n9946 ^ x379 ;
  assign n9954 = n9953 ^ n9947 ;
  assign n9955 = ~n3646 & n9954 ;
  assign n9962 = n9955 ^ n9947 ;
  assign n9961 = n9951 ^ n9948 ;
  assign n9963 = n9962 ^ n9961 ;
  assign n9964 = ~n3688 & n9963 ;
  assign n9971 = n9964 ^ n9961 ;
  assign n9965 = n9964 ^ n9963 ;
  assign n9966 = n9965 ^ n9961 ;
  assign n9956 = n9955 ^ n9954 ;
  assign n9957 = n9956 ^ n9947 ;
  assign n9958 = n9957 ^ x347 ;
  assign n9959 = ~n3724 & n9958 ;
  assign n9960 = n9959 ^ x347 ;
  assign n9967 = n9966 ^ n9960 ;
  assign n9968 = n3767 & n9967 ;
  assign n9969 = n9968 ^ n9967 ;
  assign n9970 = n9969 ^ n9960 ;
  assign n9972 = n9971 ^ n9970 ;
  assign n9973 = n3841 & n9972 ;
  assign n9984 = n9973 ^ n9970 ;
  assign n9976 = n9968 ^ n9960 ;
  assign n9977 = n9976 ^ x315 ;
  assign n9978 = ~n3803 & n9977 ;
  assign n9979 = n9978 ^ x315 ;
  assign n9974 = n9973 ^ n9972 ;
  assign n9975 = n9974 ^ n9970 ;
  assign n9980 = n9979 ^ n9975 ;
  assign n9981 = ~n3884 & n9980 ;
  assign n9982 = n9981 ^ n9980 ;
  assign n9983 = n9982 ^ n9975 ;
  assign n9985 = n9984 ^ n9983 ;
  assign n9986 = ~n3927 & n9985 ;
  assign n10001 = n9986 ^ n9983 ;
  assign n9989 = n9981 ^ n9975 ;
  assign n9990 = n9989 ^ x283 ;
  assign n9991 = ~n3959 & n9990 ;
  assign n9992 = n9991 ^ x283 ;
  assign n9987 = n9986 ^ n9985 ;
  assign n9988 = n9987 ^ n9983 ;
  assign n9993 = n9992 ^ n9988 ;
  assign n9994 = n4004 & n9993 ;
  assign n10000 = n9994 ^ n9988 ;
  assign n10002 = n10001 ^ n10000 ;
  assign n10003 = n4046 & n10002 ;
  assign n10010 = n10003 ^ n10000 ;
  assign n10004 = n10003 ^ n10002 ;
  assign n10005 = n10004 ^ n10000 ;
  assign n9995 = n9994 ^ n9993 ;
  assign n9996 = n9995 ^ n9988 ;
  assign n9997 = n9996 ^ x251 ;
  assign n9998 = ~n4083 & n9997 ;
  assign n9999 = n9998 ^ x251 ;
  assign n10006 = n10005 ^ n9999 ;
  assign n10007 = n4127 & n10006 ;
  assign n10008 = n10007 ^ n10006 ;
  assign n10009 = n10008 ^ n9999 ;
  assign n10011 = n10010 ^ n10009 ;
  assign n10012 = n4201 & n10011 ;
  assign n10023 = n10012 ^ n10009 ;
  assign n10015 = n10007 ^ n9999 ;
  assign n10016 = n10015 ^ x219 ;
  assign n10017 = ~n4163 & n10016 ;
  assign n10018 = n10017 ^ x219 ;
  assign n10013 = n10012 ^ n10011 ;
  assign n10014 = n10013 ^ n10009 ;
  assign n10019 = n10018 ^ n10014 ;
  assign n10020 = ~n4245 & n10019 ;
  assign n10021 = n10020 ^ n10019 ;
  assign n10022 = n10021 ^ n10014 ;
  assign n10024 = n10023 ^ n10022 ;
  assign n10025 = ~n4288 & n10024 ;
  assign n10040 = n10025 ^ n10022 ;
  assign n10028 = n10020 ^ n10014 ;
  assign n10029 = n10028 ^ x187 ;
  assign n10030 = ~n4320 & n10029 ;
  assign n10031 = n10030 ^ x187 ;
  assign n10026 = n10025 ^ n10024 ;
  assign n10027 = n10026 ^ n10022 ;
  assign n10032 = n10031 ^ n10027 ;
  assign n10033 = n4365 & n10032 ;
  assign n10039 = n10033 ^ n10027 ;
  assign n10041 = n10040 ^ n10039 ;
  assign n10042 = n4407 & n10041 ;
  assign n10049 = n10042 ^ n10039 ;
  assign n10043 = n10042 ^ n10041 ;
  assign n10044 = n10043 ^ n10039 ;
  assign n10034 = n10033 ^ n10032 ;
  assign n10035 = n10034 ^ n10027 ;
  assign n10036 = n10035 ^ x155 ;
  assign n10037 = ~n4444 & n10036 ;
  assign n10038 = n10037 ^ x155 ;
  assign n10045 = n10044 ^ n10038 ;
  assign n10046 = n4488 & n10045 ;
  assign n10047 = n10046 ^ n10045 ;
  assign n10048 = n10047 ^ n10038 ;
  assign n10050 = n10049 ^ n10048 ;
  assign n10051 = n4562 & n10050 ;
  assign n10062 = n10051 ^ n10048 ;
  assign n10054 = n10046 ^ n10038 ;
  assign n10055 = n10054 ^ x123 ;
  assign n10056 = ~n4524 & n10055 ;
  assign n10057 = n10056 ^ x123 ;
  assign n10052 = n10051 ^ n10050 ;
  assign n10053 = n10052 ^ n10048 ;
  assign n10058 = n10057 ^ n10053 ;
  assign n10059 = ~n4606 & n10058 ;
  assign n10060 = n10059 ^ n10058 ;
  assign n10061 = n10060 ^ n10053 ;
  assign n10063 = n10062 ^ n10061 ;
  assign n10064 = ~n4649 & n10063 ;
  assign n10079 = n10064 ^ n10061 ;
  assign n10067 = n10059 ^ n10053 ;
  assign n10068 = n10067 ^ x91 ;
  assign n10069 = ~n4681 & n10068 ;
  assign n10070 = n10069 ^ x91 ;
  assign n10065 = n10064 ^ n10063 ;
  assign n10066 = n10065 ^ n10061 ;
  assign n10071 = n10070 ^ n10066 ;
  assign n10072 = n4726 & n10071 ;
  assign n10078 = n10072 ^ n10066 ;
  assign n10080 = n10079 ^ n10078 ;
  assign n10081 = n4772 & n10080 ;
  assign n10088 = n10081 ^ n10078 ;
  assign n10082 = n10081 ^ n10080 ;
  assign n10083 = n10082 ^ n10078 ;
  assign n10073 = n10072 ^ n10071 ;
  assign n10074 = n10073 ^ n10066 ;
  assign n10075 = n10074 ^ x59 ;
  assign n10076 = ~n4806 & n10075 ;
  assign n10077 = n10076 ^ x59 ;
  assign n10084 = n10083 ^ n10077 ;
  assign n10085 = n4850 & n10084 ;
  assign n10086 = n10085 ^ n10084 ;
  assign n10087 = n10086 ^ n10077 ;
  assign n10089 = n10088 ^ n10087 ;
  assign n10090 = ~n4893 & n10089 ;
  assign n10101 = n10090 ^ n10087 ;
  assign n10093 = n10085 ^ n10077 ;
  assign n10094 = n10093 ^ x27 ;
  assign n10095 = ~n4927 & n10094 ;
  assign n10096 = n10095 ^ x27 ;
  assign n10091 = n10090 ^ n10089 ;
  assign n10092 = n10091 ^ n10087 ;
  assign n10097 = n10096 ^ n10092 ;
  assign n10098 = ~n4972 & n10097 ;
  assign n10099 = n10098 ^ n10097 ;
  assign n10100 = n10099 ^ n10092 ;
  assign n10102 = n10101 ^ n10100 ;
  assign n10103 = n5009 & n10102 ;
  assign n10104 = n10103 ^ n10102 ;
  assign n10105 = n10104 ^ n10100 ;
  assign n10106 = x508 ^ x476 ;
  assign n10107 = n3371 & n10106 ;
  assign n10114 = n10107 ^ x476 ;
  assign n10108 = n10107 ^ n10106 ;
  assign n10109 = n10108 ^ x476 ;
  assign n10110 = n10109 ^ x444 ;
  assign n10111 = n3412 & n10110 ;
  assign n10112 = n10111 ^ n10110 ;
  assign n10113 = n10112 ^ x444 ;
  assign n10115 = n10114 ^ n10113 ;
  assign n10116 = n3451 & n10115 ;
  assign n10131 = n10116 ^ n10113 ;
  assign n10119 = n10111 ^ x444 ;
  assign n10120 = n10119 ^ x412 ;
  assign n10121 = ~n3484 & n10120 ;
  assign n10122 = n10121 ^ x412 ;
  assign n10117 = n10116 ^ n10115 ;
  assign n10118 = n10117 ^ n10113 ;
  assign n10123 = n10122 ^ n10118 ;
  assign n10124 = ~n3527 & n10123 ;
  assign n10130 = n10124 ^ n10118 ;
  assign n10132 = n10131 ^ n10130 ;
  assign n10133 = ~n3570 & n10132 ;
  assign n10134 = n10133 ^ n10132 ;
  assign n10135 = n10134 ^ n10130 ;
  assign n10125 = n10124 ^ n10123 ;
  assign n10126 = n10125 ^ n10118 ;
  assign n10127 = n10126 ^ x380 ;
  assign n10128 = ~n3602 & n10127 ;
  assign n10129 = n10128 ^ x380 ;
  assign n10136 = n10135 ^ n10129 ;
  assign n10137 = ~n3646 & n10136 ;
  assign n10144 = n10137 ^ n10129 ;
  assign n10143 = n10133 ^ n10130 ;
  assign n10145 = n10144 ^ n10143 ;
  assign n10146 = ~n3688 & n10145 ;
  assign n10153 = n10146 ^ n10143 ;
  assign n10147 = n10146 ^ n10145 ;
  assign n10148 = n10147 ^ n10143 ;
  assign n10138 = n10137 ^ n10136 ;
  assign n10139 = n10138 ^ n10129 ;
  assign n10140 = n10139 ^ x348 ;
  assign n10141 = ~n3724 & n10140 ;
  assign n10142 = n10141 ^ x348 ;
  assign n10149 = n10148 ^ n10142 ;
  assign n10150 = n3767 & n10149 ;
  assign n10151 = n10150 ^ n10149 ;
  assign n10152 = n10151 ^ n10142 ;
  assign n10154 = n10153 ^ n10152 ;
  assign n10155 = n3841 & n10154 ;
  assign n10166 = n10155 ^ n10152 ;
  assign n10158 = n10150 ^ n10142 ;
  assign n10159 = n10158 ^ x316 ;
  assign n10160 = ~n3803 & n10159 ;
  assign n10161 = n10160 ^ x316 ;
  assign n10156 = n10155 ^ n10154 ;
  assign n10157 = n10156 ^ n10152 ;
  assign n10162 = n10161 ^ n10157 ;
  assign n10163 = ~n3884 & n10162 ;
  assign n10164 = n10163 ^ n10162 ;
  assign n10165 = n10164 ^ n10157 ;
  assign n10167 = n10166 ^ n10165 ;
  assign n10168 = ~n3927 & n10167 ;
  assign n10183 = n10168 ^ n10165 ;
  assign n10171 = n10163 ^ n10157 ;
  assign n10172 = n10171 ^ x284 ;
  assign n10173 = ~n3959 & n10172 ;
  assign n10174 = n10173 ^ x284 ;
  assign n10169 = n10168 ^ n10167 ;
  assign n10170 = n10169 ^ n10165 ;
  assign n10175 = n10174 ^ n10170 ;
  assign n10176 = n4004 & n10175 ;
  assign n10182 = n10176 ^ n10170 ;
  assign n10184 = n10183 ^ n10182 ;
  assign n10185 = n4046 & n10184 ;
  assign n10192 = n10185 ^ n10182 ;
  assign n10186 = n10185 ^ n10184 ;
  assign n10187 = n10186 ^ n10182 ;
  assign n10177 = n10176 ^ n10175 ;
  assign n10178 = n10177 ^ n10170 ;
  assign n10179 = n10178 ^ x252 ;
  assign n10180 = ~n4083 & n10179 ;
  assign n10181 = n10180 ^ x252 ;
  assign n10188 = n10187 ^ n10181 ;
  assign n10189 = n4127 & n10188 ;
  assign n10190 = n10189 ^ n10188 ;
  assign n10191 = n10190 ^ n10181 ;
  assign n10193 = n10192 ^ n10191 ;
  assign n10194 = n4201 & n10193 ;
  assign n10205 = n10194 ^ n10191 ;
  assign n10197 = n10189 ^ n10181 ;
  assign n10198 = n10197 ^ x220 ;
  assign n10199 = ~n4163 & n10198 ;
  assign n10200 = n10199 ^ x220 ;
  assign n10195 = n10194 ^ n10193 ;
  assign n10196 = n10195 ^ n10191 ;
  assign n10201 = n10200 ^ n10196 ;
  assign n10202 = ~n4245 & n10201 ;
  assign n10203 = n10202 ^ n10201 ;
  assign n10204 = n10203 ^ n10196 ;
  assign n10206 = n10205 ^ n10204 ;
  assign n10207 = ~n4288 & n10206 ;
  assign n10222 = n10207 ^ n10204 ;
  assign n10210 = n10202 ^ n10196 ;
  assign n10211 = n10210 ^ x188 ;
  assign n10212 = ~n4320 & n10211 ;
  assign n10213 = n10212 ^ x188 ;
  assign n10208 = n10207 ^ n10206 ;
  assign n10209 = n10208 ^ n10204 ;
  assign n10214 = n10213 ^ n10209 ;
  assign n10215 = n4365 & n10214 ;
  assign n10221 = n10215 ^ n10209 ;
  assign n10223 = n10222 ^ n10221 ;
  assign n10224 = n4407 & n10223 ;
  assign n10231 = n10224 ^ n10221 ;
  assign n10225 = n10224 ^ n10223 ;
  assign n10226 = n10225 ^ n10221 ;
  assign n10216 = n10215 ^ n10214 ;
  assign n10217 = n10216 ^ n10209 ;
  assign n10218 = n10217 ^ x156 ;
  assign n10219 = ~n4444 & n10218 ;
  assign n10220 = n10219 ^ x156 ;
  assign n10227 = n10226 ^ n10220 ;
  assign n10228 = n4488 & n10227 ;
  assign n10229 = n10228 ^ n10227 ;
  assign n10230 = n10229 ^ n10220 ;
  assign n10232 = n10231 ^ n10230 ;
  assign n10233 = n4562 & n10232 ;
  assign n10244 = n10233 ^ n10230 ;
  assign n10236 = n10228 ^ n10220 ;
  assign n10237 = n10236 ^ x124 ;
  assign n10238 = ~n4524 & n10237 ;
  assign n10239 = n10238 ^ x124 ;
  assign n10234 = n10233 ^ n10232 ;
  assign n10235 = n10234 ^ n10230 ;
  assign n10240 = n10239 ^ n10235 ;
  assign n10241 = ~n4606 & n10240 ;
  assign n10242 = n10241 ^ n10240 ;
  assign n10243 = n10242 ^ n10235 ;
  assign n10245 = n10244 ^ n10243 ;
  assign n10246 = ~n4649 & n10245 ;
  assign n10261 = n10246 ^ n10243 ;
  assign n10249 = n10241 ^ n10235 ;
  assign n10250 = n10249 ^ x92 ;
  assign n10251 = ~n4681 & n10250 ;
  assign n10252 = n10251 ^ x92 ;
  assign n10247 = n10246 ^ n10245 ;
  assign n10248 = n10247 ^ n10243 ;
  assign n10253 = n10252 ^ n10248 ;
  assign n10254 = n4726 & n10253 ;
  assign n10260 = n10254 ^ n10248 ;
  assign n10262 = n10261 ^ n10260 ;
  assign n10263 = n4772 & n10262 ;
  assign n10270 = n10263 ^ n10260 ;
  assign n10264 = n10263 ^ n10262 ;
  assign n10265 = n10264 ^ n10260 ;
  assign n10255 = n10254 ^ n10253 ;
  assign n10256 = n10255 ^ n10248 ;
  assign n10257 = n10256 ^ x60 ;
  assign n10258 = ~n4806 & n10257 ;
  assign n10259 = n10258 ^ x60 ;
  assign n10266 = n10265 ^ n10259 ;
  assign n10267 = n4850 & n10266 ;
  assign n10268 = n10267 ^ n10266 ;
  assign n10269 = n10268 ^ n10259 ;
  assign n10271 = n10270 ^ n10269 ;
  assign n10272 = ~n4893 & n10271 ;
  assign n10283 = n10272 ^ n10269 ;
  assign n10275 = n10267 ^ n10259 ;
  assign n10276 = n10275 ^ x28 ;
  assign n10277 = ~n4927 & n10276 ;
  assign n10278 = n10277 ^ x28 ;
  assign n10273 = n10272 ^ n10271 ;
  assign n10274 = n10273 ^ n10269 ;
  assign n10279 = n10278 ^ n10274 ;
  assign n10280 = ~n4972 & n10279 ;
  assign n10281 = n10280 ^ n10279 ;
  assign n10282 = n10281 ^ n10274 ;
  assign n10284 = n10283 ^ n10282 ;
  assign n10285 = n5009 & n10284 ;
  assign n10286 = n10285 ^ n10284 ;
  assign n10287 = n10286 ^ n10282 ;
  assign n10288 = x509 ^ x477 ;
  assign n10289 = n3371 & n10288 ;
  assign n10296 = n10289 ^ x477 ;
  assign n10290 = n10289 ^ n10288 ;
  assign n10291 = n10290 ^ x477 ;
  assign n10292 = n10291 ^ x445 ;
  assign n10293 = n3412 & n10292 ;
  assign n10294 = n10293 ^ n10292 ;
  assign n10295 = n10294 ^ x445 ;
  assign n10297 = n10296 ^ n10295 ;
  assign n10298 = n3451 & n10297 ;
  assign n10313 = n10298 ^ n10295 ;
  assign n10301 = n10293 ^ x445 ;
  assign n10302 = n10301 ^ x413 ;
  assign n10303 = ~n3484 & n10302 ;
  assign n10304 = n10303 ^ x413 ;
  assign n10299 = n10298 ^ n10297 ;
  assign n10300 = n10299 ^ n10295 ;
  assign n10305 = n10304 ^ n10300 ;
  assign n10306 = ~n3527 & n10305 ;
  assign n10312 = n10306 ^ n10300 ;
  assign n10314 = n10313 ^ n10312 ;
  assign n10315 = ~n3570 & n10314 ;
  assign n10316 = n10315 ^ n10314 ;
  assign n10317 = n10316 ^ n10312 ;
  assign n10307 = n10306 ^ n10305 ;
  assign n10308 = n10307 ^ n10300 ;
  assign n10309 = n10308 ^ x381 ;
  assign n10310 = ~n3602 & n10309 ;
  assign n10311 = n10310 ^ x381 ;
  assign n10318 = n10317 ^ n10311 ;
  assign n10319 = ~n3646 & n10318 ;
  assign n10326 = n10319 ^ n10311 ;
  assign n10325 = n10315 ^ n10312 ;
  assign n10327 = n10326 ^ n10325 ;
  assign n10328 = ~n3688 & n10327 ;
  assign n10335 = n10328 ^ n10325 ;
  assign n10329 = n10328 ^ n10327 ;
  assign n10330 = n10329 ^ n10325 ;
  assign n10320 = n10319 ^ n10318 ;
  assign n10321 = n10320 ^ n10311 ;
  assign n10322 = n10321 ^ x349 ;
  assign n10323 = ~n3724 & n10322 ;
  assign n10324 = n10323 ^ x349 ;
  assign n10331 = n10330 ^ n10324 ;
  assign n10332 = n3767 & n10331 ;
  assign n10333 = n10332 ^ n10331 ;
  assign n10334 = n10333 ^ n10324 ;
  assign n10336 = n10335 ^ n10334 ;
  assign n10337 = n3841 & n10336 ;
  assign n10348 = n10337 ^ n10334 ;
  assign n10340 = n10332 ^ n10324 ;
  assign n10341 = n10340 ^ x317 ;
  assign n10342 = ~n3803 & n10341 ;
  assign n10343 = n10342 ^ x317 ;
  assign n10338 = n10337 ^ n10336 ;
  assign n10339 = n10338 ^ n10334 ;
  assign n10344 = n10343 ^ n10339 ;
  assign n10345 = ~n3884 & n10344 ;
  assign n10346 = n10345 ^ n10344 ;
  assign n10347 = n10346 ^ n10339 ;
  assign n10349 = n10348 ^ n10347 ;
  assign n10350 = ~n3927 & n10349 ;
  assign n10365 = n10350 ^ n10347 ;
  assign n10353 = n10345 ^ n10339 ;
  assign n10354 = n10353 ^ x285 ;
  assign n10355 = ~n3959 & n10354 ;
  assign n10356 = n10355 ^ x285 ;
  assign n10351 = n10350 ^ n10349 ;
  assign n10352 = n10351 ^ n10347 ;
  assign n10357 = n10356 ^ n10352 ;
  assign n10358 = n4004 & n10357 ;
  assign n10364 = n10358 ^ n10352 ;
  assign n10366 = n10365 ^ n10364 ;
  assign n10367 = n4046 & n10366 ;
  assign n10374 = n10367 ^ n10364 ;
  assign n10368 = n10367 ^ n10366 ;
  assign n10369 = n10368 ^ n10364 ;
  assign n10359 = n10358 ^ n10357 ;
  assign n10360 = n10359 ^ n10352 ;
  assign n10361 = n10360 ^ x253 ;
  assign n10362 = ~n4083 & n10361 ;
  assign n10363 = n10362 ^ x253 ;
  assign n10370 = n10369 ^ n10363 ;
  assign n10371 = n4127 & n10370 ;
  assign n10372 = n10371 ^ n10370 ;
  assign n10373 = n10372 ^ n10363 ;
  assign n10375 = n10374 ^ n10373 ;
  assign n10376 = n4201 & n10375 ;
  assign n10387 = n10376 ^ n10373 ;
  assign n10379 = n10371 ^ n10363 ;
  assign n10380 = n10379 ^ x221 ;
  assign n10381 = ~n4163 & n10380 ;
  assign n10382 = n10381 ^ x221 ;
  assign n10377 = n10376 ^ n10375 ;
  assign n10378 = n10377 ^ n10373 ;
  assign n10383 = n10382 ^ n10378 ;
  assign n10384 = ~n4245 & n10383 ;
  assign n10385 = n10384 ^ n10383 ;
  assign n10386 = n10385 ^ n10378 ;
  assign n10388 = n10387 ^ n10386 ;
  assign n10389 = ~n4288 & n10388 ;
  assign n10404 = n10389 ^ n10386 ;
  assign n10392 = n10384 ^ n10378 ;
  assign n10393 = n10392 ^ x189 ;
  assign n10394 = ~n4320 & n10393 ;
  assign n10395 = n10394 ^ x189 ;
  assign n10390 = n10389 ^ n10388 ;
  assign n10391 = n10390 ^ n10386 ;
  assign n10396 = n10395 ^ n10391 ;
  assign n10397 = n4365 & n10396 ;
  assign n10403 = n10397 ^ n10391 ;
  assign n10405 = n10404 ^ n10403 ;
  assign n10406 = n4407 & n10405 ;
  assign n10413 = n10406 ^ n10403 ;
  assign n10407 = n10406 ^ n10405 ;
  assign n10408 = n10407 ^ n10403 ;
  assign n10398 = n10397 ^ n10396 ;
  assign n10399 = n10398 ^ n10391 ;
  assign n10400 = n10399 ^ x157 ;
  assign n10401 = ~n4444 & n10400 ;
  assign n10402 = n10401 ^ x157 ;
  assign n10409 = n10408 ^ n10402 ;
  assign n10410 = n4488 & n10409 ;
  assign n10411 = n10410 ^ n10409 ;
  assign n10412 = n10411 ^ n10402 ;
  assign n10414 = n10413 ^ n10412 ;
  assign n10415 = n4562 & n10414 ;
  assign n10426 = n10415 ^ n10412 ;
  assign n10418 = n10410 ^ n10402 ;
  assign n10419 = n10418 ^ x125 ;
  assign n10420 = ~n4524 & n10419 ;
  assign n10421 = n10420 ^ x125 ;
  assign n10416 = n10415 ^ n10414 ;
  assign n10417 = n10416 ^ n10412 ;
  assign n10422 = n10421 ^ n10417 ;
  assign n10423 = ~n4606 & n10422 ;
  assign n10424 = n10423 ^ n10422 ;
  assign n10425 = n10424 ^ n10417 ;
  assign n10427 = n10426 ^ n10425 ;
  assign n10428 = ~n4649 & n10427 ;
  assign n10443 = n10428 ^ n10425 ;
  assign n10431 = n10423 ^ n10417 ;
  assign n10432 = n10431 ^ x93 ;
  assign n10433 = ~n4681 & n10432 ;
  assign n10434 = n10433 ^ x93 ;
  assign n10429 = n10428 ^ n10427 ;
  assign n10430 = n10429 ^ n10425 ;
  assign n10435 = n10434 ^ n10430 ;
  assign n10436 = n4726 & n10435 ;
  assign n10442 = n10436 ^ n10430 ;
  assign n10444 = n10443 ^ n10442 ;
  assign n10445 = n4772 & n10444 ;
  assign n10452 = n10445 ^ n10442 ;
  assign n10446 = n10445 ^ n10444 ;
  assign n10447 = n10446 ^ n10442 ;
  assign n10437 = n10436 ^ n10435 ;
  assign n10438 = n10437 ^ n10430 ;
  assign n10439 = n10438 ^ x61 ;
  assign n10440 = ~n4806 & n10439 ;
  assign n10441 = n10440 ^ x61 ;
  assign n10448 = n10447 ^ n10441 ;
  assign n10449 = n4850 & n10448 ;
  assign n10450 = n10449 ^ n10448 ;
  assign n10451 = n10450 ^ n10441 ;
  assign n10453 = n10452 ^ n10451 ;
  assign n10454 = ~n4893 & n10453 ;
  assign n10465 = n10454 ^ n10451 ;
  assign n10457 = n10449 ^ n10441 ;
  assign n10458 = n10457 ^ x29 ;
  assign n10459 = ~n4927 & n10458 ;
  assign n10460 = n10459 ^ x29 ;
  assign n10455 = n10454 ^ n10453 ;
  assign n10456 = n10455 ^ n10451 ;
  assign n10461 = n10460 ^ n10456 ;
  assign n10462 = ~n4972 & n10461 ;
  assign n10463 = n10462 ^ n10461 ;
  assign n10464 = n10463 ^ n10456 ;
  assign n10466 = n10465 ^ n10464 ;
  assign n10467 = n5009 & n10466 ;
  assign n10468 = n10467 ^ n10466 ;
  assign n10469 = n10468 ^ n10464 ;
  assign n10470 = x510 ^ x478 ;
  assign n10471 = n3371 & n10470 ;
  assign n10478 = n10471 ^ x478 ;
  assign n10472 = n10471 ^ n10470 ;
  assign n10473 = n10472 ^ x478 ;
  assign n10474 = n10473 ^ x446 ;
  assign n10475 = n3412 & n10474 ;
  assign n10476 = n10475 ^ n10474 ;
  assign n10477 = n10476 ^ x446 ;
  assign n10479 = n10478 ^ n10477 ;
  assign n10480 = n3451 & n10479 ;
  assign n10495 = n10480 ^ n10477 ;
  assign n10483 = n10475 ^ x446 ;
  assign n10484 = n10483 ^ x414 ;
  assign n10485 = ~n3484 & n10484 ;
  assign n10486 = n10485 ^ x414 ;
  assign n10481 = n10480 ^ n10479 ;
  assign n10482 = n10481 ^ n10477 ;
  assign n10487 = n10486 ^ n10482 ;
  assign n10488 = ~n3527 & n10487 ;
  assign n10494 = n10488 ^ n10482 ;
  assign n10496 = n10495 ^ n10494 ;
  assign n10497 = ~n3570 & n10496 ;
  assign n10498 = n10497 ^ n10496 ;
  assign n10499 = n10498 ^ n10494 ;
  assign n10489 = n10488 ^ n10487 ;
  assign n10490 = n10489 ^ n10482 ;
  assign n10491 = n10490 ^ x382 ;
  assign n10492 = ~n3602 & n10491 ;
  assign n10493 = n10492 ^ x382 ;
  assign n10500 = n10499 ^ n10493 ;
  assign n10501 = ~n3646 & n10500 ;
  assign n10508 = n10501 ^ n10493 ;
  assign n10507 = n10497 ^ n10494 ;
  assign n10509 = n10508 ^ n10507 ;
  assign n10510 = ~n3688 & n10509 ;
  assign n10517 = n10510 ^ n10507 ;
  assign n10511 = n10510 ^ n10509 ;
  assign n10512 = n10511 ^ n10507 ;
  assign n10502 = n10501 ^ n10500 ;
  assign n10503 = n10502 ^ n10493 ;
  assign n10504 = n10503 ^ x350 ;
  assign n10505 = ~n3724 & n10504 ;
  assign n10506 = n10505 ^ x350 ;
  assign n10513 = n10512 ^ n10506 ;
  assign n10514 = n3767 & n10513 ;
  assign n10515 = n10514 ^ n10513 ;
  assign n10516 = n10515 ^ n10506 ;
  assign n10518 = n10517 ^ n10516 ;
  assign n10519 = n3841 & n10518 ;
  assign n10530 = n10519 ^ n10516 ;
  assign n10522 = n10514 ^ n10506 ;
  assign n10523 = n10522 ^ x318 ;
  assign n10524 = ~n3803 & n10523 ;
  assign n10525 = n10524 ^ x318 ;
  assign n10520 = n10519 ^ n10518 ;
  assign n10521 = n10520 ^ n10516 ;
  assign n10526 = n10525 ^ n10521 ;
  assign n10527 = ~n3884 & n10526 ;
  assign n10528 = n10527 ^ n10526 ;
  assign n10529 = n10528 ^ n10521 ;
  assign n10531 = n10530 ^ n10529 ;
  assign n10532 = ~n3927 & n10531 ;
  assign n10547 = n10532 ^ n10529 ;
  assign n10535 = n10527 ^ n10521 ;
  assign n10536 = n10535 ^ x286 ;
  assign n10537 = ~n3959 & n10536 ;
  assign n10538 = n10537 ^ x286 ;
  assign n10533 = n10532 ^ n10531 ;
  assign n10534 = n10533 ^ n10529 ;
  assign n10539 = n10538 ^ n10534 ;
  assign n10540 = n4004 & n10539 ;
  assign n10546 = n10540 ^ n10534 ;
  assign n10548 = n10547 ^ n10546 ;
  assign n10549 = n4046 & n10548 ;
  assign n10556 = n10549 ^ n10546 ;
  assign n10550 = n10549 ^ n10548 ;
  assign n10551 = n10550 ^ n10546 ;
  assign n10541 = n10540 ^ n10539 ;
  assign n10542 = n10541 ^ n10534 ;
  assign n10543 = n10542 ^ x254 ;
  assign n10544 = ~n4083 & n10543 ;
  assign n10545 = n10544 ^ x254 ;
  assign n10552 = n10551 ^ n10545 ;
  assign n10553 = n4127 & n10552 ;
  assign n10554 = n10553 ^ n10552 ;
  assign n10555 = n10554 ^ n10545 ;
  assign n10557 = n10556 ^ n10555 ;
  assign n10558 = n4201 & n10557 ;
  assign n10569 = n10558 ^ n10555 ;
  assign n10561 = n10553 ^ n10545 ;
  assign n10562 = n10561 ^ x222 ;
  assign n10563 = ~n4163 & n10562 ;
  assign n10564 = n10563 ^ x222 ;
  assign n10559 = n10558 ^ n10557 ;
  assign n10560 = n10559 ^ n10555 ;
  assign n10565 = n10564 ^ n10560 ;
  assign n10566 = ~n4245 & n10565 ;
  assign n10567 = n10566 ^ n10565 ;
  assign n10568 = n10567 ^ n10560 ;
  assign n10570 = n10569 ^ n10568 ;
  assign n10571 = ~n4288 & n10570 ;
  assign n10586 = n10571 ^ n10568 ;
  assign n10574 = n10566 ^ n10560 ;
  assign n10575 = n10574 ^ x190 ;
  assign n10576 = ~n4320 & n10575 ;
  assign n10577 = n10576 ^ x190 ;
  assign n10572 = n10571 ^ n10570 ;
  assign n10573 = n10572 ^ n10568 ;
  assign n10578 = n10577 ^ n10573 ;
  assign n10579 = n4365 & n10578 ;
  assign n10585 = n10579 ^ n10573 ;
  assign n10587 = n10586 ^ n10585 ;
  assign n10588 = n4407 & n10587 ;
  assign n10595 = n10588 ^ n10585 ;
  assign n10589 = n10588 ^ n10587 ;
  assign n10590 = n10589 ^ n10585 ;
  assign n10580 = n10579 ^ n10578 ;
  assign n10581 = n10580 ^ n10573 ;
  assign n10582 = n10581 ^ x158 ;
  assign n10583 = ~n4444 & n10582 ;
  assign n10584 = n10583 ^ x158 ;
  assign n10591 = n10590 ^ n10584 ;
  assign n10592 = n4488 & n10591 ;
  assign n10593 = n10592 ^ n10591 ;
  assign n10594 = n10593 ^ n10584 ;
  assign n10596 = n10595 ^ n10594 ;
  assign n10597 = n4562 & n10596 ;
  assign n10608 = n10597 ^ n10594 ;
  assign n10600 = n10592 ^ n10584 ;
  assign n10601 = n10600 ^ x126 ;
  assign n10602 = ~n4524 & n10601 ;
  assign n10603 = n10602 ^ x126 ;
  assign n10598 = n10597 ^ n10596 ;
  assign n10599 = n10598 ^ n10594 ;
  assign n10604 = n10603 ^ n10599 ;
  assign n10605 = ~n4606 & n10604 ;
  assign n10606 = n10605 ^ n10604 ;
  assign n10607 = n10606 ^ n10599 ;
  assign n10609 = n10608 ^ n10607 ;
  assign n10610 = ~n4649 & n10609 ;
  assign n10625 = n10610 ^ n10607 ;
  assign n10613 = n10605 ^ n10599 ;
  assign n10614 = n10613 ^ x94 ;
  assign n10615 = ~n4681 & n10614 ;
  assign n10616 = n10615 ^ x94 ;
  assign n10611 = n10610 ^ n10609 ;
  assign n10612 = n10611 ^ n10607 ;
  assign n10617 = n10616 ^ n10612 ;
  assign n10618 = n4726 & n10617 ;
  assign n10624 = n10618 ^ n10612 ;
  assign n10626 = n10625 ^ n10624 ;
  assign n10627 = n4772 & n10626 ;
  assign n10634 = n10627 ^ n10624 ;
  assign n10628 = n10627 ^ n10626 ;
  assign n10629 = n10628 ^ n10624 ;
  assign n10619 = n10618 ^ n10617 ;
  assign n10620 = n10619 ^ n10612 ;
  assign n10621 = n10620 ^ x62 ;
  assign n10622 = ~n4806 & n10621 ;
  assign n10623 = n10622 ^ x62 ;
  assign n10630 = n10629 ^ n10623 ;
  assign n10631 = n4850 & n10630 ;
  assign n10632 = n10631 ^ n10630 ;
  assign n10633 = n10632 ^ n10623 ;
  assign n10635 = n10634 ^ n10633 ;
  assign n10636 = ~n4893 & n10635 ;
  assign n10647 = n10636 ^ n10633 ;
  assign n10639 = n10631 ^ n10623 ;
  assign n10640 = n10639 ^ x30 ;
  assign n10641 = ~n4927 & n10640 ;
  assign n10642 = n10641 ^ x30 ;
  assign n10637 = n10636 ^ n10635 ;
  assign n10638 = n10637 ^ n10633 ;
  assign n10643 = n10642 ^ n10638 ;
  assign n10644 = ~n4972 & n10643 ;
  assign n10645 = n10644 ^ n10643 ;
  assign n10646 = n10645 ^ n10638 ;
  assign n10648 = n10647 ^ n10646 ;
  assign n10649 = n5009 & n10648 ;
  assign n10650 = n10649 ^ n10648 ;
  assign n10651 = n10650 ^ n10646 ;
  assign n10652 = x511 ^ x479 ;
  assign n10653 = n3371 & n10652 ;
  assign n10660 = n10653 ^ x479 ;
  assign n10654 = n10653 ^ n10652 ;
  assign n10655 = n10654 ^ x479 ;
  assign n10656 = n10655 ^ x447 ;
  assign n10657 = n3412 & n10656 ;
  assign n10658 = n10657 ^ n10656 ;
  assign n10659 = n10658 ^ x447 ;
  assign n10661 = n10660 ^ n10659 ;
  assign n10662 = n3451 & n10661 ;
  assign n10677 = n10662 ^ n10659 ;
  assign n10665 = n10657 ^ x447 ;
  assign n10666 = n10665 ^ x415 ;
  assign n10667 = ~n3484 & n10666 ;
  assign n10668 = n10667 ^ x415 ;
  assign n10663 = n10662 ^ n10661 ;
  assign n10664 = n10663 ^ n10659 ;
  assign n10669 = n10668 ^ n10664 ;
  assign n10670 = ~n3527 & n10669 ;
  assign n10676 = n10670 ^ n10664 ;
  assign n10678 = n10677 ^ n10676 ;
  assign n10679 = ~n3570 & n10678 ;
  assign n10680 = n10679 ^ n10678 ;
  assign n10681 = n10680 ^ n10676 ;
  assign n10671 = n10670 ^ n10669 ;
  assign n10672 = n10671 ^ n10664 ;
  assign n10673 = n10672 ^ x383 ;
  assign n10674 = ~n3602 & n10673 ;
  assign n10675 = n10674 ^ x383 ;
  assign n10682 = n10681 ^ n10675 ;
  assign n10683 = ~n3646 & n10682 ;
  assign n10690 = n10683 ^ n10675 ;
  assign n10689 = n10679 ^ n10676 ;
  assign n10691 = n10690 ^ n10689 ;
  assign n10692 = ~n3688 & n10691 ;
  assign n10699 = n10692 ^ n10689 ;
  assign n10693 = n10692 ^ n10691 ;
  assign n10694 = n10693 ^ n10689 ;
  assign n10684 = n10683 ^ n10682 ;
  assign n10685 = n10684 ^ n10675 ;
  assign n10686 = n10685 ^ x351 ;
  assign n10687 = ~n3724 & n10686 ;
  assign n10688 = n10687 ^ x351 ;
  assign n10695 = n10694 ^ n10688 ;
  assign n10696 = n3767 & n10695 ;
  assign n10697 = n10696 ^ n10695 ;
  assign n10698 = n10697 ^ n10688 ;
  assign n10700 = n10699 ^ n10698 ;
  assign n10701 = n3841 & n10700 ;
  assign n10712 = n10701 ^ n10698 ;
  assign n10704 = n10696 ^ n10688 ;
  assign n10705 = n10704 ^ x319 ;
  assign n10706 = ~n3803 & n10705 ;
  assign n10707 = n10706 ^ x319 ;
  assign n10702 = n10701 ^ n10700 ;
  assign n10703 = n10702 ^ n10698 ;
  assign n10708 = n10707 ^ n10703 ;
  assign n10709 = ~n3884 & n10708 ;
  assign n10710 = n10709 ^ n10708 ;
  assign n10711 = n10710 ^ n10703 ;
  assign n10713 = n10712 ^ n10711 ;
  assign n10714 = ~n3927 & n10713 ;
  assign n10729 = n10714 ^ n10711 ;
  assign n10717 = n10709 ^ n10703 ;
  assign n10718 = n10717 ^ x287 ;
  assign n10719 = ~n3959 & n10718 ;
  assign n10720 = n10719 ^ x287 ;
  assign n10715 = n10714 ^ n10713 ;
  assign n10716 = n10715 ^ n10711 ;
  assign n10721 = n10720 ^ n10716 ;
  assign n10722 = n4004 & n10721 ;
  assign n10728 = n10722 ^ n10716 ;
  assign n10730 = n10729 ^ n10728 ;
  assign n10731 = n4046 & n10730 ;
  assign n10738 = n10731 ^ n10728 ;
  assign n10732 = n10731 ^ n10730 ;
  assign n10733 = n10732 ^ n10728 ;
  assign n10723 = n10722 ^ n10721 ;
  assign n10724 = n10723 ^ n10716 ;
  assign n10725 = n10724 ^ x255 ;
  assign n10726 = ~n4083 & n10725 ;
  assign n10727 = n10726 ^ x255 ;
  assign n10734 = n10733 ^ n10727 ;
  assign n10735 = n4127 & n10734 ;
  assign n10736 = n10735 ^ n10734 ;
  assign n10737 = n10736 ^ n10727 ;
  assign n10739 = n10738 ^ n10737 ;
  assign n10740 = n4201 & n10739 ;
  assign n10751 = n10740 ^ n10737 ;
  assign n10743 = n10735 ^ n10727 ;
  assign n10744 = n10743 ^ x223 ;
  assign n10745 = ~n4163 & n10744 ;
  assign n10746 = n10745 ^ x223 ;
  assign n10741 = n10740 ^ n10739 ;
  assign n10742 = n10741 ^ n10737 ;
  assign n10747 = n10746 ^ n10742 ;
  assign n10748 = ~n4245 & n10747 ;
  assign n10749 = n10748 ^ n10747 ;
  assign n10750 = n10749 ^ n10742 ;
  assign n10752 = n10751 ^ n10750 ;
  assign n10753 = ~n4288 & n10752 ;
  assign n10768 = n10753 ^ n10750 ;
  assign n10756 = n10748 ^ n10742 ;
  assign n10757 = n10756 ^ x191 ;
  assign n10758 = ~n4320 & n10757 ;
  assign n10759 = n10758 ^ x191 ;
  assign n10754 = n10753 ^ n10752 ;
  assign n10755 = n10754 ^ n10750 ;
  assign n10760 = n10759 ^ n10755 ;
  assign n10761 = n4365 & n10760 ;
  assign n10767 = n10761 ^ n10755 ;
  assign n10769 = n10768 ^ n10767 ;
  assign n10770 = n4407 & n10769 ;
  assign n10777 = n10770 ^ n10767 ;
  assign n10771 = n10770 ^ n10769 ;
  assign n10772 = n10771 ^ n10767 ;
  assign n10762 = n10761 ^ n10760 ;
  assign n10763 = n10762 ^ n10755 ;
  assign n10764 = n10763 ^ x159 ;
  assign n10765 = ~n4444 & n10764 ;
  assign n10766 = n10765 ^ x159 ;
  assign n10773 = n10772 ^ n10766 ;
  assign n10774 = n4488 & n10773 ;
  assign n10775 = n10774 ^ n10773 ;
  assign n10776 = n10775 ^ n10766 ;
  assign n10778 = n10777 ^ n10776 ;
  assign n10779 = n4562 & n10778 ;
  assign n10790 = n10779 ^ n10776 ;
  assign n10782 = n10774 ^ n10766 ;
  assign n10783 = n10782 ^ x127 ;
  assign n10784 = ~n4524 & n10783 ;
  assign n10785 = n10784 ^ x127 ;
  assign n10780 = n10779 ^ n10778 ;
  assign n10781 = n10780 ^ n10776 ;
  assign n10786 = n10785 ^ n10781 ;
  assign n10787 = ~n4606 & n10786 ;
  assign n10788 = n10787 ^ n10786 ;
  assign n10789 = n10788 ^ n10781 ;
  assign n10791 = n10790 ^ n10789 ;
  assign n10792 = ~n4649 & n10791 ;
  assign n10807 = n10792 ^ n10789 ;
  assign n10795 = n10787 ^ n10781 ;
  assign n10796 = n10795 ^ x95 ;
  assign n10797 = ~n4681 & n10796 ;
  assign n10798 = n10797 ^ x95 ;
  assign n10793 = n10792 ^ n10791 ;
  assign n10794 = n10793 ^ n10789 ;
  assign n10799 = n10798 ^ n10794 ;
  assign n10800 = n4726 & n10799 ;
  assign n10806 = n10800 ^ n10794 ;
  assign n10808 = n10807 ^ n10806 ;
  assign n10809 = n4772 & n10808 ;
  assign n10816 = n10809 ^ n10806 ;
  assign n10810 = n10809 ^ n10808 ;
  assign n10811 = n10810 ^ n10806 ;
  assign n10801 = n10800 ^ n10799 ;
  assign n10802 = n10801 ^ n10794 ;
  assign n10803 = n10802 ^ x63 ;
  assign n10804 = ~n4806 & n10803 ;
  assign n10805 = n10804 ^ x63 ;
  assign n10812 = n10811 ^ n10805 ;
  assign n10813 = n4850 & n10812 ;
  assign n10814 = n10813 ^ n10812 ;
  assign n10815 = n10814 ^ n10805 ;
  assign n10817 = n10816 ^ n10815 ;
  assign n10818 = ~n4893 & n10817 ;
  assign n10829 = n10818 ^ n10815 ;
  assign n10821 = n10813 ^ n10805 ;
  assign n10822 = n10821 ^ x31 ;
  assign n10823 = ~n4927 & n10822 ;
  assign n10824 = n10823 ^ x31 ;
  assign n10819 = n10818 ^ n10817 ;
  assign n10820 = n10819 ^ n10815 ;
  assign n10825 = n10824 ^ n10820 ;
  assign n10826 = ~n4972 & n10825 ;
  assign n10827 = n10826 ^ n10825 ;
  assign n10828 = n10827 ^ n10820 ;
  assign n10830 = n10829 ^ n10828 ;
  assign n10831 = n5009 & n10830 ;
  assign n10832 = n10831 ^ n10830 ;
  assign n10833 = n10832 ^ n10828 ;
  assign n10834 = n5189 ^ n5186 ;
  assign n10835 = n5371 ^ n5368 ;
  assign n10836 = n5553 ^ n5550 ;
  assign n10837 = n5735 ^ n5732 ;
  assign n10838 = n5917 ^ n5914 ;
  assign n10839 = n6099 ^ n6096 ;
  assign n10840 = n6281 ^ n6278 ;
  assign n10841 = n6463 ^ n6460 ;
  assign n10842 = n6645 ^ n6642 ;
  assign n10843 = n6827 ^ n6824 ;
  assign n10844 = n7009 ^ n7006 ;
  assign n10845 = n7191 ^ n7188 ;
  assign n10846 = n7373 ^ n7370 ;
  assign n10847 = n7555 ^ n7552 ;
  assign n10848 = n7737 ^ n7734 ;
  assign n10849 = n7919 ^ n7916 ;
  assign n10850 = n8101 ^ n8098 ;
  assign n10851 = n8283 ^ n8280 ;
  assign n10852 = n8465 ^ n8462 ;
  assign n10853 = n8647 ^ n8644 ;
  assign n10854 = n8829 ^ n8826 ;
  assign n10855 = n9011 ^ n9008 ;
  assign n10856 = n9193 ^ n9190 ;
  assign n10857 = n9375 ^ n9372 ;
  assign n10858 = n9557 ^ n9554 ;
  assign n10859 = n9739 ^ n9736 ;
  assign n10860 = n9921 ^ n9918 ;
  assign n10861 = n10103 ^ n10100 ;
  assign n10862 = n10285 ^ n10282 ;
  assign n10863 = n10467 ^ n10464 ;
  assign n10864 = n10649 ^ n10646 ;
  assign n10865 = n10831 ^ n10828 ;
  assign n10866 = n5184 ^ n5176 ;
  assign n10867 = n5366 ^ n5360 ;
  assign n10868 = n5548 ^ n5542 ;
  assign n10869 = n5730 ^ n5724 ;
  assign n10870 = n5912 ^ n5906 ;
  assign n10871 = n6094 ^ n6088 ;
  assign n10872 = n6276 ^ n6270 ;
  assign n10873 = n6458 ^ n6452 ;
  assign n10874 = n6640 ^ n6634 ;
  assign n10875 = n6822 ^ n6816 ;
  assign n10876 = n7004 ^ n6998 ;
  assign n10877 = n7186 ^ n7180 ;
  assign n10878 = n7368 ^ n7362 ;
  assign n10879 = n7550 ^ n7544 ;
  assign n10880 = n7732 ^ n7726 ;
  assign n10881 = n7914 ^ n7908 ;
  assign n10882 = n8096 ^ n8090 ;
  assign n10883 = n8278 ^ n8272 ;
  assign n10884 = n8460 ^ n8454 ;
  assign n10885 = n8642 ^ n8636 ;
  assign n10886 = n8824 ^ n8818 ;
  assign n10887 = n9006 ^ n9000 ;
  assign n10888 = n9188 ^ n9182 ;
  assign n10889 = n9370 ^ n9364 ;
  assign n10890 = n9552 ^ n9546 ;
  assign n10891 = n9734 ^ n9728 ;
  assign n10892 = n9916 ^ n9910 ;
  assign n10893 = n10098 ^ n10092 ;
  assign n10894 = n10280 ^ n10274 ;
  assign n10895 = n10462 ^ n10456 ;
  assign n10896 = n10644 ^ n10638 ;
  assign n10897 = n10826 ^ n10820 ;
  assign y0 = n5191 ;
  assign y1 = n5373 ;
  assign y2 = n5555 ;
  assign y3 = n5737 ;
  assign y4 = n5919 ;
  assign y5 = n6101 ;
  assign y6 = n6283 ;
  assign y7 = n6465 ;
  assign y8 = n6647 ;
  assign y9 = n6829 ;
  assign y10 = n7011 ;
  assign y11 = n7193 ;
  assign y12 = n7375 ;
  assign y13 = n7557 ;
  assign y14 = n7739 ;
  assign y15 = n7921 ;
  assign y16 = n8103 ;
  assign y17 = n8285 ;
  assign y18 = n8467 ;
  assign y19 = n8649 ;
  assign y20 = n8831 ;
  assign y21 = n9013 ;
  assign y22 = n9195 ;
  assign y23 = n9377 ;
  assign y24 = n9559 ;
  assign y25 = n9741 ;
  assign y26 = n9923 ;
  assign y27 = n10105 ;
  assign y28 = n10287 ;
  assign y29 = n10469 ;
  assign y30 = n10651 ;
  assign y31 = n10833 ;
  assign y32 = n10834 ;
  assign y33 = n10835 ;
  assign y34 = n10836 ;
  assign y35 = n10837 ;
  assign y36 = n10838 ;
  assign y37 = n10839 ;
  assign y38 = n10840 ;
  assign y39 = n10841 ;
  assign y40 = n10842 ;
  assign y41 = n10843 ;
  assign y42 = n10844 ;
  assign y43 = n10845 ;
  assign y44 = n10846 ;
  assign y45 = n10847 ;
  assign y46 = n10848 ;
  assign y47 = n10849 ;
  assign y48 = n10850 ;
  assign y49 = n10851 ;
  assign y50 = n10852 ;
  assign y51 = n10853 ;
  assign y52 = n10854 ;
  assign y53 = n10855 ;
  assign y54 = n10856 ;
  assign y55 = n10857 ;
  assign y56 = n10858 ;
  assign y57 = n10859 ;
  assign y58 = n10860 ;
  assign y59 = n10861 ;
  assign y60 = n10862 ;
  assign y61 = n10863 ;
  assign y62 = n10864 ;
  assign y63 = n10865 ;
  assign y64 = n10866 ;
  assign y65 = n10867 ;
  assign y66 = n10868 ;
  assign y67 = n10869 ;
  assign y68 = n10870 ;
  assign y69 = n10871 ;
  assign y70 = n10872 ;
  assign y71 = n10873 ;
  assign y72 = n10874 ;
  assign y73 = n10875 ;
  assign y74 = n10876 ;
  assign y75 = n10877 ;
  assign y76 = n10878 ;
  assign y77 = n10879 ;
  assign y78 = n10880 ;
  assign y79 = n10881 ;
  assign y80 = n10882 ;
  assign y81 = n10883 ;
  assign y82 = n10884 ;
  assign y83 = n10885 ;
  assign y84 = n10886 ;
  assign y85 = n10887 ;
  assign y86 = n10888 ;
  assign y87 = n10889 ;
  assign y88 = n10890 ;
  assign y89 = n10891 ;
  assign y90 = n10892 ;
  assign y91 = n10893 ;
  assign y92 = n10894 ;
  assign y93 = n10895 ;
  assign y94 = n10896 ;
  assign y95 = n10897 ;
endmodule
