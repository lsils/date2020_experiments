module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 ;
  assign n15 = x4 & x5 ;
  assign n16 = n15 ^ x5 ;
  assign n17 = n16 ^ x4 ;
  assign n12 = x2 & x3 ;
  assign n13 = n12 ^ x3 ;
  assign n14 = n13 ^ x2 ;
  assign n18 = n17 ^ n14 ;
  assign n9 = x6 & x7 ;
  assign n10 = n9 ^ x7 ;
  assign n11 = n10 ^ x6 ;
  assign n19 = n18 ^ n11 ;
  assign n20 = x0 & x1 ;
  assign n21 = n20 ^ x1 ;
  assign n22 = n21 ^ x0 ;
  assign n23 = ~n19 & ~n22 ;
  assign n24 = n14 ^ n11 ;
  assign n25 = ~n18 & n24 ;
  assign n26 = n25 ^ n11 ;
  assign n66 = ~n23 & n26 ;
  assign n27 = n26 ^ n23 ;
  assign n67 = n66 ^ n27 ;
  assign n29 = n9 ^ x6 ;
  assign n28 = n15 ^ x4 ;
  assign n30 = n29 ^ n28 ;
  assign n31 = n12 ^ x2 ;
  assign n32 = n31 ^ n28 ;
  assign n33 = ~n30 & n32 ;
  assign n34 = n33 ^ n31 ;
  assign n35 = n31 ^ n30 ;
  assign n36 = n20 ^ x0 ;
  assign n37 = n35 & n36 ;
  assign n38 = ~n34 & ~n37 ;
  assign n39 = n38 ^ n37 ;
  assign n40 = n39 ^ n34 ;
  assign n68 = n67 ^ n40 ;
  assign n43 = n15 ^ n9 ;
  assign n44 = n43 ^ n12 ;
  assign n53 = n20 & n44 ;
  assign n50 = n15 ^ n12 ;
  assign n51 = ~n43 & n50 ;
  assign n52 = n51 ^ n12 ;
  assign n54 = n53 ^ n52 ;
  assign n46 = n16 ^ n10 ;
  assign n56 = n16 ^ n13 ;
  assign n57 = ~n46 & n56 ;
  assign n58 = n57 ^ n13 ;
  assign n47 = n46 ^ n13 ;
  assign n59 = n21 & n47 ;
  assign n60 = ~n58 & ~n59 ;
  assign n64 = ~n54 & n60 ;
  assign n41 = n40 ^ n38 ;
  assign n42 = n27 & ~n41 ;
  assign n45 = n44 ^ n20 ;
  assign n48 = n47 ^ n21 ;
  assign n49 = ~n45 & n48 ;
  assign n55 = n54 ^ n49 ;
  assign n61 = n60 ^ n49 ;
  assign n62 = ~n55 & n61 ;
  assign n63 = n42 & n62 ;
  assign n65 = n64 ^ n63 ;
  assign n69 = n68 ^ n65 ;
  assign n70 = n62 ^ n54 ;
  assign n71 = n70 ^ n38 ;
  assign n72 = ~n69 & ~n71 ;
  assign n73 = n72 ^ n70 ;
  assign y0 = n73 ;
  assign y1 = n69 ;
endmodule
