module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , y0 , y1 , y2 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 ;
  output y0 , y1 , y2 ;
  wire n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 ;
  assign n112 = x15 & x16 ;
  assign n113 = n112 ^ x16 ;
  assign n114 = x17 & n113 ;
  assign n468 = n114 ^ n113 ;
  assign n109 = x12 & x13 ;
  assign n110 = n109 ^ x13 ;
  assign n111 = x14 & n110 ;
  assign n467 = n111 ^ n110 ;
  assign n469 = n468 ^ n467 ;
  assign n116 = x9 & x10 ;
  assign n117 = n116 ^ x10 ;
  assign n118 = x11 & n117 ;
  assign n466 = n118 ^ n117 ;
  assign n475 = n467 ^ n466 ;
  assign n476 = ~n469 & n475 ;
  assign n477 = n476 ^ n466 ;
  assign n101 = x18 & x19 ;
  assign n102 = n101 ^ x19 ;
  assign n103 = x20 & n102 ;
  assign n459 = n103 ^ n102 ;
  assign n97 = x24 & x25 ;
  assign n98 = n97 ^ x25 ;
  assign n99 = x26 & n98 ;
  assign n457 = n99 ^ n98 ;
  assign n94 = x21 & x22 ;
  assign n95 = n94 ^ x22 ;
  assign n96 = x23 & n95 ;
  assign n456 = n96 ^ n95 ;
  assign n458 = n457 ^ n456 ;
  assign n464 = n459 ^ n458 ;
  assign n105 = x6 & x7 ;
  assign n106 = n105 ^ x7 ;
  assign n107 = x8 & n106 ;
  assign n463 = n107 ^ n106 ;
  assign n465 = n464 ^ n463 ;
  assign n470 = n469 ^ n466 ;
  assign n471 = n470 ^ n463 ;
  assign n472 = ~n465 & n471 ;
  assign n473 = n472 ^ n470 ;
  assign n460 = n459 ^ n456 ;
  assign n461 = ~n458 & n460 ;
  assign n462 = n461 ^ n459 ;
  assign n474 = n473 ^ n462 ;
  assign n478 = n477 ^ n474 ;
  assign n67 = x36 & x37 ;
  assign n68 = n67 ^ x37 ;
  assign n69 = x38 & n68 ;
  assign n442 = n69 ^ n68 ;
  assign n64 = x33 & x34 ;
  assign n65 = n64 ^ x34 ;
  assign n66 = x35 & n65 ;
  assign n441 = n66 ^ n65 ;
  assign n443 = n442 ^ n441 ;
  assign n71 = x30 & x31 ;
  assign n72 = n71 ^ x31 ;
  assign n73 = x32 & n72 ;
  assign n440 = n73 ^ n72 ;
  assign n449 = n441 ^ n440 ;
  assign n450 = ~n443 & n449 ;
  assign n451 = n450 ^ n440 ;
  assign n60 = x27 & x28 ;
  assign n61 = n60 ^ x28 ;
  assign n62 = x29 & n61 ;
  assign n438 = n62 ^ n61 ;
  assign n52 = x39 & x40 ;
  assign n53 = n52 ^ x40 ;
  assign n54 = x41 & n53 ;
  assign n433 = n54 ^ n53 ;
  assign n56 = x45 & x46 ;
  assign n57 = n56 ^ x46 ;
  assign n58 = x47 & n57 ;
  assign n431 = n58 ^ n57 ;
  assign n49 = x42 & x43 ;
  assign n50 = n49 ^ x43 ;
  assign n51 = x44 & n50 ;
  assign n430 = n51 ^ n50 ;
  assign n432 = n431 ^ n430 ;
  assign n437 = n433 ^ n432 ;
  assign n439 = n438 ^ n437 ;
  assign n444 = n443 ^ n440 ;
  assign n445 = n444 ^ n437 ;
  assign n446 = ~n439 & n445 ;
  assign n447 = n446 ^ n444 ;
  assign n434 = n433 ^ n430 ;
  assign n435 = ~n432 & n434 ;
  assign n436 = n435 ^ n433 ;
  assign n448 = n447 ^ n436 ;
  assign n455 = n451 ^ n448 ;
  assign n479 = n478 ^ n455 ;
  assign n481 = n470 ^ n465 ;
  assign n90 = x3 & x4 ;
  assign n91 = n90 ^ x4 ;
  assign n92 = x5 & n91 ;
  assign n480 = n92 ^ n91 ;
  assign n482 = n481 ^ n480 ;
  assign n483 = n444 ^ n439 ;
  assign n484 = n483 ^ n480 ;
  assign n485 = ~n482 & n484 ;
  assign n486 = n485 ^ n483 ;
  assign n487 = n486 ^ n455 ;
  assign n488 = ~n479 & n487 ;
  assign n489 = n488 ^ n486 ;
  assign n452 = n451 ^ n436 ;
  assign n453 = ~n448 & n452 ;
  assign n454 = n453 ^ n451 ;
  assign n490 = n489 ^ n454 ;
  assign n491 = n477 ^ n473 ;
  assign n492 = n474 & ~n491 ;
  assign n493 = n492 ^ n462 ;
  assign n494 = n493 ^ n489 ;
  assign n495 = n490 & ~n494 ;
  assign n496 = n495 ^ n454 ;
  assign n497 = n483 ^ n482 ;
  assign n147 = x0 & x1 ;
  assign n148 = n147 ^ x1 ;
  assign n149 = x2 & n148 ;
  assign n498 = n149 ^ n148 ;
  assign n499 = n497 & n498 ;
  assign n500 = n486 ^ n479 ;
  assign n501 = n499 & n500 ;
  assign n502 = n493 ^ n490 ;
  assign n503 = n501 & n502 ;
  assign n505 = ~n496 & ~n503 ;
  assign n504 = n503 ^ n496 ;
  assign n506 = n505 ^ n504 ;
  assign n161 = x41 & n52 ;
  assign n517 = n161 ^ n52 ;
  assign n159 = x47 & n56 ;
  assign n515 = n159 ^ n56 ;
  assign n158 = x44 & n49 ;
  assign n514 = n158 ^ n49 ;
  assign n516 = n515 ^ n514 ;
  assign n522 = n517 ^ n516 ;
  assign n163 = x29 & n60 ;
  assign n521 = n163 ^ n60 ;
  assign n523 = n522 ^ n521 ;
  assign n168 = x32 & n71 ;
  assign n510 = n168 ^ n71 ;
  assign n166 = x38 & n67 ;
  assign n508 = n166 ^ n67 ;
  assign n165 = x35 & n64 ;
  assign n507 = n165 ^ n64 ;
  assign n509 = n508 ^ n507 ;
  assign n524 = n510 ^ n509 ;
  assign n525 = n524 ^ n522 ;
  assign n526 = n523 & ~n525 ;
  assign n527 = n526 ^ n521 ;
  assign n518 = n517 ^ n514 ;
  assign n519 = ~n516 & n518 ;
  assign n520 = n519 ^ n517 ;
  assign n528 = n527 ^ n520 ;
  assign n511 = n510 ^ n507 ;
  assign n512 = ~n509 & n511 ;
  assign n513 = n512 ^ n510 ;
  assign n564 = n527 ^ n513 ;
  assign n565 = n528 & ~n564 ;
  assign n566 = n565 ^ n520 ;
  assign n185 = x5 & n90 ;
  assign n531 = n185 ^ n90 ;
  assign n530 = n524 ^ n523 ;
  assign n532 = n531 ^ n530 ;
  assign n195 = x17 & n112 ;
  assign n542 = n195 ^ n112 ;
  assign n194 = x14 & n109 ;
  assign n541 = n194 ^ n109 ;
  assign n543 = n542 ^ n541 ;
  assign n197 = x11 & n116 ;
  assign n540 = n197 ^ n116 ;
  assign n544 = n543 ^ n540 ;
  assign n188 = x26 & n97 ;
  assign n536 = n188 ^ n97 ;
  assign n187 = x23 & n94 ;
  assign n535 = n187 ^ n94 ;
  assign n537 = n536 ^ n535 ;
  assign n190 = x20 & n101 ;
  assign n534 = n190 ^ n101 ;
  assign n538 = n537 ^ n534 ;
  assign n192 = x8 & n105 ;
  assign n533 = n192 ^ n105 ;
  assign n539 = n538 ^ n533 ;
  assign n545 = n544 ^ n539 ;
  assign n546 = n545 ^ n531 ;
  assign n547 = n532 & ~n546 ;
  assign n548 = n547 ^ n530 ;
  assign n529 = n528 ^ n513 ;
  assign n549 = n548 ^ n529 ;
  assign n557 = n541 ^ n540 ;
  assign n558 = ~n543 & n557 ;
  assign n559 = n558 ^ n540 ;
  assign n553 = n544 ^ n538 ;
  assign n554 = n539 & ~n553 ;
  assign n555 = n554 ^ n533 ;
  assign n550 = n535 ^ n534 ;
  assign n551 = ~n537 & n550 ;
  assign n552 = n551 ^ n534 ;
  assign n556 = n555 ^ n552 ;
  assign n560 = n559 ^ n556 ;
  assign n561 = n560 ^ n529 ;
  assign n562 = ~n549 & n561 ;
  assign n563 = n562 ^ n560 ;
  assign n567 = n566 ^ n563 ;
  assign n568 = n559 ^ n555 ;
  assign n569 = n556 & ~n568 ;
  assign n570 = n569 ^ n552 ;
  assign n571 = n570 ^ n563 ;
  assign n572 = n567 & n571 ;
  assign n573 = n572 ^ n563 ;
  assign n574 = n545 ^ n532 ;
  assign n227 = x2 & n147 ;
  assign n575 = n227 ^ n147 ;
  assign n576 = n574 & n575 ;
  assign n577 = n560 ^ n549 ;
  assign n578 = n576 & n577 ;
  assign n579 = n570 ^ n567 ;
  assign n580 = n578 & n579 ;
  assign n582 = ~n573 & ~n580 ;
  assign n581 = n580 ^ n573 ;
  assign n583 = n582 ^ n581 ;
  assign n584 = n506 & n583 ;
  assign n333 = n65 ^ x33 ;
  assign n334 = x35 & ~n333 ;
  assign n597 = n334 ^ n333 ;
  assign n336 = n72 ^ x30 ;
  assign n337 = x32 & ~n336 ;
  assign n596 = n337 ^ n336 ;
  assign n598 = n597 ^ n596 ;
  assign n331 = n68 ^ x36 ;
  assign n332 = x38 & ~n331 ;
  assign n595 = n332 ^ n331 ;
  assign n604 = n596 ^ n595 ;
  assign n605 = ~n598 & n604 ;
  assign n606 = n605 ^ n595 ;
  assign n344 = n57 ^ x45 ;
  assign n345 = x47 & ~n344 ;
  assign n588 = n345 ^ n344 ;
  assign n347 = n53 ^ x39 ;
  assign n348 = x41 & ~n347 ;
  assign n586 = n348 ^ n347 ;
  assign n342 = n50 ^ x42 ;
  assign n343 = x44 & ~n342 ;
  assign n585 = n343 ^ n342 ;
  assign n587 = n586 ^ n585 ;
  assign n593 = n588 ^ n587 ;
  assign n339 = n61 ^ x27 ;
  assign n340 = x29 & ~n339 ;
  assign n592 = n340 ^ n339 ;
  assign n594 = n593 ^ n592 ;
  assign n599 = n598 ^ n595 ;
  assign n600 = n599 ^ n593 ;
  assign n601 = n594 & ~n600 ;
  assign n602 = n601 ^ n592 ;
  assign n589 = n588 ^ n585 ;
  assign n590 = ~n587 & n589 ;
  assign n591 = n590 ^ n588 ;
  assign n603 = n602 ^ n591 ;
  assign n629 = n606 ^ n603 ;
  assign n611 = n599 ^ n594 ;
  assign n367 = n91 ^ x3 ;
  assign n368 = x5 & ~n367 ;
  assign n610 = n368 ^ n367 ;
  assign n612 = n611 ^ n610 ;
  assign n375 = n117 ^ x9 ;
  assign n376 = x11 & ~n375 ;
  assign n622 = n376 ^ n375 ;
  assign n372 = n110 ^ x12 ;
  assign n373 = x14 & ~n372 ;
  assign n621 = n373 ^ n372 ;
  assign n623 = n622 ^ n621 ;
  assign n370 = n113 ^ x15 ;
  assign n371 = x17 & ~n370 ;
  assign n620 = n371 ^ n370 ;
  assign n624 = n623 ^ n620 ;
  assign n383 = n102 ^ x18 ;
  assign n384 = x20 & ~n383 ;
  assign n616 = n384 ^ n383 ;
  assign n380 = n95 ^ x21 ;
  assign n381 = x23 & ~n380 ;
  assign n615 = n381 ^ n380 ;
  assign n617 = n616 ^ n615 ;
  assign n378 = n98 ^ x24 ;
  assign n379 = x26 & ~n378 ;
  assign n614 = n379 ^ n378 ;
  assign n618 = n617 ^ n614 ;
  assign n386 = n106 ^ x6 ;
  assign n387 = x8 & ~n386 ;
  assign n613 = n387 ^ n386 ;
  assign n619 = n618 ^ n613 ;
  assign n625 = n624 ^ n619 ;
  assign n626 = n625 ^ n611 ;
  assign n627 = n612 & ~n626 ;
  assign n628 = n627 ^ n610 ;
  assign n630 = n629 ^ n628 ;
  assign n638 = n621 ^ n620 ;
  assign n639 = ~n623 & n638 ;
  assign n640 = n639 ^ n620 ;
  assign n634 = n615 ^ n614 ;
  assign n635 = ~n617 & n634 ;
  assign n636 = n635 ^ n614 ;
  assign n631 = n624 ^ n618 ;
  assign n632 = n619 & ~n631 ;
  assign n633 = n632 ^ n613 ;
  assign n637 = n636 ^ n633 ;
  assign n641 = n640 ^ n637 ;
  assign n642 = n641 ^ n629 ;
  assign n643 = n630 & ~n642 ;
  assign n644 = n643 ^ n628 ;
  assign n607 = n606 ^ n591 ;
  assign n608 = n603 & n607 ;
  assign n609 = n608 ^ n591 ;
  assign n645 = n644 ^ n609 ;
  assign n646 = n640 ^ n636 ;
  assign n647 = n637 & ~n646 ;
  assign n648 = n647 ^ n633 ;
  assign n649 = n648 ^ n644 ;
  assign n650 = n645 & ~n649 ;
  assign n651 = n650 ^ n609 ;
  assign n652 = n641 ^ n630 ;
  assign n653 = n625 ^ n612 ;
  assign n418 = n148 ^ x0 ;
  assign n419 = x2 & ~n418 ;
  assign n654 = n419 ^ n418 ;
  assign n655 = ~n653 & ~n654 ;
  assign n656 = ~n652 & n655 ;
  assign n657 = n648 ^ n645 ;
  assign n658 = n656 & ~n657 ;
  assign n660 = n651 & ~n658 ;
  assign n659 = n658 ^ n651 ;
  assign n661 = n660 ^ n659 ;
  assign n248 = n52 ^ x39 ;
  assign n249 = x41 & n248 ;
  assign n672 = n249 ^ n248 ;
  assign n251 = n56 ^ x45 ;
  assign n252 = x47 & n251 ;
  assign n670 = n252 ^ n251 ;
  assign n246 = n49 ^ x42 ;
  assign n247 = x44 & n246 ;
  assign n669 = n247 ^ n246 ;
  assign n671 = n670 ^ n669 ;
  assign n677 = n672 ^ n671 ;
  assign n257 = n60 ^ x27 ;
  assign n258 = x29 & n257 ;
  assign n676 = n258 ^ n257 ;
  assign n678 = n677 ^ n676 ;
  assign n241 = n71 ^ x30 ;
  assign n242 = x32 & n241 ;
  assign n665 = n242 ^ n241 ;
  assign n238 = n67 ^ x36 ;
  assign n239 = x38 & n238 ;
  assign n663 = n239 ^ n238 ;
  assign n236 = n64 ^ x33 ;
  assign n237 = x35 & n236 ;
  assign n662 = n237 ^ n236 ;
  assign n664 = n663 ^ n662 ;
  assign n679 = n665 ^ n664 ;
  assign n680 = n679 ^ n677 ;
  assign n681 = n678 & ~n680 ;
  assign n682 = n681 ^ n676 ;
  assign n673 = n672 ^ n669 ;
  assign n674 = ~n671 & n673 ;
  assign n675 = n674 ^ n672 ;
  assign n683 = n682 ^ n675 ;
  assign n666 = n665 ^ n662 ;
  assign n667 = ~n664 & n666 ;
  assign n668 = n667 ^ n665 ;
  assign n719 = n682 ^ n668 ;
  assign n720 = n683 & ~n719 ;
  assign n721 = n720 ^ n675 ;
  assign n268 = n90 ^ x3 ;
  assign n269 = x5 & n268 ;
  assign n686 = n269 ^ n268 ;
  assign n685 = n679 ^ n678 ;
  assign n687 = n686 ^ n685 ;
  assign n273 = n112 ^ x15 ;
  assign n274 = x17 & n273 ;
  assign n697 = n274 ^ n273 ;
  assign n271 = n109 ^ x12 ;
  assign n272 = x14 & n271 ;
  assign n696 = n272 ^ n271 ;
  assign n698 = n697 ^ n696 ;
  assign n276 = n116 ^ x9 ;
  assign n277 = x11 & n276 ;
  assign n695 = n277 ^ n276 ;
  assign n699 = n698 ^ n695 ;
  assign n281 = n97 ^ x24 ;
  assign n282 = x26 & n281 ;
  assign n691 = n282 ^ n281 ;
  assign n279 = n94 ^ x21 ;
  assign n280 = x23 & n279 ;
  assign n690 = n280 ^ n279 ;
  assign n692 = n691 ^ n690 ;
  assign n284 = n101 ^ x18 ;
  assign n285 = x20 & n284 ;
  assign n689 = n285 ^ n284 ;
  assign n693 = n692 ^ n689 ;
  assign n287 = n105 ^ x6 ;
  assign n288 = x8 & n287 ;
  assign n688 = n288 ^ n287 ;
  assign n694 = n693 ^ n688 ;
  assign n700 = n699 ^ n694 ;
  assign n701 = n700 ^ n686 ;
  assign n702 = n687 & ~n701 ;
  assign n703 = n702 ^ n685 ;
  assign n684 = n683 ^ n668 ;
  assign n704 = n703 ^ n684 ;
  assign n712 = n696 ^ n695 ;
  assign n713 = ~n698 & n712 ;
  assign n714 = n713 ^ n695 ;
  assign n708 = n699 ^ n693 ;
  assign n709 = n694 & ~n708 ;
  assign n710 = n709 ^ n688 ;
  assign n705 = n690 ^ n689 ;
  assign n706 = ~n692 & n705 ;
  assign n707 = n706 ^ n689 ;
  assign n711 = n710 ^ n707 ;
  assign n715 = n714 ^ n711 ;
  assign n716 = n715 ^ n684 ;
  assign n717 = ~n704 & n716 ;
  assign n718 = n717 ^ n715 ;
  assign n722 = n721 ^ n718 ;
  assign n723 = n714 ^ n710 ;
  assign n724 = n711 & ~n723 ;
  assign n725 = n724 ^ n707 ;
  assign n726 = n725 ^ n718 ;
  assign n727 = n722 & n726 ;
  assign n728 = n727 ^ n718 ;
  assign n729 = n700 ^ n687 ;
  assign n321 = n147 ^ x0 ;
  assign n322 = x2 & n321 ;
  assign n730 = n322 ^ n321 ;
  assign n731 = n729 & n730 ;
  assign n732 = n715 ^ n704 ;
  assign n733 = n731 & n732 ;
  assign n734 = n725 ^ n722 ;
  assign n735 = n733 & n734 ;
  assign n737 = ~n728 & ~n735 ;
  assign n736 = n735 ^ n728 ;
  assign n738 = n737 ^ n736 ;
  assign n739 = ~n661 & n738 ;
  assign n740 = n584 & ~n739 ;
  assign n741 = n740 ^ n584 ;
  assign n70 = n69 ^ n66 ;
  assign n74 = n73 ^ n70 ;
  assign n55 = n54 ^ n51 ;
  assign n59 = n58 ^ n55 ;
  assign n63 = n62 ^ n59 ;
  assign n89 = n74 ^ n63 ;
  assign n93 = n92 ^ n89 ;
  assign n115 = n114 ^ n111 ;
  assign n119 = n118 ^ n115 ;
  assign n100 = n99 ^ n96 ;
  assign n104 = n103 ^ n100 ;
  assign n108 = n107 ^ n104 ;
  assign n120 = n119 ^ n108 ;
  assign n121 = n120 ^ n89 ;
  assign n122 = n93 & ~n121 ;
  assign n123 = n122 ^ n92 ;
  assign n82 = n73 ^ n69 ;
  assign n83 = n70 & ~n82 ;
  assign n84 = n83 ^ n66 ;
  assign n78 = n58 ^ n51 ;
  assign n79 = ~n55 & n78 ;
  assign n80 = n79 ^ n58 ;
  assign n75 = n74 ^ n62 ;
  assign n76 = ~n63 & n75 ;
  assign n77 = n76 ^ n74 ;
  assign n81 = n80 ^ n77 ;
  assign n88 = n84 ^ n81 ;
  assign n124 = n123 ^ n88 ;
  assign n132 = n118 ^ n114 ;
  assign n133 = n115 & ~n132 ;
  assign n134 = n133 ^ n111 ;
  assign n128 = n103 ^ n99 ;
  assign n129 = n100 & ~n128 ;
  assign n130 = n129 ^ n96 ;
  assign n125 = n119 ^ n107 ;
  assign n126 = n108 & ~n125 ;
  assign n127 = n126 ^ n104 ;
  assign n131 = n130 ^ n127 ;
  assign n135 = n134 ^ n131 ;
  assign n136 = n135 ^ n88 ;
  assign n137 = n124 & ~n136 ;
  assign n138 = n137 ^ n123 ;
  assign n85 = n84 ^ n80 ;
  assign n86 = n81 & ~n85 ;
  assign n87 = n86 ^ n77 ;
  assign n139 = n138 ^ n87 ;
  assign n140 = n134 ^ n130 ;
  assign n141 = n131 & ~n140 ;
  assign n142 = n141 ^ n127 ;
  assign n143 = n142 ^ n87 ;
  assign n144 = ~n139 & n143 ;
  assign n145 = n144 ^ n142 ;
  assign n146 = n142 ^ n139 ;
  assign n150 = n120 ^ n93 ;
  assign n151 = n149 & n150 ;
  assign n152 = n135 ^ n124 ;
  assign n153 = n151 & n152 ;
  assign n154 = n146 & n153 ;
  assign n156 = ~n145 & ~n154 ;
  assign n155 = n154 ^ n145 ;
  assign n157 = n156 ^ n155 ;
  assign n167 = n166 ^ n165 ;
  assign n169 = n168 ^ n167 ;
  assign n160 = n159 ^ n158 ;
  assign n162 = n161 ^ n160 ;
  assign n164 = n163 ^ n162 ;
  assign n184 = n169 ^ n164 ;
  assign n186 = n185 ^ n184 ;
  assign n196 = n195 ^ n194 ;
  assign n198 = n197 ^ n196 ;
  assign n189 = n188 ^ n187 ;
  assign n191 = n190 ^ n189 ;
  assign n193 = n192 ^ n191 ;
  assign n199 = n198 ^ n193 ;
  assign n200 = n199 ^ n185 ;
  assign n201 = n186 & ~n200 ;
  assign n202 = n201 ^ n184 ;
  assign n177 = n168 ^ n166 ;
  assign n178 = n167 & ~n177 ;
  assign n179 = n178 ^ n165 ;
  assign n173 = n161 ^ n159 ;
  assign n174 = ~n160 & n173 ;
  assign n175 = n174 ^ n161 ;
  assign n170 = n169 ^ n163 ;
  assign n171 = ~n164 & n170 ;
  assign n172 = n171 ^ n169 ;
  assign n176 = n175 ^ n172 ;
  assign n183 = n179 ^ n176 ;
  assign n203 = n202 ^ n183 ;
  assign n211 = n197 ^ n195 ;
  assign n212 = n196 & ~n211 ;
  assign n213 = n212 ^ n194 ;
  assign n207 = n198 ^ n191 ;
  assign n208 = ~n193 & n207 ;
  assign n209 = n208 ^ n198 ;
  assign n204 = n190 ^ n188 ;
  assign n205 = n189 & ~n204 ;
  assign n206 = n205 ^ n187 ;
  assign n210 = n209 ^ n206 ;
  assign n214 = n213 ^ n210 ;
  assign n215 = n214 ^ n183 ;
  assign n216 = n203 & ~n215 ;
  assign n217 = n216 ^ n202 ;
  assign n180 = n179 ^ n175 ;
  assign n181 = n176 & ~n180 ;
  assign n182 = n181 ^ n172 ;
  assign n218 = n217 ^ n182 ;
  assign n219 = n213 ^ n206 ;
  assign n220 = ~n210 & n219 ;
  assign n221 = n220 ^ n213 ;
  assign n222 = n221 ^ n182 ;
  assign n223 = n218 & n222 ;
  assign n224 = n223 ^ n182 ;
  assign n225 = n221 ^ n218 ;
  assign n226 = n214 ^ n203 ;
  assign n228 = n199 ^ n186 ;
  assign n229 = n227 & n228 ;
  assign n230 = n226 & n229 ;
  assign n231 = n225 & n230 ;
  assign n233 = ~n224 & ~n231 ;
  assign n232 = n231 ^ n224 ;
  assign n234 = n233 ^ n232 ;
  assign n235 = n157 & n234 ;
  assign n240 = n239 ^ n237 ;
  assign n256 = n242 ^ n240 ;
  assign n259 = n258 ^ n256 ;
  assign n250 = n249 ^ n247 ;
  assign n260 = n252 ^ n250 ;
  assign n261 = n260 ^ n256 ;
  assign n262 = n259 & ~n261 ;
  assign n263 = n262 ^ n258 ;
  assign n253 = n252 ^ n247 ;
  assign n254 = n250 & ~n253 ;
  assign n255 = n254 ^ n249 ;
  assign n264 = n263 ^ n255 ;
  assign n243 = n242 ^ n237 ;
  assign n244 = ~n240 & n243 ;
  assign n245 = n244 ^ n242 ;
  assign n310 = n255 ^ n245 ;
  assign n311 = ~n264 & n310 ;
  assign n312 = n311 ^ n245 ;
  assign n266 = n260 ^ n258 ;
  assign n267 = n266 ^ n256 ;
  assign n270 = n269 ^ n267 ;
  assign n283 = n282 ^ n280 ;
  assign n286 = n285 ^ n283 ;
  assign n289 = n288 ^ n286 ;
  assign n275 = n274 ^ n272 ;
  assign n278 = n277 ^ n275 ;
  assign n290 = n289 ^ n278 ;
  assign n291 = n290 ^ n267 ;
  assign n292 = n270 & ~n291 ;
  assign n293 = n292 ^ n269 ;
  assign n265 = n264 ^ n245 ;
  assign n294 = n293 ^ n265 ;
  assign n303 = n277 ^ n272 ;
  assign n304 = ~n275 & n303 ;
  assign n305 = n304 ^ n277 ;
  assign n298 = n288 ^ n278 ;
  assign n299 = n286 ^ n278 ;
  assign n300 = n298 & ~n299 ;
  assign n301 = n300 ^ n288 ;
  assign n295 = n285 ^ n280 ;
  assign n296 = ~n283 & n295 ;
  assign n297 = n296 ^ n285 ;
  assign n302 = n301 ^ n297 ;
  assign n306 = n305 ^ n302 ;
  assign n307 = n306 ^ n293 ;
  assign n308 = n294 & ~n307 ;
  assign n309 = n308 ^ n265 ;
  assign n313 = n312 ^ n309 ;
  assign n314 = n305 ^ n301 ;
  assign n315 = n302 & ~n314 ;
  assign n316 = n315 ^ n297 ;
  assign n317 = n316 ^ n312 ;
  assign n318 = n313 & ~n317 ;
  assign n319 = n318 ^ n309 ;
  assign n320 = n316 ^ n313 ;
  assign n323 = n290 ^ n270 ;
  assign n324 = n322 & n323 ;
  assign n325 = n306 ^ n294 ;
  assign n326 = n324 & n325 ;
  assign n327 = n320 & n326 ;
  assign n329 = ~n319 & ~n327 ;
  assign n328 = n327 ^ n319 ;
  assign n330 = n329 ^ n328 ;
  assign n346 = n345 ^ n343 ;
  assign n349 = n348 ^ n346 ;
  assign n365 = n349 ^ n340 ;
  assign n335 = n334 ^ n332 ;
  assign n338 = n337 ^ n335 ;
  assign n366 = n365 ^ n338 ;
  assign n369 = n368 ^ n366 ;
  assign n382 = n381 ^ n379 ;
  assign n385 = n384 ^ n382 ;
  assign n388 = n387 ^ n385 ;
  assign n374 = n373 ^ n371 ;
  assign n377 = n376 ^ n374 ;
  assign n389 = n388 ^ n377 ;
  assign n390 = n389 ^ n366 ;
  assign n391 = n369 & ~n390 ;
  assign n392 = n391 ^ n368 ;
  assign n357 = n337 ^ n334 ;
  assign n358 = n337 ^ n332 ;
  assign n359 = ~n357 & n358 ;
  assign n360 = n359 ^ n332 ;
  assign n353 = n348 ^ n343 ;
  assign n354 = n346 & ~n353 ;
  assign n355 = n354 ^ n345 ;
  assign n341 = n340 ^ n338 ;
  assign n350 = n349 ^ n338 ;
  assign n351 = n341 & ~n350 ;
  assign n352 = n351 ^ n340 ;
  assign n356 = n355 ^ n352 ;
  assign n364 = n360 ^ n356 ;
  assign n393 = n392 ^ n364 ;
  assign n402 = n376 ^ n373 ;
  assign n403 = n374 & ~n402 ;
  assign n404 = n403 ^ n371 ;
  assign n397 = n387 ^ n377 ;
  assign n398 = n385 ^ n377 ;
  assign n399 = n397 & ~n398 ;
  assign n400 = n399 ^ n387 ;
  assign n394 = n384 ^ n381 ;
  assign n395 = n382 & ~n394 ;
  assign n396 = n395 ^ n379 ;
  assign n401 = n400 ^ n396 ;
  assign n405 = n404 ^ n401 ;
  assign n406 = n405 ^ n364 ;
  assign n407 = n393 & ~n406 ;
  assign n408 = n407 ^ n392 ;
  assign n361 = n360 ^ n355 ;
  assign n362 = n356 & ~n361 ;
  assign n363 = n362 ^ n352 ;
  assign n409 = n408 ^ n363 ;
  assign n410 = n404 ^ n396 ;
  assign n411 = ~n401 & n410 ;
  assign n412 = n411 ^ n404 ;
  assign n413 = n412 ^ n363 ;
  assign n414 = n409 & n413 ;
  assign n415 = n414 ^ n363 ;
  assign n416 = n412 ^ n409 ;
  assign n417 = n405 ^ n393 ;
  assign n420 = n389 ^ n369 ;
  assign n421 = n419 & n420 ;
  assign n422 = n417 & n421 ;
  assign n423 = n416 & n422 ;
  assign n425 = ~n415 & ~n423 ;
  assign n424 = n423 ^ n415 ;
  assign n426 = n425 ^ n424 ;
  assign n427 = n330 & n426 ;
  assign n428 = n235 & ~n427 ;
  assign n429 = n428 ^ n235 ;
  assign n742 = n741 ^ n429 ;
  assign n827 = n329 & n425 ;
  assign n828 = n827 ^ n427 ;
  assign n829 = n156 & n233 ;
  assign n830 = ~n828 & ~n829 ;
  assign n831 = n830 ^ n427 ;
  assign n832 = n235 & n831 ;
  assign n833 = n832 ^ n427 ;
  assign n834 = n828 ^ n428 ;
  assign n835 = n834 ^ n829 ;
  assign n836 = n835 ^ n832 ;
  assign n863 = n326 ^ n320 ;
  assign n862 = n422 ^ n416 ;
  assign n864 = n863 ^ n862 ;
  assign n865 = n426 ^ n330 ;
  assign n866 = n424 ^ n328 ;
  assign n868 = n323 ^ n322 ;
  assign n869 = n420 ^ n419 ;
  assign n870 = ~n868 & n869 ;
  assign n867 = n325 ^ n324 ;
  assign n871 = n870 ^ n867 ;
  assign n872 = n421 ^ n417 ;
  assign n873 = n872 ^ n870 ;
  assign n874 = ~n871 & ~n873 ;
  assign n875 = n874 ^ n867 ;
  assign n876 = n875 ^ n862 ;
  assign n877 = ~n864 & n876 ;
  assign n878 = n877 ^ n863 ;
  assign n879 = n878 ^ n328 ;
  assign n880 = ~n866 & ~n879 ;
  assign n881 = n880 ^ n424 ;
  assign n882 = n881 ^ n330 ;
  assign n883 = ~n865 & ~n882 ;
  assign n884 = n883 ^ n426 ;
  assign n885 = n864 & ~n884 ;
  assign n886 = n885 ^ n863 ;
  assign n838 = n230 ^ n225 ;
  assign n837 = n153 ^ n146 ;
  assign n839 = n838 ^ n837 ;
  assign n840 = n234 ^ n157 ;
  assign n841 = n232 ^ n155 ;
  assign n843 = n229 ^ n226 ;
  assign n842 = n152 ^ n151 ;
  assign n844 = n843 ^ n842 ;
  assign n845 = n228 ^ n227 ;
  assign n846 = n150 ^ n149 ;
  assign n847 = ~n845 & n846 ;
  assign n848 = n847 ^ n842 ;
  assign n849 = ~n844 & ~n848 ;
  assign n850 = n849 ^ n843 ;
  assign n851 = n850 ^ n838 ;
  assign n852 = ~n839 & n851 ;
  assign n853 = n852 ^ n838 ;
  assign n854 = n853 ^ n232 ;
  assign n855 = ~n841 & ~n854 ;
  assign n856 = n855 ^ n155 ;
  assign n857 = n856 ^ n234 ;
  assign n858 = ~n840 & ~n857 ;
  assign n859 = n858 ^ n157 ;
  assign n860 = n839 & ~n859 ;
  assign n861 = n860 ^ n838 ;
  assign n887 = n886 ^ n861 ;
  assign n890 = n872 ^ n867 ;
  assign n891 = n884 & n890 ;
  assign n892 = n891 ^ n872 ;
  assign n888 = n844 & ~n859 ;
  assign n889 = n888 ^ n843 ;
  assign n893 = n892 ^ n889 ;
  assign n894 = n846 ^ n845 ;
  assign n895 = ~n859 & n894 ;
  assign n896 = n895 ^ n845 ;
  assign n897 = n869 ^ n868 ;
  assign n898 = ~n884 & n897 ;
  assign n899 = n898 ^ n868 ;
  assign n900 = ~n896 & n899 ;
  assign n901 = n900 ^ n892 ;
  assign n902 = ~n893 & n901 ;
  assign n903 = n902 ^ n892 ;
  assign n904 = n903 ^ n886 ;
  assign n905 = ~n887 & n904 ;
  assign n906 = n905 ^ n886 ;
  assign n907 = ~n836 & ~n906 ;
  assign n908 = ~n833 & ~n907 ;
  assign n909 = n829 ^ n235 ;
  assign n910 = n909 ^ n828 ;
  assign n911 = n910 ^ n828 ;
  assign n912 = ~n428 & n911 ;
  assign n913 = n912 ^ n828 ;
  assign n914 = ~n908 & n913 ;
  assign n915 = n914 ^ n828 ;
  assign n745 = n660 & n737 ;
  assign n746 = n745 ^ n739 ;
  assign n743 = n505 & n582 ;
  assign n744 = n743 ^ n584 ;
  assign n747 = n746 ^ n744 ;
  assign n773 = n738 ^ n661 ;
  assign n774 = n736 ^ n659 ;
  assign n784 = n657 ^ n656 ;
  assign n776 = n655 ^ n652 ;
  assign n775 = n732 ^ n731 ;
  assign n777 = n776 ^ n775 ;
  assign n778 = n730 ^ n729 ;
  assign n779 = n654 ^ n653 ;
  assign n780 = ~n778 & n779 ;
  assign n781 = n780 ^ n776 ;
  assign n782 = ~n777 & ~n781 ;
  assign n783 = n782 ^ n780 ;
  assign n785 = n784 ^ n783 ;
  assign n786 = n734 ^ n733 ;
  assign n787 = n786 ^ n783 ;
  assign n788 = ~n785 & n787 ;
  assign n789 = n788 ^ n784 ;
  assign n790 = n789 ^ n659 ;
  assign n791 = n774 & ~n790 ;
  assign n792 = n791 ^ n736 ;
  assign n793 = n792 ^ n738 ;
  assign n794 = n773 & n793 ;
  assign n795 = n794 ^ n661 ;
  assign n796 = n786 ^ n784 ;
  assign n797 = ~n795 & ~n796 ;
  assign n798 = n797 ^ n784 ;
  assign n749 = n579 ^ n578 ;
  assign n748 = n502 ^ n501 ;
  assign n750 = n749 ^ n748 ;
  assign n751 = n583 ^ n506 ;
  assign n752 = n581 ^ n504 ;
  assign n754 = n500 ^ n499 ;
  assign n753 = n577 ^ n576 ;
  assign n755 = n754 ^ n753 ;
  assign n756 = n575 ^ n574 ;
  assign n757 = n498 ^ n497 ;
  assign n758 = ~n756 & n757 ;
  assign n759 = n758 ^ n754 ;
  assign n760 = n755 & n759 ;
  assign n761 = n760 ^ n758 ;
  assign n762 = n761 ^ n748 ;
  assign n763 = ~n750 & ~n762 ;
  assign n764 = n763 ^ n749 ;
  assign n765 = n764 ^ n581 ;
  assign n766 = ~n752 & ~n765 ;
  assign n767 = n766 ^ n504 ;
  assign n768 = n767 ^ n583 ;
  assign n769 = ~n751 & ~n768 ;
  assign n770 = n769 ^ n506 ;
  assign n771 = n750 & ~n770 ;
  assign n772 = n771 ^ n749 ;
  assign n799 = n798 ^ n772 ;
  assign n802 = n757 ^ n756 ;
  assign n803 = ~n770 & n802 ;
  assign n804 = n803 ^ n756 ;
  assign n805 = n779 ^ n778 ;
  assign n806 = n795 & n805 ;
  assign n807 = n806 ^ n778 ;
  assign n808 = ~n804 & n807 ;
  assign n800 = n755 & n770 ;
  assign n801 = n800 ^ n754 ;
  assign n809 = n808 ^ n801 ;
  assign n810 = ~n777 & ~n795 ;
  assign n811 = n810 ^ n776 ;
  assign n812 = n811 ^ n808 ;
  assign n813 = ~n809 & ~n812 ;
  assign n814 = n813 ^ n808 ;
  assign n815 = n814 ^ n798 ;
  assign n816 = n799 & n815 ;
  assign n817 = n816 ^ n772 ;
  assign n818 = n817 ^ n746 ;
  assign n819 = ~n747 & ~n818 ;
  assign n820 = n819 ^ n746 ;
  assign n821 = n741 ^ n739 ;
  assign n822 = n820 & ~n821 ;
  assign n823 = ~n740 & n744 ;
  assign n824 = n823 ^ n746 ;
  assign n825 = ~n822 & n824 ;
  assign n826 = n825 ^ n746 ;
  assign n916 = n915 ^ n826 ;
  assign n920 = ~n740 & ~n822 ;
  assign n921 = ~n799 & ~n920 ;
  assign n922 = n921 ^ n772 ;
  assign n917 = ~n428 & ~n908 ;
  assign n918 = n887 & n917 ;
  assign n919 = n918 ^ n886 ;
  assign n923 = n922 ^ n919 ;
  assign n926 = n811 ^ n801 ;
  assign n927 = n920 & ~n926 ;
  assign n928 = n927 ^ n811 ;
  assign n924 = n893 & n917 ;
  assign n925 = n924 ^ n892 ;
  assign n929 = n928 ^ n925 ;
  assign n930 = n899 ^ n896 ;
  assign n931 = ~n917 & n930 ;
  assign n932 = n931 ^ n896 ;
  assign n933 = n807 ^ n804 ;
  assign n934 = ~n920 & n933 ;
  assign n935 = n934 ^ n804 ;
  assign n936 = ~n932 & n935 ;
  assign n937 = n936 ^ n925 ;
  assign n938 = n929 & ~n937 ;
  assign n939 = n938 ^ n925 ;
  assign n940 = n939 ^ n919 ;
  assign n941 = ~n923 & n940 ;
  assign n942 = n941 ^ n919 ;
  assign n943 = n942 ^ n826 ;
  assign n944 = ~n916 & n943 ;
  assign n945 = n944 ^ n915 ;
  assign n946 = n945 ^ n429 ;
  assign n947 = ~n742 & n946 ;
  assign n948 = n947 ^ n741 ;
  assign n952 = n884 ^ n859 ;
  assign n953 = ~n917 & n952 ;
  assign n954 = n953 ^ n859 ;
  assign n949 = n795 ^ n770 ;
  assign n950 = ~n920 & ~n949 ;
  assign n951 = n950 ^ n770 ;
  assign n955 = n954 ^ n951 ;
  assign n956 = n948 & n955 ;
  assign n957 = n956 ^ n951 ;
  assign n958 = n920 ^ n917 ;
  assign n959 = ~n948 & n958 ;
  assign n960 = n959 ^ n917 ;
  assign y0 = n957 ;
  assign y1 = n960 ;
  assign y2 = n948 ;
endmodule
