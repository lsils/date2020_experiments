module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 ;
  assign n3180 = x526 ^ x14 ;
  assign n3179 = x527 ^ x15 ;
  assign n3181 = n3180 ^ n3179 ;
  assign n3178 = x528 ^ x16 ;
  assign n3209 = n3180 ^ n3178 ;
  assign n3210 = n3181 & ~n3209 ;
  assign n3211 = n3210 ^ n3179 ;
  assign n3183 = x522 ^ x10 ;
  assign n3182 = n3181 ^ n3178 ;
  assign n3184 = n3183 ^ n3182 ;
  assign n3176 = x525 ^ x13 ;
  assign n3174 = x523 ^ x11 ;
  assign n3173 = x524 ^ x12 ;
  assign n3175 = n3174 ^ n3173 ;
  assign n3177 = n3176 ^ n3175 ;
  assign n3206 = n3183 ^ n3177 ;
  assign n3207 = n3184 & ~n3206 ;
  assign n3208 = n3207 ^ n3182 ;
  assign n3212 = n3211 ^ n3208 ;
  assign n3203 = n3176 ^ n3174 ;
  assign n3204 = n3175 & ~n3203 ;
  assign n3205 = n3204 ^ n3173 ;
  assign n3229 = n3211 ^ n3205 ;
  assign n3230 = n3212 & ~n3229 ;
  assign n3231 = n3230 ^ n3208 ;
  assign n3185 = n3184 ^ n3177 ;
  assign n3172 = x514 ^ x2 ;
  assign n3186 = n3185 ^ n3172 ;
  assign n3169 = x515 ^ x3 ;
  assign n3167 = x521 ^ x9 ;
  assign n3165 = x519 ^ x7 ;
  assign n3164 = x520 ^ x8 ;
  assign n3166 = n3165 ^ n3164 ;
  assign n3168 = n3167 ^ n3166 ;
  assign n3170 = n3169 ^ n3168 ;
  assign n3162 = x518 ^ x6 ;
  assign n3160 = x516 ^ x4 ;
  assign n3159 = x517 ^ x5 ;
  assign n3161 = n3160 ^ n3159 ;
  assign n3163 = n3162 ^ n3161 ;
  assign n3171 = n3170 ^ n3163 ;
  assign n3214 = n3185 ^ n3171 ;
  assign n3215 = n3186 & ~n3214 ;
  assign n3216 = n3215 ^ n3172 ;
  assign n3213 = n3212 ^ n3205 ;
  assign n3217 = n3216 ^ n3213 ;
  assign n3199 = n3162 ^ n3160 ;
  assign n3200 = n3161 & ~n3199 ;
  assign n3201 = n3200 ^ n3159 ;
  assign n3195 = n3168 ^ n3163 ;
  assign n3196 = ~n3170 & n3195 ;
  assign n3197 = n3196 ^ n3163 ;
  assign n3192 = n3167 ^ n3165 ;
  assign n3193 = n3166 & ~n3192 ;
  assign n3194 = n3193 ^ n3164 ;
  assign n3198 = n3197 ^ n3194 ;
  assign n3202 = n3201 ^ n3198 ;
  assign n3226 = n3213 ^ n3202 ;
  assign n3227 = n3217 & ~n3226 ;
  assign n3228 = n3227 ^ n3216 ;
  assign n3232 = n3231 ^ n3228 ;
  assign n3223 = n3201 ^ n3197 ;
  assign n3224 = n3198 & ~n3223 ;
  assign n3225 = n3224 ^ n3194 ;
  assign n3238 = n3231 ^ n3225 ;
  assign n3239 = n3232 & ~n3238 ;
  assign n3240 = n3239 ^ n3228 ;
  assign n3157 = x513 ^ x1 ;
  assign n3126 = x533 ^ x21 ;
  assign n3124 = x531 ^ x19 ;
  assign n3123 = x532 ^ x20 ;
  assign n3125 = n3124 ^ n3123 ;
  assign n3127 = n3126 ^ n3125 ;
  assign n3121 = x530 ^ x18 ;
  assign n3119 = x536 ^ x24 ;
  assign n3117 = x534 ^ x22 ;
  assign n3116 = x535 ^ x23 ;
  assign n3118 = n3117 ^ n3116 ;
  assign n3120 = n3119 ^ n3118 ;
  assign n3122 = n3121 ^ n3120 ;
  assign n3128 = n3127 ^ n3122 ;
  assign n3114 = x529 ^ x17 ;
  assign n3100 = x540 ^ x28 ;
  assign n3098 = x538 ^ x26 ;
  assign n3097 = x539 ^ x27 ;
  assign n3099 = n3098 ^ n3097 ;
  assign n3101 = n3100 ^ n3099 ;
  assign n3090 = x543 ^ x31 ;
  assign n3088 = x542 ^ x30 ;
  assign n3087 = x541 ^ x29 ;
  assign n3089 = n3088 ^ n3087 ;
  assign n3095 = n3090 ^ n3089 ;
  assign n3094 = x537 ^ x25 ;
  assign n3096 = n3095 ^ n3094 ;
  assign n3113 = n3101 ^ n3096 ;
  assign n3115 = n3114 ^ n3113 ;
  assign n3156 = n3128 ^ n3115 ;
  assign n3158 = n3157 ^ n3156 ;
  assign n3187 = n3186 ^ n3171 ;
  assign n3188 = n3187 ^ n3157 ;
  assign n3189 = n3158 & ~n3188 ;
  assign n3190 = n3189 ^ n3156 ;
  assign n3140 = n3126 ^ n3124 ;
  assign n3141 = n3125 & ~n3140 ;
  assign n3142 = n3141 ^ n3123 ;
  assign n3136 = n3119 ^ n3117 ;
  assign n3137 = n3118 & ~n3136 ;
  assign n3138 = n3137 ^ n3116 ;
  assign n3133 = n3127 ^ n3121 ;
  assign n3134 = n3122 & ~n3133 ;
  assign n3135 = n3134 ^ n3120 ;
  assign n3139 = n3138 ^ n3135 ;
  assign n3143 = n3142 ^ n3139 ;
  assign n3129 = n3128 ^ n3114 ;
  assign n3130 = n3115 & ~n3129 ;
  assign n3131 = n3130 ^ n3113 ;
  assign n3106 = n3100 ^ n3098 ;
  assign n3107 = n3099 & ~n3106 ;
  assign n3108 = n3107 ^ n3097 ;
  assign n3102 = n3101 ^ n3095 ;
  assign n3103 = n3096 & ~n3102 ;
  assign n3104 = n3103 ^ n3094 ;
  assign n3091 = n3090 ^ n3088 ;
  assign n3092 = n3089 & ~n3091 ;
  assign n3093 = n3092 ^ n3087 ;
  assign n3105 = n3104 ^ n3093 ;
  assign n3112 = n3108 ^ n3105 ;
  assign n3132 = n3131 ^ n3112 ;
  assign n3155 = n3143 ^ n3132 ;
  assign n3191 = n3190 ^ n3155 ;
  assign n3218 = n3217 ^ n3202 ;
  assign n3219 = n3218 ^ n3155 ;
  assign n3220 = n3191 & ~n3219 ;
  assign n3221 = n3220 ^ n3190 ;
  assign n3148 = n3142 ^ n3138 ;
  assign n3149 = n3139 & ~n3148 ;
  assign n3150 = n3149 ^ n3135 ;
  assign n3144 = n3143 ^ n3112 ;
  assign n3145 = n3132 & ~n3144 ;
  assign n3146 = n3145 ^ n3131 ;
  assign n3109 = n3108 ^ n3104 ;
  assign n3110 = n3105 & ~n3109 ;
  assign n3111 = n3110 ^ n3093 ;
  assign n3147 = n3146 ^ n3111 ;
  assign n3154 = n3150 ^ n3147 ;
  assign n3222 = n3221 ^ n3154 ;
  assign n3233 = n3232 ^ n3225 ;
  assign n3234 = n3233 ^ n3221 ;
  assign n3235 = n3222 & ~n3234 ;
  assign n3236 = n3235 ^ n3154 ;
  assign n3151 = n3150 ^ n3146 ;
  assign n3152 = n3147 & ~n3151 ;
  assign n3153 = n3152 ^ n3111 ;
  assign n3237 = n3236 ^ n3153 ;
  assign n3241 = n3240 ^ n3237 ;
  assign n3242 = n3218 ^ n3191 ;
  assign n3243 = n3187 ^ n3158 ;
  assign n3244 = x512 ^ x0 ;
  assign n3245 = n3243 & n3244 ;
  assign n3246 = n3242 & n3245 ;
  assign n3247 = n3233 ^ n3222 ;
  assign n3248 = n3246 & n3247 ;
  assign n3249 = n3241 & n3248 ;
  assign n3250 = n3240 ^ n3153 ;
  assign n3251 = ~n3237 & n3250 ;
  assign n3252 = n3251 ^ n3240 ;
  assign n3253 = n3249 & n3252 ;
  assign n643 = x514 ^ x34 ;
  assign n640 = x522 ^ x42 ;
  assign n638 = x528 ^ x48 ;
  assign n636 = x526 ^ x46 ;
  assign n635 = x527 ^ x47 ;
  assign n637 = n636 ^ n635 ;
  assign n639 = n638 ^ n637 ;
  assign n641 = n640 ^ n639 ;
  assign n633 = x525 ^ x45 ;
  assign n631 = x523 ^ x43 ;
  assign n630 = x524 ^ x44 ;
  assign n632 = n631 ^ n630 ;
  assign n634 = n633 ^ n632 ;
  assign n642 = n641 ^ n634 ;
  assign n644 = n643 ^ n642 ;
  assign n627 = x515 ^ x35 ;
  assign n625 = x521 ^ x41 ;
  assign n623 = x519 ^ x39 ;
  assign n622 = x520 ^ x40 ;
  assign n624 = n623 ^ n622 ;
  assign n626 = n625 ^ n624 ;
  assign n628 = n627 ^ n626 ;
  assign n620 = x518 ^ x38 ;
  assign n618 = x516 ^ x36 ;
  assign n617 = x517 ^ x37 ;
  assign n619 = n618 ^ n617 ;
  assign n621 = n620 ^ n619 ;
  assign n629 = n628 ^ n621 ;
  assign n672 = n643 ^ n629 ;
  assign n673 = n644 & ~n672 ;
  assign n674 = n673 ^ n642 ;
  assign n668 = n633 ^ n631 ;
  assign n669 = n632 & ~n668 ;
  assign n670 = n669 ^ n630 ;
  assign n664 = n638 ^ n636 ;
  assign n665 = n637 & ~n664 ;
  assign n666 = n665 ^ n635 ;
  assign n661 = n639 ^ n634 ;
  assign n662 = ~n641 & n661 ;
  assign n663 = n662 ^ n634 ;
  assign n667 = n666 ^ n663 ;
  assign n671 = n670 ^ n667 ;
  assign n675 = n674 ^ n671 ;
  assign n657 = n620 ^ n618 ;
  assign n658 = n619 & ~n657 ;
  assign n659 = n658 ^ n617 ;
  assign n653 = n626 ^ n621 ;
  assign n654 = ~n628 & n653 ;
  assign n655 = n654 ^ n621 ;
  assign n650 = n625 ^ n623 ;
  assign n651 = n624 & ~n650 ;
  assign n652 = n651 ^ n622 ;
  assign n656 = n655 ^ n652 ;
  assign n660 = n659 ^ n656 ;
  assign n687 = n674 ^ n660 ;
  assign n688 = n675 & ~n687 ;
  assign n689 = n688 ^ n671 ;
  assign n684 = n670 ^ n666 ;
  assign n685 = n667 & ~n684 ;
  assign n686 = n685 ^ n663 ;
  assign n690 = n689 ^ n686 ;
  assign n681 = n659 ^ n655 ;
  assign n682 = n656 & ~n681 ;
  assign n683 = n682 ^ n652 ;
  assign n696 = n686 ^ n683 ;
  assign n697 = ~n690 & n696 ;
  assign n698 = n697 ^ n683 ;
  assign n615 = x513 ^ x33 ;
  assign n581 = x533 ^ x53 ;
  assign n579 = x531 ^ x51 ;
  assign n578 = x532 ^ x52 ;
  assign n580 = n579 ^ n578 ;
  assign n582 = n581 ^ n580 ;
  assign n576 = x530 ^ x50 ;
  assign n574 = x536 ^ x56 ;
  assign n572 = x534 ^ x54 ;
  assign n571 = x535 ^ x55 ;
  assign n573 = n572 ^ n571 ;
  assign n575 = n574 ^ n573 ;
  assign n577 = n576 ^ n575 ;
  assign n583 = n582 ^ n577 ;
  assign n554 = x538 ^ x58 ;
  assign n553 = x539 ^ x59 ;
  assign n555 = n554 ^ n553 ;
  assign n552 = x540 ^ x60 ;
  assign n556 = n555 ^ n552 ;
  assign n550 = x537 ^ x57 ;
  assign n547 = x541 ^ x61 ;
  assign n546 = x542 ^ x62 ;
  assign n548 = n547 ^ n546 ;
  assign n545 = x543 ^ x63 ;
  assign n549 = n548 ^ n545 ;
  assign n551 = n550 ^ n549 ;
  assign n569 = n556 ^ n551 ;
  assign n568 = x529 ^ x49 ;
  assign n570 = n569 ^ n568 ;
  assign n614 = n583 ^ n570 ;
  assign n616 = n615 ^ n614 ;
  assign n645 = n644 ^ n629 ;
  assign n646 = n645 ^ n615 ;
  assign n647 = n616 & ~n646 ;
  assign n648 = n647 ^ n614 ;
  assign n595 = n581 ^ n579 ;
  assign n596 = n580 & ~n595 ;
  assign n597 = n596 ^ n578 ;
  assign n591 = n574 ^ n572 ;
  assign n592 = n573 & ~n591 ;
  assign n593 = n592 ^ n571 ;
  assign n588 = n582 ^ n576 ;
  assign n589 = n577 & ~n588 ;
  assign n590 = n589 ^ n575 ;
  assign n594 = n593 ^ n590 ;
  assign n598 = n597 ^ n594 ;
  assign n584 = n583 ^ n569 ;
  assign n585 = n570 & ~n584 ;
  assign n586 = n585 ^ n568 ;
  assign n564 = n553 ^ n552 ;
  assign n565 = ~n555 & n564 ;
  assign n566 = n565 ^ n552 ;
  assign n560 = n546 ^ n545 ;
  assign n561 = ~n548 & n560 ;
  assign n562 = n561 ^ n545 ;
  assign n557 = n556 ^ n550 ;
  assign n558 = n551 & ~n557 ;
  assign n559 = n558 ^ n549 ;
  assign n563 = n562 ^ n559 ;
  assign n567 = n566 ^ n563 ;
  assign n587 = n586 ^ n567 ;
  assign n613 = n598 ^ n587 ;
  assign n649 = n648 ^ n613 ;
  assign n676 = n675 ^ n660 ;
  assign n677 = n676 ^ n613 ;
  assign n678 = n649 & ~n677 ;
  assign n679 = n678 ^ n648 ;
  assign n606 = n597 ^ n593 ;
  assign n607 = n594 & ~n606 ;
  assign n608 = n607 ^ n590 ;
  assign n602 = n566 ^ n562 ;
  assign n603 = n563 & ~n602 ;
  assign n604 = n603 ^ n559 ;
  assign n599 = n598 ^ n586 ;
  assign n600 = n587 & ~n599 ;
  assign n601 = n600 ^ n567 ;
  assign n605 = n604 ^ n601 ;
  assign n612 = n608 ^ n605 ;
  assign n680 = n679 ^ n612 ;
  assign n691 = n690 ^ n683 ;
  assign n692 = n691 ^ n679 ;
  assign n693 = n680 & ~n692 ;
  assign n694 = n693 ^ n612 ;
  assign n609 = n608 ^ n604 ;
  assign n610 = n605 & ~n609 ;
  assign n611 = n610 ^ n601 ;
  assign n695 = n694 ^ n611 ;
  assign n699 = n698 ^ n695 ;
  assign n700 = n645 ^ n616 ;
  assign n701 = x512 ^ x32 ;
  assign n702 = n700 & n701 ;
  assign n703 = n676 ^ n649 ;
  assign n704 = n702 & n703 ;
  assign n705 = n691 ^ n680 ;
  assign n706 = n704 & n705 ;
  assign n707 = n699 & n706 ;
  assign n708 = n698 ^ n694 ;
  assign n709 = n695 & ~n708 ;
  assign n710 = n709 ^ n611 ;
  assign n711 = n707 & n710 ;
  assign n810 = x514 ^ x66 ;
  assign n807 = x522 ^ x74 ;
  assign n805 = x528 ^ x80 ;
  assign n803 = x526 ^ x78 ;
  assign n802 = x527 ^ x79 ;
  assign n804 = n803 ^ n802 ;
  assign n806 = n805 ^ n804 ;
  assign n808 = n807 ^ n806 ;
  assign n800 = x525 ^ x77 ;
  assign n798 = x523 ^ x75 ;
  assign n797 = x524 ^ x76 ;
  assign n799 = n798 ^ n797 ;
  assign n801 = n800 ^ n799 ;
  assign n809 = n808 ^ n801 ;
  assign n811 = n810 ^ n809 ;
  assign n794 = x515 ^ x67 ;
  assign n792 = x521 ^ x73 ;
  assign n790 = x519 ^ x71 ;
  assign n789 = x520 ^ x72 ;
  assign n791 = n790 ^ n789 ;
  assign n793 = n792 ^ n791 ;
  assign n795 = n794 ^ n793 ;
  assign n787 = x518 ^ x70 ;
  assign n785 = x516 ^ x68 ;
  assign n784 = x517 ^ x69 ;
  assign n786 = n785 ^ n784 ;
  assign n788 = n787 ^ n786 ;
  assign n796 = n795 ^ n788 ;
  assign n839 = n810 ^ n796 ;
  assign n840 = n811 & ~n839 ;
  assign n841 = n840 ^ n809 ;
  assign n835 = n800 ^ n798 ;
  assign n836 = n799 & ~n835 ;
  assign n837 = n836 ^ n797 ;
  assign n831 = n805 ^ n803 ;
  assign n832 = n804 & ~n831 ;
  assign n833 = n832 ^ n802 ;
  assign n828 = n806 ^ n801 ;
  assign n829 = ~n808 & n828 ;
  assign n830 = n829 ^ n801 ;
  assign n834 = n833 ^ n830 ;
  assign n838 = n837 ^ n834 ;
  assign n842 = n841 ^ n838 ;
  assign n824 = n787 ^ n785 ;
  assign n825 = n786 & ~n824 ;
  assign n826 = n825 ^ n784 ;
  assign n820 = n793 ^ n788 ;
  assign n821 = ~n795 & n820 ;
  assign n822 = n821 ^ n788 ;
  assign n817 = n792 ^ n790 ;
  assign n818 = n791 & ~n817 ;
  assign n819 = n818 ^ n789 ;
  assign n823 = n822 ^ n819 ;
  assign n827 = n826 ^ n823 ;
  assign n854 = n841 ^ n827 ;
  assign n855 = n842 & ~n854 ;
  assign n856 = n855 ^ n838 ;
  assign n851 = n837 ^ n833 ;
  assign n852 = n834 & ~n851 ;
  assign n853 = n852 ^ n830 ;
  assign n857 = n856 ^ n853 ;
  assign n848 = n826 ^ n822 ;
  assign n849 = n823 & ~n848 ;
  assign n850 = n849 ^ n819 ;
  assign n863 = n853 ^ n850 ;
  assign n864 = ~n857 & n863 ;
  assign n865 = n864 ^ n850 ;
  assign n782 = x513 ^ x65 ;
  assign n748 = x533 ^ x85 ;
  assign n746 = x531 ^ x83 ;
  assign n745 = x532 ^ x84 ;
  assign n747 = n746 ^ n745 ;
  assign n749 = n748 ^ n747 ;
  assign n743 = x530 ^ x82 ;
  assign n741 = x536 ^ x88 ;
  assign n739 = x534 ^ x86 ;
  assign n738 = x535 ^ x87 ;
  assign n740 = n739 ^ n738 ;
  assign n742 = n741 ^ n740 ;
  assign n744 = n743 ^ n742 ;
  assign n750 = n749 ^ n744 ;
  assign n721 = x538 ^ x90 ;
  assign n720 = x539 ^ x91 ;
  assign n722 = n721 ^ n720 ;
  assign n719 = x540 ^ x92 ;
  assign n723 = n722 ^ n719 ;
  assign n717 = x537 ^ x89 ;
  assign n714 = x541 ^ x93 ;
  assign n713 = x542 ^ x94 ;
  assign n715 = n714 ^ n713 ;
  assign n712 = x543 ^ x95 ;
  assign n716 = n715 ^ n712 ;
  assign n718 = n717 ^ n716 ;
  assign n736 = n723 ^ n718 ;
  assign n735 = x529 ^ x81 ;
  assign n737 = n736 ^ n735 ;
  assign n781 = n750 ^ n737 ;
  assign n783 = n782 ^ n781 ;
  assign n812 = n811 ^ n796 ;
  assign n813 = n812 ^ n782 ;
  assign n814 = n783 & ~n813 ;
  assign n815 = n814 ^ n781 ;
  assign n762 = n748 ^ n746 ;
  assign n763 = n747 & ~n762 ;
  assign n764 = n763 ^ n745 ;
  assign n758 = n741 ^ n739 ;
  assign n759 = n740 & ~n758 ;
  assign n760 = n759 ^ n738 ;
  assign n755 = n749 ^ n743 ;
  assign n756 = n744 & ~n755 ;
  assign n757 = n756 ^ n742 ;
  assign n761 = n760 ^ n757 ;
  assign n765 = n764 ^ n761 ;
  assign n751 = n750 ^ n736 ;
  assign n752 = n737 & ~n751 ;
  assign n753 = n752 ^ n735 ;
  assign n731 = n720 ^ n719 ;
  assign n732 = ~n722 & n731 ;
  assign n733 = n732 ^ n719 ;
  assign n727 = n713 ^ n712 ;
  assign n728 = ~n715 & n727 ;
  assign n729 = n728 ^ n712 ;
  assign n724 = n723 ^ n717 ;
  assign n725 = n718 & ~n724 ;
  assign n726 = n725 ^ n716 ;
  assign n730 = n729 ^ n726 ;
  assign n734 = n733 ^ n730 ;
  assign n754 = n753 ^ n734 ;
  assign n780 = n765 ^ n754 ;
  assign n816 = n815 ^ n780 ;
  assign n843 = n842 ^ n827 ;
  assign n844 = n843 ^ n780 ;
  assign n845 = n816 & ~n844 ;
  assign n846 = n845 ^ n815 ;
  assign n773 = n764 ^ n760 ;
  assign n774 = n761 & ~n773 ;
  assign n775 = n774 ^ n757 ;
  assign n769 = n733 ^ n729 ;
  assign n770 = n730 & ~n769 ;
  assign n771 = n770 ^ n726 ;
  assign n766 = n765 ^ n753 ;
  assign n767 = n754 & ~n766 ;
  assign n768 = n767 ^ n734 ;
  assign n772 = n771 ^ n768 ;
  assign n779 = n775 ^ n772 ;
  assign n847 = n846 ^ n779 ;
  assign n858 = n857 ^ n850 ;
  assign n859 = n858 ^ n846 ;
  assign n860 = n847 & ~n859 ;
  assign n861 = n860 ^ n779 ;
  assign n776 = n775 ^ n771 ;
  assign n777 = n772 & ~n776 ;
  assign n778 = n777 ^ n768 ;
  assign n862 = n861 ^ n778 ;
  assign n866 = n865 ^ n862 ;
  assign n867 = n812 ^ n783 ;
  assign n868 = x512 ^ x64 ;
  assign n869 = n867 & n868 ;
  assign n870 = n843 ^ n816 ;
  assign n871 = n869 & n870 ;
  assign n872 = n858 ^ n847 ;
  assign n873 = n871 & n872 ;
  assign n874 = n866 & n873 ;
  assign n875 = n865 ^ n861 ;
  assign n876 = n862 & ~n875 ;
  assign n877 = n876 ^ n778 ;
  assign n878 = n874 & n877 ;
  assign n977 = x514 ^ x98 ;
  assign n974 = x522 ^ x106 ;
  assign n972 = x528 ^ x112 ;
  assign n970 = x526 ^ x110 ;
  assign n969 = x527 ^ x111 ;
  assign n971 = n970 ^ n969 ;
  assign n973 = n972 ^ n971 ;
  assign n975 = n974 ^ n973 ;
  assign n967 = x525 ^ x109 ;
  assign n965 = x523 ^ x107 ;
  assign n964 = x524 ^ x108 ;
  assign n966 = n965 ^ n964 ;
  assign n968 = n967 ^ n966 ;
  assign n976 = n975 ^ n968 ;
  assign n978 = n977 ^ n976 ;
  assign n961 = x515 ^ x99 ;
  assign n959 = x521 ^ x105 ;
  assign n957 = x519 ^ x103 ;
  assign n956 = x520 ^ x104 ;
  assign n958 = n957 ^ n956 ;
  assign n960 = n959 ^ n958 ;
  assign n962 = n961 ^ n960 ;
  assign n954 = x518 ^ x102 ;
  assign n952 = x516 ^ x100 ;
  assign n951 = x517 ^ x101 ;
  assign n953 = n952 ^ n951 ;
  assign n955 = n954 ^ n953 ;
  assign n963 = n962 ^ n955 ;
  assign n1006 = n977 ^ n963 ;
  assign n1007 = n978 & ~n1006 ;
  assign n1008 = n1007 ^ n976 ;
  assign n1002 = n967 ^ n965 ;
  assign n1003 = n966 & ~n1002 ;
  assign n1004 = n1003 ^ n964 ;
  assign n998 = n972 ^ n970 ;
  assign n999 = n971 & ~n998 ;
  assign n1000 = n999 ^ n969 ;
  assign n995 = n973 ^ n968 ;
  assign n996 = ~n975 & n995 ;
  assign n997 = n996 ^ n968 ;
  assign n1001 = n1000 ^ n997 ;
  assign n1005 = n1004 ^ n1001 ;
  assign n1009 = n1008 ^ n1005 ;
  assign n991 = n954 ^ n952 ;
  assign n992 = n953 & ~n991 ;
  assign n993 = n992 ^ n951 ;
  assign n987 = n960 ^ n955 ;
  assign n988 = ~n962 & n987 ;
  assign n989 = n988 ^ n955 ;
  assign n984 = n959 ^ n957 ;
  assign n985 = n958 & ~n984 ;
  assign n986 = n985 ^ n956 ;
  assign n990 = n989 ^ n986 ;
  assign n994 = n993 ^ n990 ;
  assign n1021 = n1008 ^ n994 ;
  assign n1022 = n1009 & ~n1021 ;
  assign n1023 = n1022 ^ n1005 ;
  assign n1018 = n1004 ^ n1000 ;
  assign n1019 = n1001 & ~n1018 ;
  assign n1020 = n1019 ^ n997 ;
  assign n1024 = n1023 ^ n1020 ;
  assign n1015 = n993 ^ n989 ;
  assign n1016 = n990 & ~n1015 ;
  assign n1017 = n1016 ^ n986 ;
  assign n1030 = n1020 ^ n1017 ;
  assign n1031 = ~n1024 & n1030 ;
  assign n1032 = n1031 ^ n1017 ;
  assign n949 = x513 ^ x97 ;
  assign n915 = x533 ^ x117 ;
  assign n913 = x531 ^ x115 ;
  assign n912 = x532 ^ x116 ;
  assign n914 = n913 ^ n912 ;
  assign n916 = n915 ^ n914 ;
  assign n910 = x530 ^ x114 ;
  assign n908 = x536 ^ x120 ;
  assign n906 = x534 ^ x118 ;
  assign n905 = x535 ^ x119 ;
  assign n907 = n906 ^ n905 ;
  assign n909 = n908 ^ n907 ;
  assign n911 = n910 ^ n909 ;
  assign n917 = n916 ^ n911 ;
  assign n888 = x538 ^ x122 ;
  assign n887 = x539 ^ x123 ;
  assign n889 = n888 ^ n887 ;
  assign n886 = x540 ^ x124 ;
  assign n890 = n889 ^ n886 ;
  assign n884 = x537 ^ x121 ;
  assign n881 = x541 ^ x125 ;
  assign n880 = x542 ^ x126 ;
  assign n882 = n881 ^ n880 ;
  assign n879 = x543 ^ x127 ;
  assign n883 = n882 ^ n879 ;
  assign n885 = n884 ^ n883 ;
  assign n903 = n890 ^ n885 ;
  assign n902 = x529 ^ x113 ;
  assign n904 = n903 ^ n902 ;
  assign n948 = n917 ^ n904 ;
  assign n950 = n949 ^ n948 ;
  assign n979 = n978 ^ n963 ;
  assign n980 = n979 ^ n949 ;
  assign n981 = n950 & ~n980 ;
  assign n982 = n981 ^ n948 ;
  assign n929 = n915 ^ n913 ;
  assign n930 = n914 & ~n929 ;
  assign n931 = n930 ^ n912 ;
  assign n925 = n908 ^ n906 ;
  assign n926 = n907 & ~n925 ;
  assign n927 = n926 ^ n905 ;
  assign n922 = n916 ^ n910 ;
  assign n923 = n911 & ~n922 ;
  assign n924 = n923 ^ n909 ;
  assign n928 = n927 ^ n924 ;
  assign n932 = n931 ^ n928 ;
  assign n918 = n917 ^ n903 ;
  assign n919 = n904 & ~n918 ;
  assign n920 = n919 ^ n902 ;
  assign n898 = n887 ^ n886 ;
  assign n899 = ~n889 & n898 ;
  assign n900 = n899 ^ n886 ;
  assign n894 = n880 ^ n879 ;
  assign n895 = ~n882 & n894 ;
  assign n896 = n895 ^ n879 ;
  assign n891 = n890 ^ n884 ;
  assign n892 = n885 & ~n891 ;
  assign n893 = n892 ^ n883 ;
  assign n897 = n896 ^ n893 ;
  assign n901 = n900 ^ n897 ;
  assign n921 = n920 ^ n901 ;
  assign n947 = n932 ^ n921 ;
  assign n983 = n982 ^ n947 ;
  assign n1010 = n1009 ^ n994 ;
  assign n1011 = n1010 ^ n947 ;
  assign n1012 = n983 & ~n1011 ;
  assign n1013 = n1012 ^ n982 ;
  assign n940 = n931 ^ n927 ;
  assign n941 = n928 & ~n940 ;
  assign n942 = n941 ^ n924 ;
  assign n936 = n900 ^ n896 ;
  assign n937 = n897 & ~n936 ;
  assign n938 = n937 ^ n893 ;
  assign n933 = n932 ^ n920 ;
  assign n934 = n921 & ~n933 ;
  assign n935 = n934 ^ n901 ;
  assign n939 = n938 ^ n935 ;
  assign n946 = n942 ^ n939 ;
  assign n1014 = n1013 ^ n946 ;
  assign n1025 = n1024 ^ n1017 ;
  assign n1026 = n1025 ^ n1013 ;
  assign n1027 = n1014 & ~n1026 ;
  assign n1028 = n1027 ^ n946 ;
  assign n943 = n942 ^ n938 ;
  assign n944 = n939 & ~n943 ;
  assign n945 = n944 ^ n935 ;
  assign n1029 = n1028 ^ n945 ;
  assign n1033 = n1032 ^ n1029 ;
  assign n1034 = n1010 ^ n983 ;
  assign n1035 = n979 ^ n950 ;
  assign n1036 = x512 ^ x96 ;
  assign n1037 = n1035 & n1036 ;
  assign n1038 = n1034 & n1037 ;
  assign n1039 = n1025 ^ n1014 ;
  assign n1040 = n1038 & n1039 ;
  assign n1041 = n1033 & n1040 ;
  assign n1042 = n1032 ^ n1028 ;
  assign n1043 = n1029 & ~n1042 ;
  assign n1044 = n1043 ^ n945 ;
  assign n1045 = n1041 & n1044 ;
  assign n1144 = x514 ^ x130 ;
  assign n1141 = x522 ^ x138 ;
  assign n1139 = x528 ^ x144 ;
  assign n1137 = x526 ^ x142 ;
  assign n1136 = x527 ^ x143 ;
  assign n1138 = n1137 ^ n1136 ;
  assign n1140 = n1139 ^ n1138 ;
  assign n1142 = n1141 ^ n1140 ;
  assign n1134 = x525 ^ x141 ;
  assign n1132 = x523 ^ x139 ;
  assign n1131 = x524 ^ x140 ;
  assign n1133 = n1132 ^ n1131 ;
  assign n1135 = n1134 ^ n1133 ;
  assign n1143 = n1142 ^ n1135 ;
  assign n1145 = n1144 ^ n1143 ;
  assign n1128 = x515 ^ x131 ;
  assign n1126 = x521 ^ x137 ;
  assign n1124 = x519 ^ x135 ;
  assign n1123 = x520 ^ x136 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1127 = n1126 ^ n1125 ;
  assign n1129 = n1128 ^ n1127 ;
  assign n1121 = x518 ^ x134 ;
  assign n1119 = x516 ^ x132 ;
  assign n1118 = x517 ^ x133 ;
  assign n1120 = n1119 ^ n1118 ;
  assign n1122 = n1121 ^ n1120 ;
  assign n1130 = n1129 ^ n1122 ;
  assign n1173 = n1144 ^ n1130 ;
  assign n1174 = n1145 & ~n1173 ;
  assign n1175 = n1174 ^ n1143 ;
  assign n1169 = n1134 ^ n1132 ;
  assign n1170 = n1133 & ~n1169 ;
  assign n1171 = n1170 ^ n1131 ;
  assign n1165 = n1139 ^ n1137 ;
  assign n1166 = n1138 & ~n1165 ;
  assign n1167 = n1166 ^ n1136 ;
  assign n1162 = n1140 ^ n1135 ;
  assign n1163 = ~n1142 & n1162 ;
  assign n1164 = n1163 ^ n1135 ;
  assign n1168 = n1167 ^ n1164 ;
  assign n1172 = n1171 ^ n1168 ;
  assign n1176 = n1175 ^ n1172 ;
  assign n1158 = n1121 ^ n1119 ;
  assign n1159 = n1120 & ~n1158 ;
  assign n1160 = n1159 ^ n1118 ;
  assign n1154 = n1127 ^ n1122 ;
  assign n1155 = ~n1129 & n1154 ;
  assign n1156 = n1155 ^ n1122 ;
  assign n1151 = n1126 ^ n1124 ;
  assign n1152 = n1125 & ~n1151 ;
  assign n1153 = n1152 ^ n1123 ;
  assign n1157 = n1156 ^ n1153 ;
  assign n1161 = n1160 ^ n1157 ;
  assign n1188 = n1175 ^ n1161 ;
  assign n1189 = n1176 & ~n1188 ;
  assign n1190 = n1189 ^ n1172 ;
  assign n1185 = n1171 ^ n1167 ;
  assign n1186 = n1168 & ~n1185 ;
  assign n1187 = n1186 ^ n1164 ;
  assign n1191 = n1190 ^ n1187 ;
  assign n1182 = n1160 ^ n1156 ;
  assign n1183 = n1157 & ~n1182 ;
  assign n1184 = n1183 ^ n1153 ;
  assign n1197 = n1187 ^ n1184 ;
  assign n1198 = ~n1191 & n1197 ;
  assign n1199 = n1198 ^ n1184 ;
  assign n1116 = x513 ^ x129 ;
  assign n1082 = x533 ^ x149 ;
  assign n1080 = x531 ^ x147 ;
  assign n1079 = x532 ^ x148 ;
  assign n1081 = n1080 ^ n1079 ;
  assign n1083 = n1082 ^ n1081 ;
  assign n1077 = x530 ^ x146 ;
  assign n1075 = x536 ^ x152 ;
  assign n1073 = x534 ^ x150 ;
  assign n1072 = x535 ^ x151 ;
  assign n1074 = n1073 ^ n1072 ;
  assign n1076 = n1075 ^ n1074 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1084 = n1083 ^ n1078 ;
  assign n1055 = x538 ^ x154 ;
  assign n1054 = x539 ^ x155 ;
  assign n1056 = n1055 ^ n1054 ;
  assign n1053 = x540 ^ x156 ;
  assign n1057 = n1056 ^ n1053 ;
  assign n1051 = x537 ^ x153 ;
  assign n1048 = x541 ^ x157 ;
  assign n1047 = x542 ^ x158 ;
  assign n1049 = n1048 ^ n1047 ;
  assign n1046 = x543 ^ x159 ;
  assign n1050 = n1049 ^ n1046 ;
  assign n1052 = n1051 ^ n1050 ;
  assign n1070 = n1057 ^ n1052 ;
  assign n1069 = x529 ^ x145 ;
  assign n1071 = n1070 ^ n1069 ;
  assign n1115 = n1084 ^ n1071 ;
  assign n1117 = n1116 ^ n1115 ;
  assign n1146 = n1145 ^ n1130 ;
  assign n1147 = n1146 ^ n1116 ;
  assign n1148 = n1117 & ~n1147 ;
  assign n1149 = n1148 ^ n1115 ;
  assign n1096 = n1082 ^ n1080 ;
  assign n1097 = n1081 & ~n1096 ;
  assign n1098 = n1097 ^ n1079 ;
  assign n1092 = n1075 ^ n1073 ;
  assign n1093 = n1074 & ~n1092 ;
  assign n1094 = n1093 ^ n1072 ;
  assign n1089 = n1083 ^ n1077 ;
  assign n1090 = n1078 & ~n1089 ;
  assign n1091 = n1090 ^ n1076 ;
  assign n1095 = n1094 ^ n1091 ;
  assign n1099 = n1098 ^ n1095 ;
  assign n1085 = n1084 ^ n1070 ;
  assign n1086 = n1071 & ~n1085 ;
  assign n1087 = n1086 ^ n1069 ;
  assign n1065 = n1054 ^ n1053 ;
  assign n1066 = ~n1056 & n1065 ;
  assign n1067 = n1066 ^ n1053 ;
  assign n1061 = n1047 ^ n1046 ;
  assign n1062 = ~n1049 & n1061 ;
  assign n1063 = n1062 ^ n1046 ;
  assign n1058 = n1057 ^ n1051 ;
  assign n1059 = n1052 & ~n1058 ;
  assign n1060 = n1059 ^ n1050 ;
  assign n1064 = n1063 ^ n1060 ;
  assign n1068 = n1067 ^ n1064 ;
  assign n1088 = n1087 ^ n1068 ;
  assign n1114 = n1099 ^ n1088 ;
  assign n1150 = n1149 ^ n1114 ;
  assign n1177 = n1176 ^ n1161 ;
  assign n1178 = n1177 ^ n1114 ;
  assign n1179 = n1150 & ~n1178 ;
  assign n1180 = n1179 ^ n1149 ;
  assign n1107 = n1098 ^ n1094 ;
  assign n1108 = n1095 & ~n1107 ;
  assign n1109 = n1108 ^ n1091 ;
  assign n1103 = n1067 ^ n1063 ;
  assign n1104 = n1064 & ~n1103 ;
  assign n1105 = n1104 ^ n1060 ;
  assign n1100 = n1099 ^ n1087 ;
  assign n1101 = n1088 & ~n1100 ;
  assign n1102 = n1101 ^ n1068 ;
  assign n1106 = n1105 ^ n1102 ;
  assign n1113 = n1109 ^ n1106 ;
  assign n1181 = n1180 ^ n1113 ;
  assign n1192 = n1191 ^ n1184 ;
  assign n1193 = n1192 ^ n1180 ;
  assign n1194 = n1181 & ~n1193 ;
  assign n1195 = n1194 ^ n1113 ;
  assign n1110 = n1109 ^ n1105 ;
  assign n1111 = n1106 & ~n1110 ;
  assign n1112 = n1111 ^ n1102 ;
  assign n1196 = n1195 ^ n1112 ;
  assign n1200 = n1199 ^ n1196 ;
  assign n1201 = n1177 ^ n1150 ;
  assign n1202 = n1146 ^ n1117 ;
  assign n1203 = x512 ^ x128 ;
  assign n1204 = n1202 & n1203 ;
  assign n1205 = n1201 & n1204 ;
  assign n1206 = n1192 ^ n1181 ;
  assign n1207 = n1205 & n1206 ;
  assign n1208 = n1200 & n1207 ;
  assign n1209 = n1199 ^ n1195 ;
  assign n1210 = n1196 & ~n1209 ;
  assign n1211 = n1210 ^ n1112 ;
  assign n1212 = n1208 & n1211 ;
  assign n1311 = x514 ^ x162 ;
  assign n1308 = x522 ^ x170 ;
  assign n1306 = x528 ^ x176 ;
  assign n1304 = x526 ^ x174 ;
  assign n1303 = x527 ^ x175 ;
  assign n1305 = n1304 ^ n1303 ;
  assign n1307 = n1306 ^ n1305 ;
  assign n1309 = n1308 ^ n1307 ;
  assign n1301 = x525 ^ x173 ;
  assign n1299 = x523 ^ x171 ;
  assign n1298 = x524 ^ x172 ;
  assign n1300 = n1299 ^ n1298 ;
  assign n1302 = n1301 ^ n1300 ;
  assign n1310 = n1309 ^ n1302 ;
  assign n1312 = n1311 ^ n1310 ;
  assign n1295 = x515 ^ x163 ;
  assign n1293 = x521 ^ x169 ;
  assign n1291 = x519 ^ x167 ;
  assign n1290 = x520 ^ x168 ;
  assign n1292 = n1291 ^ n1290 ;
  assign n1294 = n1293 ^ n1292 ;
  assign n1296 = n1295 ^ n1294 ;
  assign n1288 = x518 ^ x166 ;
  assign n1286 = x516 ^ x164 ;
  assign n1285 = x517 ^ x165 ;
  assign n1287 = n1286 ^ n1285 ;
  assign n1289 = n1288 ^ n1287 ;
  assign n1297 = n1296 ^ n1289 ;
  assign n1340 = n1311 ^ n1297 ;
  assign n1341 = n1312 & ~n1340 ;
  assign n1342 = n1341 ^ n1310 ;
  assign n1336 = n1301 ^ n1299 ;
  assign n1337 = n1300 & ~n1336 ;
  assign n1338 = n1337 ^ n1298 ;
  assign n1332 = n1306 ^ n1304 ;
  assign n1333 = n1305 & ~n1332 ;
  assign n1334 = n1333 ^ n1303 ;
  assign n1329 = n1307 ^ n1302 ;
  assign n1330 = ~n1309 & n1329 ;
  assign n1331 = n1330 ^ n1302 ;
  assign n1335 = n1334 ^ n1331 ;
  assign n1339 = n1338 ^ n1335 ;
  assign n1343 = n1342 ^ n1339 ;
  assign n1325 = n1288 ^ n1286 ;
  assign n1326 = n1287 & ~n1325 ;
  assign n1327 = n1326 ^ n1285 ;
  assign n1321 = n1294 ^ n1289 ;
  assign n1322 = ~n1296 & n1321 ;
  assign n1323 = n1322 ^ n1289 ;
  assign n1318 = n1293 ^ n1291 ;
  assign n1319 = n1292 & ~n1318 ;
  assign n1320 = n1319 ^ n1290 ;
  assign n1324 = n1323 ^ n1320 ;
  assign n1328 = n1327 ^ n1324 ;
  assign n1355 = n1342 ^ n1328 ;
  assign n1356 = n1343 & ~n1355 ;
  assign n1357 = n1356 ^ n1339 ;
  assign n1352 = n1338 ^ n1334 ;
  assign n1353 = n1335 & ~n1352 ;
  assign n1354 = n1353 ^ n1331 ;
  assign n1358 = n1357 ^ n1354 ;
  assign n1349 = n1327 ^ n1323 ;
  assign n1350 = n1324 & ~n1349 ;
  assign n1351 = n1350 ^ n1320 ;
  assign n1364 = n1354 ^ n1351 ;
  assign n1365 = ~n1358 & n1364 ;
  assign n1366 = n1365 ^ n1351 ;
  assign n1283 = x513 ^ x161 ;
  assign n1249 = x533 ^ x181 ;
  assign n1247 = x531 ^ x179 ;
  assign n1246 = x532 ^ x180 ;
  assign n1248 = n1247 ^ n1246 ;
  assign n1250 = n1249 ^ n1248 ;
  assign n1244 = x530 ^ x178 ;
  assign n1242 = x536 ^ x184 ;
  assign n1240 = x534 ^ x182 ;
  assign n1239 = x535 ^ x183 ;
  assign n1241 = n1240 ^ n1239 ;
  assign n1243 = n1242 ^ n1241 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1251 = n1250 ^ n1245 ;
  assign n1222 = x538 ^ x186 ;
  assign n1221 = x539 ^ x187 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1220 = x540 ^ x188 ;
  assign n1224 = n1223 ^ n1220 ;
  assign n1218 = x537 ^ x185 ;
  assign n1215 = x541 ^ x189 ;
  assign n1214 = x542 ^ x190 ;
  assign n1216 = n1215 ^ n1214 ;
  assign n1213 = x543 ^ x191 ;
  assign n1217 = n1216 ^ n1213 ;
  assign n1219 = n1218 ^ n1217 ;
  assign n1237 = n1224 ^ n1219 ;
  assign n1236 = x529 ^ x177 ;
  assign n1238 = n1237 ^ n1236 ;
  assign n1282 = n1251 ^ n1238 ;
  assign n1284 = n1283 ^ n1282 ;
  assign n1313 = n1312 ^ n1297 ;
  assign n1314 = n1313 ^ n1283 ;
  assign n1315 = n1284 & ~n1314 ;
  assign n1316 = n1315 ^ n1282 ;
  assign n1263 = n1249 ^ n1247 ;
  assign n1264 = n1248 & ~n1263 ;
  assign n1265 = n1264 ^ n1246 ;
  assign n1259 = n1242 ^ n1240 ;
  assign n1260 = n1241 & ~n1259 ;
  assign n1261 = n1260 ^ n1239 ;
  assign n1256 = n1250 ^ n1244 ;
  assign n1257 = n1245 & ~n1256 ;
  assign n1258 = n1257 ^ n1243 ;
  assign n1262 = n1261 ^ n1258 ;
  assign n1266 = n1265 ^ n1262 ;
  assign n1252 = n1251 ^ n1237 ;
  assign n1253 = n1238 & ~n1252 ;
  assign n1254 = n1253 ^ n1236 ;
  assign n1232 = n1221 ^ n1220 ;
  assign n1233 = ~n1223 & n1232 ;
  assign n1234 = n1233 ^ n1220 ;
  assign n1228 = n1214 ^ n1213 ;
  assign n1229 = ~n1216 & n1228 ;
  assign n1230 = n1229 ^ n1213 ;
  assign n1225 = n1224 ^ n1218 ;
  assign n1226 = n1219 & ~n1225 ;
  assign n1227 = n1226 ^ n1217 ;
  assign n1231 = n1230 ^ n1227 ;
  assign n1235 = n1234 ^ n1231 ;
  assign n1255 = n1254 ^ n1235 ;
  assign n1281 = n1266 ^ n1255 ;
  assign n1317 = n1316 ^ n1281 ;
  assign n1344 = n1343 ^ n1328 ;
  assign n1345 = n1344 ^ n1281 ;
  assign n1346 = n1317 & ~n1345 ;
  assign n1347 = n1346 ^ n1316 ;
  assign n1274 = n1265 ^ n1261 ;
  assign n1275 = n1262 & ~n1274 ;
  assign n1276 = n1275 ^ n1258 ;
  assign n1270 = n1234 ^ n1230 ;
  assign n1271 = n1231 & ~n1270 ;
  assign n1272 = n1271 ^ n1227 ;
  assign n1267 = n1266 ^ n1254 ;
  assign n1268 = n1255 & ~n1267 ;
  assign n1269 = n1268 ^ n1235 ;
  assign n1273 = n1272 ^ n1269 ;
  assign n1280 = n1276 ^ n1273 ;
  assign n1348 = n1347 ^ n1280 ;
  assign n1359 = n1358 ^ n1351 ;
  assign n1360 = n1359 ^ n1347 ;
  assign n1361 = n1348 & ~n1360 ;
  assign n1362 = n1361 ^ n1280 ;
  assign n1277 = n1276 ^ n1272 ;
  assign n1278 = n1273 & ~n1277 ;
  assign n1279 = n1278 ^ n1269 ;
  assign n1363 = n1362 ^ n1279 ;
  assign n1367 = n1366 ^ n1363 ;
  assign n1368 = n1344 ^ n1317 ;
  assign n1369 = n1313 ^ n1284 ;
  assign n1370 = x512 ^ x160 ;
  assign n1371 = n1369 & n1370 ;
  assign n1372 = n1368 & n1371 ;
  assign n1373 = n1359 ^ n1348 ;
  assign n1374 = n1372 & n1373 ;
  assign n1375 = n1367 & n1374 ;
  assign n1376 = n1366 ^ n1362 ;
  assign n1377 = n1363 & ~n1376 ;
  assign n1378 = n1377 ^ n1279 ;
  assign n1379 = n1375 & n1378 ;
  assign n1478 = x514 ^ x194 ;
  assign n1475 = x522 ^ x202 ;
  assign n1473 = x528 ^ x208 ;
  assign n1471 = x526 ^ x206 ;
  assign n1470 = x527 ^ x207 ;
  assign n1472 = n1471 ^ n1470 ;
  assign n1474 = n1473 ^ n1472 ;
  assign n1476 = n1475 ^ n1474 ;
  assign n1468 = x525 ^ x205 ;
  assign n1466 = x523 ^ x203 ;
  assign n1465 = x524 ^ x204 ;
  assign n1467 = n1466 ^ n1465 ;
  assign n1469 = n1468 ^ n1467 ;
  assign n1477 = n1476 ^ n1469 ;
  assign n1479 = n1478 ^ n1477 ;
  assign n1462 = x515 ^ x195 ;
  assign n1460 = x521 ^ x201 ;
  assign n1458 = x519 ^ x199 ;
  assign n1457 = x520 ^ x200 ;
  assign n1459 = n1458 ^ n1457 ;
  assign n1461 = n1460 ^ n1459 ;
  assign n1463 = n1462 ^ n1461 ;
  assign n1455 = x518 ^ x198 ;
  assign n1453 = x516 ^ x196 ;
  assign n1452 = x517 ^ x197 ;
  assign n1454 = n1453 ^ n1452 ;
  assign n1456 = n1455 ^ n1454 ;
  assign n1464 = n1463 ^ n1456 ;
  assign n1507 = n1478 ^ n1464 ;
  assign n1508 = n1479 & ~n1507 ;
  assign n1509 = n1508 ^ n1477 ;
  assign n1503 = n1468 ^ n1466 ;
  assign n1504 = n1467 & ~n1503 ;
  assign n1505 = n1504 ^ n1465 ;
  assign n1499 = n1473 ^ n1471 ;
  assign n1500 = n1472 & ~n1499 ;
  assign n1501 = n1500 ^ n1470 ;
  assign n1496 = n1474 ^ n1469 ;
  assign n1497 = ~n1476 & n1496 ;
  assign n1498 = n1497 ^ n1469 ;
  assign n1502 = n1501 ^ n1498 ;
  assign n1506 = n1505 ^ n1502 ;
  assign n1510 = n1509 ^ n1506 ;
  assign n1492 = n1455 ^ n1453 ;
  assign n1493 = n1454 & ~n1492 ;
  assign n1494 = n1493 ^ n1452 ;
  assign n1488 = n1461 ^ n1456 ;
  assign n1489 = ~n1463 & n1488 ;
  assign n1490 = n1489 ^ n1456 ;
  assign n1485 = n1460 ^ n1458 ;
  assign n1486 = n1459 & ~n1485 ;
  assign n1487 = n1486 ^ n1457 ;
  assign n1491 = n1490 ^ n1487 ;
  assign n1495 = n1494 ^ n1491 ;
  assign n1522 = n1509 ^ n1495 ;
  assign n1523 = n1510 & ~n1522 ;
  assign n1524 = n1523 ^ n1506 ;
  assign n1519 = n1505 ^ n1501 ;
  assign n1520 = n1502 & ~n1519 ;
  assign n1521 = n1520 ^ n1498 ;
  assign n1525 = n1524 ^ n1521 ;
  assign n1516 = n1494 ^ n1490 ;
  assign n1517 = n1491 & ~n1516 ;
  assign n1518 = n1517 ^ n1487 ;
  assign n1531 = n1521 ^ n1518 ;
  assign n1532 = ~n1525 & n1531 ;
  assign n1533 = n1532 ^ n1518 ;
  assign n1450 = x513 ^ x193 ;
  assign n1416 = x533 ^ x213 ;
  assign n1414 = x531 ^ x211 ;
  assign n1413 = x532 ^ x212 ;
  assign n1415 = n1414 ^ n1413 ;
  assign n1417 = n1416 ^ n1415 ;
  assign n1411 = x530 ^ x210 ;
  assign n1409 = x536 ^ x216 ;
  assign n1407 = x534 ^ x214 ;
  assign n1406 = x535 ^ x215 ;
  assign n1408 = n1407 ^ n1406 ;
  assign n1410 = n1409 ^ n1408 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1418 = n1417 ^ n1412 ;
  assign n1389 = x538 ^ x218 ;
  assign n1388 = x539 ^ x219 ;
  assign n1390 = n1389 ^ n1388 ;
  assign n1387 = x540 ^ x220 ;
  assign n1391 = n1390 ^ n1387 ;
  assign n1385 = x537 ^ x217 ;
  assign n1382 = x541 ^ x221 ;
  assign n1381 = x542 ^ x222 ;
  assign n1383 = n1382 ^ n1381 ;
  assign n1380 = x543 ^ x223 ;
  assign n1384 = n1383 ^ n1380 ;
  assign n1386 = n1385 ^ n1384 ;
  assign n1404 = n1391 ^ n1386 ;
  assign n1403 = x529 ^ x209 ;
  assign n1405 = n1404 ^ n1403 ;
  assign n1449 = n1418 ^ n1405 ;
  assign n1451 = n1450 ^ n1449 ;
  assign n1480 = n1479 ^ n1464 ;
  assign n1481 = n1480 ^ n1450 ;
  assign n1482 = n1451 & ~n1481 ;
  assign n1483 = n1482 ^ n1449 ;
  assign n1430 = n1416 ^ n1414 ;
  assign n1431 = n1415 & ~n1430 ;
  assign n1432 = n1431 ^ n1413 ;
  assign n1426 = n1409 ^ n1407 ;
  assign n1427 = n1408 & ~n1426 ;
  assign n1428 = n1427 ^ n1406 ;
  assign n1423 = n1417 ^ n1411 ;
  assign n1424 = n1412 & ~n1423 ;
  assign n1425 = n1424 ^ n1410 ;
  assign n1429 = n1428 ^ n1425 ;
  assign n1433 = n1432 ^ n1429 ;
  assign n1419 = n1418 ^ n1404 ;
  assign n1420 = n1405 & ~n1419 ;
  assign n1421 = n1420 ^ n1403 ;
  assign n1399 = n1388 ^ n1387 ;
  assign n1400 = ~n1390 & n1399 ;
  assign n1401 = n1400 ^ n1387 ;
  assign n1395 = n1381 ^ n1380 ;
  assign n1396 = ~n1383 & n1395 ;
  assign n1397 = n1396 ^ n1380 ;
  assign n1392 = n1391 ^ n1385 ;
  assign n1393 = n1386 & ~n1392 ;
  assign n1394 = n1393 ^ n1384 ;
  assign n1398 = n1397 ^ n1394 ;
  assign n1402 = n1401 ^ n1398 ;
  assign n1422 = n1421 ^ n1402 ;
  assign n1448 = n1433 ^ n1422 ;
  assign n1484 = n1483 ^ n1448 ;
  assign n1511 = n1510 ^ n1495 ;
  assign n1512 = n1511 ^ n1448 ;
  assign n1513 = n1484 & ~n1512 ;
  assign n1514 = n1513 ^ n1483 ;
  assign n1441 = n1432 ^ n1428 ;
  assign n1442 = n1429 & ~n1441 ;
  assign n1443 = n1442 ^ n1425 ;
  assign n1437 = n1401 ^ n1397 ;
  assign n1438 = n1398 & ~n1437 ;
  assign n1439 = n1438 ^ n1394 ;
  assign n1434 = n1433 ^ n1421 ;
  assign n1435 = n1422 & ~n1434 ;
  assign n1436 = n1435 ^ n1402 ;
  assign n1440 = n1439 ^ n1436 ;
  assign n1447 = n1443 ^ n1440 ;
  assign n1515 = n1514 ^ n1447 ;
  assign n1526 = n1525 ^ n1518 ;
  assign n1527 = n1526 ^ n1514 ;
  assign n1528 = n1515 & ~n1527 ;
  assign n1529 = n1528 ^ n1447 ;
  assign n1444 = n1443 ^ n1439 ;
  assign n1445 = n1440 & ~n1444 ;
  assign n1446 = n1445 ^ n1436 ;
  assign n1530 = n1529 ^ n1446 ;
  assign n1534 = n1533 ^ n1530 ;
  assign n1535 = n1511 ^ n1484 ;
  assign n1536 = n1480 ^ n1451 ;
  assign n1537 = x512 ^ x192 ;
  assign n1538 = n1536 & n1537 ;
  assign n1539 = n1535 & n1538 ;
  assign n1540 = n1526 ^ n1515 ;
  assign n1541 = n1539 & n1540 ;
  assign n1542 = n1534 & n1541 ;
  assign n1543 = n1533 ^ n1529 ;
  assign n1544 = n1530 & ~n1543 ;
  assign n1545 = n1544 ^ n1446 ;
  assign n1546 = n1542 & n1545 ;
  assign n1645 = x514 ^ x226 ;
  assign n1642 = x522 ^ x234 ;
  assign n1640 = x528 ^ x240 ;
  assign n1638 = x526 ^ x238 ;
  assign n1637 = x527 ^ x239 ;
  assign n1639 = n1638 ^ n1637 ;
  assign n1641 = n1640 ^ n1639 ;
  assign n1643 = n1642 ^ n1641 ;
  assign n1635 = x525 ^ x237 ;
  assign n1633 = x523 ^ x235 ;
  assign n1632 = x524 ^ x236 ;
  assign n1634 = n1633 ^ n1632 ;
  assign n1636 = n1635 ^ n1634 ;
  assign n1644 = n1643 ^ n1636 ;
  assign n1646 = n1645 ^ n1644 ;
  assign n1629 = x515 ^ x227 ;
  assign n1627 = x521 ^ x233 ;
  assign n1625 = x519 ^ x231 ;
  assign n1624 = x520 ^ x232 ;
  assign n1626 = n1625 ^ n1624 ;
  assign n1628 = n1627 ^ n1626 ;
  assign n1630 = n1629 ^ n1628 ;
  assign n1622 = x518 ^ x230 ;
  assign n1620 = x516 ^ x228 ;
  assign n1619 = x517 ^ x229 ;
  assign n1621 = n1620 ^ n1619 ;
  assign n1623 = n1622 ^ n1621 ;
  assign n1631 = n1630 ^ n1623 ;
  assign n1674 = n1645 ^ n1631 ;
  assign n1675 = n1646 & ~n1674 ;
  assign n1676 = n1675 ^ n1644 ;
  assign n1670 = n1635 ^ n1633 ;
  assign n1671 = n1634 & ~n1670 ;
  assign n1672 = n1671 ^ n1632 ;
  assign n1666 = n1640 ^ n1638 ;
  assign n1667 = n1639 & ~n1666 ;
  assign n1668 = n1667 ^ n1637 ;
  assign n1663 = n1641 ^ n1636 ;
  assign n1664 = ~n1643 & n1663 ;
  assign n1665 = n1664 ^ n1636 ;
  assign n1669 = n1668 ^ n1665 ;
  assign n1673 = n1672 ^ n1669 ;
  assign n1677 = n1676 ^ n1673 ;
  assign n1659 = n1622 ^ n1620 ;
  assign n1660 = n1621 & ~n1659 ;
  assign n1661 = n1660 ^ n1619 ;
  assign n1655 = n1628 ^ n1623 ;
  assign n1656 = ~n1630 & n1655 ;
  assign n1657 = n1656 ^ n1623 ;
  assign n1652 = n1627 ^ n1625 ;
  assign n1653 = n1626 & ~n1652 ;
  assign n1654 = n1653 ^ n1624 ;
  assign n1658 = n1657 ^ n1654 ;
  assign n1662 = n1661 ^ n1658 ;
  assign n1689 = n1676 ^ n1662 ;
  assign n1690 = n1677 & ~n1689 ;
  assign n1691 = n1690 ^ n1673 ;
  assign n1686 = n1672 ^ n1668 ;
  assign n1687 = n1669 & ~n1686 ;
  assign n1688 = n1687 ^ n1665 ;
  assign n1692 = n1691 ^ n1688 ;
  assign n1683 = n1661 ^ n1657 ;
  assign n1684 = n1658 & ~n1683 ;
  assign n1685 = n1684 ^ n1654 ;
  assign n1698 = n1688 ^ n1685 ;
  assign n1699 = ~n1692 & n1698 ;
  assign n1700 = n1699 ^ n1685 ;
  assign n1617 = x513 ^ x225 ;
  assign n1583 = x533 ^ x245 ;
  assign n1581 = x531 ^ x243 ;
  assign n1580 = x532 ^ x244 ;
  assign n1582 = n1581 ^ n1580 ;
  assign n1584 = n1583 ^ n1582 ;
  assign n1578 = x530 ^ x242 ;
  assign n1576 = x536 ^ x248 ;
  assign n1574 = x534 ^ x246 ;
  assign n1573 = x535 ^ x247 ;
  assign n1575 = n1574 ^ n1573 ;
  assign n1577 = n1576 ^ n1575 ;
  assign n1579 = n1578 ^ n1577 ;
  assign n1585 = n1584 ^ n1579 ;
  assign n1556 = x538 ^ x250 ;
  assign n1555 = x539 ^ x251 ;
  assign n1557 = n1556 ^ n1555 ;
  assign n1554 = x540 ^ x252 ;
  assign n1558 = n1557 ^ n1554 ;
  assign n1552 = x537 ^ x249 ;
  assign n1549 = x541 ^ x253 ;
  assign n1548 = x542 ^ x254 ;
  assign n1550 = n1549 ^ n1548 ;
  assign n1547 = x543 ^ x255 ;
  assign n1551 = n1550 ^ n1547 ;
  assign n1553 = n1552 ^ n1551 ;
  assign n1571 = n1558 ^ n1553 ;
  assign n1570 = x529 ^ x241 ;
  assign n1572 = n1571 ^ n1570 ;
  assign n1616 = n1585 ^ n1572 ;
  assign n1618 = n1617 ^ n1616 ;
  assign n1647 = n1646 ^ n1631 ;
  assign n1648 = n1647 ^ n1617 ;
  assign n1649 = n1618 & ~n1648 ;
  assign n1650 = n1649 ^ n1616 ;
  assign n1597 = n1583 ^ n1581 ;
  assign n1598 = n1582 & ~n1597 ;
  assign n1599 = n1598 ^ n1580 ;
  assign n1593 = n1576 ^ n1574 ;
  assign n1594 = n1575 & ~n1593 ;
  assign n1595 = n1594 ^ n1573 ;
  assign n1590 = n1584 ^ n1578 ;
  assign n1591 = n1579 & ~n1590 ;
  assign n1592 = n1591 ^ n1577 ;
  assign n1596 = n1595 ^ n1592 ;
  assign n1600 = n1599 ^ n1596 ;
  assign n1586 = n1585 ^ n1571 ;
  assign n1587 = n1572 & ~n1586 ;
  assign n1588 = n1587 ^ n1570 ;
  assign n1566 = n1555 ^ n1554 ;
  assign n1567 = ~n1557 & n1566 ;
  assign n1568 = n1567 ^ n1554 ;
  assign n1562 = n1548 ^ n1547 ;
  assign n1563 = ~n1550 & n1562 ;
  assign n1564 = n1563 ^ n1547 ;
  assign n1559 = n1558 ^ n1552 ;
  assign n1560 = n1553 & ~n1559 ;
  assign n1561 = n1560 ^ n1551 ;
  assign n1565 = n1564 ^ n1561 ;
  assign n1569 = n1568 ^ n1565 ;
  assign n1589 = n1588 ^ n1569 ;
  assign n1615 = n1600 ^ n1589 ;
  assign n1651 = n1650 ^ n1615 ;
  assign n1678 = n1677 ^ n1662 ;
  assign n1679 = n1678 ^ n1615 ;
  assign n1680 = n1651 & ~n1679 ;
  assign n1681 = n1680 ^ n1650 ;
  assign n1608 = n1599 ^ n1595 ;
  assign n1609 = n1596 & ~n1608 ;
  assign n1610 = n1609 ^ n1592 ;
  assign n1604 = n1568 ^ n1564 ;
  assign n1605 = n1565 & ~n1604 ;
  assign n1606 = n1605 ^ n1561 ;
  assign n1601 = n1600 ^ n1588 ;
  assign n1602 = n1589 & ~n1601 ;
  assign n1603 = n1602 ^ n1569 ;
  assign n1607 = n1606 ^ n1603 ;
  assign n1614 = n1610 ^ n1607 ;
  assign n1682 = n1681 ^ n1614 ;
  assign n1693 = n1692 ^ n1685 ;
  assign n1694 = n1693 ^ n1681 ;
  assign n1695 = n1682 & ~n1694 ;
  assign n1696 = n1695 ^ n1614 ;
  assign n1611 = n1610 ^ n1606 ;
  assign n1612 = n1607 & ~n1611 ;
  assign n1613 = n1612 ^ n1603 ;
  assign n1697 = n1696 ^ n1613 ;
  assign n1701 = n1700 ^ n1697 ;
  assign n1702 = n1678 ^ n1651 ;
  assign n1703 = n1647 ^ n1618 ;
  assign n1704 = x512 ^ x224 ;
  assign n1705 = n1703 & n1704 ;
  assign n1706 = n1702 & n1705 ;
  assign n1707 = n1693 ^ n1682 ;
  assign n1708 = n1706 & n1707 ;
  assign n1709 = n1701 & n1708 ;
  assign n1710 = n1700 ^ n1696 ;
  assign n1711 = n1697 & ~n1710 ;
  assign n1712 = n1711 ^ n1613 ;
  assign n1713 = n1709 & n1712 ;
  assign n1812 = x514 ^ x258 ;
  assign n1809 = x522 ^ x266 ;
  assign n1807 = x528 ^ x272 ;
  assign n1805 = x526 ^ x270 ;
  assign n1804 = x527 ^ x271 ;
  assign n1806 = n1805 ^ n1804 ;
  assign n1808 = n1807 ^ n1806 ;
  assign n1810 = n1809 ^ n1808 ;
  assign n1802 = x525 ^ x269 ;
  assign n1800 = x523 ^ x267 ;
  assign n1799 = x524 ^ x268 ;
  assign n1801 = n1800 ^ n1799 ;
  assign n1803 = n1802 ^ n1801 ;
  assign n1811 = n1810 ^ n1803 ;
  assign n1813 = n1812 ^ n1811 ;
  assign n1796 = x515 ^ x259 ;
  assign n1794 = x521 ^ x265 ;
  assign n1792 = x519 ^ x263 ;
  assign n1791 = x520 ^ x264 ;
  assign n1793 = n1792 ^ n1791 ;
  assign n1795 = n1794 ^ n1793 ;
  assign n1797 = n1796 ^ n1795 ;
  assign n1789 = x518 ^ x262 ;
  assign n1787 = x516 ^ x260 ;
  assign n1786 = x517 ^ x261 ;
  assign n1788 = n1787 ^ n1786 ;
  assign n1790 = n1789 ^ n1788 ;
  assign n1798 = n1797 ^ n1790 ;
  assign n1841 = n1812 ^ n1798 ;
  assign n1842 = n1813 & ~n1841 ;
  assign n1843 = n1842 ^ n1811 ;
  assign n1837 = n1802 ^ n1800 ;
  assign n1838 = n1801 & ~n1837 ;
  assign n1839 = n1838 ^ n1799 ;
  assign n1833 = n1807 ^ n1805 ;
  assign n1834 = n1806 & ~n1833 ;
  assign n1835 = n1834 ^ n1804 ;
  assign n1830 = n1808 ^ n1803 ;
  assign n1831 = ~n1810 & n1830 ;
  assign n1832 = n1831 ^ n1803 ;
  assign n1836 = n1835 ^ n1832 ;
  assign n1840 = n1839 ^ n1836 ;
  assign n1844 = n1843 ^ n1840 ;
  assign n1826 = n1789 ^ n1787 ;
  assign n1827 = n1788 & ~n1826 ;
  assign n1828 = n1827 ^ n1786 ;
  assign n1822 = n1795 ^ n1790 ;
  assign n1823 = ~n1797 & n1822 ;
  assign n1824 = n1823 ^ n1790 ;
  assign n1819 = n1794 ^ n1792 ;
  assign n1820 = n1793 & ~n1819 ;
  assign n1821 = n1820 ^ n1791 ;
  assign n1825 = n1824 ^ n1821 ;
  assign n1829 = n1828 ^ n1825 ;
  assign n1856 = n1843 ^ n1829 ;
  assign n1857 = n1844 & ~n1856 ;
  assign n1858 = n1857 ^ n1840 ;
  assign n1853 = n1839 ^ n1835 ;
  assign n1854 = n1836 & ~n1853 ;
  assign n1855 = n1854 ^ n1832 ;
  assign n1859 = n1858 ^ n1855 ;
  assign n1850 = n1828 ^ n1824 ;
  assign n1851 = n1825 & ~n1850 ;
  assign n1852 = n1851 ^ n1821 ;
  assign n1865 = n1855 ^ n1852 ;
  assign n1866 = ~n1859 & n1865 ;
  assign n1867 = n1866 ^ n1852 ;
  assign n1784 = x513 ^ x257 ;
  assign n1750 = x533 ^ x277 ;
  assign n1748 = x531 ^ x275 ;
  assign n1747 = x532 ^ x276 ;
  assign n1749 = n1748 ^ n1747 ;
  assign n1751 = n1750 ^ n1749 ;
  assign n1745 = x530 ^ x274 ;
  assign n1743 = x536 ^ x280 ;
  assign n1741 = x534 ^ x278 ;
  assign n1740 = x535 ^ x279 ;
  assign n1742 = n1741 ^ n1740 ;
  assign n1744 = n1743 ^ n1742 ;
  assign n1746 = n1745 ^ n1744 ;
  assign n1752 = n1751 ^ n1746 ;
  assign n1723 = x538 ^ x282 ;
  assign n1722 = x539 ^ x283 ;
  assign n1724 = n1723 ^ n1722 ;
  assign n1721 = x540 ^ x284 ;
  assign n1725 = n1724 ^ n1721 ;
  assign n1719 = x537 ^ x281 ;
  assign n1716 = x541 ^ x285 ;
  assign n1715 = x542 ^ x286 ;
  assign n1717 = n1716 ^ n1715 ;
  assign n1714 = x543 ^ x287 ;
  assign n1718 = n1717 ^ n1714 ;
  assign n1720 = n1719 ^ n1718 ;
  assign n1738 = n1725 ^ n1720 ;
  assign n1737 = x529 ^ x273 ;
  assign n1739 = n1738 ^ n1737 ;
  assign n1783 = n1752 ^ n1739 ;
  assign n1785 = n1784 ^ n1783 ;
  assign n1814 = n1813 ^ n1798 ;
  assign n1815 = n1814 ^ n1784 ;
  assign n1816 = n1785 & ~n1815 ;
  assign n1817 = n1816 ^ n1783 ;
  assign n1764 = n1750 ^ n1748 ;
  assign n1765 = n1749 & ~n1764 ;
  assign n1766 = n1765 ^ n1747 ;
  assign n1760 = n1743 ^ n1741 ;
  assign n1761 = n1742 & ~n1760 ;
  assign n1762 = n1761 ^ n1740 ;
  assign n1757 = n1751 ^ n1745 ;
  assign n1758 = n1746 & ~n1757 ;
  assign n1759 = n1758 ^ n1744 ;
  assign n1763 = n1762 ^ n1759 ;
  assign n1767 = n1766 ^ n1763 ;
  assign n1753 = n1752 ^ n1738 ;
  assign n1754 = n1739 & ~n1753 ;
  assign n1755 = n1754 ^ n1737 ;
  assign n1733 = n1722 ^ n1721 ;
  assign n1734 = ~n1724 & n1733 ;
  assign n1735 = n1734 ^ n1721 ;
  assign n1729 = n1715 ^ n1714 ;
  assign n1730 = ~n1717 & n1729 ;
  assign n1731 = n1730 ^ n1714 ;
  assign n1726 = n1725 ^ n1719 ;
  assign n1727 = n1720 & ~n1726 ;
  assign n1728 = n1727 ^ n1718 ;
  assign n1732 = n1731 ^ n1728 ;
  assign n1736 = n1735 ^ n1732 ;
  assign n1756 = n1755 ^ n1736 ;
  assign n1782 = n1767 ^ n1756 ;
  assign n1818 = n1817 ^ n1782 ;
  assign n1845 = n1844 ^ n1829 ;
  assign n1846 = n1845 ^ n1782 ;
  assign n1847 = n1818 & ~n1846 ;
  assign n1848 = n1847 ^ n1817 ;
  assign n1775 = n1766 ^ n1762 ;
  assign n1776 = n1763 & ~n1775 ;
  assign n1777 = n1776 ^ n1759 ;
  assign n1771 = n1735 ^ n1731 ;
  assign n1772 = n1732 & ~n1771 ;
  assign n1773 = n1772 ^ n1728 ;
  assign n1768 = n1767 ^ n1755 ;
  assign n1769 = n1756 & ~n1768 ;
  assign n1770 = n1769 ^ n1736 ;
  assign n1774 = n1773 ^ n1770 ;
  assign n1781 = n1777 ^ n1774 ;
  assign n1849 = n1848 ^ n1781 ;
  assign n1860 = n1859 ^ n1852 ;
  assign n1861 = n1860 ^ n1848 ;
  assign n1862 = n1849 & ~n1861 ;
  assign n1863 = n1862 ^ n1781 ;
  assign n1778 = n1777 ^ n1773 ;
  assign n1779 = n1774 & ~n1778 ;
  assign n1780 = n1779 ^ n1770 ;
  assign n1864 = n1863 ^ n1780 ;
  assign n1868 = n1867 ^ n1864 ;
  assign n1869 = n1845 ^ n1818 ;
  assign n1870 = n1814 ^ n1785 ;
  assign n1871 = x512 ^ x256 ;
  assign n1872 = n1870 & n1871 ;
  assign n1873 = n1869 & n1872 ;
  assign n1874 = n1860 ^ n1849 ;
  assign n1875 = n1873 & n1874 ;
  assign n1876 = n1868 & n1875 ;
  assign n1877 = n1867 ^ n1863 ;
  assign n1878 = n1864 & ~n1877 ;
  assign n1879 = n1878 ^ n1780 ;
  assign n1880 = n1876 & n1879 ;
  assign n1979 = x514 ^ x290 ;
  assign n1976 = x522 ^ x298 ;
  assign n1974 = x528 ^ x304 ;
  assign n1972 = x526 ^ x302 ;
  assign n1971 = x527 ^ x303 ;
  assign n1973 = n1972 ^ n1971 ;
  assign n1975 = n1974 ^ n1973 ;
  assign n1977 = n1976 ^ n1975 ;
  assign n1969 = x525 ^ x301 ;
  assign n1967 = x523 ^ x299 ;
  assign n1966 = x524 ^ x300 ;
  assign n1968 = n1967 ^ n1966 ;
  assign n1970 = n1969 ^ n1968 ;
  assign n1978 = n1977 ^ n1970 ;
  assign n1980 = n1979 ^ n1978 ;
  assign n1963 = x515 ^ x291 ;
  assign n1961 = x521 ^ x297 ;
  assign n1959 = x519 ^ x295 ;
  assign n1958 = x520 ^ x296 ;
  assign n1960 = n1959 ^ n1958 ;
  assign n1962 = n1961 ^ n1960 ;
  assign n1964 = n1963 ^ n1962 ;
  assign n1956 = x518 ^ x294 ;
  assign n1954 = x516 ^ x292 ;
  assign n1953 = x517 ^ x293 ;
  assign n1955 = n1954 ^ n1953 ;
  assign n1957 = n1956 ^ n1955 ;
  assign n1965 = n1964 ^ n1957 ;
  assign n2008 = n1979 ^ n1965 ;
  assign n2009 = n1980 & ~n2008 ;
  assign n2010 = n2009 ^ n1978 ;
  assign n2004 = n1969 ^ n1967 ;
  assign n2005 = n1968 & ~n2004 ;
  assign n2006 = n2005 ^ n1966 ;
  assign n2000 = n1974 ^ n1972 ;
  assign n2001 = n1973 & ~n2000 ;
  assign n2002 = n2001 ^ n1971 ;
  assign n1997 = n1975 ^ n1970 ;
  assign n1998 = ~n1977 & n1997 ;
  assign n1999 = n1998 ^ n1970 ;
  assign n2003 = n2002 ^ n1999 ;
  assign n2007 = n2006 ^ n2003 ;
  assign n2011 = n2010 ^ n2007 ;
  assign n1993 = n1956 ^ n1954 ;
  assign n1994 = n1955 & ~n1993 ;
  assign n1995 = n1994 ^ n1953 ;
  assign n1989 = n1962 ^ n1957 ;
  assign n1990 = ~n1964 & n1989 ;
  assign n1991 = n1990 ^ n1957 ;
  assign n1986 = n1961 ^ n1959 ;
  assign n1987 = n1960 & ~n1986 ;
  assign n1988 = n1987 ^ n1958 ;
  assign n1992 = n1991 ^ n1988 ;
  assign n1996 = n1995 ^ n1992 ;
  assign n2023 = n2010 ^ n1996 ;
  assign n2024 = n2011 & ~n2023 ;
  assign n2025 = n2024 ^ n2007 ;
  assign n2020 = n2006 ^ n2002 ;
  assign n2021 = n2003 & ~n2020 ;
  assign n2022 = n2021 ^ n1999 ;
  assign n2026 = n2025 ^ n2022 ;
  assign n2017 = n1995 ^ n1991 ;
  assign n2018 = n1992 & ~n2017 ;
  assign n2019 = n2018 ^ n1988 ;
  assign n2032 = n2022 ^ n2019 ;
  assign n2033 = ~n2026 & n2032 ;
  assign n2034 = n2033 ^ n2019 ;
  assign n1951 = x513 ^ x289 ;
  assign n1917 = x533 ^ x309 ;
  assign n1915 = x531 ^ x307 ;
  assign n1914 = x532 ^ x308 ;
  assign n1916 = n1915 ^ n1914 ;
  assign n1918 = n1917 ^ n1916 ;
  assign n1912 = x530 ^ x306 ;
  assign n1910 = x536 ^ x312 ;
  assign n1908 = x534 ^ x310 ;
  assign n1907 = x535 ^ x311 ;
  assign n1909 = n1908 ^ n1907 ;
  assign n1911 = n1910 ^ n1909 ;
  assign n1913 = n1912 ^ n1911 ;
  assign n1919 = n1918 ^ n1913 ;
  assign n1890 = x538 ^ x314 ;
  assign n1889 = x539 ^ x315 ;
  assign n1891 = n1890 ^ n1889 ;
  assign n1888 = x540 ^ x316 ;
  assign n1892 = n1891 ^ n1888 ;
  assign n1886 = x537 ^ x313 ;
  assign n1883 = x541 ^ x317 ;
  assign n1882 = x542 ^ x318 ;
  assign n1884 = n1883 ^ n1882 ;
  assign n1881 = x543 ^ x319 ;
  assign n1885 = n1884 ^ n1881 ;
  assign n1887 = n1886 ^ n1885 ;
  assign n1905 = n1892 ^ n1887 ;
  assign n1904 = x529 ^ x305 ;
  assign n1906 = n1905 ^ n1904 ;
  assign n1950 = n1919 ^ n1906 ;
  assign n1952 = n1951 ^ n1950 ;
  assign n1981 = n1980 ^ n1965 ;
  assign n1982 = n1981 ^ n1951 ;
  assign n1983 = n1952 & ~n1982 ;
  assign n1984 = n1983 ^ n1950 ;
  assign n1931 = n1917 ^ n1915 ;
  assign n1932 = n1916 & ~n1931 ;
  assign n1933 = n1932 ^ n1914 ;
  assign n1927 = n1910 ^ n1908 ;
  assign n1928 = n1909 & ~n1927 ;
  assign n1929 = n1928 ^ n1907 ;
  assign n1924 = n1918 ^ n1912 ;
  assign n1925 = n1913 & ~n1924 ;
  assign n1926 = n1925 ^ n1911 ;
  assign n1930 = n1929 ^ n1926 ;
  assign n1934 = n1933 ^ n1930 ;
  assign n1920 = n1919 ^ n1905 ;
  assign n1921 = n1906 & ~n1920 ;
  assign n1922 = n1921 ^ n1904 ;
  assign n1900 = n1889 ^ n1888 ;
  assign n1901 = ~n1891 & n1900 ;
  assign n1902 = n1901 ^ n1888 ;
  assign n1896 = n1882 ^ n1881 ;
  assign n1897 = ~n1884 & n1896 ;
  assign n1898 = n1897 ^ n1881 ;
  assign n1893 = n1892 ^ n1886 ;
  assign n1894 = n1887 & ~n1893 ;
  assign n1895 = n1894 ^ n1885 ;
  assign n1899 = n1898 ^ n1895 ;
  assign n1903 = n1902 ^ n1899 ;
  assign n1923 = n1922 ^ n1903 ;
  assign n1949 = n1934 ^ n1923 ;
  assign n1985 = n1984 ^ n1949 ;
  assign n2012 = n2011 ^ n1996 ;
  assign n2013 = n2012 ^ n1949 ;
  assign n2014 = n1985 & ~n2013 ;
  assign n2015 = n2014 ^ n1984 ;
  assign n1942 = n1933 ^ n1929 ;
  assign n1943 = n1930 & ~n1942 ;
  assign n1944 = n1943 ^ n1926 ;
  assign n1938 = n1902 ^ n1898 ;
  assign n1939 = n1899 & ~n1938 ;
  assign n1940 = n1939 ^ n1895 ;
  assign n1935 = n1934 ^ n1922 ;
  assign n1936 = n1923 & ~n1935 ;
  assign n1937 = n1936 ^ n1903 ;
  assign n1941 = n1940 ^ n1937 ;
  assign n1948 = n1944 ^ n1941 ;
  assign n2016 = n2015 ^ n1948 ;
  assign n2027 = n2026 ^ n2019 ;
  assign n2028 = n2027 ^ n2015 ;
  assign n2029 = n2016 & ~n2028 ;
  assign n2030 = n2029 ^ n1948 ;
  assign n1945 = n1944 ^ n1940 ;
  assign n1946 = n1941 & ~n1945 ;
  assign n1947 = n1946 ^ n1937 ;
  assign n2031 = n2030 ^ n1947 ;
  assign n2035 = n2034 ^ n2031 ;
  assign n2036 = n2012 ^ n1985 ;
  assign n2037 = n1981 ^ n1952 ;
  assign n2038 = x512 ^ x288 ;
  assign n2039 = n2037 & n2038 ;
  assign n2040 = n2036 & n2039 ;
  assign n2041 = n2027 ^ n2016 ;
  assign n2042 = n2040 & n2041 ;
  assign n2043 = n2035 & n2042 ;
  assign n2044 = n2034 ^ n2030 ;
  assign n2045 = n2031 & ~n2044 ;
  assign n2046 = n2045 ^ n1947 ;
  assign n2047 = n2043 & n2046 ;
  assign n2146 = x514 ^ x322 ;
  assign n2143 = x522 ^ x330 ;
  assign n2141 = x528 ^ x336 ;
  assign n2139 = x526 ^ x334 ;
  assign n2138 = x527 ^ x335 ;
  assign n2140 = n2139 ^ n2138 ;
  assign n2142 = n2141 ^ n2140 ;
  assign n2144 = n2143 ^ n2142 ;
  assign n2136 = x525 ^ x333 ;
  assign n2134 = x523 ^ x331 ;
  assign n2133 = x524 ^ x332 ;
  assign n2135 = n2134 ^ n2133 ;
  assign n2137 = n2136 ^ n2135 ;
  assign n2145 = n2144 ^ n2137 ;
  assign n2147 = n2146 ^ n2145 ;
  assign n2130 = x515 ^ x323 ;
  assign n2128 = x521 ^ x329 ;
  assign n2126 = x519 ^ x327 ;
  assign n2125 = x520 ^ x328 ;
  assign n2127 = n2126 ^ n2125 ;
  assign n2129 = n2128 ^ n2127 ;
  assign n2131 = n2130 ^ n2129 ;
  assign n2123 = x518 ^ x326 ;
  assign n2121 = x516 ^ x324 ;
  assign n2120 = x517 ^ x325 ;
  assign n2122 = n2121 ^ n2120 ;
  assign n2124 = n2123 ^ n2122 ;
  assign n2132 = n2131 ^ n2124 ;
  assign n2175 = n2146 ^ n2132 ;
  assign n2176 = n2147 & ~n2175 ;
  assign n2177 = n2176 ^ n2145 ;
  assign n2171 = n2136 ^ n2134 ;
  assign n2172 = n2135 & ~n2171 ;
  assign n2173 = n2172 ^ n2133 ;
  assign n2167 = n2141 ^ n2139 ;
  assign n2168 = n2140 & ~n2167 ;
  assign n2169 = n2168 ^ n2138 ;
  assign n2164 = n2142 ^ n2137 ;
  assign n2165 = ~n2144 & n2164 ;
  assign n2166 = n2165 ^ n2137 ;
  assign n2170 = n2169 ^ n2166 ;
  assign n2174 = n2173 ^ n2170 ;
  assign n2178 = n2177 ^ n2174 ;
  assign n2160 = n2123 ^ n2121 ;
  assign n2161 = n2122 & ~n2160 ;
  assign n2162 = n2161 ^ n2120 ;
  assign n2156 = n2129 ^ n2124 ;
  assign n2157 = ~n2131 & n2156 ;
  assign n2158 = n2157 ^ n2124 ;
  assign n2153 = n2128 ^ n2126 ;
  assign n2154 = n2127 & ~n2153 ;
  assign n2155 = n2154 ^ n2125 ;
  assign n2159 = n2158 ^ n2155 ;
  assign n2163 = n2162 ^ n2159 ;
  assign n2190 = n2177 ^ n2163 ;
  assign n2191 = n2178 & ~n2190 ;
  assign n2192 = n2191 ^ n2174 ;
  assign n2187 = n2173 ^ n2169 ;
  assign n2188 = n2170 & ~n2187 ;
  assign n2189 = n2188 ^ n2166 ;
  assign n2193 = n2192 ^ n2189 ;
  assign n2184 = n2162 ^ n2158 ;
  assign n2185 = n2159 & ~n2184 ;
  assign n2186 = n2185 ^ n2155 ;
  assign n2199 = n2189 ^ n2186 ;
  assign n2200 = ~n2193 & n2199 ;
  assign n2201 = n2200 ^ n2186 ;
  assign n2118 = x513 ^ x321 ;
  assign n2084 = x533 ^ x341 ;
  assign n2082 = x531 ^ x339 ;
  assign n2081 = x532 ^ x340 ;
  assign n2083 = n2082 ^ n2081 ;
  assign n2085 = n2084 ^ n2083 ;
  assign n2079 = x530 ^ x338 ;
  assign n2077 = x536 ^ x344 ;
  assign n2075 = x534 ^ x342 ;
  assign n2074 = x535 ^ x343 ;
  assign n2076 = n2075 ^ n2074 ;
  assign n2078 = n2077 ^ n2076 ;
  assign n2080 = n2079 ^ n2078 ;
  assign n2086 = n2085 ^ n2080 ;
  assign n2057 = x538 ^ x346 ;
  assign n2056 = x539 ^ x347 ;
  assign n2058 = n2057 ^ n2056 ;
  assign n2055 = x540 ^ x348 ;
  assign n2059 = n2058 ^ n2055 ;
  assign n2053 = x537 ^ x345 ;
  assign n2050 = x541 ^ x349 ;
  assign n2049 = x542 ^ x350 ;
  assign n2051 = n2050 ^ n2049 ;
  assign n2048 = x543 ^ x351 ;
  assign n2052 = n2051 ^ n2048 ;
  assign n2054 = n2053 ^ n2052 ;
  assign n2072 = n2059 ^ n2054 ;
  assign n2071 = x529 ^ x337 ;
  assign n2073 = n2072 ^ n2071 ;
  assign n2117 = n2086 ^ n2073 ;
  assign n2119 = n2118 ^ n2117 ;
  assign n2148 = n2147 ^ n2132 ;
  assign n2149 = n2148 ^ n2118 ;
  assign n2150 = n2119 & ~n2149 ;
  assign n2151 = n2150 ^ n2117 ;
  assign n2098 = n2084 ^ n2082 ;
  assign n2099 = n2083 & ~n2098 ;
  assign n2100 = n2099 ^ n2081 ;
  assign n2094 = n2077 ^ n2075 ;
  assign n2095 = n2076 & ~n2094 ;
  assign n2096 = n2095 ^ n2074 ;
  assign n2091 = n2085 ^ n2079 ;
  assign n2092 = n2080 & ~n2091 ;
  assign n2093 = n2092 ^ n2078 ;
  assign n2097 = n2096 ^ n2093 ;
  assign n2101 = n2100 ^ n2097 ;
  assign n2087 = n2086 ^ n2072 ;
  assign n2088 = n2073 & ~n2087 ;
  assign n2089 = n2088 ^ n2071 ;
  assign n2067 = n2056 ^ n2055 ;
  assign n2068 = ~n2058 & n2067 ;
  assign n2069 = n2068 ^ n2055 ;
  assign n2063 = n2049 ^ n2048 ;
  assign n2064 = ~n2051 & n2063 ;
  assign n2065 = n2064 ^ n2048 ;
  assign n2060 = n2059 ^ n2053 ;
  assign n2061 = n2054 & ~n2060 ;
  assign n2062 = n2061 ^ n2052 ;
  assign n2066 = n2065 ^ n2062 ;
  assign n2070 = n2069 ^ n2066 ;
  assign n2090 = n2089 ^ n2070 ;
  assign n2116 = n2101 ^ n2090 ;
  assign n2152 = n2151 ^ n2116 ;
  assign n2179 = n2178 ^ n2163 ;
  assign n2180 = n2179 ^ n2116 ;
  assign n2181 = n2152 & ~n2180 ;
  assign n2182 = n2181 ^ n2151 ;
  assign n2109 = n2100 ^ n2096 ;
  assign n2110 = n2097 & ~n2109 ;
  assign n2111 = n2110 ^ n2093 ;
  assign n2105 = n2069 ^ n2065 ;
  assign n2106 = n2066 & ~n2105 ;
  assign n2107 = n2106 ^ n2062 ;
  assign n2102 = n2101 ^ n2089 ;
  assign n2103 = n2090 & ~n2102 ;
  assign n2104 = n2103 ^ n2070 ;
  assign n2108 = n2107 ^ n2104 ;
  assign n2115 = n2111 ^ n2108 ;
  assign n2183 = n2182 ^ n2115 ;
  assign n2194 = n2193 ^ n2186 ;
  assign n2195 = n2194 ^ n2182 ;
  assign n2196 = n2183 & ~n2195 ;
  assign n2197 = n2196 ^ n2115 ;
  assign n2112 = n2111 ^ n2107 ;
  assign n2113 = n2108 & ~n2112 ;
  assign n2114 = n2113 ^ n2104 ;
  assign n2198 = n2197 ^ n2114 ;
  assign n2202 = n2201 ^ n2198 ;
  assign n2203 = n2179 ^ n2152 ;
  assign n2204 = n2148 ^ n2119 ;
  assign n2205 = x512 ^ x320 ;
  assign n2206 = n2204 & n2205 ;
  assign n2207 = n2203 & n2206 ;
  assign n2208 = n2194 ^ n2183 ;
  assign n2209 = n2207 & n2208 ;
  assign n2210 = n2202 & n2209 ;
  assign n2211 = n2201 ^ n2197 ;
  assign n2212 = n2198 & ~n2211 ;
  assign n2213 = n2212 ^ n2114 ;
  assign n2214 = n2210 & n2213 ;
  assign n2313 = x514 ^ x354 ;
  assign n2310 = x522 ^ x362 ;
  assign n2308 = x528 ^ x368 ;
  assign n2306 = x526 ^ x366 ;
  assign n2305 = x527 ^ x367 ;
  assign n2307 = n2306 ^ n2305 ;
  assign n2309 = n2308 ^ n2307 ;
  assign n2311 = n2310 ^ n2309 ;
  assign n2303 = x525 ^ x365 ;
  assign n2301 = x523 ^ x363 ;
  assign n2300 = x524 ^ x364 ;
  assign n2302 = n2301 ^ n2300 ;
  assign n2304 = n2303 ^ n2302 ;
  assign n2312 = n2311 ^ n2304 ;
  assign n2314 = n2313 ^ n2312 ;
  assign n2297 = x515 ^ x355 ;
  assign n2295 = x521 ^ x361 ;
  assign n2293 = x519 ^ x359 ;
  assign n2292 = x520 ^ x360 ;
  assign n2294 = n2293 ^ n2292 ;
  assign n2296 = n2295 ^ n2294 ;
  assign n2298 = n2297 ^ n2296 ;
  assign n2290 = x518 ^ x358 ;
  assign n2288 = x516 ^ x356 ;
  assign n2287 = x517 ^ x357 ;
  assign n2289 = n2288 ^ n2287 ;
  assign n2291 = n2290 ^ n2289 ;
  assign n2299 = n2298 ^ n2291 ;
  assign n2342 = n2313 ^ n2299 ;
  assign n2343 = n2314 & ~n2342 ;
  assign n2344 = n2343 ^ n2312 ;
  assign n2338 = n2303 ^ n2301 ;
  assign n2339 = n2302 & ~n2338 ;
  assign n2340 = n2339 ^ n2300 ;
  assign n2334 = n2308 ^ n2306 ;
  assign n2335 = n2307 & ~n2334 ;
  assign n2336 = n2335 ^ n2305 ;
  assign n2331 = n2309 ^ n2304 ;
  assign n2332 = ~n2311 & n2331 ;
  assign n2333 = n2332 ^ n2304 ;
  assign n2337 = n2336 ^ n2333 ;
  assign n2341 = n2340 ^ n2337 ;
  assign n2345 = n2344 ^ n2341 ;
  assign n2327 = n2290 ^ n2288 ;
  assign n2328 = n2289 & ~n2327 ;
  assign n2329 = n2328 ^ n2287 ;
  assign n2323 = n2296 ^ n2291 ;
  assign n2324 = ~n2298 & n2323 ;
  assign n2325 = n2324 ^ n2291 ;
  assign n2320 = n2295 ^ n2293 ;
  assign n2321 = n2294 & ~n2320 ;
  assign n2322 = n2321 ^ n2292 ;
  assign n2326 = n2325 ^ n2322 ;
  assign n2330 = n2329 ^ n2326 ;
  assign n2357 = n2344 ^ n2330 ;
  assign n2358 = n2345 & ~n2357 ;
  assign n2359 = n2358 ^ n2341 ;
  assign n2354 = n2340 ^ n2336 ;
  assign n2355 = n2337 & ~n2354 ;
  assign n2356 = n2355 ^ n2333 ;
  assign n2360 = n2359 ^ n2356 ;
  assign n2351 = n2329 ^ n2325 ;
  assign n2352 = n2326 & ~n2351 ;
  assign n2353 = n2352 ^ n2322 ;
  assign n2366 = n2356 ^ n2353 ;
  assign n2367 = ~n2360 & n2366 ;
  assign n2368 = n2367 ^ n2353 ;
  assign n2285 = x513 ^ x353 ;
  assign n2251 = x533 ^ x373 ;
  assign n2249 = x531 ^ x371 ;
  assign n2248 = x532 ^ x372 ;
  assign n2250 = n2249 ^ n2248 ;
  assign n2252 = n2251 ^ n2250 ;
  assign n2246 = x530 ^ x370 ;
  assign n2244 = x536 ^ x376 ;
  assign n2242 = x534 ^ x374 ;
  assign n2241 = x535 ^ x375 ;
  assign n2243 = n2242 ^ n2241 ;
  assign n2245 = n2244 ^ n2243 ;
  assign n2247 = n2246 ^ n2245 ;
  assign n2253 = n2252 ^ n2247 ;
  assign n2224 = x538 ^ x378 ;
  assign n2223 = x539 ^ x379 ;
  assign n2225 = n2224 ^ n2223 ;
  assign n2222 = x540 ^ x380 ;
  assign n2226 = n2225 ^ n2222 ;
  assign n2220 = x537 ^ x377 ;
  assign n2217 = x541 ^ x381 ;
  assign n2216 = x542 ^ x382 ;
  assign n2218 = n2217 ^ n2216 ;
  assign n2215 = x543 ^ x383 ;
  assign n2219 = n2218 ^ n2215 ;
  assign n2221 = n2220 ^ n2219 ;
  assign n2239 = n2226 ^ n2221 ;
  assign n2238 = x529 ^ x369 ;
  assign n2240 = n2239 ^ n2238 ;
  assign n2284 = n2253 ^ n2240 ;
  assign n2286 = n2285 ^ n2284 ;
  assign n2315 = n2314 ^ n2299 ;
  assign n2316 = n2315 ^ n2285 ;
  assign n2317 = n2286 & ~n2316 ;
  assign n2318 = n2317 ^ n2284 ;
  assign n2265 = n2251 ^ n2249 ;
  assign n2266 = n2250 & ~n2265 ;
  assign n2267 = n2266 ^ n2248 ;
  assign n2261 = n2244 ^ n2242 ;
  assign n2262 = n2243 & ~n2261 ;
  assign n2263 = n2262 ^ n2241 ;
  assign n2258 = n2252 ^ n2246 ;
  assign n2259 = n2247 & ~n2258 ;
  assign n2260 = n2259 ^ n2245 ;
  assign n2264 = n2263 ^ n2260 ;
  assign n2268 = n2267 ^ n2264 ;
  assign n2254 = n2253 ^ n2239 ;
  assign n2255 = n2240 & ~n2254 ;
  assign n2256 = n2255 ^ n2238 ;
  assign n2234 = n2223 ^ n2222 ;
  assign n2235 = ~n2225 & n2234 ;
  assign n2236 = n2235 ^ n2222 ;
  assign n2230 = n2216 ^ n2215 ;
  assign n2231 = ~n2218 & n2230 ;
  assign n2232 = n2231 ^ n2215 ;
  assign n2227 = n2226 ^ n2220 ;
  assign n2228 = n2221 & ~n2227 ;
  assign n2229 = n2228 ^ n2219 ;
  assign n2233 = n2232 ^ n2229 ;
  assign n2237 = n2236 ^ n2233 ;
  assign n2257 = n2256 ^ n2237 ;
  assign n2283 = n2268 ^ n2257 ;
  assign n2319 = n2318 ^ n2283 ;
  assign n2346 = n2345 ^ n2330 ;
  assign n2347 = n2346 ^ n2283 ;
  assign n2348 = n2319 & ~n2347 ;
  assign n2349 = n2348 ^ n2318 ;
  assign n2276 = n2267 ^ n2263 ;
  assign n2277 = n2264 & ~n2276 ;
  assign n2278 = n2277 ^ n2260 ;
  assign n2272 = n2236 ^ n2232 ;
  assign n2273 = n2233 & ~n2272 ;
  assign n2274 = n2273 ^ n2229 ;
  assign n2269 = n2268 ^ n2256 ;
  assign n2270 = n2257 & ~n2269 ;
  assign n2271 = n2270 ^ n2237 ;
  assign n2275 = n2274 ^ n2271 ;
  assign n2282 = n2278 ^ n2275 ;
  assign n2350 = n2349 ^ n2282 ;
  assign n2361 = n2360 ^ n2353 ;
  assign n2362 = n2361 ^ n2349 ;
  assign n2363 = n2350 & ~n2362 ;
  assign n2364 = n2363 ^ n2282 ;
  assign n2279 = n2278 ^ n2274 ;
  assign n2280 = n2275 & ~n2279 ;
  assign n2281 = n2280 ^ n2271 ;
  assign n2365 = n2364 ^ n2281 ;
  assign n2369 = n2368 ^ n2365 ;
  assign n2370 = n2346 ^ n2319 ;
  assign n2371 = n2315 ^ n2286 ;
  assign n2372 = x512 ^ x352 ;
  assign n2373 = n2371 & n2372 ;
  assign n2374 = n2370 & n2373 ;
  assign n2375 = n2361 ^ n2350 ;
  assign n2376 = n2374 & n2375 ;
  assign n2377 = n2369 & n2376 ;
  assign n2378 = n2368 ^ n2364 ;
  assign n2379 = n2365 & ~n2378 ;
  assign n2380 = n2379 ^ n2281 ;
  assign n2381 = n2377 & n2380 ;
  assign n2480 = x514 ^ x418 ;
  assign n2477 = x522 ^ x426 ;
  assign n2475 = x528 ^ x432 ;
  assign n2473 = x526 ^ x430 ;
  assign n2472 = x527 ^ x431 ;
  assign n2474 = n2473 ^ n2472 ;
  assign n2476 = n2475 ^ n2474 ;
  assign n2478 = n2477 ^ n2476 ;
  assign n2470 = x525 ^ x429 ;
  assign n2468 = x523 ^ x427 ;
  assign n2467 = x524 ^ x428 ;
  assign n2469 = n2468 ^ n2467 ;
  assign n2471 = n2470 ^ n2469 ;
  assign n2479 = n2478 ^ n2471 ;
  assign n2481 = n2480 ^ n2479 ;
  assign n2464 = x515 ^ x419 ;
  assign n2462 = x521 ^ x425 ;
  assign n2460 = x519 ^ x423 ;
  assign n2459 = x520 ^ x424 ;
  assign n2461 = n2460 ^ n2459 ;
  assign n2463 = n2462 ^ n2461 ;
  assign n2465 = n2464 ^ n2463 ;
  assign n2457 = x518 ^ x422 ;
  assign n2455 = x516 ^ x420 ;
  assign n2454 = x517 ^ x421 ;
  assign n2456 = n2455 ^ n2454 ;
  assign n2458 = n2457 ^ n2456 ;
  assign n2466 = n2465 ^ n2458 ;
  assign n2509 = n2480 ^ n2466 ;
  assign n2510 = n2481 & ~n2509 ;
  assign n2511 = n2510 ^ n2479 ;
  assign n2505 = n2470 ^ n2468 ;
  assign n2506 = n2469 & ~n2505 ;
  assign n2507 = n2506 ^ n2467 ;
  assign n2501 = n2475 ^ n2473 ;
  assign n2502 = n2474 & ~n2501 ;
  assign n2503 = n2502 ^ n2472 ;
  assign n2498 = n2476 ^ n2471 ;
  assign n2499 = ~n2478 & n2498 ;
  assign n2500 = n2499 ^ n2471 ;
  assign n2504 = n2503 ^ n2500 ;
  assign n2508 = n2507 ^ n2504 ;
  assign n2512 = n2511 ^ n2508 ;
  assign n2494 = n2457 ^ n2455 ;
  assign n2495 = n2456 & ~n2494 ;
  assign n2496 = n2495 ^ n2454 ;
  assign n2490 = n2463 ^ n2458 ;
  assign n2491 = ~n2465 & n2490 ;
  assign n2492 = n2491 ^ n2458 ;
  assign n2487 = n2462 ^ n2460 ;
  assign n2488 = n2461 & ~n2487 ;
  assign n2489 = n2488 ^ n2459 ;
  assign n2493 = n2492 ^ n2489 ;
  assign n2497 = n2496 ^ n2493 ;
  assign n2524 = n2511 ^ n2497 ;
  assign n2525 = n2512 & ~n2524 ;
  assign n2526 = n2525 ^ n2508 ;
  assign n2521 = n2507 ^ n2503 ;
  assign n2522 = n2504 & ~n2521 ;
  assign n2523 = n2522 ^ n2500 ;
  assign n2527 = n2526 ^ n2523 ;
  assign n2518 = n2496 ^ n2492 ;
  assign n2519 = n2493 & ~n2518 ;
  assign n2520 = n2519 ^ n2489 ;
  assign n2533 = n2523 ^ n2520 ;
  assign n2534 = ~n2527 & n2533 ;
  assign n2535 = n2534 ^ n2520 ;
  assign n2452 = x513 ^ x417 ;
  assign n2418 = x533 ^ x437 ;
  assign n2416 = x531 ^ x435 ;
  assign n2415 = x532 ^ x436 ;
  assign n2417 = n2416 ^ n2415 ;
  assign n2419 = n2418 ^ n2417 ;
  assign n2413 = x530 ^ x434 ;
  assign n2411 = x536 ^ x440 ;
  assign n2409 = x534 ^ x438 ;
  assign n2408 = x535 ^ x439 ;
  assign n2410 = n2409 ^ n2408 ;
  assign n2412 = n2411 ^ n2410 ;
  assign n2414 = n2413 ^ n2412 ;
  assign n2420 = n2419 ^ n2414 ;
  assign n2391 = x538 ^ x442 ;
  assign n2390 = x539 ^ x443 ;
  assign n2392 = n2391 ^ n2390 ;
  assign n2389 = x540 ^ x444 ;
  assign n2393 = n2392 ^ n2389 ;
  assign n2387 = x537 ^ x441 ;
  assign n2384 = x541 ^ x445 ;
  assign n2383 = x542 ^ x446 ;
  assign n2385 = n2384 ^ n2383 ;
  assign n2382 = x543 ^ x447 ;
  assign n2386 = n2385 ^ n2382 ;
  assign n2388 = n2387 ^ n2386 ;
  assign n2406 = n2393 ^ n2388 ;
  assign n2405 = x529 ^ x433 ;
  assign n2407 = n2406 ^ n2405 ;
  assign n2451 = n2420 ^ n2407 ;
  assign n2453 = n2452 ^ n2451 ;
  assign n2482 = n2481 ^ n2466 ;
  assign n2483 = n2482 ^ n2452 ;
  assign n2484 = n2453 & ~n2483 ;
  assign n2485 = n2484 ^ n2451 ;
  assign n2432 = n2418 ^ n2416 ;
  assign n2433 = n2417 & ~n2432 ;
  assign n2434 = n2433 ^ n2415 ;
  assign n2428 = n2411 ^ n2409 ;
  assign n2429 = n2410 & ~n2428 ;
  assign n2430 = n2429 ^ n2408 ;
  assign n2425 = n2419 ^ n2413 ;
  assign n2426 = n2414 & ~n2425 ;
  assign n2427 = n2426 ^ n2412 ;
  assign n2431 = n2430 ^ n2427 ;
  assign n2435 = n2434 ^ n2431 ;
  assign n2421 = n2420 ^ n2406 ;
  assign n2422 = n2407 & ~n2421 ;
  assign n2423 = n2422 ^ n2405 ;
  assign n2401 = n2390 ^ n2389 ;
  assign n2402 = ~n2392 & n2401 ;
  assign n2403 = n2402 ^ n2389 ;
  assign n2397 = n2383 ^ n2382 ;
  assign n2398 = ~n2385 & n2397 ;
  assign n2399 = n2398 ^ n2382 ;
  assign n2394 = n2393 ^ n2387 ;
  assign n2395 = n2388 & ~n2394 ;
  assign n2396 = n2395 ^ n2386 ;
  assign n2400 = n2399 ^ n2396 ;
  assign n2404 = n2403 ^ n2400 ;
  assign n2424 = n2423 ^ n2404 ;
  assign n2450 = n2435 ^ n2424 ;
  assign n2486 = n2485 ^ n2450 ;
  assign n2513 = n2512 ^ n2497 ;
  assign n2514 = n2513 ^ n2450 ;
  assign n2515 = n2486 & ~n2514 ;
  assign n2516 = n2515 ^ n2485 ;
  assign n2443 = n2434 ^ n2430 ;
  assign n2444 = n2431 & ~n2443 ;
  assign n2445 = n2444 ^ n2427 ;
  assign n2439 = n2403 ^ n2399 ;
  assign n2440 = n2400 & ~n2439 ;
  assign n2441 = n2440 ^ n2396 ;
  assign n2436 = n2435 ^ n2423 ;
  assign n2437 = n2424 & ~n2436 ;
  assign n2438 = n2437 ^ n2404 ;
  assign n2442 = n2441 ^ n2438 ;
  assign n2449 = n2445 ^ n2442 ;
  assign n2517 = n2516 ^ n2449 ;
  assign n2528 = n2527 ^ n2520 ;
  assign n2529 = n2528 ^ n2516 ;
  assign n2530 = n2517 & ~n2529 ;
  assign n2531 = n2530 ^ n2449 ;
  assign n2446 = n2445 ^ n2441 ;
  assign n2447 = n2442 & ~n2446 ;
  assign n2448 = n2447 ^ n2438 ;
  assign n2532 = n2531 ^ n2448 ;
  assign n2536 = n2535 ^ n2532 ;
  assign n2537 = n2513 ^ n2486 ;
  assign n2538 = n2482 ^ n2453 ;
  assign n2539 = x512 ^ x416 ;
  assign n2540 = n2538 & n2539 ;
  assign n2541 = n2537 & n2540 ;
  assign n2542 = n2528 ^ n2517 ;
  assign n2543 = n2541 & n2542 ;
  assign n2544 = n2536 & n2543 ;
  assign n2545 = n2535 ^ n2531 ;
  assign n2546 = n2532 & ~n2545 ;
  assign n2547 = n2546 ^ n2448 ;
  assign n2548 = n2544 & n2547 ;
  assign n2624 = x536 ^ x472 ;
  assign n2622 = x535 ^ x471 ;
  assign n2621 = x534 ^ x470 ;
  assign n2623 = n2622 ^ n2621 ;
  assign n2629 = n2624 ^ n2623 ;
  assign n2628 = x530 ^ x466 ;
  assign n2630 = n2629 ^ n2628 ;
  assign n2617 = x533 ^ x469 ;
  assign n2615 = x531 ^ x467 ;
  assign n2614 = x532 ^ x468 ;
  assign n2616 = n2615 ^ n2614 ;
  assign n2631 = n2617 ^ n2616 ;
  assign n2632 = n2631 ^ n2629 ;
  assign n2633 = n2630 & ~n2632 ;
  assign n2634 = n2633 ^ n2628 ;
  assign n2625 = n2624 ^ n2622 ;
  assign n2626 = n2623 & ~n2625 ;
  assign n2627 = n2626 ^ n2621 ;
  assign n2635 = n2634 ^ n2627 ;
  assign n2618 = n2617 ^ n2615 ;
  assign n2619 = n2616 & ~n2618 ;
  assign n2620 = n2619 ^ n2614 ;
  assign n2688 = n2634 ^ n2620 ;
  assign n2689 = n2635 & n2688 ;
  assign n2690 = n2689 ^ n2634 ;
  assign n2649 = x539 ^ x475 ;
  assign n2648 = x538 ^ x474 ;
  assign n2650 = n2649 ^ n2648 ;
  assign n2647 = x540 ^ x476 ;
  assign n2651 = n2650 ^ n2647 ;
  assign n2640 = x543 ^ x479 ;
  assign n2638 = x542 ^ x478 ;
  assign n2637 = x541 ^ x477 ;
  assign n2639 = n2638 ^ n2637 ;
  assign n2645 = n2640 ^ n2639 ;
  assign n2644 = x537 ^ x473 ;
  assign n2646 = n2645 ^ n2644 ;
  assign n2661 = n2651 ^ n2646 ;
  assign n2660 = x529 ^ x465 ;
  assign n2662 = n2661 ^ n2660 ;
  assign n2663 = n2631 ^ n2630 ;
  assign n2664 = n2663 ^ n2660 ;
  assign n2665 = ~n2662 & n2664 ;
  assign n2666 = n2665 ^ n2663 ;
  assign n2656 = n2649 ^ n2647 ;
  assign n2657 = n2650 & ~n2656 ;
  assign n2658 = n2657 ^ n2648 ;
  assign n2652 = n2651 ^ n2644 ;
  assign n2653 = ~n2646 & n2652 ;
  assign n2654 = n2653 ^ n2651 ;
  assign n2641 = n2640 ^ n2638 ;
  assign n2642 = n2639 & ~n2641 ;
  assign n2643 = n2642 ^ n2637 ;
  assign n2655 = n2654 ^ n2643 ;
  assign n2659 = n2658 ^ n2655 ;
  assign n2667 = n2666 ^ n2659 ;
  assign n2636 = n2635 ^ n2620 ;
  assign n2684 = n2659 ^ n2636 ;
  assign n2685 = ~n2667 & n2684 ;
  assign n2686 = n2685 ^ n2636 ;
  assign n2681 = n2658 ^ n2643 ;
  assign n2682 = ~n2655 & n2681 ;
  assign n2683 = n2682 ^ n2658 ;
  assign n2687 = n2686 ^ n2683 ;
  assign n2691 = n2690 ^ n2687 ;
  assign n2670 = n2663 ^ n2662 ;
  assign n2669 = x513 ^ x449 ;
  assign n2671 = n2670 ^ n2669 ;
  assign n2585 = x518 ^ x454 ;
  assign n2583 = x516 ^ x452 ;
  assign n2582 = x517 ^ x453 ;
  assign n2584 = n2583 ^ n2582 ;
  assign n2586 = n2585 ^ n2584 ;
  assign n2580 = x515 ^ x451 ;
  assign n2575 = x521 ^ x457 ;
  assign n2573 = x519 ^ x455 ;
  assign n2572 = x520 ^ x456 ;
  assign n2574 = n2573 ^ n2572 ;
  assign n2579 = n2575 ^ n2574 ;
  assign n2581 = n2580 ^ n2579 ;
  assign n2599 = n2586 ^ n2581 ;
  assign n2559 = x525 ^ x461 ;
  assign n2557 = x523 ^ x459 ;
  assign n2556 = x524 ^ x460 ;
  assign n2558 = n2557 ^ n2556 ;
  assign n2560 = n2559 ^ n2558 ;
  assign n2554 = x522 ^ x458 ;
  assign n2552 = x528 ^ x464 ;
  assign n2550 = x526 ^ x462 ;
  assign n2549 = x527 ^ x463 ;
  assign n2551 = n2550 ^ n2549 ;
  assign n2553 = n2552 ^ n2551 ;
  assign n2555 = n2554 ^ n2553 ;
  assign n2597 = n2560 ^ n2555 ;
  assign n2596 = x514 ^ x450 ;
  assign n2598 = n2597 ^ n2596 ;
  assign n2672 = n2599 ^ n2598 ;
  assign n2673 = n2672 ^ n2670 ;
  assign n2674 = n2671 & ~n2673 ;
  assign n2675 = n2674 ^ n2669 ;
  assign n2668 = n2667 ^ n2636 ;
  assign n2676 = n2675 ^ n2668 ;
  assign n2600 = n2599 ^ n2597 ;
  assign n2601 = n2598 & ~n2600 ;
  assign n2602 = n2601 ^ n2596 ;
  assign n2591 = n2585 ^ n2583 ;
  assign n2592 = n2584 & ~n2591 ;
  assign n2593 = n2592 ^ n2582 ;
  assign n2587 = n2586 ^ n2579 ;
  assign n2588 = ~n2581 & n2587 ;
  assign n2589 = n2588 ^ n2586 ;
  assign n2576 = n2575 ^ n2573 ;
  assign n2577 = n2574 & ~n2576 ;
  assign n2578 = n2577 ^ n2572 ;
  assign n2590 = n2589 ^ n2578 ;
  assign n2594 = n2593 ^ n2590 ;
  assign n2568 = n2559 ^ n2557 ;
  assign n2569 = n2558 & ~n2568 ;
  assign n2570 = n2569 ^ n2556 ;
  assign n2564 = n2552 ^ n2550 ;
  assign n2565 = n2551 & ~n2564 ;
  assign n2566 = n2565 ^ n2549 ;
  assign n2561 = n2560 ^ n2553 ;
  assign n2562 = ~n2555 & n2561 ;
  assign n2563 = n2562 ^ n2560 ;
  assign n2567 = n2566 ^ n2563 ;
  assign n2571 = n2570 ^ n2567 ;
  assign n2595 = n2594 ^ n2571 ;
  assign n2677 = n2602 ^ n2595 ;
  assign n2678 = n2677 ^ n2668 ;
  assign n2679 = n2676 & ~n2678 ;
  assign n2680 = n2679 ^ n2675 ;
  assign n2692 = n2691 ^ n2680 ;
  assign n2610 = n2593 ^ n2589 ;
  assign n2611 = n2590 & n2610 ;
  assign n2612 = n2611 ^ n2589 ;
  assign n2606 = n2570 ^ n2566 ;
  assign n2607 = n2567 & ~n2606 ;
  assign n2608 = n2607 ^ n2563 ;
  assign n2603 = n2602 ^ n2571 ;
  assign n2604 = ~n2595 & n2603 ;
  assign n2605 = n2604 ^ n2602 ;
  assign n2609 = n2608 ^ n2605 ;
  assign n2613 = n2612 ^ n2609 ;
  assign n2693 = n2692 ^ n2613 ;
  assign n2694 = n2677 ^ n2676 ;
  assign n2695 = x512 ^ x448 ;
  assign n2696 = n2672 ^ n2671 ;
  assign n2697 = n2695 & n2696 ;
  assign n2698 = n2694 & n2697 ;
  assign n2699 = n2693 & n2698 ;
  assign n2706 = n2680 ^ n2613 ;
  assign n2707 = ~n2692 & n2706 ;
  assign n2708 = n2707 ^ n2613 ;
  assign n2703 = n2690 ^ n2686 ;
  assign n2704 = n2687 & ~n2703 ;
  assign n2705 = n2704 ^ n2683 ;
  assign n2709 = n2708 ^ n2705 ;
  assign n2700 = n2612 ^ n2608 ;
  assign n2701 = n2609 & ~n2700 ;
  assign n2702 = n2701 ^ n2605 ;
  assign n2710 = n2709 ^ n2702 ;
  assign n2711 = n2699 & n2710 ;
  assign n2712 = n2708 ^ n2702 ;
  assign n2713 = n2709 & ~n2712 ;
  assign n2714 = n2713 ^ n2705 ;
  assign n2716 = ~n2711 & ~n2714 ;
  assign n2715 = n2714 ^ n2711 ;
  assign n2717 = n2716 ^ n2715 ;
  assign n2793 = x534 ^ x502 ;
  assign n2792 = x535 ^ x503 ;
  assign n2794 = n2793 ^ n2792 ;
  assign n2791 = x536 ^ x504 ;
  assign n2801 = n2793 ^ n2791 ;
  assign n2802 = n2794 & ~n2801 ;
  assign n2803 = n2802 ^ n2792 ;
  assign n2795 = n2794 ^ n2791 ;
  assign n2790 = x530 ^ x498 ;
  assign n2796 = n2795 ^ n2790 ;
  assign n2786 = x533 ^ x501 ;
  assign n2784 = x531 ^ x499 ;
  assign n2783 = x532 ^ x500 ;
  assign n2785 = n2784 ^ n2783 ;
  assign n2797 = n2786 ^ n2785 ;
  assign n2798 = n2797 ^ n2795 ;
  assign n2799 = n2796 & ~n2798 ;
  assign n2800 = n2799 ^ n2790 ;
  assign n2804 = n2803 ^ n2800 ;
  assign n2787 = n2786 ^ n2784 ;
  assign n2788 = n2785 & ~n2787 ;
  assign n2789 = n2788 ^ n2783 ;
  assign n2857 = n2803 ^ n2789 ;
  assign n2858 = n2804 & ~n2857 ;
  assign n2859 = n2858 ^ n2800 ;
  assign n2830 = x529 ^ x497 ;
  assign n2816 = x540 ^ x508 ;
  assign n2814 = x538 ^ x506 ;
  assign n2813 = x539 ^ x507 ;
  assign n2815 = n2814 ^ n2813 ;
  assign n2817 = n2816 ^ n2815 ;
  assign n2810 = x543 ^ x511 ;
  assign n2808 = x541 ^ x509 ;
  assign n2807 = x542 ^ x510 ;
  assign n2809 = n2808 ^ n2807 ;
  assign n2811 = n2810 ^ n2809 ;
  assign n2806 = x537 ^ x505 ;
  assign n2812 = n2811 ^ n2806 ;
  assign n2829 = n2817 ^ n2812 ;
  assign n2831 = n2830 ^ n2829 ;
  assign n2832 = n2797 ^ n2796 ;
  assign n2833 = n2832 ^ n2830 ;
  assign n2834 = n2831 & ~n2833 ;
  assign n2835 = n2834 ^ n2829 ;
  assign n2825 = n2816 ^ n2814 ;
  assign n2826 = n2815 & ~n2825 ;
  assign n2827 = n2826 ^ n2813 ;
  assign n2821 = n2810 ^ n2808 ;
  assign n2822 = n2809 & ~n2821 ;
  assign n2823 = n2822 ^ n2807 ;
  assign n2818 = n2817 ^ n2811 ;
  assign n2819 = n2812 & ~n2818 ;
  assign n2820 = n2819 ^ n2806 ;
  assign n2824 = n2823 ^ n2820 ;
  assign n2828 = n2827 ^ n2824 ;
  assign n2836 = n2835 ^ n2828 ;
  assign n2805 = n2804 ^ n2789 ;
  assign n2853 = n2835 ^ n2805 ;
  assign n2854 = ~n2836 & n2853 ;
  assign n2855 = n2854 ^ n2805 ;
  assign n2850 = n2827 ^ n2823 ;
  assign n2851 = n2824 & ~n2850 ;
  assign n2852 = n2851 ^ n2820 ;
  assign n2856 = n2855 ^ n2852 ;
  assign n2860 = n2859 ^ n2856 ;
  assign n2839 = x513 ^ x481 ;
  assign n2838 = n2832 ^ n2831 ;
  assign n2840 = n2839 ^ n2838 ;
  assign n2754 = x515 ^ x483 ;
  assign n2752 = x521 ^ x489 ;
  assign n2750 = x519 ^ x487 ;
  assign n2749 = x520 ^ x488 ;
  assign n2751 = n2750 ^ n2749 ;
  assign n2753 = n2752 ^ n2751 ;
  assign n2755 = n2754 ^ n2753 ;
  assign n2747 = x518 ^ x486 ;
  assign n2745 = x516 ^ x484 ;
  assign n2744 = x517 ^ x485 ;
  assign n2746 = n2745 ^ n2744 ;
  assign n2748 = n2747 ^ n2746 ;
  assign n2756 = n2755 ^ n2748 ;
  assign n2728 = x525 ^ x493 ;
  assign n2726 = x523 ^ x491 ;
  assign n2725 = x524 ^ x492 ;
  assign n2727 = n2726 ^ n2725 ;
  assign n2729 = n2728 ^ n2727 ;
  assign n2723 = x522 ^ x490 ;
  assign n2721 = x528 ^ x496 ;
  assign n2719 = x526 ^ x494 ;
  assign n2718 = x527 ^ x495 ;
  assign n2720 = n2719 ^ n2718 ;
  assign n2722 = n2721 ^ n2720 ;
  assign n2724 = n2723 ^ n2722 ;
  assign n2742 = n2729 ^ n2724 ;
  assign n2741 = x514 ^ x482 ;
  assign n2743 = n2742 ^ n2741 ;
  assign n2841 = n2756 ^ n2743 ;
  assign n2842 = n2841 ^ n2839 ;
  assign n2843 = n2840 & ~n2842 ;
  assign n2844 = n2843 ^ n2838 ;
  assign n2837 = n2836 ^ n2805 ;
  assign n2845 = n2844 ^ n2837 ;
  assign n2768 = n2747 ^ n2745 ;
  assign n2769 = n2746 & ~n2768 ;
  assign n2770 = n2769 ^ n2744 ;
  assign n2764 = n2753 ^ n2748 ;
  assign n2765 = ~n2755 & n2764 ;
  assign n2766 = n2765 ^ n2748 ;
  assign n2761 = n2752 ^ n2750 ;
  assign n2762 = n2751 & ~n2761 ;
  assign n2763 = n2762 ^ n2749 ;
  assign n2767 = n2766 ^ n2763 ;
  assign n2771 = n2770 ^ n2767 ;
  assign n2757 = n2756 ^ n2742 ;
  assign n2758 = n2743 & ~n2757 ;
  assign n2759 = n2758 ^ n2741 ;
  assign n2737 = n2728 ^ n2726 ;
  assign n2738 = n2727 & ~n2737 ;
  assign n2739 = n2738 ^ n2725 ;
  assign n2733 = n2721 ^ n2719 ;
  assign n2734 = n2720 & ~n2733 ;
  assign n2735 = n2734 ^ n2718 ;
  assign n2730 = n2729 ^ n2722 ;
  assign n2731 = ~n2724 & n2730 ;
  assign n2732 = n2731 ^ n2729 ;
  assign n2736 = n2735 ^ n2732 ;
  assign n2740 = n2739 ^ n2736 ;
  assign n2760 = n2759 ^ n2740 ;
  assign n2846 = n2771 ^ n2760 ;
  assign n2847 = n2846 ^ n2837 ;
  assign n2848 = n2845 & ~n2847 ;
  assign n2849 = n2848 ^ n2844 ;
  assign n2861 = n2860 ^ n2849 ;
  assign n2779 = n2770 ^ n2766 ;
  assign n2780 = n2767 & ~n2779 ;
  assign n2781 = n2780 ^ n2763 ;
  assign n2775 = n2739 ^ n2735 ;
  assign n2776 = n2736 & ~n2775 ;
  assign n2777 = n2776 ^ n2732 ;
  assign n2772 = n2771 ^ n2740 ;
  assign n2773 = n2760 & ~n2772 ;
  assign n2774 = n2773 ^ n2759 ;
  assign n2778 = n2777 ^ n2774 ;
  assign n2782 = n2781 ^ n2778 ;
  assign n2862 = n2861 ^ n2782 ;
  assign n2863 = n2841 ^ n2840 ;
  assign n2864 = x512 ^ x480 ;
  assign n2865 = n2863 & n2864 ;
  assign n2866 = n2846 ^ n2845 ;
  assign n2867 = n2865 & n2866 ;
  assign n2868 = n2862 & n2867 ;
  assign n2875 = n2849 ^ n2782 ;
  assign n2876 = ~n2861 & n2875 ;
  assign n2877 = n2876 ^ n2782 ;
  assign n2872 = n2859 ^ n2852 ;
  assign n2873 = n2856 & n2872 ;
  assign n2874 = n2873 ^ n2852 ;
  assign n2878 = n2877 ^ n2874 ;
  assign n2869 = n2781 ^ n2777 ;
  assign n2870 = n2778 & ~n2869 ;
  assign n2871 = n2870 ^ n2774 ;
  assign n2879 = n2878 ^ n2871 ;
  assign n2880 = n2868 & n2879 ;
  assign n2881 = n2877 ^ n2871 ;
  assign n2882 = n2878 & ~n2881 ;
  assign n2883 = n2882 ^ n2874 ;
  assign n2885 = ~n2880 & ~n2883 ;
  assign n2884 = n2883 ^ n2880 ;
  assign n2886 = n2885 ^ n2884 ;
  assign n2888 = ~n2717 & n2886 ;
  assign n2887 = n2886 ^ n2717 ;
  assign n2889 = n2888 ^ n2887 ;
  assign n2890 = n2889 ^ n2886 ;
  assign n2891 = n2548 & ~n2890 ;
  assign n2990 = x514 ^ x386 ;
  assign n2987 = x522 ^ x394 ;
  assign n2985 = x528 ^ x400 ;
  assign n2983 = x526 ^ x398 ;
  assign n2982 = x527 ^ x399 ;
  assign n2984 = n2983 ^ n2982 ;
  assign n2986 = n2985 ^ n2984 ;
  assign n2988 = n2987 ^ n2986 ;
  assign n2980 = x525 ^ x397 ;
  assign n2978 = x523 ^ x395 ;
  assign n2977 = x524 ^ x396 ;
  assign n2979 = n2978 ^ n2977 ;
  assign n2981 = n2980 ^ n2979 ;
  assign n2989 = n2988 ^ n2981 ;
  assign n2991 = n2990 ^ n2989 ;
  assign n2974 = x515 ^ x387 ;
  assign n2972 = x521 ^ x393 ;
  assign n2970 = x519 ^ x391 ;
  assign n2969 = x520 ^ x392 ;
  assign n2971 = n2970 ^ n2969 ;
  assign n2973 = n2972 ^ n2971 ;
  assign n2975 = n2974 ^ n2973 ;
  assign n2967 = x518 ^ x390 ;
  assign n2965 = x516 ^ x388 ;
  assign n2964 = x517 ^ x389 ;
  assign n2966 = n2965 ^ n2964 ;
  assign n2968 = n2967 ^ n2966 ;
  assign n2976 = n2975 ^ n2968 ;
  assign n3019 = n2990 ^ n2976 ;
  assign n3020 = n2991 & ~n3019 ;
  assign n3021 = n3020 ^ n2989 ;
  assign n3015 = n2980 ^ n2978 ;
  assign n3016 = n2979 & ~n3015 ;
  assign n3017 = n3016 ^ n2977 ;
  assign n3011 = n2985 ^ n2983 ;
  assign n3012 = n2984 & ~n3011 ;
  assign n3013 = n3012 ^ n2982 ;
  assign n3008 = n2986 ^ n2981 ;
  assign n3009 = ~n2988 & n3008 ;
  assign n3010 = n3009 ^ n2981 ;
  assign n3014 = n3013 ^ n3010 ;
  assign n3018 = n3017 ^ n3014 ;
  assign n3022 = n3021 ^ n3018 ;
  assign n3004 = n2967 ^ n2965 ;
  assign n3005 = n2966 & ~n3004 ;
  assign n3006 = n3005 ^ n2964 ;
  assign n3000 = n2973 ^ n2968 ;
  assign n3001 = ~n2975 & n3000 ;
  assign n3002 = n3001 ^ n2968 ;
  assign n2997 = n2972 ^ n2970 ;
  assign n2998 = n2971 & ~n2997 ;
  assign n2999 = n2998 ^ n2969 ;
  assign n3003 = n3002 ^ n2999 ;
  assign n3007 = n3006 ^ n3003 ;
  assign n3034 = n3021 ^ n3007 ;
  assign n3035 = n3022 & ~n3034 ;
  assign n3036 = n3035 ^ n3018 ;
  assign n3031 = n3017 ^ n3013 ;
  assign n3032 = n3014 & ~n3031 ;
  assign n3033 = n3032 ^ n3010 ;
  assign n3037 = n3036 ^ n3033 ;
  assign n3028 = n3006 ^ n3002 ;
  assign n3029 = n3003 & ~n3028 ;
  assign n3030 = n3029 ^ n2999 ;
  assign n3043 = n3033 ^ n3030 ;
  assign n3044 = ~n3037 & n3043 ;
  assign n3045 = n3044 ^ n3030 ;
  assign n2962 = x513 ^ x385 ;
  assign n2928 = x533 ^ x405 ;
  assign n2926 = x531 ^ x403 ;
  assign n2925 = x532 ^ x404 ;
  assign n2927 = n2926 ^ n2925 ;
  assign n2929 = n2928 ^ n2927 ;
  assign n2923 = x530 ^ x402 ;
  assign n2921 = x536 ^ x408 ;
  assign n2919 = x534 ^ x406 ;
  assign n2918 = x535 ^ x407 ;
  assign n2920 = n2919 ^ n2918 ;
  assign n2922 = n2921 ^ n2920 ;
  assign n2924 = n2923 ^ n2922 ;
  assign n2930 = n2929 ^ n2924 ;
  assign n2901 = x538 ^ x410 ;
  assign n2900 = x539 ^ x411 ;
  assign n2902 = n2901 ^ n2900 ;
  assign n2899 = x540 ^ x412 ;
  assign n2903 = n2902 ^ n2899 ;
  assign n2897 = x537 ^ x409 ;
  assign n2894 = x541 ^ x413 ;
  assign n2893 = x542 ^ x414 ;
  assign n2895 = n2894 ^ n2893 ;
  assign n2892 = x543 ^ x415 ;
  assign n2896 = n2895 ^ n2892 ;
  assign n2898 = n2897 ^ n2896 ;
  assign n2916 = n2903 ^ n2898 ;
  assign n2915 = x529 ^ x401 ;
  assign n2917 = n2916 ^ n2915 ;
  assign n2961 = n2930 ^ n2917 ;
  assign n2963 = n2962 ^ n2961 ;
  assign n2992 = n2991 ^ n2976 ;
  assign n2993 = n2992 ^ n2962 ;
  assign n2994 = n2963 & ~n2993 ;
  assign n2995 = n2994 ^ n2961 ;
  assign n2942 = n2928 ^ n2926 ;
  assign n2943 = n2927 & ~n2942 ;
  assign n2944 = n2943 ^ n2925 ;
  assign n2938 = n2921 ^ n2919 ;
  assign n2939 = n2920 & ~n2938 ;
  assign n2940 = n2939 ^ n2918 ;
  assign n2935 = n2929 ^ n2923 ;
  assign n2936 = n2924 & ~n2935 ;
  assign n2937 = n2936 ^ n2922 ;
  assign n2941 = n2940 ^ n2937 ;
  assign n2945 = n2944 ^ n2941 ;
  assign n2931 = n2930 ^ n2916 ;
  assign n2932 = n2917 & ~n2931 ;
  assign n2933 = n2932 ^ n2915 ;
  assign n2911 = n2900 ^ n2899 ;
  assign n2912 = ~n2902 & n2911 ;
  assign n2913 = n2912 ^ n2899 ;
  assign n2907 = n2893 ^ n2892 ;
  assign n2908 = ~n2895 & n2907 ;
  assign n2909 = n2908 ^ n2892 ;
  assign n2904 = n2903 ^ n2897 ;
  assign n2905 = n2898 & ~n2904 ;
  assign n2906 = n2905 ^ n2896 ;
  assign n2910 = n2909 ^ n2906 ;
  assign n2914 = n2913 ^ n2910 ;
  assign n2934 = n2933 ^ n2914 ;
  assign n2960 = n2945 ^ n2934 ;
  assign n2996 = n2995 ^ n2960 ;
  assign n3023 = n3022 ^ n3007 ;
  assign n3024 = n3023 ^ n2960 ;
  assign n3025 = n2996 & ~n3024 ;
  assign n3026 = n3025 ^ n2995 ;
  assign n2953 = n2944 ^ n2940 ;
  assign n2954 = n2941 & ~n2953 ;
  assign n2955 = n2954 ^ n2937 ;
  assign n2949 = n2913 ^ n2909 ;
  assign n2950 = n2910 & ~n2949 ;
  assign n2951 = n2950 ^ n2906 ;
  assign n2946 = n2945 ^ n2933 ;
  assign n2947 = n2934 & ~n2946 ;
  assign n2948 = n2947 ^ n2914 ;
  assign n2952 = n2951 ^ n2948 ;
  assign n2959 = n2955 ^ n2952 ;
  assign n3027 = n3026 ^ n2959 ;
  assign n3038 = n3037 ^ n3030 ;
  assign n3039 = n3038 ^ n3026 ;
  assign n3040 = n3027 & ~n3039 ;
  assign n3041 = n3040 ^ n2959 ;
  assign n2956 = n2955 ^ n2951 ;
  assign n2957 = n2952 & ~n2956 ;
  assign n2958 = n2957 ^ n2948 ;
  assign n3042 = n3041 ^ n2958 ;
  assign n3046 = n3045 ^ n3042 ;
  assign n3047 = n3023 ^ n2996 ;
  assign n3048 = n2992 ^ n2963 ;
  assign n3049 = x512 ^ x384 ;
  assign n3050 = n3048 & n3049 ;
  assign n3051 = n3047 & n3050 ;
  assign n3052 = n3038 ^ n3027 ;
  assign n3053 = n3051 & n3052 ;
  assign n3054 = n3046 & n3053 ;
  assign n3055 = n3045 ^ n3041 ;
  assign n3056 = n3042 & ~n3055 ;
  assign n3057 = n3056 ^ n2958 ;
  assign n3058 = n3054 & n3057 ;
  assign n3059 = n2891 & ~n3058 ;
  assign n3060 = n3059 ^ n2891 ;
  assign n3061 = n2381 & n3060 ;
  assign n3063 = ~n2214 & n3061 ;
  assign n3062 = n3061 ^ n2214 ;
  assign n3064 = n3063 ^ n3062 ;
  assign n3065 = n3064 ^ n2214 ;
  assign n3066 = n2047 & n3065 ;
  assign n3068 = ~n1880 & n3066 ;
  assign n3067 = n3066 ^ n1880 ;
  assign n3069 = n3068 ^ n3067 ;
  assign n3070 = n3069 ^ n1880 ;
  assign n3071 = n1713 & n3070 ;
  assign n3073 = ~n1546 & n3071 ;
  assign n3072 = n3071 ^ n1546 ;
  assign n3074 = n3073 ^ n3072 ;
  assign n3075 = n3074 ^ n1546 ;
  assign n3076 = n1379 & n3075 ;
  assign n3078 = ~n1212 & n3076 ;
  assign n3077 = n3076 ^ n1212 ;
  assign n3079 = n3078 ^ n3077 ;
  assign n3080 = n3079 ^ n1212 ;
  assign n3081 = n1045 & n3080 ;
  assign n3083 = ~n878 & n3081 ;
  assign n3082 = n3081 ^ n878 ;
  assign n3084 = n3083 ^ n3082 ;
  assign n3085 = n3084 ^ n878 ;
  assign n3086 = n711 & n3085 ;
  assign n3254 = n3253 ^ n3086 ;
  assign n3763 = n3252 ^ n3249 ;
  assign n3269 = n2547 ^ n2544 ;
  assign n3267 = ~n2716 & ~n2885 ;
  assign n3268 = n3267 ^ n2890 ;
  assign n3270 = n3269 ^ n3268 ;
  assign n3271 = n2890 ^ n2548 ;
  assign n3330 = n3269 ^ n2548 ;
  assign n3274 = n2879 ^ n2868 ;
  assign n3273 = n2710 ^ n2699 ;
  assign n3275 = n3274 ^ n3273 ;
  assign n3276 = n2884 ^ n2715 ;
  assign n3286 = n2698 ^ n2693 ;
  assign n3278 = n2866 ^ n2865 ;
  assign n3277 = n2697 ^ n2694 ;
  assign n3279 = n3278 ^ n3277 ;
  assign n3280 = n2864 ^ n2863 ;
  assign n3281 = n2696 ^ n2695 ;
  assign n3282 = ~n3280 & n3281 ;
  assign n3283 = n3282 ^ n3277 ;
  assign n3284 = n3279 & n3283 ;
  assign n3285 = n3284 ^ n3282 ;
  assign n3287 = n3286 ^ n3285 ;
  assign n3288 = n2867 ^ n2862 ;
  assign n3289 = n3288 ^ n3285 ;
  assign n3290 = n3287 & n3289 ;
  assign n3291 = n3290 ^ n3286 ;
  assign n3292 = n3291 ^ n3273 ;
  assign n3293 = n3291 ^ n3274 ;
  assign n3294 = n3292 & n3293 ;
  assign n3295 = n3294 ^ n3273 ;
  assign n3296 = n3295 ^ n2884 ;
  assign n3297 = ~n3276 & ~n3296 ;
  assign n3298 = n3297 ^ n2884 ;
  assign n3299 = n3298 ^ n2886 ;
  assign n3300 = ~n2887 & n3299 ;
  assign n3301 = n3300 ^ n2717 ;
  assign n3302 = n3275 & ~n3301 ;
  assign n3303 = n3302 ^ n3273 ;
  assign n3272 = n2543 ^ n2536 ;
  assign n3304 = n3303 ^ n3272 ;
  assign n3308 = n2542 ^ n2541 ;
  assign n3305 = n3288 ^ n3286 ;
  assign n3306 = ~n3301 & n3305 ;
  assign n3307 = n3306 ^ n3286 ;
  assign n3309 = n3308 ^ n3307 ;
  assign n3312 = n2540 ^ n2537 ;
  assign n3310 = n3279 & ~n3301 ;
  assign n3311 = n3310 ^ n3277 ;
  assign n3313 = n3312 ^ n3311 ;
  assign n3314 = n2539 ^ n2538 ;
  assign n3315 = n3281 ^ n3280 ;
  assign n3316 = n3301 & n3315 ;
  assign n3317 = n3316 ^ n3280 ;
  assign n3318 = n3314 & ~n3317 ;
  assign n3319 = n3318 ^ n3311 ;
  assign n3320 = ~n3313 & ~n3319 ;
  assign n3321 = n3320 ^ n3311 ;
  assign n3322 = n3321 ^ n3307 ;
  assign n3323 = ~n3309 & n3322 ;
  assign n3324 = n3323 ^ n3307 ;
  assign n3325 = n3324 ^ n3272 ;
  assign n3326 = ~n3304 & ~n3325 ;
  assign n3327 = n3326 ^ n3272 ;
  assign n3328 = n3327 ^ n3268 ;
  assign n3329 = n3270 & ~n3328 ;
  assign n3331 = n3330 ^ n3329 ;
  assign n3332 = n3271 & ~n3331 ;
  assign n3333 = n3332 ^ n2890 ;
  assign n3334 = ~n3270 & n3333 ;
  assign n3335 = n3334 ^ n3269 ;
  assign n3266 = n3057 ^ n3054 ;
  assign n3336 = n3335 ^ n3266 ;
  assign n3337 = ~n3266 & n3335 ;
  assign n3338 = n3337 ^ n3059 ;
  assign n3339 = n3337 ^ n3336 ;
  assign n3341 = n3304 & n3333 ;
  assign n3342 = n3341 ^ n3272 ;
  assign n3340 = n3053 ^ n3046 ;
  assign n3343 = n3342 ^ n3340 ;
  assign n3346 = n3052 ^ n3051 ;
  assign n3344 = n3309 & n3333 ;
  assign n3345 = n3344 ^ n3308 ;
  assign n3347 = n3346 ^ n3345 ;
  assign n3350 = n3050 ^ n3047 ;
  assign n3348 = n3313 & n3333 ;
  assign n3349 = n3348 ^ n3312 ;
  assign n3351 = n3350 ^ n3349 ;
  assign n3352 = n3049 ^ n3048 ;
  assign n3353 = n3317 ^ n3314 ;
  assign n3354 = n3333 & n3353 ;
  assign n3355 = n3354 ^ n3314 ;
  assign n3356 = n3352 & ~n3355 ;
  assign n3357 = n3356 ^ n3349 ;
  assign n3358 = ~n3351 & ~n3357 ;
  assign n3359 = n3358 ^ n3349 ;
  assign n3360 = n3359 ^ n3345 ;
  assign n3361 = ~n3347 & n3360 ;
  assign n3362 = n3361 ^ n3345 ;
  assign n3363 = n3362 ^ n3340 ;
  assign n3364 = ~n3343 & ~n3363 ;
  assign n3365 = n3364 ^ n3340 ;
  assign n3366 = ~n3339 & ~n3365 ;
  assign n3367 = ~n3338 & ~n3366 ;
  assign n3368 = n3060 ^ n3058 ;
  assign n3369 = ~n3367 & ~n3368 ;
  assign n3370 = n3336 & n3369 ;
  assign n3371 = n3370 ^ n3335 ;
  assign n3265 = n2380 ^ n2377 ;
  assign n3372 = n3371 ^ n3265 ;
  assign n3373 = n3060 ^ n2381 ;
  assign n3402 = n3265 ^ n2381 ;
  assign n3375 = n3343 & ~n3369 ;
  assign n3376 = n3375 ^ n3340 ;
  assign n3374 = n2376 ^ n2369 ;
  assign n3377 = n3376 ^ n3374 ;
  assign n3380 = n2375 ^ n2374 ;
  assign n3378 = n3347 & ~n3369 ;
  assign n3379 = n3378 ^ n3346 ;
  assign n3381 = n3380 ^ n3379 ;
  assign n3384 = n2373 ^ n2370 ;
  assign n3382 = n3351 & ~n3369 ;
  assign n3383 = n3382 ^ n3350 ;
  assign n3385 = n3384 ^ n3383 ;
  assign n3386 = n2372 ^ n2371 ;
  assign n3387 = n3355 ^ n3352 ;
  assign n3388 = ~n3369 & n3387 ;
  assign n3389 = n3388 ^ n3352 ;
  assign n3390 = n3386 & ~n3389 ;
  assign n3391 = n3390 ^ n3383 ;
  assign n3392 = ~n3385 & ~n3391 ;
  assign n3393 = n3392 ^ n3383 ;
  assign n3394 = n3393 ^ n3379 ;
  assign n3395 = ~n3381 & n3394 ;
  assign n3396 = n3395 ^ n3379 ;
  assign n3397 = n3396 ^ n3374 ;
  assign n3398 = ~n3377 & ~n3397 ;
  assign n3399 = n3398 ^ n3374 ;
  assign n3400 = n3399 ^ n3371 ;
  assign n3401 = ~n3372 & n3400 ;
  assign n3403 = n3402 ^ n3401 ;
  assign n3404 = ~n3373 & ~n3403 ;
  assign n3405 = n3404 ^ n3060 ;
  assign n3406 = n3372 & n3405 ;
  assign n3407 = n3406 ^ n3371 ;
  assign n3264 = n2213 ^ n2210 ;
  assign n3408 = n3407 ^ n3264 ;
  assign n3409 = ~n3264 & n3407 ;
  assign n3410 = n3409 ^ n3063 ;
  assign n3411 = n3409 ^ n3408 ;
  assign n3413 = n3377 & ~n3405 ;
  assign n3414 = n3413 ^ n3374 ;
  assign n3412 = n2209 ^ n2202 ;
  assign n3415 = n3414 ^ n3412 ;
  assign n3418 = n2208 ^ n2207 ;
  assign n3416 = n3381 & ~n3405 ;
  assign n3417 = n3416 ^ n3380 ;
  assign n3419 = n3418 ^ n3417 ;
  assign n3422 = n2206 ^ n2203 ;
  assign n3420 = n3385 & ~n3405 ;
  assign n3421 = n3420 ^ n3384 ;
  assign n3423 = n3422 ^ n3421 ;
  assign n3424 = n2205 ^ n2204 ;
  assign n3425 = n3389 ^ n3386 ;
  assign n3426 = ~n3405 & n3425 ;
  assign n3427 = n3426 ^ n3386 ;
  assign n3428 = n3424 & ~n3427 ;
  assign n3429 = n3428 ^ n3421 ;
  assign n3430 = ~n3423 & ~n3429 ;
  assign n3431 = n3430 ^ n3421 ;
  assign n3432 = n3431 ^ n3417 ;
  assign n3433 = ~n3419 & n3432 ;
  assign n3434 = n3433 ^ n3417 ;
  assign n3435 = n3434 ^ n3412 ;
  assign n3436 = ~n3415 & ~n3435 ;
  assign n3437 = n3436 ^ n3412 ;
  assign n3438 = ~n3411 & ~n3437 ;
  assign n3439 = ~n3410 & ~n3438 ;
  assign n3440 = ~n3064 & ~n3439 ;
  assign n3441 = n3408 & n3440 ;
  assign n3442 = n3441 ^ n3407 ;
  assign n3263 = n2046 ^ n2043 ;
  assign n3443 = n3442 ^ n3263 ;
  assign n3444 = n3065 ^ n2047 ;
  assign n3473 = n3263 ^ n2047 ;
  assign n3446 = n3415 & ~n3440 ;
  assign n3447 = n3446 ^ n3412 ;
  assign n3445 = n2042 ^ n2035 ;
  assign n3448 = n3447 ^ n3445 ;
  assign n3451 = n2041 ^ n2040 ;
  assign n3449 = n3419 & ~n3440 ;
  assign n3450 = n3449 ^ n3418 ;
  assign n3452 = n3451 ^ n3450 ;
  assign n3455 = n2039 ^ n2036 ;
  assign n3453 = n3423 & ~n3440 ;
  assign n3454 = n3453 ^ n3422 ;
  assign n3456 = n3455 ^ n3454 ;
  assign n3457 = n2038 ^ n2037 ;
  assign n3458 = n3427 ^ n3424 ;
  assign n3459 = ~n3440 & n3458 ;
  assign n3460 = n3459 ^ n3424 ;
  assign n3461 = n3457 & ~n3460 ;
  assign n3462 = n3461 ^ n3454 ;
  assign n3463 = ~n3456 & ~n3462 ;
  assign n3464 = n3463 ^ n3454 ;
  assign n3465 = n3464 ^ n3450 ;
  assign n3466 = ~n3452 & n3465 ;
  assign n3467 = n3466 ^ n3450 ;
  assign n3468 = n3467 ^ n3445 ;
  assign n3469 = ~n3448 & ~n3468 ;
  assign n3470 = n3469 ^ n3445 ;
  assign n3471 = n3470 ^ n3442 ;
  assign n3472 = ~n3443 & n3471 ;
  assign n3474 = n3473 ^ n3472 ;
  assign n3475 = ~n3444 & ~n3474 ;
  assign n3476 = n3475 ^ n3065 ;
  assign n3477 = n3443 & n3476 ;
  assign n3478 = n3477 ^ n3442 ;
  assign n3262 = n1879 ^ n1876 ;
  assign n3479 = n3478 ^ n3262 ;
  assign n3480 = ~n3262 & n3478 ;
  assign n3481 = n3480 ^ n3068 ;
  assign n3482 = n3480 ^ n3479 ;
  assign n3484 = n3448 & ~n3476 ;
  assign n3485 = n3484 ^ n3445 ;
  assign n3483 = n1875 ^ n1868 ;
  assign n3486 = n3485 ^ n3483 ;
  assign n3489 = n1874 ^ n1873 ;
  assign n3487 = n3452 & ~n3476 ;
  assign n3488 = n3487 ^ n3451 ;
  assign n3490 = n3489 ^ n3488 ;
  assign n3493 = n1872 ^ n1869 ;
  assign n3491 = n3456 & ~n3476 ;
  assign n3492 = n3491 ^ n3455 ;
  assign n3494 = n3493 ^ n3492 ;
  assign n3495 = n1871 ^ n1870 ;
  assign n3496 = n3460 ^ n3457 ;
  assign n3497 = ~n3476 & n3496 ;
  assign n3498 = n3497 ^ n3457 ;
  assign n3499 = n3495 & ~n3498 ;
  assign n3500 = n3499 ^ n3492 ;
  assign n3501 = ~n3494 & ~n3500 ;
  assign n3502 = n3501 ^ n3492 ;
  assign n3503 = n3502 ^ n3488 ;
  assign n3504 = ~n3490 & n3503 ;
  assign n3505 = n3504 ^ n3488 ;
  assign n3506 = n3505 ^ n3483 ;
  assign n3507 = ~n3486 & ~n3506 ;
  assign n3508 = n3507 ^ n3483 ;
  assign n3509 = ~n3482 & ~n3508 ;
  assign n3510 = ~n3481 & ~n3509 ;
  assign n3511 = ~n3069 & ~n3510 ;
  assign n3512 = n3479 & n3511 ;
  assign n3513 = n3512 ^ n3478 ;
  assign n3261 = n1712 ^ n1709 ;
  assign n3514 = n3513 ^ n3261 ;
  assign n3515 = n3070 ^ n1713 ;
  assign n3544 = n3261 ^ n1713 ;
  assign n3517 = n3486 & ~n3511 ;
  assign n3518 = n3517 ^ n3483 ;
  assign n3516 = n1708 ^ n1701 ;
  assign n3519 = n3518 ^ n3516 ;
  assign n3522 = n1707 ^ n1706 ;
  assign n3520 = n3490 & ~n3511 ;
  assign n3521 = n3520 ^ n3489 ;
  assign n3523 = n3522 ^ n3521 ;
  assign n3526 = n1705 ^ n1702 ;
  assign n3524 = n3494 & ~n3511 ;
  assign n3525 = n3524 ^ n3493 ;
  assign n3527 = n3526 ^ n3525 ;
  assign n3528 = n1704 ^ n1703 ;
  assign n3529 = n3498 ^ n3495 ;
  assign n3530 = ~n3511 & n3529 ;
  assign n3531 = n3530 ^ n3495 ;
  assign n3532 = n3528 & ~n3531 ;
  assign n3533 = n3532 ^ n3525 ;
  assign n3534 = ~n3527 & ~n3533 ;
  assign n3535 = n3534 ^ n3525 ;
  assign n3536 = n3535 ^ n3521 ;
  assign n3537 = ~n3523 & n3536 ;
  assign n3538 = n3537 ^ n3521 ;
  assign n3539 = n3538 ^ n3516 ;
  assign n3540 = ~n3519 & ~n3539 ;
  assign n3541 = n3540 ^ n3516 ;
  assign n3542 = n3541 ^ n3513 ;
  assign n3543 = ~n3514 & n3542 ;
  assign n3545 = n3544 ^ n3543 ;
  assign n3546 = ~n3515 & ~n3545 ;
  assign n3547 = n3546 ^ n3070 ;
  assign n3548 = n3514 & n3547 ;
  assign n3549 = n3548 ^ n3513 ;
  assign n3260 = n1545 ^ n1542 ;
  assign n3550 = n3549 ^ n3260 ;
  assign n3551 = ~n3260 & n3549 ;
  assign n3552 = n3551 ^ n3073 ;
  assign n3553 = n3551 ^ n3550 ;
  assign n3555 = n3519 & ~n3547 ;
  assign n3556 = n3555 ^ n3516 ;
  assign n3554 = n1541 ^ n1534 ;
  assign n3557 = n3556 ^ n3554 ;
  assign n3560 = n1540 ^ n1539 ;
  assign n3558 = n3523 & ~n3547 ;
  assign n3559 = n3558 ^ n3522 ;
  assign n3561 = n3560 ^ n3559 ;
  assign n3564 = n1538 ^ n1535 ;
  assign n3562 = n3527 & ~n3547 ;
  assign n3563 = n3562 ^ n3526 ;
  assign n3565 = n3564 ^ n3563 ;
  assign n3566 = n1537 ^ n1536 ;
  assign n3567 = n3531 ^ n3528 ;
  assign n3568 = ~n3547 & n3567 ;
  assign n3569 = n3568 ^ n3528 ;
  assign n3570 = n3566 & ~n3569 ;
  assign n3571 = n3570 ^ n3563 ;
  assign n3572 = ~n3565 & ~n3571 ;
  assign n3573 = n3572 ^ n3563 ;
  assign n3574 = n3573 ^ n3559 ;
  assign n3575 = ~n3561 & n3574 ;
  assign n3576 = n3575 ^ n3559 ;
  assign n3577 = n3576 ^ n3554 ;
  assign n3578 = ~n3557 & ~n3577 ;
  assign n3579 = n3578 ^ n3554 ;
  assign n3580 = ~n3553 & ~n3579 ;
  assign n3581 = ~n3552 & ~n3580 ;
  assign n3582 = ~n3074 & ~n3581 ;
  assign n3583 = n3550 & n3582 ;
  assign n3584 = n3583 ^ n3549 ;
  assign n3259 = n1378 ^ n1375 ;
  assign n3585 = n3584 ^ n3259 ;
  assign n3586 = n3075 ^ n1379 ;
  assign n3615 = n3259 ^ n1379 ;
  assign n3588 = n3557 & ~n3582 ;
  assign n3589 = n3588 ^ n3554 ;
  assign n3587 = n1374 ^ n1367 ;
  assign n3590 = n3589 ^ n3587 ;
  assign n3593 = n1373 ^ n1372 ;
  assign n3591 = n3561 & ~n3582 ;
  assign n3592 = n3591 ^ n3560 ;
  assign n3594 = n3593 ^ n3592 ;
  assign n3597 = n1371 ^ n1368 ;
  assign n3595 = n3565 & ~n3582 ;
  assign n3596 = n3595 ^ n3564 ;
  assign n3598 = n3597 ^ n3596 ;
  assign n3599 = n1370 ^ n1369 ;
  assign n3600 = n3569 ^ n3566 ;
  assign n3601 = ~n3582 & n3600 ;
  assign n3602 = n3601 ^ n3566 ;
  assign n3603 = n3599 & ~n3602 ;
  assign n3604 = n3603 ^ n3596 ;
  assign n3605 = ~n3598 & ~n3604 ;
  assign n3606 = n3605 ^ n3596 ;
  assign n3607 = n3606 ^ n3592 ;
  assign n3608 = ~n3594 & n3607 ;
  assign n3609 = n3608 ^ n3592 ;
  assign n3610 = n3609 ^ n3587 ;
  assign n3611 = ~n3590 & ~n3610 ;
  assign n3612 = n3611 ^ n3587 ;
  assign n3613 = n3612 ^ n3584 ;
  assign n3614 = ~n3585 & n3613 ;
  assign n3616 = n3615 ^ n3614 ;
  assign n3617 = ~n3586 & ~n3616 ;
  assign n3618 = n3617 ^ n3075 ;
  assign n3619 = n3585 & n3618 ;
  assign n3620 = n3619 ^ n3584 ;
  assign n3258 = n1211 ^ n1208 ;
  assign n3621 = n3620 ^ n3258 ;
  assign n3622 = ~n3258 & n3620 ;
  assign n3623 = n3622 ^ n3078 ;
  assign n3624 = n3622 ^ n3621 ;
  assign n3626 = n3590 & ~n3618 ;
  assign n3627 = n3626 ^ n3587 ;
  assign n3625 = n1207 ^ n1200 ;
  assign n3628 = n3627 ^ n3625 ;
  assign n3631 = n1206 ^ n1205 ;
  assign n3629 = n3594 & ~n3618 ;
  assign n3630 = n3629 ^ n3593 ;
  assign n3632 = n3631 ^ n3630 ;
  assign n3635 = n1204 ^ n1201 ;
  assign n3633 = n3598 & ~n3618 ;
  assign n3634 = n3633 ^ n3597 ;
  assign n3636 = n3635 ^ n3634 ;
  assign n3637 = n1203 ^ n1202 ;
  assign n3638 = n3602 ^ n3599 ;
  assign n3639 = ~n3618 & n3638 ;
  assign n3640 = n3639 ^ n3599 ;
  assign n3641 = n3637 & ~n3640 ;
  assign n3642 = n3641 ^ n3634 ;
  assign n3643 = ~n3636 & ~n3642 ;
  assign n3644 = n3643 ^ n3634 ;
  assign n3645 = n3644 ^ n3630 ;
  assign n3646 = ~n3632 & n3645 ;
  assign n3647 = n3646 ^ n3630 ;
  assign n3648 = n3647 ^ n3625 ;
  assign n3649 = ~n3628 & ~n3648 ;
  assign n3650 = n3649 ^ n3625 ;
  assign n3651 = ~n3624 & ~n3650 ;
  assign n3652 = ~n3623 & ~n3651 ;
  assign n3653 = ~n3079 & ~n3652 ;
  assign n3654 = n3621 & n3653 ;
  assign n3655 = n3654 ^ n3620 ;
  assign n3257 = n1044 ^ n1041 ;
  assign n3656 = n3655 ^ n3257 ;
  assign n3657 = n3080 ^ n1045 ;
  assign n3686 = n3257 ^ n1045 ;
  assign n3659 = n3628 & ~n3653 ;
  assign n3660 = n3659 ^ n3625 ;
  assign n3658 = n1040 ^ n1033 ;
  assign n3661 = n3660 ^ n3658 ;
  assign n3664 = n1039 ^ n1038 ;
  assign n3662 = n3632 & ~n3653 ;
  assign n3663 = n3662 ^ n3631 ;
  assign n3665 = n3664 ^ n3663 ;
  assign n3668 = n1037 ^ n1034 ;
  assign n3666 = n3636 & ~n3653 ;
  assign n3667 = n3666 ^ n3635 ;
  assign n3669 = n3668 ^ n3667 ;
  assign n3670 = n1036 ^ n1035 ;
  assign n3671 = n3640 ^ n3637 ;
  assign n3672 = ~n3653 & n3671 ;
  assign n3673 = n3672 ^ n3637 ;
  assign n3674 = n3670 & ~n3673 ;
  assign n3675 = n3674 ^ n3667 ;
  assign n3676 = ~n3669 & ~n3675 ;
  assign n3677 = n3676 ^ n3667 ;
  assign n3678 = n3677 ^ n3663 ;
  assign n3679 = ~n3665 & n3678 ;
  assign n3680 = n3679 ^ n3663 ;
  assign n3681 = n3680 ^ n3658 ;
  assign n3682 = ~n3661 & ~n3681 ;
  assign n3683 = n3682 ^ n3658 ;
  assign n3684 = n3683 ^ n3655 ;
  assign n3685 = ~n3656 & n3684 ;
  assign n3687 = n3686 ^ n3685 ;
  assign n3688 = ~n3657 & ~n3687 ;
  assign n3689 = n3688 ^ n3080 ;
  assign n3690 = n3656 & n3689 ;
  assign n3691 = n3690 ^ n3655 ;
  assign n3256 = n877 ^ n874 ;
  assign n3692 = n3691 ^ n3256 ;
  assign n3693 = ~n3256 & n3691 ;
  assign n3694 = n3693 ^ n3083 ;
  assign n3695 = n3693 ^ n3692 ;
  assign n3697 = n3661 & ~n3689 ;
  assign n3698 = n3697 ^ n3658 ;
  assign n3696 = n873 ^ n866 ;
  assign n3699 = n3698 ^ n3696 ;
  assign n3702 = n872 ^ n871 ;
  assign n3700 = n3665 & ~n3689 ;
  assign n3701 = n3700 ^ n3664 ;
  assign n3703 = n3702 ^ n3701 ;
  assign n3706 = n870 ^ n869 ;
  assign n3704 = n3669 & ~n3689 ;
  assign n3705 = n3704 ^ n3668 ;
  assign n3707 = n3706 ^ n3705 ;
  assign n3708 = n868 ^ n867 ;
  assign n3709 = n3673 ^ n3670 ;
  assign n3710 = ~n3689 & n3709 ;
  assign n3711 = n3710 ^ n3670 ;
  assign n3712 = n3708 & ~n3711 ;
  assign n3713 = n3712 ^ n3705 ;
  assign n3714 = ~n3707 & ~n3713 ;
  assign n3715 = n3714 ^ n3705 ;
  assign n3716 = n3715 ^ n3701 ;
  assign n3717 = ~n3703 & n3716 ;
  assign n3718 = n3717 ^ n3701 ;
  assign n3719 = n3718 ^ n3696 ;
  assign n3720 = ~n3699 & ~n3719 ;
  assign n3721 = n3720 ^ n3696 ;
  assign n3722 = ~n3695 & ~n3721 ;
  assign n3723 = ~n3694 & ~n3722 ;
  assign n3724 = ~n3084 & ~n3723 ;
  assign n3725 = n3692 & n3724 ;
  assign n3726 = n3725 ^ n3691 ;
  assign n3255 = n710 ^ n707 ;
  assign n3727 = n3726 ^ n3255 ;
  assign n3728 = n3085 ^ n711 ;
  assign n3757 = n3255 ^ n711 ;
  assign n3730 = n3699 & ~n3724 ;
  assign n3731 = n3730 ^ n3696 ;
  assign n3729 = n706 ^ n699 ;
  assign n3732 = n3731 ^ n3729 ;
  assign n3735 = n705 ^ n704 ;
  assign n3733 = n3703 & ~n3724 ;
  assign n3734 = n3733 ^ n3702 ;
  assign n3736 = n3735 ^ n3734 ;
  assign n3738 = n3707 & ~n3724 ;
  assign n3739 = n3738 ^ n3706 ;
  assign n3737 = n703 ^ n702 ;
  assign n3740 = n3739 ^ n3737 ;
  assign n3741 = n701 ^ n700 ;
  assign n3742 = n3711 ^ n3708 ;
  assign n3743 = ~n3724 & n3742 ;
  assign n3744 = n3743 ^ n3708 ;
  assign n3745 = n3741 & ~n3744 ;
  assign n3746 = n3745 ^ n3737 ;
  assign n3747 = ~n3740 & n3746 ;
  assign n3748 = n3747 ^ n3737 ;
  assign n3749 = n3748 ^ n3734 ;
  assign n3750 = ~n3736 & ~n3749 ;
  assign n3751 = n3750 ^ n3734 ;
  assign n3752 = n3751 ^ n3729 ;
  assign n3753 = ~n3732 & ~n3752 ;
  assign n3754 = n3753 ^ n3729 ;
  assign n3755 = n3754 ^ n3726 ;
  assign n3756 = ~n3727 & n3755 ;
  assign n3758 = n3757 ^ n3756 ;
  assign n3759 = ~n3728 & ~n3758 ;
  assign n3760 = n3759 ^ n3085 ;
  assign n3761 = n3727 & ~n3760 ;
  assign n3762 = n3761 ^ n3255 ;
  assign n3764 = n3763 ^ n3762 ;
  assign n3766 = n3732 & ~n3760 ;
  assign n3767 = n3766 ^ n3729 ;
  assign n3765 = n3248 ^ n3241 ;
  assign n3768 = n3767 ^ n3765 ;
  assign n3771 = n3247 ^ n3246 ;
  assign n3769 = n3736 & ~n3760 ;
  assign n3770 = n3769 ^ n3735 ;
  assign n3772 = n3771 ^ n3770 ;
  assign n3775 = n3245 ^ n3242 ;
  assign n3773 = n3740 & n3760 ;
  assign n3774 = n3773 ^ n3739 ;
  assign n3776 = n3775 ^ n3774 ;
  assign n3777 = n3244 ^ n3243 ;
  assign n3778 = n3744 ^ n3741 ;
  assign n3779 = n3760 & n3778 ;
  assign n3780 = n3779 ^ n3744 ;
  assign n3781 = n3777 & ~n3780 ;
  assign n3782 = n3781 ^ n3774 ;
  assign n3783 = ~n3776 & ~n3782 ;
  assign n3784 = n3783 ^ n3774 ;
  assign n3785 = n3784 ^ n3770 ;
  assign n3786 = ~n3772 & n3785 ;
  assign n3787 = n3786 ^ n3770 ;
  assign n3788 = n3787 ^ n3767 ;
  assign n3789 = ~n3768 & n3788 ;
  assign n3790 = n3789 ^ n3767 ;
  assign n3791 = n3790 ^ n3763 ;
  assign n3792 = ~n3764 & n3791 ;
  assign n3793 = n3792 ^ n3762 ;
  assign n3794 = n3793 ^ n3086 ;
  assign n3795 = ~n3254 & ~n3794 ;
  assign n3796 = n3795 ^ n3253 ;
  assign n3797 = x480 ^ x448 ;
  assign n3798 = ~n3301 & n3797 ;
  assign n3799 = n3798 ^ x448 ;
  assign n3800 = n3799 ^ x416 ;
  assign n3801 = n3333 & n3800 ;
  assign n3802 = n3801 ^ x416 ;
  assign n3803 = n3802 ^ x384 ;
  assign n3804 = ~n3369 & n3803 ;
  assign n3805 = n3804 ^ x384 ;
  assign n3806 = n3805 ^ x352 ;
  assign n3807 = ~n3405 & n3806 ;
  assign n3808 = n3807 ^ x352 ;
  assign n3809 = n3808 ^ x320 ;
  assign n3810 = ~n3440 & n3809 ;
  assign n3811 = n3810 ^ x320 ;
  assign n3812 = n3811 ^ x288 ;
  assign n3813 = ~n3476 & n3812 ;
  assign n3814 = n3813 ^ x288 ;
  assign n3815 = n3814 ^ x256 ;
  assign n3816 = ~n3511 & n3815 ;
  assign n3817 = n3816 ^ x256 ;
  assign n3818 = n3817 ^ x224 ;
  assign n3819 = ~n3547 & n3818 ;
  assign n3820 = n3819 ^ x224 ;
  assign n3821 = n3820 ^ x192 ;
  assign n3822 = ~n3582 & n3821 ;
  assign n3823 = n3822 ^ x192 ;
  assign n3824 = n3823 ^ x160 ;
  assign n3825 = ~n3618 & n3824 ;
  assign n3826 = n3825 ^ x160 ;
  assign n3827 = n3826 ^ x128 ;
  assign n3828 = ~n3653 & n3827 ;
  assign n3829 = n3828 ^ x128 ;
  assign n3830 = n3829 ^ x96 ;
  assign n3831 = ~n3689 & n3830 ;
  assign n3832 = n3831 ^ x96 ;
  assign n3833 = n3832 ^ x64 ;
  assign n3834 = ~n3724 & n3833 ;
  assign n3835 = n3834 ^ x64 ;
  assign n3836 = n3835 ^ x32 ;
  assign n3837 = ~n3760 & n3836 ;
  assign n3838 = n3837 ^ x32 ;
  assign n3839 = n3838 ^ x0 ;
  assign n3840 = n3796 & n3839 ;
  assign n3841 = n3840 ^ x0 ;
  assign n3842 = x481 ^ x449 ;
  assign n3843 = ~n3301 & n3842 ;
  assign n3844 = n3843 ^ x449 ;
  assign n3845 = n3844 ^ x417 ;
  assign n3846 = n3333 & n3845 ;
  assign n3847 = n3846 ^ x417 ;
  assign n3848 = n3847 ^ x385 ;
  assign n3849 = ~n3369 & n3848 ;
  assign n3850 = n3849 ^ x385 ;
  assign n3851 = n3850 ^ x353 ;
  assign n3852 = ~n3405 & n3851 ;
  assign n3853 = n3852 ^ x353 ;
  assign n3854 = n3853 ^ x321 ;
  assign n3855 = ~n3440 & n3854 ;
  assign n3856 = n3855 ^ x321 ;
  assign n3857 = n3856 ^ x289 ;
  assign n3858 = ~n3476 & n3857 ;
  assign n3859 = n3858 ^ x289 ;
  assign n3860 = n3859 ^ x257 ;
  assign n3861 = ~n3511 & n3860 ;
  assign n3862 = n3861 ^ x257 ;
  assign n3863 = n3862 ^ x225 ;
  assign n3864 = ~n3547 & n3863 ;
  assign n3865 = n3864 ^ x225 ;
  assign n3866 = n3865 ^ x193 ;
  assign n3867 = ~n3582 & n3866 ;
  assign n3868 = n3867 ^ x193 ;
  assign n3869 = n3868 ^ x161 ;
  assign n3870 = ~n3618 & n3869 ;
  assign n3871 = n3870 ^ x161 ;
  assign n3872 = n3871 ^ x129 ;
  assign n3873 = ~n3653 & n3872 ;
  assign n3874 = n3873 ^ x129 ;
  assign n3875 = n3874 ^ x97 ;
  assign n3876 = ~n3689 & n3875 ;
  assign n3877 = n3876 ^ x97 ;
  assign n3878 = n3877 ^ x65 ;
  assign n3879 = ~n3724 & n3878 ;
  assign n3880 = n3879 ^ x65 ;
  assign n3881 = n3880 ^ x33 ;
  assign n3882 = ~n3760 & n3881 ;
  assign n3883 = n3882 ^ x33 ;
  assign n3884 = n3883 ^ x1 ;
  assign n3885 = n3796 & n3884 ;
  assign n3886 = n3885 ^ x1 ;
  assign n3887 = x482 ^ x450 ;
  assign n3888 = ~n3301 & n3887 ;
  assign n3889 = n3888 ^ x450 ;
  assign n3890 = n3889 ^ x418 ;
  assign n3891 = n3333 & n3890 ;
  assign n3892 = n3891 ^ x418 ;
  assign n3893 = n3892 ^ x386 ;
  assign n3894 = ~n3369 & n3893 ;
  assign n3895 = n3894 ^ x386 ;
  assign n3896 = n3895 ^ x354 ;
  assign n3897 = ~n3405 & n3896 ;
  assign n3898 = n3897 ^ x354 ;
  assign n3899 = n3898 ^ x322 ;
  assign n3900 = ~n3440 & n3899 ;
  assign n3901 = n3900 ^ x322 ;
  assign n3902 = n3901 ^ x290 ;
  assign n3903 = ~n3476 & n3902 ;
  assign n3904 = n3903 ^ x290 ;
  assign n3905 = n3904 ^ x258 ;
  assign n3906 = ~n3511 & n3905 ;
  assign n3907 = n3906 ^ x258 ;
  assign n3908 = n3907 ^ x226 ;
  assign n3909 = ~n3547 & n3908 ;
  assign n3910 = n3909 ^ x226 ;
  assign n3911 = n3910 ^ x194 ;
  assign n3912 = ~n3582 & n3911 ;
  assign n3913 = n3912 ^ x194 ;
  assign n3914 = n3913 ^ x162 ;
  assign n3915 = ~n3618 & n3914 ;
  assign n3916 = n3915 ^ x162 ;
  assign n3917 = n3916 ^ x130 ;
  assign n3918 = ~n3653 & n3917 ;
  assign n3919 = n3918 ^ x130 ;
  assign n3920 = n3919 ^ x98 ;
  assign n3921 = ~n3689 & n3920 ;
  assign n3922 = n3921 ^ x98 ;
  assign n3923 = n3922 ^ x66 ;
  assign n3924 = ~n3724 & n3923 ;
  assign n3925 = n3924 ^ x66 ;
  assign n3926 = n3925 ^ x34 ;
  assign n3927 = ~n3760 & n3926 ;
  assign n3928 = n3927 ^ x34 ;
  assign n3929 = n3928 ^ x2 ;
  assign n3930 = n3796 & n3929 ;
  assign n3931 = n3930 ^ x2 ;
  assign n3932 = x483 ^ x451 ;
  assign n3933 = ~n3301 & n3932 ;
  assign n3934 = n3933 ^ x451 ;
  assign n3935 = n3934 ^ x419 ;
  assign n3936 = n3333 & n3935 ;
  assign n3937 = n3936 ^ x419 ;
  assign n3938 = n3937 ^ x387 ;
  assign n3939 = ~n3369 & n3938 ;
  assign n3940 = n3939 ^ x387 ;
  assign n3941 = n3940 ^ x355 ;
  assign n3942 = ~n3405 & n3941 ;
  assign n3943 = n3942 ^ x355 ;
  assign n3944 = n3943 ^ x323 ;
  assign n3945 = ~n3440 & n3944 ;
  assign n3946 = n3945 ^ x323 ;
  assign n3947 = n3946 ^ x291 ;
  assign n3948 = ~n3476 & n3947 ;
  assign n3949 = n3948 ^ x291 ;
  assign n3950 = n3949 ^ x259 ;
  assign n3951 = ~n3511 & n3950 ;
  assign n3952 = n3951 ^ x259 ;
  assign n3953 = n3952 ^ x227 ;
  assign n3954 = ~n3547 & n3953 ;
  assign n3955 = n3954 ^ x227 ;
  assign n3956 = n3955 ^ x195 ;
  assign n3957 = ~n3582 & n3956 ;
  assign n3958 = n3957 ^ x195 ;
  assign n3959 = n3958 ^ x163 ;
  assign n3960 = ~n3618 & n3959 ;
  assign n3961 = n3960 ^ x163 ;
  assign n3962 = n3961 ^ x131 ;
  assign n3963 = ~n3653 & n3962 ;
  assign n3964 = n3963 ^ x131 ;
  assign n3965 = n3964 ^ x99 ;
  assign n3966 = ~n3689 & n3965 ;
  assign n3967 = n3966 ^ x99 ;
  assign n3968 = n3967 ^ x67 ;
  assign n3969 = ~n3724 & n3968 ;
  assign n3970 = n3969 ^ x67 ;
  assign n3971 = n3970 ^ x35 ;
  assign n3972 = ~n3760 & n3971 ;
  assign n3973 = n3972 ^ x35 ;
  assign n3974 = n3973 ^ x3 ;
  assign n3975 = n3796 & n3974 ;
  assign n3976 = n3975 ^ x3 ;
  assign n3977 = x484 ^ x452 ;
  assign n3978 = ~n3301 & n3977 ;
  assign n3979 = n3978 ^ x452 ;
  assign n3980 = n3979 ^ x420 ;
  assign n3981 = n3333 & n3980 ;
  assign n3982 = n3981 ^ x420 ;
  assign n3983 = n3982 ^ x388 ;
  assign n3984 = ~n3369 & n3983 ;
  assign n3985 = n3984 ^ x388 ;
  assign n3986 = n3985 ^ x356 ;
  assign n3987 = ~n3405 & n3986 ;
  assign n3988 = n3987 ^ x356 ;
  assign n3989 = n3988 ^ x324 ;
  assign n3990 = ~n3440 & n3989 ;
  assign n3991 = n3990 ^ x324 ;
  assign n3992 = n3991 ^ x292 ;
  assign n3993 = ~n3476 & n3992 ;
  assign n3994 = n3993 ^ x292 ;
  assign n3995 = n3994 ^ x260 ;
  assign n3996 = ~n3511 & n3995 ;
  assign n3997 = n3996 ^ x260 ;
  assign n3998 = n3997 ^ x228 ;
  assign n3999 = ~n3547 & n3998 ;
  assign n4000 = n3999 ^ x228 ;
  assign n4001 = n4000 ^ x196 ;
  assign n4002 = ~n3582 & n4001 ;
  assign n4003 = n4002 ^ x196 ;
  assign n4004 = n4003 ^ x164 ;
  assign n4005 = ~n3618 & n4004 ;
  assign n4006 = n4005 ^ x164 ;
  assign n4007 = n4006 ^ x132 ;
  assign n4008 = ~n3653 & n4007 ;
  assign n4009 = n4008 ^ x132 ;
  assign n4010 = n4009 ^ x100 ;
  assign n4011 = ~n3689 & n4010 ;
  assign n4012 = n4011 ^ x100 ;
  assign n4013 = n4012 ^ x68 ;
  assign n4014 = ~n3724 & n4013 ;
  assign n4015 = n4014 ^ x68 ;
  assign n4016 = n4015 ^ x36 ;
  assign n4017 = ~n3760 & n4016 ;
  assign n4018 = n4017 ^ x36 ;
  assign n4019 = n4018 ^ x4 ;
  assign n4020 = n3796 & n4019 ;
  assign n4021 = n4020 ^ x4 ;
  assign n4022 = x485 ^ x453 ;
  assign n4023 = ~n3301 & n4022 ;
  assign n4024 = n4023 ^ x453 ;
  assign n4025 = n4024 ^ x421 ;
  assign n4026 = n3333 & n4025 ;
  assign n4027 = n4026 ^ x421 ;
  assign n4028 = n4027 ^ x389 ;
  assign n4029 = ~n3369 & n4028 ;
  assign n4030 = n4029 ^ x389 ;
  assign n4031 = n4030 ^ x357 ;
  assign n4032 = ~n3405 & n4031 ;
  assign n4033 = n4032 ^ x357 ;
  assign n4034 = n4033 ^ x325 ;
  assign n4035 = ~n3440 & n4034 ;
  assign n4036 = n4035 ^ x325 ;
  assign n4037 = n4036 ^ x293 ;
  assign n4038 = ~n3476 & n4037 ;
  assign n4039 = n4038 ^ x293 ;
  assign n4040 = n4039 ^ x261 ;
  assign n4041 = ~n3511 & n4040 ;
  assign n4042 = n4041 ^ x261 ;
  assign n4043 = n4042 ^ x229 ;
  assign n4044 = ~n3547 & n4043 ;
  assign n4045 = n4044 ^ x229 ;
  assign n4046 = n4045 ^ x197 ;
  assign n4047 = ~n3582 & n4046 ;
  assign n4048 = n4047 ^ x197 ;
  assign n4049 = n4048 ^ x165 ;
  assign n4050 = ~n3618 & n4049 ;
  assign n4051 = n4050 ^ x165 ;
  assign n4052 = n4051 ^ x133 ;
  assign n4053 = ~n3653 & n4052 ;
  assign n4054 = n4053 ^ x133 ;
  assign n4055 = n4054 ^ x101 ;
  assign n4056 = ~n3689 & n4055 ;
  assign n4057 = n4056 ^ x101 ;
  assign n4058 = n4057 ^ x69 ;
  assign n4059 = ~n3724 & n4058 ;
  assign n4060 = n4059 ^ x69 ;
  assign n4061 = n4060 ^ x37 ;
  assign n4062 = ~n3760 & n4061 ;
  assign n4063 = n4062 ^ x37 ;
  assign n4064 = n4063 ^ x5 ;
  assign n4065 = n3796 & n4064 ;
  assign n4066 = n4065 ^ x5 ;
  assign n4067 = x486 ^ x454 ;
  assign n4068 = ~n3301 & n4067 ;
  assign n4069 = n4068 ^ x454 ;
  assign n4070 = n4069 ^ x422 ;
  assign n4071 = n3333 & n4070 ;
  assign n4072 = n4071 ^ x422 ;
  assign n4073 = n4072 ^ x390 ;
  assign n4074 = ~n3369 & n4073 ;
  assign n4075 = n4074 ^ x390 ;
  assign n4076 = n4075 ^ x358 ;
  assign n4077 = ~n3405 & n4076 ;
  assign n4078 = n4077 ^ x358 ;
  assign n4079 = n4078 ^ x326 ;
  assign n4080 = ~n3440 & n4079 ;
  assign n4081 = n4080 ^ x326 ;
  assign n4082 = n4081 ^ x294 ;
  assign n4083 = ~n3476 & n4082 ;
  assign n4084 = n4083 ^ x294 ;
  assign n4085 = n4084 ^ x262 ;
  assign n4086 = ~n3511 & n4085 ;
  assign n4087 = n4086 ^ x262 ;
  assign n4088 = n4087 ^ x230 ;
  assign n4089 = ~n3547 & n4088 ;
  assign n4090 = n4089 ^ x230 ;
  assign n4091 = n4090 ^ x198 ;
  assign n4092 = ~n3582 & n4091 ;
  assign n4093 = n4092 ^ x198 ;
  assign n4094 = n4093 ^ x166 ;
  assign n4095 = ~n3618 & n4094 ;
  assign n4096 = n4095 ^ x166 ;
  assign n4097 = n4096 ^ x134 ;
  assign n4098 = ~n3653 & n4097 ;
  assign n4099 = n4098 ^ x134 ;
  assign n4100 = n4099 ^ x102 ;
  assign n4101 = ~n3689 & n4100 ;
  assign n4102 = n4101 ^ x102 ;
  assign n4103 = n4102 ^ x70 ;
  assign n4104 = ~n3724 & n4103 ;
  assign n4105 = n4104 ^ x70 ;
  assign n4106 = n4105 ^ x38 ;
  assign n4107 = ~n3760 & n4106 ;
  assign n4108 = n4107 ^ x38 ;
  assign n4109 = n4108 ^ x6 ;
  assign n4110 = n3796 & n4109 ;
  assign n4111 = n4110 ^ x6 ;
  assign n4112 = x487 ^ x455 ;
  assign n4113 = ~n3301 & n4112 ;
  assign n4114 = n4113 ^ x455 ;
  assign n4115 = n4114 ^ x423 ;
  assign n4116 = n3333 & n4115 ;
  assign n4117 = n4116 ^ x423 ;
  assign n4118 = n4117 ^ x391 ;
  assign n4119 = ~n3369 & n4118 ;
  assign n4120 = n4119 ^ x391 ;
  assign n4121 = n4120 ^ x359 ;
  assign n4122 = ~n3405 & n4121 ;
  assign n4123 = n4122 ^ x359 ;
  assign n4124 = n4123 ^ x327 ;
  assign n4125 = ~n3440 & n4124 ;
  assign n4126 = n4125 ^ x327 ;
  assign n4127 = n4126 ^ x295 ;
  assign n4128 = ~n3476 & n4127 ;
  assign n4129 = n4128 ^ x295 ;
  assign n4130 = n4129 ^ x263 ;
  assign n4131 = ~n3511 & n4130 ;
  assign n4132 = n4131 ^ x263 ;
  assign n4133 = n4132 ^ x231 ;
  assign n4134 = ~n3547 & n4133 ;
  assign n4135 = n4134 ^ x231 ;
  assign n4136 = n4135 ^ x199 ;
  assign n4137 = ~n3582 & n4136 ;
  assign n4138 = n4137 ^ x199 ;
  assign n4139 = n4138 ^ x167 ;
  assign n4140 = ~n3618 & n4139 ;
  assign n4141 = n4140 ^ x167 ;
  assign n4142 = n4141 ^ x135 ;
  assign n4143 = ~n3653 & n4142 ;
  assign n4144 = n4143 ^ x135 ;
  assign n4145 = n4144 ^ x103 ;
  assign n4146 = ~n3689 & n4145 ;
  assign n4147 = n4146 ^ x103 ;
  assign n4148 = n4147 ^ x71 ;
  assign n4149 = ~n3724 & n4148 ;
  assign n4150 = n4149 ^ x71 ;
  assign n4151 = n4150 ^ x39 ;
  assign n4152 = ~n3760 & n4151 ;
  assign n4153 = n4152 ^ x39 ;
  assign n4154 = n4153 ^ x7 ;
  assign n4155 = n3796 & n4154 ;
  assign n4156 = n4155 ^ x7 ;
  assign n4157 = x488 ^ x456 ;
  assign n4158 = ~n3301 & n4157 ;
  assign n4159 = n4158 ^ x456 ;
  assign n4160 = n4159 ^ x424 ;
  assign n4161 = n3333 & n4160 ;
  assign n4162 = n4161 ^ x424 ;
  assign n4163 = n4162 ^ x392 ;
  assign n4164 = ~n3369 & n4163 ;
  assign n4165 = n4164 ^ x392 ;
  assign n4166 = n4165 ^ x360 ;
  assign n4167 = ~n3405 & n4166 ;
  assign n4168 = n4167 ^ x360 ;
  assign n4169 = n4168 ^ x328 ;
  assign n4170 = ~n3440 & n4169 ;
  assign n4171 = n4170 ^ x328 ;
  assign n4172 = n4171 ^ x296 ;
  assign n4173 = ~n3476 & n4172 ;
  assign n4174 = n4173 ^ x296 ;
  assign n4175 = n4174 ^ x264 ;
  assign n4176 = ~n3511 & n4175 ;
  assign n4177 = n4176 ^ x264 ;
  assign n4178 = n4177 ^ x232 ;
  assign n4179 = ~n3547 & n4178 ;
  assign n4180 = n4179 ^ x232 ;
  assign n4181 = n4180 ^ x200 ;
  assign n4182 = ~n3582 & n4181 ;
  assign n4183 = n4182 ^ x200 ;
  assign n4184 = n4183 ^ x168 ;
  assign n4185 = ~n3618 & n4184 ;
  assign n4186 = n4185 ^ x168 ;
  assign n4187 = n4186 ^ x136 ;
  assign n4188 = ~n3653 & n4187 ;
  assign n4189 = n4188 ^ x136 ;
  assign n4190 = n4189 ^ x104 ;
  assign n4191 = ~n3689 & n4190 ;
  assign n4192 = n4191 ^ x104 ;
  assign n4193 = n4192 ^ x72 ;
  assign n4194 = ~n3724 & n4193 ;
  assign n4195 = n4194 ^ x72 ;
  assign n4196 = n4195 ^ x40 ;
  assign n4197 = ~n3760 & n4196 ;
  assign n4198 = n4197 ^ x40 ;
  assign n4199 = n4198 ^ x8 ;
  assign n4200 = n3796 & n4199 ;
  assign n4201 = n4200 ^ x8 ;
  assign n4202 = x489 ^ x457 ;
  assign n4203 = ~n3301 & n4202 ;
  assign n4204 = n4203 ^ x457 ;
  assign n4205 = n4204 ^ x425 ;
  assign n4206 = n3333 & n4205 ;
  assign n4207 = n4206 ^ x425 ;
  assign n4208 = n4207 ^ x393 ;
  assign n4209 = ~n3369 & n4208 ;
  assign n4210 = n4209 ^ x393 ;
  assign n4211 = n4210 ^ x361 ;
  assign n4212 = ~n3405 & n4211 ;
  assign n4213 = n4212 ^ x361 ;
  assign n4214 = n4213 ^ x329 ;
  assign n4215 = ~n3440 & n4214 ;
  assign n4216 = n4215 ^ x329 ;
  assign n4217 = n4216 ^ x297 ;
  assign n4218 = ~n3476 & n4217 ;
  assign n4219 = n4218 ^ x297 ;
  assign n4220 = n4219 ^ x265 ;
  assign n4221 = ~n3511 & n4220 ;
  assign n4222 = n4221 ^ x265 ;
  assign n4223 = n4222 ^ x233 ;
  assign n4224 = ~n3547 & n4223 ;
  assign n4225 = n4224 ^ x233 ;
  assign n4226 = n4225 ^ x201 ;
  assign n4227 = ~n3582 & n4226 ;
  assign n4228 = n4227 ^ x201 ;
  assign n4229 = n4228 ^ x169 ;
  assign n4230 = ~n3618 & n4229 ;
  assign n4231 = n4230 ^ x169 ;
  assign n4232 = n4231 ^ x137 ;
  assign n4233 = ~n3653 & n4232 ;
  assign n4234 = n4233 ^ x137 ;
  assign n4235 = n4234 ^ x105 ;
  assign n4236 = ~n3689 & n4235 ;
  assign n4237 = n4236 ^ x105 ;
  assign n4238 = n4237 ^ x73 ;
  assign n4239 = ~n3724 & n4238 ;
  assign n4240 = n4239 ^ x73 ;
  assign n4241 = n4240 ^ x41 ;
  assign n4242 = ~n3760 & n4241 ;
  assign n4243 = n4242 ^ x41 ;
  assign n4244 = n4243 ^ x9 ;
  assign n4245 = n3796 & n4244 ;
  assign n4246 = n4245 ^ x9 ;
  assign n4247 = x490 ^ x458 ;
  assign n4248 = ~n3301 & n4247 ;
  assign n4249 = n4248 ^ x458 ;
  assign n4250 = n4249 ^ x426 ;
  assign n4251 = n3333 & n4250 ;
  assign n4252 = n4251 ^ x426 ;
  assign n4253 = n4252 ^ x394 ;
  assign n4254 = ~n3369 & n4253 ;
  assign n4255 = n4254 ^ x394 ;
  assign n4256 = n4255 ^ x362 ;
  assign n4257 = ~n3405 & n4256 ;
  assign n4258 = n4257 ^ x362 ;
  assign n4259 = n4258 ^ x330 ;
  assign n4260 = ~n3440 & n4259 ;
  assign n4261 = n4260 ^ x330 ;
  assign n4262 = n4261 ^ x298 ;
  assign n4263 = ~n3476 & n4262 ;
  assign n4264 = n4263 ^ x298 ;
  assign n4265 = n4264 ^ x266 ;
  assign n4266 = ~n3511 & n4265 ;
  assign n4267 = n4266 ^ x266 ;
  assign n4268 = n4267 ^ x234 ;
  assign n4269 = ~n3547 & n4268 ;
  assign n4270 = n4269 ^ x234 ;
  assign n4271 = n4270 ^ x202 ;
  assign n4272 = ~n3582 & n4271 ;
  assign n4273 = n4272 ^ x202 ;
  assign n4274 = n4273 ^ x170 ;
  assign n4275 = ~n3618 & n4274 ;
  assign n4276 = n4275 ^ x170 ;
  assign n4277 = n4276 ^ x138 ;
  assign n4278 = ~n3653 & n4277 ;
  assign n4279 = n4278 ^ x138 ;
  assign n4280 = n4279 ^ x106 ;
  assign n4281 = ~n3689 & n4280 ;
  assign n4282 = n4281 ^ x106 ;
  assign n4283 = n4282 ^ x74 ;
  assign n4284 = ~n3724 & n4283 ;
  assign n4285 = n4284 ^ x74 ;
  assign n4286 = n4285 ^ x42 ;
  assign n4287 = ~n3760 & n4286 ;
  assign n4288 = n4287 ^ x42 ;
  assign n4289 = n4288 ^ x10 ;
  assign n4290 = n3796 & n4289 ;
  assign n4291 = n4290 ^ x10 ;
  assign n4292 = x491 ^ x459 ;
  assign n4293 = ~n3301 & n4292 ;
  assign n4294 = n4293 ^ x459 ;
  assign n4295 = n4294 ^ x427 ;
  assign n4296 = n3333 & n4295 ;
  assign n4297 = n4296 ^ x427 ;
  assign n4298 = n4297 ^ x395 ;
  assign n4299 = ~n3369 & n4298 ;
  assign n4300 = n4299 ^ x395 ;
  assign n4301 = n4300 ^ x363 ;
  assign n4302 = ~n3405 & n4301 ;
  assign n4303 = n4302 ^ x363 ;
  assign n4304 = n4303 ^ x331 ;
  assign n4305 = ~n3440 & n4304 ;
  assign n4306 = n4305 ^ x331 ;
  assign n4307 = n4306 ^ x299 ;
  assign n4308 = ~n3476 & n4307 ;
  assign n4309 = n4308 ^ x299 ;
  assign n4310 = n4309 ^ x267 ;
  assign n4311 = ~n3511 & n4310 ;
  assign n4312 = n4311 ^ x267 ;
  assign n4313 = n4312 ^ x235 ;
  assign n4314 = ~n3547 & n4313 ;
  assign n4315 = n4314 ^ x235 ;
  assign n4316 = n4315 ^ x203 ;
  assign n4317 = ~n3582 & n4316 ;
  assign n4318 = n4317 ^ x203 ;
  assign n4319 = n4318 ^ x171 ;
  assign n4320 = ~n3618 & n4319 ;
  assign n4321 = n4320 ^ x171 ;
  assign n4322 = n4321 ^ x139 ;
  assign n4323 = ~n3653 & n4322 ;
  assign n4324 = n4323 ^ x139 ;
  assign n4325 = n4324 ^ x107 ;
  assign n4326 = ~n3689 & n4325 ;
  assign n4327 = n4326 ^ x107 ;
  assign n4328 = n4327 ^ x75 ;
  assign n4329 = ~n3724 & n4328 ;
  assign n4330 = n4329 ^ x75 ;
  assign n4331 = n4330 ^ x43 ;
  assign n4332 = ~n3760 & n4331 ;
  assign n4333 = n4332 ^ x43 ;
  assign n4334 = n4333 ^ x11 ;
  assign n4335 = n3796 & n4334 ;
  assign n4336 = n4335 ^ x11 ;
  assign n4337 = x492 ^ x460 ;
  assign n4338 = ~n3301 & n4337 ;
  assign n4339 = n4338 ^ x460 ;
  assign n4340 = n4339 ^ x428 ;
  assign n4341 = n3333 & n4340 ;
  assign n4342 = n4341 ^ x428 ;
  assign n4343 = n4342 ^ x396 ;
  assign n4344 = ~n3369 & n4343 ;
  assign n4345 = n4344 ^ x396 ;
  assign n4346 = n4345 ^ x364 ;
  assign n4347 = ~n3405 & n4346 ;
  assign n4348 = n4347 ^ x364 ;
  assign n4349 = n4348 ^ x332 ;
  assign n4350 = ~n3440 & n4349 ;
  assign n4351 = n4350 ^ x332 ;
  assign n4352 = n4351 ^ x300 ;
  assign n4353 = ~n3476 & n4352 ;
  assign n4354 = n4353 ^ x300 ;
  assign n4355 = n4354 ^ x268 ;
  assign n4356 = ~n3511 & n4355 ;
  assign n4357 = n4356 ^ x268 ;
  assign n4358 = n4357 ^ x236 ;
  assign n4359 = ~n3547 & n4358 ;
  assign n4360 = n4359 ^ x236 ;
  assign n4361 = n4360 ^ x204 ;
  assign n4362 = ~n3582 & n4361 ;
  assign n4363 = n4362 ^ x204 ;
  assign n4364 = n4363 ^ x172 ;
  assign n4365 = ~n3618 & n4364 ;
  assign n4366 = n4365 ^ x172 ;
  assign n4367 = n4366 ^ x140 ;
  assign n4368 = ~n3653 & n4367 ;
  assign n4369 = n4368 ^ x140 ;
  assign n4370 = n4369 ^ x108 ;
  assign n4371 = ~n3689 & n4370 ;
  assign n4372 = n4371 ^ x108 ;
  assign n4373 = n4372 ^ x76 ;
  assign n4374 = ~n3724 & n4373 ;
  assign n4375 = n4374 ^ x76 ;
  assign n4376 = n4375 ^ x44 ;
  assign n4377 = ~n3760 & n4376 ;
  assign n4378 = n4377 ^ x44 ;
  assign n4379 = n4378 ^ x12 ;
  assign n4380 = n3796 & n4379 ;
  assign n4381 = n4380 ^ x12 ;
  assign n4382 = x493 ^ x461 ;
  assign n4383 = ~n3301 & n4382 ;
  assign n4384 = n4383 ^ x461 ;
  assign n4385 = n4384 ^ x429 ;
  assign n4386 = n3333 & n4385 ;
  assign n4387 = n4386 ^ x429 ;
  assign n4388 = n4387 ^ x397 ;
  assign n4389 = ~n3369 & n4388 ;
  assign n4390 = n4389 ^ x397 ;
  assign n4391 = n4390 ^ x365 ;
  assign n4392 = ~n3405 & n4391 ;
  assign n4393 = n4392 ^ x365 ;
  assign n4394 = n4393 ^ x333 ;
  assign n4395 = ~n3440 & n4394 ;
  assign n4396 = n4395 ^ x333 ;
  assign n4397 = n4396 ^ x301 ;
  assign n4398 = ~n3476 & n4397 ;
  assign n4399 = n4398 ^ x301 ;
  assign n4400 = n4399 ^ x269 ;
  assign n4401 = ~n3511 & n4400 ;
  assign n4402 = n4401 ^ x269 ;
  assign n4403 = n4402 ^ x237 ;
  assign n4404 = ~n3547 & n4403 ;
  assign n4405 = n4404 ^ x237 ;
  assign n4406 = n4405 ^ x205 ;
  assign n4407 = ~n3582 & n4406 ;
  assign n4408 = n4407 ^ x205 ;
  assign n4409 = n4408 ^ x173 ;
  assign n4410 = ~n3618 & n4409 ;
  assign n4411 = n4410 ^ x173 ;
  assign n4412 = n4411 ^ x141 ;
  assign n4413 = ~n3653 & n4412 ;
  assign n4414 = n4413 ^ x141 ;
  assign n4415 = n4414 ^ x109 ;
  assign n4416 = ~n3689 & n4415 ;
  assign n4417 = n4416 ^ x109 ;
  assign n4418 = n4417 ^ x77 ;
  assign n4419 = ~n3724 & n4418 ;
  assign n4420 = n4419 ^ x77 ;
  assign n4421 = n4420 ^ x45 ;
  assign n4422 = ~n3760 & n4421 ;
  assign n4423 = n4422 ^ x45 ;
  assign n4424 = n4423 ^ x13 ;
  assign n4425 = n3796 & n4424 ;
  assign n4426 = n4425 ^ x13 ;
  assign n4427 = x494 ^ x462 ;
  assign n4428 = ~n3301 & n4427 ;
  assign n4429 = n4428 ^ x462 ;
  assign n4430 = n4429 ^ x430 ;
  assign n4431 = n3333 & n4430 ;
  assign n4432 = n4431 ^ x430 ;
  assign n4433 = n4432 ^ x398 ;
  assign n4434 = ~n3369 & n4433 ;
  assign n4435 = n4434 ^ x398 ;
  assign n4436 = n4435 ^ x366 ;
  assign n4437 = ~n3405 & n4436 ;
  assign n4438 = n4437 ^ x366 ;
  assign n4439 = n4438 ^ x334 ;
  assign n4440 = ~n3440 & n4439 ;
  assign n4441 = n4440 ^ x334 ;
  assign n4442 = n4441 ^ x302 ;
  assign n4443 = ~n3476 & n4442 ;
  assign n4444 = n4443 ^ x302 ;
  assign n4445 = n4444 ^ x270 ;
  assign n4446 = ~n3511 & n4445 ;
  assign n4447 = n4446 ^ x270 ;
  assign n4448 = n4447 ^ x238 ;
  assign n4449 = ~n3547 & n4448 ;
  assign n4450 = n4449 ^ x238 ;
  assign n4451 = n4450 ^ x206 ;
  assign n4452 = ~n3582 & n4451 ;
  assign n4453 = n4452 ^ x206 ;
  assign n4454 = n4453 ^ x174 ;
  assign n4455 = ~n3618 & n4454 ;
  assign n4456 = n4455 ^ x174 ;
  assign n4457 = n4456 ^ x142 ;
  assign n4458 = ~n3653 & n4457 ;
  assign n4459 = n4458 ^ x142 ;
  assign n4460 = n4459 ^ x110 ;
  assign n4461 = ~n3689 & n4460 ;
  assign n4462 = n4461 ^ x110 ;
  assign n4463 = n4462 ^ x78 ;
  assign n4464 = ~n3724 & n4463 ;
  assign n4465 = n4464 ^ x78 ;
  assign n4466 = n4465 ^ x46 ;
  assign n4467 = ~n3760 & n4466 ;
  assign n4468 = n4467 ^ x46 ;
  assign n4469 = n4468 ^ x14 ;
  assign n4470 = n3796 & n4469 ;
  assign n4471 = n4470 ^ x14 ;
  assign n4472 = x495 ^ x463 ;
  assign n4473 = ~n3301 & n4472 ;
  assign n4474 = n4473 ^ x463 ;
  assign n4475 = n4474 ^ x431 ;
  assign n4476 = n3333 & n4475 ;
  assign n4477 = n4476 ^ x431 ;
  assign n4478 = n4477 ^ x399 ;
  assign n4479 = ~n3369 & n4478 ;
  assign n4480 = n4479 ^ x399 ;
  assign n4481 = n4480 ^ x367 ;
  assign n4482 = ~n3405 & n4481 ;
  assign n4483 = n4482 ^ x367 ;
  assign n4484 = n4483 ^ x335 ;
  assign n4485 = ~n3440 & n4484 ;
  assign n4486 = n4485 ^ x335 ;
  assign n4487 = n4486 ^ x303 ;
  assign n4488 = ~n3476 & n4487 ;
  assign n4489 = n4488 ^ x303 ;
  assign n4490 = n4489 ^ x271 ;
  assign n4491 = ~n3511 & n4490 ;
  assign n4492 = n4491 ^ x271 ;
  assign n4493 = n4492 ^ x239 ;
  assign n4494 = ~n3547 & n4493 ;
  assign n4495 = n4494 ^ x239 ;
  assign n4496 = n4495 ^ x207 ;
  assign n4497 = ~n3582 & n4496 ;
  assign n4498 = n4497 ^ x207 ;
  assign n4499 = n4498 ^ x175 ;
  assign n4500 = ~n3618 & n4499 ;
  assign n4501 = n4500 ^ x175 ;
  assign n4502 = n4501 ^ x143 ;
  assign n4503 = ~n3653 & n4502 ;
  assign n4504 = n4503 ^ x143 ;
  assign n4505 = n4504 ^ x111 ;
  assign n4506 = ~n3689 & n4505 ;
  assign n4507 = n4506 ^ x111 ;
  assign n4508 = n4507 ^ x79 ;
  assign n4509 = ~n3724 & n4508 ;
  assign n4510 = n4509 ^ x79 ;
  assign n4511 = n4510 ^ x47 ;
  assign n4512 = ~n3760 & n4511 ;
  assign n4513 = n4512 ^ x47 ;
  assign n4514 = n4513 ^ x15 ;
  assign n4515 = n3796 & n4514 ;
  assign n4516 = n4515 ^ x15 ;
  assign n4517 = x496 ^ x464 ;
  assign n4518 = ~n3301 & n4517 ;
  assign n4519 = n4518 ^ x464 ;
  assign n4520 = n4519 ^ x432 ;
  assign n4521 = n3333 & n4520 ;
  assign n4522 = n4521 ^ x432 ;
  assign n4523 = n4522 ^ x400 ;
  assign n4524 = ~n3369 & n4523 ;
  assign n4525 = n4524 ^ x400 ;
  assign n4526 = n4525 ^ x368 ;
  assign n4527 = ~n3405 & n4526 ;
  assign n4528 = n4527 ^ x368 ;
  assign n4529 = n4528 ^ x336 ;
  assign n4530 = ~n3440 & n4529 ;
  assign n4531 = n4530 ^ x336 ;
  assign n4532 = n4531 ^ x304 ;
  assign n4533 = ~n3476 & n4532 ;
  assign n4534 = n4533 ^ x304 ;
  assign n4535 = n4534 ^ x272 ;
  assign n4536 = ~n3511 & n4535 ;
  assign n4537 = n4536 ^ x272 ;
  assign n4538 = n4537 ^ x240 ;
  assign n4539 = ~n3547 & n4538 ;
  assign n4540 = n4539 ^ x240 ;
  assign n4541 = n4540 ^ x208 ;
  assign n4542 = ~n3582 & n4541 ;
  assign n4543 = n4542 ^ x208 ;
  assign n4544 = n4543 ^ x176 ;
  assign n4545 = ~n3618 & n4544 ;
  assign n4546 = n4545 ^ x176 ;
  assign n4547 = n4546 ^ x144 ;
  assign n4548 = ~n3653 & n4547 ;
  assign n4549 = n4548 ^ x144 ;
  assign n4550 = n4549 ^ x112 ;
  assign n4551 = ~n3689 & n4550 ;
  assign n4552 = n4551 ^ x112 ;
  assign n4553 = n4552 ^ x80 ;
  assign n4554 = ~n3724 & n4553 ;
  assign n4555 = n4554 ^ x80 ;
  assign n4556 = n4555 ^ x48 ;
  assign n4557 = ~n3760 & n4556 ;
  assign n4558 = n4557 ^ x48 ;
  assign n4559 = n4558 ^ x16 ;
  assign n4560 = n3796 & n4559 ;
  assign n4561 = n4560 ^ x16 ;
  assign n4562 = x497 ^ x465 ;
  assign n4563 = ~n3301 & n4562 ;
  assign n4564 = n4563 ^ x465 ;
  assign n4565 = n4564 ^ x433 ;
  assign n4566 = n3333 & n4565 ;
  assign n4567 = n4566 ^ x433 ;
  assign n4568 = n4567 ^ x401 ;
  assign n4569 = ~n3369 & n4568 ;
  assign n4570 = n4569 ^ x401 ;
  assign n4571 = n4570 ^ x369 ;
  assign n4572 = ~n3405 & n4571 ;
  assign n4573 = n4572 ^ x369 ;
  assign n4574 = n4573 ^ x337 ;
  assign n4575 = ~n3440 & n4574 ;
  assign n4576 = n4575 ^ x337 ;
  assign n4577 = n4576 ^ x305 ;
  assign n4578 = ~n3476 & n4577 ;
  assign n4579 = n4578 ^ x305 ;
  assign n4580 = n4579 ^ x273 ;
  assign n4581 = ~n3511 & n4580 ;
  assign n4582 = n4581 ^ x273 ;
  assign n4583 = n4582 ^ x241 ;
  assign n4584 = ~n3547 & n4583 ;
  assign n4585 = n4584 ^ x241 ;
  assign n4586 = n4585 ^ x209 ;
  assign n4587 = ~n3582 & n4586 ;
  assign n4588 = n4587 ^ x209 ;
  assign n4589 = n4588 ^ x177 ;
  assign n4590 = ~n3618 & n4589 ;
  assign n4591 = n4590 ^ x177 ;
  assign n4592 = n4591 ^ x145 ;
  assign n4593 = ~n3653 & n4592 ;
  assign n4594 = n4593 ^ x145 ;
  assign n4595 = n4594 ^ x113 ;
  assign n4596 = ~n3689 & n4595 ;
  assign n4597 = n4596 ^ x113 ;
  assign n4598 = n4597 ^ x81 ;
  assign n4599 = ~n3724 & n4598 ;
  assign n4600 = n4599 ^ x81 ;
  assign n4601 = n4600 ^ x49 ;
  assign n4602 = ~n3760 & n4601 ;
  assign n4603 = n4602 ^ x49 ;
  assign n4604 = n4603 ^ x17 ;
  assign n4605 = n3796 & n4604 ;
  assign n4606 = n4605 ^ x17 ;
  assign n4607 = x498 ^ x466 ;
  assign n4608 = ~n3301 & n4607 ;
  assign n4609 = n4608 ^ x466 ;
  assign n4610 = n4609 ^ x434 ;
  assign n4611 = n3333 & n4610 ;
  assign n4612 = n4611 ^ x434 ;
  assign n4613 = n4612 ^ x402 ;
  assign n4614 = ~n3369 & n4613 ;
  assign n4615 = n4614 ^ x402 ;
  assign n4616 = n4615 ^ x370 ;
  assign n4617 = ~n3405 & n4616 ;
  assign n4618 = n4617 ^ x370 ;
  assign n4619 = n4618 ^ x338 ;
  assign n4620 = ~n3440 & n4619 ;
  assign n4621 = n4620 ^ x338 ;
  assign n4622 = n4621 ^ x306 ;
  assign n4623 = ~n3476 & n4622 ;
  assign n4624 = n4623 ^ x306 ;
  assign n4625 = n4624 ^ x274 ;
  assign n4626 = ~n3511 & n4625 ;
  assign n4627 = n4626 ^ x274 ;
  assign n4628 = n4627 ^ x242 ;
  assign n4629 = ~n3547 & n4628 ;
  assign n4630 = n4629 ^ x242 ;
  assign n4631 = n4630 ^ x210 ;
  assign n4632 = ~n3582 & n4631 ;
  assign n4633 = n4632 ^ x210 ;
  assign n4634 = n4633 ^ x178 ;
  assign n4635 = ~n3618 & n4634 ;
  assign n4636 = n4635 ^ x178 ;
  assign n4637 = n4636 ^ x146 ;
  assign n4638 = ~n3653 & n4637 ;
  assign n4639 = n4638 ^ x146 ;
  assign n4640 = n4639 ^ x114 ;
  assign n4641 = ~n3689 & n4640 ;
  assign n4642 = n4641 ^ x114 ;
  assign n4643 = n4642 ^ x82 ;
  assign n4644 = ~n3724 & n4643 ;
  assign n4645 = n4644 ^ x82 ;
  assign n4646 = n4645 ^ x50 ;
  assign n4647 = ~n3760 & n4646 ;
  assign n4648 = n4647 ^ x50 ;
  assign n4649 = n4648 ^ x18 ;
  assign n4650 = n3796 & n4649 ;
  assign n4651 = n4650 ^ x18 ;
  assign n4652 = x499 ^ x467 ;
  assign n4653 = ~n3301 & n4652 ;
  assign n4654 = n4653 ^ x467 ;
  assign n4655 = n4654 ^ x435 ;
  assign n4656 = n3333 & n4655 ;
  assign n4657 = n4656 ^ x435 ;
  assign n4658 = n4657 ^ x403 ;
  assign n4659 = ~n3369 & n4658 ;
  assign n4660 = n4659 ^ x403 ;
  assign n4661 = n4660 ^ x371 ;
  assign n4662 = ~n3405 & n4661 ;
  assign n4663 = n4662 ^ x371 ;
  assign n4664 = n4663 ^ x339 ;
  assign n4665 = ~n3440 & n4664 ;
  assign n4666 = n4665 ^ x339 ;
  assign n4667 = n4666 ^ x307 ;
  assign n4668 = ~n3476 & n4667 ;
  assign n4669 = n4668 ^ x307 ;
  assign n4670 = n4669 ^ x275 ;
  assign n4671 = ~n3511 & n4670 ;
  assign n4672 = n4671 ^ x275 ;
  assign n4673 = n4672 ^ x243 ;
  assign n4674 = ~n3547 & n4673 ;
  assign n4675 = n4674 ^ x243 ;
  assign n4676 = n4675 ^ x211 ;
  assign n4677 = ~n3582 & n4676 ;
  assign n4678 = n4677 ^ x211 ;
  assign n4679 = n4678 ^ x179 ;
  assign n4680 = ~n3618 & n4679 ;
  assign n4681 = n4680 ^ x179 ;
  assign n4682 = n4681 ^ x147 ;
  assign n4683 = ~n3653 & n4682 ;
  assign n4684 = n4683 ^ x147 ;
  assign n4685 = n4684 ^ x115 ;
  assign n4686 = ~n3689 & n4685 ;
  assign n4687 = n4686 ^ x115 ;
  assign n4688 = n4687 ^ x83 ;
  assign n4689 = ~n3724 & n4688 ;
  assign n4690 = n4689 ^ x83 ;
  assign n4691 = n4690 ^ x51 ;
  assign n4692 = ~n3760 & n4691 ;
  assign n4693 = n4692 ^ x51 ;
  assign n4694 = n4693 ^ x19 ;
  assign n4695 = n3796 & n4694 ;
  assign n4696 = n4695 ^ x19 ;
  assign n4697 = x500 ^ x468 ;
  assign n4698 = ~n3301 & n4697 ;
  assign n4699 = n4698 ^ x468 ;
  assign n4700 = n4699 ^ x436 ;
  assign n4701 = n3333 & n4700 ;
  assign n4702 = n4701 ^ x436 ;
  assign n4703 = n4702 ^ x404 ;
  assign n4704 = ~n3369 & n4703 ;
  assign n4705 = n4704 ^ x404 ;
  assign n4706 = n4705 ^ x372 ;
  assign n4707 = ~n3405 & n4706 ;
  assign n4708 = n4707 ^ x372 ;
  assign n4709 = n4708 ^ x340 ;
  assign n4710 = ~n3440 & n4709 ;
  assign n4711 = n4710 ^ x340 ;
  assign n4712 = n4711 ^ x308 ;
  assign n4713 = ~n3476 & n4712 ;
  assign n4714 = n4713 ^ x308 ;
  assign n4715 = n4714 ^ x276 ;
  assign n4716 = ~n3511 & n4715 ;
  assign n4717 = n4716 ^ x276 ;
  assign n4718 = n4717 ^ x244 ;
  assign n4719 = ~n3547 & n4718 ;
  assign n4720 = n4719 ^ x244 ;
  assign n4721 = n4720 ^ x212 ;
  assign n4722 = ~n3582 & n4721 ;
  assign n4723 = n4722 ^ x212 ;
  assign n4724 = n4723 ^ x180 ;
  assign n4725 = ~n3618 & n4724 ;
  assign n4726 = n4725 ^ x180 ;
  assign n4727 = n4726 ^ x148 ;
  assign n4728 = ~n3653 & n4727 ;
  assign n4729 = n4728 ^ x148 ;
  assign n4730 = n4729 ^ x116 ;
  assign n4731 = ~n3689 & n4730 ;
  assign n4732 = n4731 ^ x116 ;
  assign n4733 = n4732 ^ x84 ;
  assign n4734 = ~n3724 & n4733 ;
  assign n4735 = n4734 ^ x84 ;
  assign n4736 = n4735 ^ x52 ;
  assign n4737 = ~n3760 & n4736 ;
  assign n4738 = n4737 ^ x52 ;
  assign n4739 = n4738 ^ x20 ;
  assign n4740 = n3796 & n4739 ;
  assign n4741 = n4740 ^ x20 ;
  assign n4742 = x501 ^ x469 ;
  assign n4743 = ~n3301 & n4742 ;
  assign n4744 = n4743 ^ x469 ;
  assign n4745 = n4744 ^ x437 ;
  assign n4746 = n3333 & n4745 ;
  assign n4747 = n4746 ^ x437 ;
  assign n4748 = n4747 ^ x405 ;
  assign n4749 = ~n3369 & n4748 ;
  assign n4750 = n4749 ^ x405 ;
  assign n4751 = n4750 ^ x373 ;
  assign n4752 = ~n3405 & n4751 ;
  assign n4753 = n4752 ^ x373 ;
  assign n4754 = n4753 ^ x341 ;
  assign n4755 = ~n3440 & n4754 ;
  assign n4756 = n4755 ^ x341 ;
  assign n4757 = n4756 ^ x309 ;
  assign n4758 = ~n3476 & n4757 ;
  assign n4759 = n4758 ^ x309 ;
  assign n4760 = n4759 ^ x277 ;
  assign n4761 = ~n3511 & n4760 ;
  assign n4762 = n4761 ^ x277 ;
  assign n4763 = n4762 ^ x245 ;
  assign n4764 = ~n3547 & n4763 ;
  assign n4765 = n4764 ^ x245 ;
  assign n4766 = n4765 ^ x213 ;
  assign n4767 = ~n3582 & n4766 ;
  assign n4768 = n4767 ^ x213 ;
  assign n4769 = n4768 ^ x181 ;
  assign n4770 = ~n3618 & n4769 ;
  assign n4771 = n4770 ^ x181 ;
  assign n4772 = n4771 ^ x149 ;
  assign n4773 = ~n3653 & n4772 ;
  assign n4774 = n4773 ^ x149 ;
  assign n4775 = n4774 ^ x117 ;
  assign n4776 = ~n3689 & n4775 ;
  assign n4777 = n4776 ^ x117 ;
  assign n4778 = n4777 ^ x85 ;
  assign n4779 = ~n3724 & n4778 ;
  assign n4780 = n4779 ^ x85 ;
  assign n4781 = n4780 ^ x53 ;
  assign n4782 = ~n3760 & n4781 ;
  assign n4783 = n4782 ^ x53 ;
  assign n4784 = n4783 ^ x21 ;
  assign n4785 = n3796 & n4784 ;
  assign n4786 = n4785 ^ x21 ;
  assign n4787 = x502 ^ x470 ;
  assign n4788 = ~n3301 & n4787 ;
  assign n4789 = n4788 ^ x470 ;
  assign n4790 = n4789 ^ x438 ;
  assign n4791 = n3333 & n4790 ;
  assign n4792 = n4791 ^ x438 ;
  assign n4793 = n4792 ^ x406 ;
  assign n4794 = ~n3369 & n4793 ;
  assign n4795 = n4794 ^ x406 ;
  assign n4796 = n4795 ^ x374 ;
  assign n4797 = ~n3405 & n4796 ;
  assign n4798 = n4797 ^ x374 ;
  assign n4799 = n4798 ^ x342 ;
  assign n4800 = ~n3440 & n4799 ;
  assign n4801 = n4800 ^ x342 ;
  assign n4802 = n4801 ^ x310 ;
  assign n4803 = ~n3476 & n4802 ;
  assign n4804 = n4803 ^ x310 ;
  assign n4805 = n4804 ^ x278 ;
  assign n4806 = ~n3511 & n4805 ;
  assign n4807 = n4806 ^ x278 ;
  assign n4808 = n4807 ^ x246 ;
  assign n4809 = ~n3547 & n4808 ;
  assign n4810 = n4809 ^ x246 ;
  assign n4811 = n4810 ^ x214 ;
  assign n4812 = ~n3582 & n4811 ;
  assign n4813 = n4812 ^ x214 ;
  assign n4814 = n4813 ^ x182 ;
  assign n4815 = ~n3618 & n4814 ;
  assign n4816 = n4815 ^ x182 ;
  assign n4817 = n4816 ^ x150 ;
  assign n4818 = ~n3653 & n4817 ;
  assign n4819 = n4818 ^ x150 ;
  assign n4820 = n4819 ^ x118 ;
  assign n4821 = ~n3689 & n4820 ;
  assign n4822 = n4821 ^ x118 ;
  assign n4823 = n4822 ^ x86 ;
  assign n4824 = ~n3724 & n4823 ;
  assign n4825 = n4824 ^ x86 ;
  assign n4826 = n4825 ^ x54 ;
  assign n4827 = ~n3760 & n4826 ;
  assign n4828 = n4827 ^ x54 ;
  assign n4829 = n4828 ^ x22 ;
  assign n4830 = n3796 & n4829 ;
  assign n4831 = n4830 ^ x22 ;
  assign n4832 = x503 ^ x471 ;
  assign n4833 = ~n3301 & n4832 ;
  assign n4834 = n4833 ^ x471 ;
  assign n4835 = n4834 ^ x439 ;
  assign n4836 = n3333 & n4835 ;
  assign n4837 = n4836 ^ x439 ;
  assign n4838 = n4837 ^ x407 ;
  assign n4839 = ~n3369 & n4838 ;
  assign n4840 = n4839 ^ x407 ;
  assign n4841 = n4840 ^ x375 ;
  assign n4842 = ~n3405 & n4841 ;
  assign n4843 = n4842 ^ x375 ;
  assign n4844 = n4843 ^ x343 ;
  assign n4845 = ~n3440 & n4844 ;
  assign n4846 = n4845 ^ x343 ;
  assign n4847 = n4846 ^ x311 ;
  assign n4848 = ~n3476 & n4847 ;
  assign n4849 = n4848 ^ x311 ;
  assign n4850 = n4849 ^ x279 ;
  assign n4851 = ~n3511 & n4850 ;
  assign n4852 = n4851 ^ x279 ;
  assign n4853 = n4852 ^ x247 ;
  assign n4854 = ~n3547 & n4853 ;
  assign n4855 = n4854 ^ x247 ;
  assign n4856 = n4855 ^ x215 ;
  assign n4857 = ~n3582 & n4856 ;
  assign n4858 = n4857 ^ x215 ;
  assign n4859 = n4858 ^ x183 ;
  assign n4860 = ~n3618 & n4859 ;
  assign n4861 = n4860 ^ x183 ;
  assign n4862 = n4861 ^ x151 ;
  assign n4863 = ~n3653 & n4862 ;
  assign n4864 = n4863 ^ x151 ;
  assign n4865 = n4864 ^ x119 ;
  assign n4866 = ~n3689 & n4865 ;
  assign n4867 = n4866 ^ x119 ;
  assign n4868 = n4867 ^ x87 ;
  assign n4869 = ~n3724 & n4868 ;
  assign n4870 = n4869 ^ x87 ;
  assign n4871 = n4870 ^ x55 ;
  assign n4872 = ~n3760 & n4871 ;
  assign n4873 = n4872 ^ x55 ;
  assign n4874 = n4873 ^ x23 ;
  assign n4875 = n3796 & n4874 ;
  assign n4876 = n4875 ^ x23 ;
  assign n4877 = x504 ^ x472 ;
  assign n4878 = ~n3301 & n4877 ;
  assign n4879 = n4878 ^ x472 ;
  assign n4880 = n4879 ^ x440 ;
  assign n4881 = n3333 & n4880 ;
  assign n4882 = n4881 ^ x440 ;
  assign n4883 = n4882 ^ x408 ;
  assign n4884 = ~n3369 & n4883 ;
  assign n4885 = n4884 ^ x408 ;
  assign n4886 = n4885 ^ x376 ;
  assign n4887 = ~n3405 & n4886 ;
  assign n4888 = n4887 ^ x376 ;
  assign n4889 = n4888 ^ x344 ;
  assign n4890 = ~n3440 & n4889 ;
  assign n4891 = n4890 ^ x344 ;
  assign n4892 = n4891 ^ x312 ;
  assign n4893 = ~n3476 & n4892 ;
  assign n4894 = n4893 ^ x312 ;
  assign n4895 = n4894 ^ x280 ;
  assign n4896 = ~n3511 & n4895 ;
  assign n4897 = n4896 ^ x280 ;
  assign n4898 = n4897 ^ x248 ;
  assign n4899 = ~n3547 & n4898 ;
  assign n4900 = n4899 ^ x248 ;
  assign n4901 = n4900 ^ x216 ;
  assign n4902 = ~n3582 & n4901 ;
  assign n4903 = n4902 ^ x216 ;
  assign n4904 = n4903 ^ x184 ;
  assign n4905 = ~n3618 & n4904 ;
  assign n4906 = n4905 ^ x184 ;
  assign n4907 = n4906 ^ x152 ;
  assign n4908 = ~n3653 & n4907 ;
  assign n4909 = n4908 ^ x152 ;
  assign n4910 = n4909 ^ x120 ;
  assign n4911 = ~n3689 & n4910 ;
  assign n4912 = n4911 ^ x120 ;
  assign n4913 = n4912 ^ x88 ;
  assign n4914 = ~n3724 & n4913 ;
  assign n4915 = n4914 ^ x88 ;
  assign n4916 = n4915 ^ x56 ;
  assign n4917 = ~n3760 & n4916 ;
  assign n4918 = n4917 ^ x56 ;
  assign n4919 = n4918 ^ x24 ;
  assign n4920 = n3796 & n4919 ;
  assign n4921 = n4920 ^ x24 ;
  assign n4922 = x505 ^ x473 ;
  assign n4923 = ~n3301 & n4922 ;
  assign n4924 = n4923 ^ x473 ;
  assign n4925 = n4924 ^ x441 ;
  assign n4926 = n3333 & n4925 ;
  assign n4927 = n4926 ^ x441 ;
  assign n4928 = n4927 ^ x409 ;
  assign n4929 = ~n3369 & n4928 ;
  assign n4930 = n4929 ^ x409 ;
  assign n4931 = n4930 ^ x377 ;
  assign n4932 = ~n3405 & n4931 ;
  assign n4933 = n4932 ^ x377 ;
  assign n4934 = n4933 ^ x345 ;
  assign n4935 = ~n3440 & n4934 ;
  assign n4936 = n4935 ^ x345 ;
  assign n4937 = n4936 ^ x313 ;
  assign n4938 = ~n3476 & n4937 ;
  assign n4939 = n4938 ^ x313 ;
  assign n4940 = n4939 ^ x281 ;
  assign n4941 = ~n3511 & n4940 ;
  assign n4942 = n4941 ^ x281 ;
  assign n4943 = n4942 ^ x249 ;
  assign n4944 = ~n3547 & n4943 ;
  assign n4945 = n4944 ^ x249 ;
  assign n4946 = n4945 ^ x217 ;
  assign n4947 = ~n3582 & n4946 ;
  assign n4948 = n4947 ^ x217 ;
  assign n4949 = n4948 ^ x185 ;
  assign n4950 = ~n3618 & n4949 ;
  assign n4951 = n4950 ^ x185 ;
  assign n4952 = n4951 ^ x153 ;
  assign n4953 = ~n3653 & n4952 ;
  assign n4954 = n4953 ^ x153 ;
  assign n4955 = n4954 ^ x121 ;
  assign n4956 = ~n3689 & n4955 ;
  assign n4957 = n4956 ^ x121 ;
  assign n4958 = n4957 ^ x89 ;
  assign n4959 = ~n3724 & n4958 ;
  assign n4960 = n4959 ^ x89 ;
  assign n4961 = n4960 ^ x57 ;
  assign n4962 = ~n3760 & n4961 ;
  assign n4963 = n4962 ^ x57 ;
  assign n4964 = n4963 ^ x25 ;
  assign n4965 = n3796 & n4964 ;
  assign n4966 = n4965 ^ x25 ;
  assign n4967 = x506 ^ x474 ;
  assign n4968 = ~n3301 & n4967 ;
  assign n4969 = n4968 ^ x474 ;
  assign n4970 = n4969 ^ x442 ;
  assign n4971 = n3333 & n4970 ;
  assign n4972 = n4971 ^ x442 ;
  assign n4973 = n4972 ^ x410 ;
  assign n4974 = ~n3369 & n4973 ;
  assign n4975 = n4974 ^ x410 ;
  assign n4976 = n4975 ^ x378 ;
  assign n4977 = ~n3405 & n4976 ;
  assign n4978 = n4977 ^ x378 ;
  assign n4979 = n4978 ^ x346 ;
  assign n4980 = ~n3440 & n4979 ;
  assign n4981 = n4980 ^ x346 ;
  assign n4982 = n4981 ^ x314 ;
  assign n4983 = ~n3476 & n4982 ;
  assign n4984 = n4983 ^ x314 ;
  assign n4985 = n4984 ^ x282 ;
  assign n4986 = ~n3511 & n4985 ;
  assign n4987 = n4986 ^ x282 ;
  assign n4988 = n4987 ^ x250 ;
  assign n4989 = ~n3547 & n4988 ;
  assign n4990 = n4989 ^ x250 ;
  assign n4991 = n4990 ^ x218 ;
  assign n4992 = ~n3582 & n4991 ;
  assign n4993 = n4992 ^ x218 ;
  assign n4994 = n4993 ^ x186 ;
  assign n4995 = ~n3618 & n4994 ;
  assign n4996 = n4995 ^ x186 ;
  assign n4997 = n4996 ^ x154 ;
  assign n4998 = ~n3653 & n4997 ;
  assign n4999 = n4998 ^ x154 ;
  assign n5000 = n4999 ^ x122 ;
  assign n5001 = ~n3689 & n5000 ;
  assign n5002 = n5001 ^ x122 ;
  assign n5003 = n5002 ^ x90 ;
  assign n5004 = ~n3724 & n5003 ;
  assign n5005 = n5004 ^ x90 ;
  assign n5006 = n5005 ^ x58 ;
  assign n5007 = ~n3760 & n5006 ;
  assign n5008 = n5007 ^ x58 ;
  assign n5009 = n5008 ^ x26 ;
  assign n5010 = n3796 & n5009 ;
  assign n5011 = n5010 ^ x26 ;
  assign n5012 = x507 ^ x475 ;
  assign n5013 = ~n3301 & n5012 ;
  assign n5014 = n5013 ^ x475 ;
  assign n5015 = n5014 ^ x443 ;
  assign n5016 = n3333 & n5015 ;
  assign n5017 = n5016 ^ x443 ;
  assign n5018 = n5017 ^ x411 ;
  assign n5019 = ~n3369 & n5018 ;
  assign n5020 = n5019 ^ x411 ;
  assign n5021 = n5020 ^ x379 ;
  assign n5022 = ~n3405 & n5021 ;
  assign n5023 = n5022 ^ x379 ;
  assign n5024 = n5023 ^ x347 ;
  assign n5025 = ~n3440 & n5024 ;
  assign n5026 = n5025 ^ x347 ;
  assign n5027 = n5026 ^ x315 ;
  assign n5028 = ~n3476 & n5027 ;
  assign n5029 = n5028 ^ x315 ;
  assign n5030 = n5029 ^ x283 ;
  assign n5031 = ~n3511 & n5030 ;
  assign n5032 = n5031 ^ x283 ;
  assign n5033 = n5032 ^ x251 ;
  assign n5034 = ~n3547 & n5033 ;
  assign n5035 = n5034 ^ x251 ;
  assign n5036 = n5035 ^ x219 ;
  assign n5037 = ~n3582 & n5036 ;
  assign n5038 = n5037 ^ x219 ;
  assign n5039 = n5038 ^ x187 ;
  assign n5040 = ~n3618 & n5039 ;
  assign n5041 = n5040 ^ x187 ;
  assign n5042 = n5041 ^ x155 ;
  assign n5043 = ~n3653 & n5042 ;
  assign n5044 = n5043 ^ x155 ;
  assign n5045 = n5044 ^ x123 ;
  assign n5046 = ~n3689 & n5045 ;
  assign n5047 = n5046 ^ x123 ;
  assign n5048 = n5047 ^ x91 ;
  assign n5049 = ~n3724 & n5048 ;
  assign n5050 = n5049 ^ x91 ;
  assign n5051 = n5050 ^ x59 ;
  assign n5052 = ~n3760 & n5051 ;
  assign n5053 = n5052 ^ x59 ;
  assign n5054 = n5053 ^ x27 ;
  assign n5055 = n3796 & n5054 ;
  assign n5056 = n5055 ^ x27 ;
  assign n5057 = x508 ^ x476 ;
  assign n5058 = ~n3301 & n5057 ;
  assign n5059 = n5058 ^ x476 ;
  assign n5060 = n5059 ^ x444 ;
  assign n5061 = n3333 & n5060 ;
  assign n5062 = n5061 ^ x444 ;
  assign n5063 = n5062 ^ x412 ;
  assign n5064 = ~n3369 & n5063 ;
  assign n5065 = n5064 ^ x412 ;
  assign n5066 = n5065 ^ x380 ;
  assign n5067 = ~n3405 & n5066 ;
  assign n5068 = n5067 ^ x380 ;
  assign n5069 = n5068 ^ x348 ;
  assign n5070 = ~n3440 & n5069 ;
  assign n5071 = n5070 ^ x348 ;
  assign n5072 = n5071 ^ x316 ;
  assign n5073 = ~n3476 & n5072 ;
  assign n5074 = n5073 ^ x316 ;
  assign n5075 = n5074 ^ x284 ;
  assign n5076 = ~n3511 & n5075 ;
  assign n5077 = n5076 ^ x284 ;
  assign n5078 = n5077 ^ x252 ;
  assign n5079 = ~n3547 & n5078 ;
  assign n5080 = n5079 ^ x252 ;
  assign n5081 = n5080 ^ x220 ;
  assign n5082 = ~n3582 & n5081 ;
  assign n5083 = n5082 ^ x220 ;
  assign n5084 = n5083 ^ x188 ;
  assign n5085 = ~n3618 & n5084 ;
  assign n5086 = n5085 ^ x188 ;
  assign n5087 = n5086 ^ x156 ;
  assign n5088 = ~n3653 & n5087 ;
  assign n5089 = n5088 ^ x156 ;
  assign n5090 = n5089 ^ x124 ;
  assign n5091 = ~n3689 & n5090 ;
  assign n5092 = n5091 ^ x124 ;
  assign n5093 = n5092 ^ x92 ;
  assign n5094 = ~n3724 & n5093 ;
  assign n5095 = n5094 ^ x92 ;
  assign n5096 = n5095 ^ x60 ;
  assign n5097 = ~n3760 & n5096 ;
  assign n5098 = n5097 ^ x60 ;
  assign n5099 = n5098 ^ x28 ;
  assign n5100 = n3796 & n5099 ;
  assign n5101 = n5100 ^ x28 ;
  assign n5102 = x509 ^ x477 ;
  assign n5103 = ~n3301 & n5102 ;
  assign n5104 = n5103 ^ x477 ;
  assign n5105 = n5104 ^ x445 ;
  assign n5106 = n3333 & n5105 ;
  assign n5107 = n5106 ^ x445 ;
  assign n5108 = n5107 ^ x413 ;
  assign n5109 = ~n3369 & n5108 ;
  assign n5110 = n5109 ^ x413 ;
  assign n5111 = n5110 ^ x381 ;
  assign n5112 = ~n3405 & n5111 ;
  assign n5113 = n5112 ^ x381 ;
  assign n5114 = n5113 ^ x349 ;
  assign n5115 = ~n3440 & n5114 ;
  assign n5116 = n5115 ^ x349 ;
  assign n5117 = n5116 ^ x317 ;
  assign n5118 = ~n3476 & n5117 ;
  assign n5119 = n5118 ^ x317 ;
  assign n5120 = n5119 ^ x285 ;
  assign n5121 = ~n3511 & n5120 ;
  assign n5122 = n5121 ^ x285 ;
  assign n5123 = n5122 ^ x253 ;
  assign n5124 = ~n3547 & n5123 ;
  assign n5125 = n5124 ^ x253 ;
  assign n5126 = n5125 ^ x221 ;
  assign n5127 = ~n3582 & n5126 ;
  assign n5128 = n5127 ^ x221 ;
  assign n5129 = n5128 ^ x189 ;
  assign n5130 = ~n3618 & n5129 ;
  assign n5131 = n5130 ^ x189 ;
  assign n5132 = n5131 ^ x157 ;
  assign n5133 = ~n3653 & n5132 ;
  assign n5134 = n5133 ^ x157 ;
  assign n5135 = n5134 ^ x125 ;
  assign n5136 = ~n3689 & n5135 ;
  assign n5137 = n5136 ^ x125 ;
  assign n5138 = n5137 ^ x93 ;
  assign n5139 = ~n3724 & n5138 ;
  assign n5140 = n5139 ^ x93 ;
  assign n5141 = n5140 ^ x61 ;
  assign n5142 = ~n3760 & n5141 ;
  assign n5143 = n5142 ^ x61 ;
  assign n5144 = n5143 ^ x29 ;
  assign n5145 = n3796 & n5144 ;
  assign n5146 = n5145 ^ x29 ;
  assign n5147 = x510 ^ x478 ;
  assign n5148 = ~n3301 & n5147 ;
  assign n5149 = n5148 ^ x478 ;
  assign n5150 = n5149 ^ x446 ;
  assign n5151 = n3333 & n5150 ;
  assign n5152 = n5151 ^ x446 ;
  assign n5153 = n5152 ^ x414 ;
  assign n5154 = ~n3369 & n5153 ;
  assign n5155 = n5154 ^ x414 ;
  assign n5156 = n5155 ^ x382 ;
  assign n5157 = ~n3405 & n5156 ;
  assign n5158 = n5157 ^ x382 ;
  assign n5159 = n5158 ^ x350 ;
  assign n5160 = ~n3440 & n5159 ;
  assign n5161 = n5160 ^ x350 ;
  assign n5162 = n5161 ^ x318 ;
  assign n5163 = ~n3476 & n5162 ;
  assign n5164 = n5163 ^ x318 ;
  assign n5165 = n5164 ^ x286 ;
  assign n5166 = ~n3511 & n5165 ;
  assign n5167 = n5166 ^ x286 ;
  assign n5168 = n5167 ^ x254 ;
  assign n5169 = ~n3547 & n5168 ;
  assign n5170 = n5169 ^ x254 ;
  assign n5171 = n5170 ^ x222 ;
  assign n5172 = ~n3582 & n5171 ;
  assign n5173 = n5172 ^ x222 ;
  assign n5174 = n5173 ^ x190 ;
  assign n5175 = ~n3618 & n5174 ;
  assign n5176 = n5175 ^ x190 ;
  assign n5177 = n5176 ^ x158 ;
  assign n5178 = ~n3653 & n5177 ;
  assign n5179 = n5178 ^ x158 ;
  assign n5180 = n5179 ^ x126 ;
  assign n5181 = ~n3689 & n5180 ;
  assign n5182 = n5181 ^ x126 ;
  assign n5183 = n5182 ^ x94 ;
  assign n5184 = ~n3724 & n5183 ;
  assign n5185 = n5184 ^ x94 ;
  assign n5186 = n5185 ^ x62 ;
  assign n5187 = ~n3760 & n5186 ;
  assign n5188 = n5187 ^ x62 ;
  assign n5189 = n5188 ^ x30 ;
  assign n5190 = n3796 & n5189 ;
  assign n5191 = n5190 ^ x30 ;
  assign n5192 = x511 ^ x479 ;
  assign n5193 = ~n3301 & n5192 ;
  assign n5194 = n5193 ^ x479 ;
  assign n5195 = n5194 ^ x447 ;
  assign n5196 = n3333 & n5195 ;
  assign n5197 = n5196 ^ x447 ;
  assign n5198 = n5197 ^ x415 ;
  assign n5199 = ~n3369 & n5198 ;
  assign n5200 = n5199 ^ x415 ;
  assign n5201 = n5200 ^ x383 ;
  assign n5202 = ~n3405 & n5201 ;
  assign n5203 = n5202 ^ x383 ;
  assign n5204 = n5203 ^ x351 ;
  assign n5205 = ~n3440 & n5204 ;
  assign n5206 = n5205 ^ x351 ;
  assign n5207 = n5206 ^ x319 ;
  assign n5208 = ~n3476 & n5207 ;
  assign n5209 = n5208 ^ x319 ;
  assign n5210 = n5209 ^ x287 ;
  assign n5211 = ~n3511 & n5210 ;
  assign n5212 = n5211 ^ x287 ;
  assign n5213 = n5212 ^ x255 ;
  assign n5214 = ~n3547 & n5213 ;
  assign n5215 = n5214 ^ x255 ;
  assign n5216 = n5215 ^ x223 ;
  assign n5217 = ~n3582 & n5216 ;
  assign n5218 = n5217 ^ x223 ;
  assign n5219 = n5218 ^ x191 ;
  assign n5220 = ~n3618 & n5219 ;
  assign n5221 = n5220 ^ x191 ;
  assign n5222 = n5221 ^ x159 ;
  assign n5223 = ~n3653 & n5222 ;
  assign n5224 = n5223 ^ x159 ;
  assign n5225 = n5224 ^ x127 ;
  assign n5226 = ~n3689 & n5225 ;
  assign n5227 = n5226 ^ x127 ;
  assign n5228 = n5227 ^ x95 ;
  assign n5229 = ~n3724 & n5228 ;
  assign n5230 = n5229 ^ x95 ;
  assign n5231 = n5230 ^ x63 ;
  assign n5232 = ~n3760 & n5231 ;
  assign n5233 = n5232 ^ x63 ;
  assign n5234 = n5233 ^ x31 ;
  assign n5235 = n3796 & n5234 ;
  assign n5236 = n5235 ^ x31 ;
  assign y0 = n3841 ;
  assign y1 = n3886 ;
  assign y2 = n3931 ;
  assign y3 = n3976 ;
  assign y4 = n4021 ;
  assign y5 = n4066 ;
  assign y6 = n4111 ;
  assign y7 = n4156 ;
  assign y8 = n4201 ;
  assign y9 = n4246 ;
  assign y10 = n4291 ;
  assign y11 = n4336 ;
  assign y12 = n4381 ;
  assign y13 = n4426 ;
  assign y14 = n4471 ;
  assign y15 = n4516 ;
  assign y16 = n4561 ;
  assign y17 = n4606 ;
  assign y18 = n4651 ;
  assign y19 = n4696 ;
  assign y20 = n4741 ;
  assign y21 = n4786 ;
  assign y22 = n4831 ;
  assign y23 = n4876 ;
  assign y24 = n4921 ;
  assign y25 = n4966 ;
  assign y26 = n5011 ;
  assign y27 = n5056 ;
  assign y28 = n5101 ;
  assign y29 = n5146 ;
  assign y30 = n5191 ;
  assign y31 = n5236 ;
endmodule
