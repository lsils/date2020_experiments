// Benchmark "knn_comb_BMR_2_8" written by ABC on Tue Nov 26 14:01:11 2019

module knn_comb_BMR_2_8 ( 
    \p_input[0] , \p_input[1] , \p_input[2] , \p_input[3] , \p_input[4] ,
    \p_input[5] , \p_input[6] , \p_input[7] , \p_input[8] , \p_input[9] ,
    \p_input[10] , \p_input[11] , \p_input[12] , \p_input[13] ,
    \p_input[14] , \p_input[15] , \p_input[16] , \p_input[17] ,
    \p_input[18] , \p_input[19] , \p_input[20] , \p_input[21] ,
    \p_input[22] , \p_input[23] , \p_input[24] , \p_input[25] ,
    \p_input[26] , \p_input[27] , \p_input[28] , \p_input[29] ,
    \p_input[30] , \p_input[31] , \p_input[32] , \p_input[33] ,
    \p_input[34] , \p_input[35] , \p_input[36] , \p_input[37] ,
    \p_input[38] , \p_input[39] , \p_input[40] , \p_input[41] ,
    \p_input[42] , \p_input[43] , \p_input[44] , \p_input[45] ,
    \p_input[46] , \p_input[47] , \p_input[48] , \p_input[49] ,
    \p_input[50] , \p_input[51] , \p_input[52] , \p_input[53] ,
    \p_input[54] , \p_input[55] , \p_input[56] , \p_input[57] ,
    \p_input[58] , \p_input[59] , \p_input[60] , \p_input[61] ,
    \p_input[62] , \p_input[63] , \p_input[64] , \p_input[65] ,
    \p_input[66] , \p_input[67] , \p_input[68] , \p_input[69] ,
    \p_input[70] , \p_input[71] , \p_input[72] , \p_input[73] ,
    \p_input[74] , \p_input[75] , \p_input[76] , \p_input[77] ,
    \p_input[78] , \p_input[79] , \p_input[80] , \p_input[81] ,
    \p_input[82] , \p_input[83] , \p_input[84] , \p_input[85] ,
    \p_input[86] , \p_input[87] , \p_input[88] , \p_input[89] ,
    \p_input[90] , \p_input[91] , \p_input[92] , \p_input[93] ,
    \p_input[94] , \p_input[95] , \p_input[96] , \p_input[97] ,
    \p_input[98] , \p_input[99] , \p_input[100] , \p_input[101] ,
    \p_input[102] , \p_input[103] , \p_input[104] , \p_input[105] ,
    \p_input[106] , \p_input[107] , \p_input[108] , \p_input[109] ,
    \p_input[110] , \p_input[111] , \p_input[112] , \p_input[113] ,
    \p_input[114] , \p_input[115] , \p_input[116] , \p_input[117] ,
    \p_input[118] , \p_input[119] , \p_input[120] , \p_input[121] ,
    \p_input[122] , \p_input[123] , \p_input[124] , \p_input[125] ,
    \p_input[126] , \p_input[127] , \p_input[128] , \p_input[129] ,
    \p_input[130] , \p_input[131] , \p_input[132] , \p_input[133] ,
    \p_input[134] , \p_input[135] , \p_input[136] , \p_input[137] ,
    \p_input[138] , \p_input[139] , \p_input[140] , \p_input[141] ,
    \p_input[142] , \p_input[143] , \p_input[144] , \p_input[145] ,
    \p_input[146] , \p_input[147] , \p_input[148] , \p_input[149] ,
    \p_input[150] , \p_input[151] , \p_input[152] , \p_input[153] ,
    \p_input[154] , \p_input[155] , \p_input[156] , \p_input[157] ,
    \p_input[158] , \p_input[159] , \p_input[160] , \p_input[161] ,
    \p_input[162] , \p_input[163] , \p_input[164] , \p_input[165] ,
    \p_input[166] , \p_input[167] , \p_input[168] , \p_input[169] ,
    \p_input[170] , \p_input[171] , \p_input[172] , \p_input[173] ,
    \p_input[174] , \p_input[175] , \p_input[176] , \p_input[177] ,
    \p_input[178] , \p_input[179] , \p_input[180] , \p_input[181] ,
    \p_input[182] , \p_input[183] , \p_input[184] , \p_input[185] ,
    \p_input[186] , \p_input[187] , \p_input[188] , \p_input[189] ,
    \p_input[190] , \p_input[191] , \p_input[192] , \p_input[193] ,
    \p_input[194] , \p_input[195] , \p_input[196] , \p_input[197] ,
    \p_input[198] , \p_input[199] , \p_input[200] , \p_input[201] ,
    \p_input[202] , \p_input[203] , \p_input[204] , \p_input[205] ,
    \p_input[206] , \p_input[207] , \p_input[208] , \p_input[209] ,
    \p_input[210] , \p_input[211] , \p_input[212] , \p_input[213] ,
    \p_input[214] , \p_input[215] , \p_input[216] , \p_input[217] ,
    \p_input[218] , \p_input[219] , \p_input[220] , \p_input[221] ,
    \p_input[222] , \p_input[223] , \p_input[224] , \p_input[225] ,
    \p_input[226] , \p_input[227] , \p_input[228] , \p_input[229] ,
    \p_input[230] , \p_input[231] , \p_input[232] , \p_input[233] ,
    \p_input[234] , \p_input[235] , \p_input[236] , \p_input[237] ,
    \p_input[238] , \p_input[239] , \p_input[240] , \p_input[241] ,
    \p_input[242] , \p_input[243] , \p_input[244] , \p_input[245] ,
    \p_input[246] , \p_input[247] , \p_input[248] , \p_input[249] ,
    \p_input[250] , \p_input[251] , \p_input[252] , \p_input[253] ,
    \p_input[254] , \p_input[255] , \p_input[256] , \p_input[257] ,
    \p_input[258] , \p_input[259] , \p_input[260] , \p_input[261] ,
    \p_input[262] , \p_input[263] , \p_input[264] , \p_input[265] ,
    \p_input[266] , \p_input[267] , \p_input[268] , \p_input[269] ,
    \p_input[270] , \p_input[271] , \p_input[272] , \p_input[273] ,
    \p_input[274] , \p_input[275] , \p_input[276] , \p_input[277] ,
    \p_input[278] , \p_input[279] , \p_input[280] , \p_input[281] ,
    \p_input[282] , \p_input[283] , \p_input[284] , \p_input[285] ,
    \p_input[286] , \p_input[287] ,
    \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] , \o[8] ,
    \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] , \o[16] ,
    \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] , \o[24] ,
    \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] , \o[32] ,
    \o[33] , \o[34] , \o[35] , \o[36] , \o[37] , \o[38] , \o[39] , \o[40] ,
    \o[41] , \o[42] , \o[43] , \o[44] , \o[45] , \o[46] , \o[47] , \o[48] ,
    \o[49] , \o[50] , \o[51] , \o[52] , \o[53] , \o[54] , \o[55] , \o[56] ,
    \o[57] , \o[58] , \o[59] , \o[60] , \o[61] , \o[62] , \o[63]   );
  input  \p_input[0] , \p_input[1] , \p_input[2] , \p_input[3] ,
    \p_input[4] , \p_input[5] , \p_input[6] , \p_input[7] , \p_input[8] ,
    \p_input[9] , \p_input[10] , \p_input[11] , \p_input[12] ,
    \p_input[13] , \p_input[14] , \p_input[15] , \p_input[16] ,
    \p_input[17] , \p_input[18] , \p_input[19] , \p_input[20] ,
    \p_input[21] , \p_input[22] , \p_input[23] , \p_input[24] ,
    \p_input[25] , \p_input[26] , \p_input[27] , \p_input[28] ,
    \p_input[29] , \p_input[30] , \p_input[31] , \p_input[32] ,
    \p_input[33] , \p_input[34] , \p_input[35] , \p_input[36] ,
    \p_input[37] , \p_input[38] , \p_input[39] , \p_input[40] ,
    \p_input[41] , \p_input[42] , \p_input[43] , \p_input[44] ,
    \p_input[45] , \p_input[46] , \p_input[47] , \p_input[48] ,
    \p_input[49] , \p_input[50] , \p_input[51] , \p_input[52] ,
    \p_input[53] , \p_input[54] , \p_input[55] , \p_input[56] ,
    \p_input[57] , \p_input[58] , \p_input[59] , \p_input[60] ,
    \p_input[61] , \p_input[62] , \p_input[63] , \p_input[64] ,
    \p_input[65] , \p_input[66] , \p_input[67] , \p_input[68] ,
    \p_input[69] , \p_input[70] , \p_input[71] , \p_input[72] ,
    \p_input[73] , \p_input[74] , \p_input[75] , \p_input[76] ,
    \p_input[77] , \p_input[78] , \p_input[79] , \p_input[80] ,
    \p_input[81] , \p_input[82] , \p_input[83] , \p_input[84] ,
    \p_input[85] , \p_input[86] , \p_input[87] , \p_input[88] ,
    \p_input[89] , \p_input[90] , \p_input[91] , \p_input[92] ,
    \p_input[93] , \p_input[94] , \p_input[95] , \p_input[96] ,
    \p_input[97] , \p_input[98] , \p_input[99] , \p_input[100] ,
    \p_input[101] , \p_input[102] , \p_input[103] , \p_input[104] ,
    \p_input[105] , \p_input[106] , \p_input[107] , \p_input[108] ,
    \p_input[109] , \p_input[110] , \p_input[111] , \p_input[112] ,
    \p_input[113] , \p_input[114] , \p_input[115] , \p_input[116] ,
    \p_input[117] , \p_input[118] , \p_input[119] , \p_input[120] ,
    \p_input[121] , \p_input[122] , \p_input[123] , \p_input[124] ,
    \p_input[125] , \p_input[126] , \p_input[127] , \p_input[128] ,
    \p_input[129] , \p_input[130] , \p_input[131] , \p_input[132] ,
    \p_input[133] , \p_input[134] , \p_input[135] , \p_input[136] ,
    \p_input[137] , \p_input[138] , \p_input[139] , \p_input[140] ,
    \p_input[141] , \p_input[142] , \p_input[143] , \p_input[144] ,
    \p_input[145] , \p_input[146] , \p_input[147] , \p_input[148] ,
    \p_input[149] , \p_input[150] , \p_input[151] , \p_input[152] ,
    \p_input[153] , \p_input[154] , \p_input[155] , \p_input[156] ,
    \p_input[157] , \p_input[158] , \p_input[159] , \p_input[160] ,
    \p_input[161] , \p_input[162] , \p_input[163] , \p_input[164] ,
    \p_input[165] , \p_input[166] , \p_input[167] , \p_input[168] ,
    \p_input[169] , \p_input[170] , \p_input[171] , \p_input[172] ,
    \p_input[173] , \p_input[174] , \p_input[175] , \p_input[176] ,
    \p_input[177] , \p_input[178] , \p_input[179] , \p_input[180] ,
    \p_input[181] , \p_input[182] , \p_input[183] , \p_input[184] ,
    \p_input[185] , \p_input[186] , \p_input[187] , \p_input[188] ,
    \p_input[189] , \p_input[190] , \p_input[191] , \p_input[192] ,
    \p_input[193] , \p_input[194] , \p_input[195] , \p_input[196] ,
    \p_input[197] , \p_input[198] , \p_input[199] , \p_input[200] ,
    \p_input[201] , \p_input[202] , \p_input[203] , \p_input[204] ,
    \p_input[205] , \p_input[206] , \p_input[207] , \p_input[208] ,
    \p_input[209] , \p_input[210] , \p_input[211] , \p_input[212] ,
    \p_input[213] , \p_input[214] , \p_input[215] , \p_input[216] ,
    \p_input[217] , \p_input[218] , \p_input[219] , \p_input[220] ,
    \p_input[221] , \p_input[222] , \p_input[223] , \p_input[224] ,
    \p_input[225] , \p_input[226] , \p_input[227] , \p_input[228] ,
    \p_input[229] , \p_input[230] , \p_input[231] , \p_input[232] ,
    \p_input[233] , \p_input[234] , \p_input[235] , \p_input[236] ,
    \p_input[237] , \p_input[238] , \p_input[239] , \p_input[240] ,
    \p_input[241] , \p_input[242] , \p_input[243] , \p_input[244] ,
    \p_input[245] , \p_input[246] , \p_input[247] , \p_input[248] ,
    \p_input[249] , \p_input[250] , \p_input[251] , \p_input[252] ,
    \p_input[253] , \p_input[254] , \p_input[255] , \p_input[256] ,
    \p_input[257] , \p_input[258] , \p_input[259] , \p_input[260] ,
    \p_input[261] , \p_input[262] , \p_input[263] , \p_input[264] ,
    \p_input[265] , \p_input[266] , \p_input[267] , \p_input[268] ,
    \p_input[269] , \p_input[270] , \p_input[271] , \p_input[272] ,
    \p_input[273] , \p_input[274] , \p_input[275] , \p_input[276] ,
    \p_input[277] , \p_input[278] , \p_input[279] , \p_input[280] ,
    \p_input[281] , \p_input[282] , \p_input[283] , \p_input[284] ,
    \p_input[285] , \p_input[286] , \p_input[287] ;
  output \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] ,
    \o[8] , \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] ,
    \o[16] , \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] ,
    \o[24] , \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] ,
    \o[32] , \o[33] , \o[34] , \o[35] , \o[36] , \o[37] , \o[38] , \o[39] ,
    \o[40] , \o[41] , \o[42] , \o[43] , \o[44] , \o[45] , \o[46] , \o[47] ,
    \o[48] , \o[49] , \o[50] , \o[51] , \o[52] , \o[53] , \o[54] , \o[55] ,
    \o[56] , \o[57] , \o[58] , \o[59] , \o[60] , \o[61] , \o[62] , \o[63] ;
  wire new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_,
    new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_,
    new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_,
    new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_,
    new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_,
    new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_,
    new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_,
    new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_,
    new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_,
    new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_,
    new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_,
    new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_,
    new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_,
    new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_,
    new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_,
    new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_,
    new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_,
    new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_,
    new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_,
    new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_,
    new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_,
    new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_,
    new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_,
    new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_,
    new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_,
    new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_,
    new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_,
    new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_,
    new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_,
    new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_,
    new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_,
    new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_,
    new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_,
    new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_,
    new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_,
    new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_,
    new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_,
    new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_,
    new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_,
    new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_,
    new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_,
    new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_,
    new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_,
    new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_,
    new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_,
    new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_,
    new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_,
    new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_,
    new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_,
    new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_,
    new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_,
    new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_,
    new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_,
    new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_,
    new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_,
    new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_,
    new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_,
    new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_,
    new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_,
    new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_,
    new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_,
    new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_,
    new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_,
    new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_,
    new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_,
    new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_,
    new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_,
    new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_,
    new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_,
    new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_,
    new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_,
    new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_,
    new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_,
    new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_,
    new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_,
    new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_,
    new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_,
    new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_,
    new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_,
    new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_,
    new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_,
    new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_,
    new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_,
    new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_,
    new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_,
    new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_,
    new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_,
    new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_,
    new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_,
    new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_,
    new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_,
    new_n3451_, new_n3452_, new_n3453_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_,
    new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_,
    new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_,
    new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_,
    new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_,
    new_n3567_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3626_, new_n3627_, new_n3628_,
    new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_,
    new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_,
    new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_,
    new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_,
    new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_,
    new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_,
    new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_,
    new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_,
    new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_,
    new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_,
    new_n3793_, new_n3794_, new_n3795_, new_n3797_, new_n3798_, new_n3799_,
    new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_, new_n3805_,
    new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_, new_n3811_,
    new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_, new_n3817_,
    new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_, new_n3823_,
    new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_, new_n3829_,
    new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_, new_n3835_,
    new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_, new_n3841_,
    new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_, new_n3847_,
    new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_, new_n3854_,
    new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_,
    new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_,
    new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_,
    new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_,
    new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_,
    new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_,
    new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_,
    new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_,
    new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_,
    new_n3909_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3968_, new_n3969_, new_n3970_,
    new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_,
    new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_,
    new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_,
    new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_,
    new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_,
    new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_,
    new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_,
    new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_,
    new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_,
    new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_,
    new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_,
    new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_,
    new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_,
    new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4139_, new_n4140_, new_n4141_,
    new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_,
    new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_,
    new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4159_,
    new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_, new_n4165_,
    new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_, new_n4171_,
    new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_, new_n4177_,
    new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_, new_n4183_,
    new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4196_,
    new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_,
    new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_,
    new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_,
    new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_,
    new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_,
    new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_,
    new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_,
    new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_,
    new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_,
    new_n4251_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4310_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_,
    new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_,
    new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_,
    new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_,
    new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_,
    new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_,
    new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_,
    new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_,
    new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_,
    new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_,
    new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_,
    new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_,
    new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_,
    new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_,
    new_n4477_, new_n4478_, new_n4479_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_,
    new_n4502_, new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_,
    new_n4508_, new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_,
    new_n4514_, new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_,
    new_n4520_, new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_,
    new_n4526_, new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_,
    new_n4532_, new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_,
    new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_,
    new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_,
    new_n4593_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4652_, new_n4653_, new_n4654_,
    new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_,
    new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_,
    new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_,
    new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_,
    new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_,
    new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_,
    new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_,
    new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_,
    new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_, new_n4782_,
    new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_,
    new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_,
    new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_,
    new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_,
    new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_,
    new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_,
    new_n4819_, new_n4820_, new_n4821_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4880_,
    new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_,
    new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_,
    new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_,
    new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_,
    new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_,
    new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_,
    new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_,
    new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_,
    new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_,
    new_n4935_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4994_, new_n4995_, new_n4996_,
    new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_,
    new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_,
    new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_,
    new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_,
    new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_,
    new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_,
    new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_,
    new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_,
    new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5108_, new_n5109_, new_n5111_, new_n5112_, new_n5114_,
    new_n5115_, new_n5117_, new_n5118_, new_n5120_, new_n5121_, new_n5123_,
    new_n5124_, new_n5126_, new_n5127_, new_n5129_, new_n5130_, new_n5132_,
    new_n5133_, new_n5135_, new_n5136_, new_n5138_, new_n5139_, new_n5141_,
    new_n5142_, new_n5144_, new_n5145_, new_n5147_, new_n5148_, new_n5150_,
    new_n5151_, new_n5153_, new_n5154_, new_n5156_, new_n5157_, new_n5159_,
    new_n5160_, new_n5162_, new_n5163_, new_n5165_, new_n5166_, new_n5168_,
    new_n5169_, new_n5171_, new_n5172_, new_n5174_, new_n5175_, new_n5177_,
    new_n5178_, new_n5180_, new_n5181_, new_n5183_, new_n5184_, new_n5186_,
    new_n5187_, new_n5189_, new_n5190_, new_n5192_, new_n5193_, new_n5195_,
    new_n5196_, new_n5198_, new_n5199_, new_n5201_, new_n5202_;
  assign new_n353_ = ~\p_input[30]  & ~\p_input[286] ;
  assign new_n354_ = \p_input[30]  & \p_input[286] ;
  assign new_n355_ = ~new_n353_ & ~new_n354_;
  assign new_n356_ = ~\p_input[29]  & ~\p_input[285] ;
  assign new_n357_ = \p_input[29]  & \p_input[285] ;
  assign new_n358_ = ~new_n356_ & ~new_n357_;
  assign new_n359_ = new_n355_ & new_n358_;
  assign new_n360_ = ~new_n355_ & ~new_n358_;
  assign new_n361_ = ~new_n359_ & ~new_n360_;
  assign new_n362_ = ~\p_input[31]  & ~\p_input[287] ;
  assign new_n363_ = \p_input[31]  & \p_input[287] ;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign new_n365_ = ~new_n361_ & ~new_n364_;
  assign new_n366_ = new_n361_ & new_n364_;
  assign new_n367_ = ~new_n365_ & ~new_n366_;
  assign new_n368_ = ~\p_input[25]  & ~\p_input[281] ;
  assign new_n369_ = \p_input[25]  & \p_input[281] ;
  assign new_n370_ = ~new_n368_ & ~new_n369_;
  assign new_n371_ = ~new_n367_ & ~new_n370_;
  assign new_n372_ = new_n367_ & new_n370_;
  assign new_n373_ = ~new_n371_ & ~new_n372_;
  assign new_n374_ = ~\p_input[27]  & ~\p_input[283] ;
  assign new_n375_ = \p_input[27]  & \p_input[283] ;
  assign new_n376_ = ~new_n374_ & ~new_n375_;
  assign new_n377_ = ~\p_input[26]  & ~\p_input[282] ;
  assign new_n378_ = \p_input[26]  & \p_input[282] ;
  assign new_n379_ = ~new_n377_ & ~new_n378_;
  assign new_n380_ = ~new_n376_ & ~new_n379_;
  assign new_n381_ = new_n376_ & new_n379_;
  assign new_n382_ = ~new_n380_ & ~new_n381_;
  assign new_n383_ = ~\p_input[28]  & ~\p_input[284] ;
  assign new_n384_ = \p_input[28]  & \p_input[284] ;
  assign new_n385_ = ~new_n383_ & ~new_n384_;
  assign new_n386_ = ~new_n382_ & ~new_n385_;
  assign new_n387_ = new_n382_ & new_n385_;
  assign new_n388_ = ~new_n386_ & ~new_n387_;
  assign new_n389_ = new_n373_ & ~new_n388_;
  assign new_n390_ = ~new_n371_ & ~new_n389_;
  assign new_n391_ = ~new_n359_ & ~new_n366_;
  assign new_n392_ = ~new_n390_ & new_n391_;
  assign new_n393_ = new_n390_ & ~new_n391_;
  assign new_n394_ = ~new_n392_ & ~new_n393_;
  assign new_n395_ = ~new_n381_ & ~new_n387_;
  assign new_n396_ = new_n394_ & new_n395_;
  assign new_n397_ = ~new_n392_ & ~new_n396_;
  assign new_n398_ = ~new_n394_ & ~new_n395_;
  assign new_n399_ = ~new_n396_ & ~new_n398_;
  assign new_n400_ = ~new_n373_ & new_n388_;
  assign new_n401_ = ~new_n389_ & ~new_n400_;
  assign new_n402_ = ~\p_input[17]  & ~\p_input[273] ;
  assign new_n403_ = \p_input[17]  & \p_input[273] ;
  assign new_n404_ = ~new_n402_ & ~new_n403_;
  assign new_n405_ = new_n401_ & ~new_n404_;
  assign new_n406_ = ~\p_input[23]  & ~\p_input[279] ;
  assign new_n407_ = \p_input[23]  & \p_input[279] ;
  assign new_n408_ = ~new_n406_ & ~new_n407_;
  assign new_n409_ = ~\p_input[22]  & ~\p_input[278] ;
  assign new_n410_ = \p_input[22]  & \p_input[278] ;
  assign new_n411_ = ~new_n409_ & ~new_n410_;
  assign new_n412_ = ~new_n408_ & ~new_n411_;
  assign new_n413_ = new_n408_ & new_n411_;
  assign new_n414_ = ~new_n412_ & ~new_n413_;
  assign new_n415_ = ~\p_input[24]  & ~\p_input[280] ;
  assign new_n416_ = \p_input[24]  & \p_input[280] ;
  assign new_n417_ = ~new_n415_ & ~new_n416_;
  assign new_n418_ = ~new_n414_ & ~new_n417_;
  assign new_n419_ = new_n414_ & new_n417_;
  assign new_n420_ = ~new_n418_ & ~new_n419_;
  assign new_n421_ = ~\p_input[18]  & ~\p_input[274] ;
  assign new_n422_ = \p_input[18]  & \p_input[274] ;
  assign new_n423_ = ~new_n421_ & ~new_n422_;
  assign new_n424_ = ~new_n420_ & ~new_n423_;
  assign new_n425_ = new_n420_ & new_n423_;
  assign new_n426_ = ~new_n424_ & ~new_n425_;
  assign new_n427_ = ~\p_input[20]  & ~\p_input[276] ;
  assign new_n428_ = \p_input[20]  & \p_input[276] ;
  assign new_n429_ = ~new_n427_ & ~new_n428_;
  assign new_n430_ = ~\p_input[19]  & ~\p_input[275] ;
  assign new_n431_ = \p_input[19]  & \p_input[275] ;
  assign new_n432_ = ~new_n430_ & ~new_n431_;
  assign new_n433_ = ~new_n429_ & ~new_n432_;
  assign new_n434_ = new_n429_ & new_n432_;
  assign new_n435_ = ~new_n433_ & ~new_n434_;
  assign new_n436_ = ~\p_input[21]  & ~\p_input[277] ;
  assign new_n437_ = \p_input[21]  & \p_input[277] ;
  assign new_n438_ = ~new_n436_ & ~new_n437_;
  assign new_n439_ = ~new_n435_ & ~new_n438_;
  assign new_n440_ = new_n435_ & new_n438_;
  assign new_n441_ = ~new_n439_ & ~new_n440_;
  assign new_n442_ = new_n426_ & ~new_n441_;
  assign new_n443_ = ~new_n426_ & new_n441_;
  assign new_n444_ = ~new_n442_ & ~new_n443_;
  assign new_n445_ = ~new_n401_ & new_n404_;
  assign new_n446_ = ~new_n405_ & ~new_n445_;
  assign new_n447_ = new_n444_ & new_n446_;
  assign new_n448_ = ~new_n405_ & ~new_n447_;
  assign new_n449_ = new_n399_ & ~new_n448_;
  assign new_n450_ = ~new_n424_ & ~new_n442_;
  assign new_n451_ = ~new_n413_ & ~new_n419_;
  assign new_n452_ = ~new_n450_ & new_n451_;
  assign new_n453_ = new_n450_ & ~new_n451_;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_ = ~new_n434_ & ~new_n440_;
  assign new_n456_ = new_n454_ & new_n455_;
  assign new_n457_ = ~new_n454_ & ~new_n455_;
  assign new_n458_ = ~new_n456_ & ~new_n457_;
  assign new_n459_ = ~new_n399_ & new_n448_;
  assign new_n460_ = ~new_n449_ & ~new_n459_;
  assign new_n461_ = new_n458_ & new_n460_;
  assign new_n462_ = ~new_n449_ & ~new_n461_;
  assign new_n463_ = ~new_n397_ & ~new_n462_;
  assign new_n464_ = new_n397_ & new_n462_;
  assign new_n465_ = ~new_n463_ & ~new_n464_;
  assign new_n466_ = ~new_n452_ & ~new_n456_;
  assign new_n467_ = new_n465_ & ~new_n466_;
  assign new_n468_ = ~new_n463_ & ~new_n467_;
  assign new_n469_ = ~new_n465_ & new_n466_;
  assign new_n470_ = ~new_n467_ & ~new_n469_;
  assign new_n471_ = ~new_n458_ & ~new_n460_;
  assign new_n472_ = ~new_n461_ & ~new_n471_;
  assign new_n473_ = ~new_n444_ & ~new_n446_;
  assign new_n474_ = ~new_n447_ & ~new_n473_;
  assign new_n475_ = ~\p_input[1]  & ~\p_input[257] ;
  assign new_n476_ = \p_input[1]  & \p_input[257] ;
  assign new_n477_ = ~new_n475_ & ~new_n476_;
  assign new_n478_ = new_n474_ & ~new_n477_;
  assign new_n479_ = ~\p_input[8]  & ~\p_input[264] ;
  assign new_n480_ = \p_input[8]  & \p_input[264] ;
  assign new_n481_ = ~new_n479_ & ~new_n480_;
  assign new_n482_ = ~\p_input[7]  & ~\p_input[263] ;
  assign new_n483_ = \p_input[7]  & \p_input[263] ;
  assign new_n484_ = ~new_n482_ & ~new_n483_;
  assign new_n485_ = ~new_n481_ & ~new_n484_;
  assign new_n486_ = new_n481_ & new_n484_;
  assign new_n487_ = ~new_n485_ & ~new_n486_;
  assign new_n488_ = ~\p_input[9]  & ~\p_input[265] ;
  assign new_n489_ = \p_input[9]  & \p_input[265] ;
  assign new_n490_ = ~new_n488_ & ~new_n489_;
  assign new_n491_ = ~new_n487_ & ~new_n490_;
  assign new_n492_ = new_n487_ & new_n490_;
  assign new_n493_ = ~new_n491_ & ~new_n492_;
  assign new_n494_ = ~\p_input[3]  & ~\p_input[259] ;
  assign new_n495_ = \p_input[3]  & \p_input[259] ;
  assign new_n496_ = ~new_n494_ & ~new_n495_;
  assign new_n497_ = ~new_n493_ & ~new_n496_;
  assign new_n498_ = new_n493_ & new_n496_;
  assign new_n499_ = ~new_n497_ & ~new_n498_;
  assign new_n500_ = ~\p_input[5]  & ~\p_input[261] ;
  assign new_n501_ = \p_input[5]  & \p_input[261] ;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = ~\p_input[4]  & ~\p_input[260] ;
  assign new_n504_ = \p_input[4]  & \p_input[260] ;
  assign new_n505_ = ~new_n503_ & ~new_n504_;
  assign new_n506_ = ~new_n502_ & ~new_n505_;
  assign new_n507_ = new_n502_ & new_n505_;
  assign new_n508_ = ~new_n506_ & ~new_n507_;
  assign new_n509_ = ~\p_input[6]  & ~\p_input[262] ;
  assign new_n510_ = \p_input[6]  & \p_input[262] ;
  assign new_n511_ = ~new_n509_ & ~new_n510_;
  assign new_n512_ = ~new_n508_ & ~new_n511_;
  assign new_n513_ = new_n508_ & new_n511_;
  assign new_n514_ = ~new_n512_ & ~new_n513_;
  assign new_n515_ = new_n499_ & ~new_n514_;
  assign new_n516_ = ~new_n499_ & new_n514_;
  assign new_n517_ = ~new_n515_ & ~new_n516_;
  assign new_n518_ = ~\p_input[15]  & ~\p_input[271] ;
  assign new_n519_ = \p_input[15]  & \p_input[271] ;
  assign new_n520_ = ~new_n518_ & ~new_n519_;
  assign new_n521_ = ~\p_input[14]  & ~\p_input[270] ;
  assign new_n522_ = \p_input[14]  & \p_input[270] ;
  assign new_n523_ = ~new_n521_ & ~new_n522_;
  assign new_n524_ = ~new_n520_ & ~new_n523_;
  assign new_n525_ = new_n520_ & new_n523_;
  assign new_n526_ = ~new_n524_ & ~new_n525_;
  assign new_n527_ = ~\p_input[16]  & ~\p_input[272] ;
  assign new_n528_ = \p_input[16]  & \p_input[272] ;
  assign new_n529_ = ~new_n527_ & ~new_n528_;
  assign new_n530_ = ~new_n526_ & ~new_n529_;
  assign new_n531_ = new_n526_ & new_n529_;
  assign new_n532_ = ~new_n530_ & ~new_n531_;
  assign new_n533_ = ~\p_input[10]  & ~\p_input[266] ;
  assign new_n534_ = \p_input[10]  & \p_input[266] ;
  assign new_n535_ = ~new_n533_ & ~new_n534_;
  assign new_n536_ = ~new_n532_ & ~new_n535_;
  assign new_n537_ = new_n532_ & new_n535_;
  assign new_n538_ = ~new_n536_ & ~new_n537_;
  assign new_n539_ = ~\p_input[12]  & ~\p_input[268] ;
  assign new_n540_ = \p_input[12]  & \p_input[268] ;
  assign new_n541_ = ~new_n539_ & ~new_n540_;
  assign new_n542_ = ~\p_input[11]  & ~\p_input[267] ;
  assign new_n543_ = \p_input[11]  & \p_input[267] ;
  assign new_n544_ = ~new_n542_ & ~new_n543_;
  assign new_n545_ = ~new_n541_ & ~new_n544_;
  assign new_n546_ = new_n541_ & new_n544_;
  assign new_n547_ = ~new_n545_ & ~new_n546_;
  assign new_n548_ = ~\p_input[13]  & ~\p_input[269] ;
  assign new_n549_ = \p_input[13]  & \p_input[269] ;
  assign new_n550_ = ~new_n548_ & ~new_n549_;
  assign new_n551_ = ~new_n547_ & ~new_n550_;
  assign new_n552_ = new_n547_ & new_n550_;
  assign new_n553_ = ~new_n551_ & ~new_n552_;
  assign new_n554_ = new_n538_ & ~new_n553_;
  assign new_n555_ = ~new_n538_ & new_n553_;
  assign new_n556_ = ~new_n554_ & ~new_n555_;
  assign new_n557_ = ~\p_input[2]  & ~\p_input[258] ;
  assign new_n558_ = \p_input[2]  & \p_input[258] ;
  assign new_n559_ = ~new_n557_ & ~new_n558_;
  assign new_n560_ = new_n556_ & ~new_n559_;
  assign new_n561_ = ~new_n556_ & new_n559_;
  assign new_n562_ = ~new_n560_ & ~new_n561_;
  assign new_n563_ = new_n517_ & new_n562_;
  assign new_n564_ = ~new_n517_ & ~new_n562_;
  assign new_n565_ = ~new_n563_ & ~new_n564_;
  assign new_n566_ = ~new_n474_ & new_n477_;
  assign new_n567_ = ~new_n478_ & ~new_n566_;
  assign new_n568_ = new_n565_ & new_n567_;
  assign new_n569_ = ~new_n478_ & ~new_n568_;
  assign new_n570_ = new_n472_ & ~new_n569_;
  assign new_n571_ = ~new_n497_ & ~new_n515_;
  assign new_n572_ = ~new_n486_ & ~new_n492_;
  assign new_n573_ = ~new_n571_ & new_n572_;
  assign new_n574_ = new_n571_ & ~new_n572_;
  assign new_n575_ = ~new_n573_ & ~new_n574_;
  assign new_n576_ = ~new_n507_ & ~new_n513_;
  assign new_n577_ = new_n575_ & new_n576_;
  assign new_n578_ = ~new_n575_ & ~new_n576_;
  assign new_n579_ = ~new_n577_ & ~new_n578_;
  assign new_n580_ = ~new_n536_ & ~new_n554_;
  assign new_n581_ = ~new_n525_ & ~new_n531_;
  assign new_n582_ = ~new_n580_ & new_n581_;
  assign new_n583_ = new_n580_ & ~new_n581_;
  assign new_n584_ = ~new_n582_ & ~new_n583_;
  assign new_n585_ = ~new_n546_ & ~new_n552_;
  assign new_n586_ = new_n584_ & new_n585_;
  assign new_n587_ = ~new_n584_ & ~new_n585_;
  assign new_n588_ = ~new_n586_ & ~new_n587_;
  assign new_n589_ = ~new_n560_ & ~new_n563_;
  assign new_n590_ = new_n588_ & ~new_n589_;
  assign new_n591_ = ~new_n588_ & new_n589_;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign new_n593_ = new_n579_ & new_n592_;
  assign new_n594_ = ~new_n579_ & ~new_n592_;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign new_n596_ = ~new_n472_ & new_n569_;
  assign new_n597_ = ~new_n570_ & ~new_n596_;
  assign new_n598_ = new_n595_ & new_n597_;
  assign new_n599_ = ~new_n570_ & ~new_n598_;
  assign new_n600_ = new_n470_ & ~new_n599_;
  assign new_n601_ = ~new_n582_ & ~new_n586_;
  assign new_n602_ = ~new_n590_ & ~new_n593_;
  assign new_n603_ = ~new_n601_ & ~new_n602_;
  assign new_n604_ = new_n601_ & new_n602_;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = ~new_n573_ & ~new_n577_;
  assign new_n607_ = new_n605_ & ~new_n606_;
  assign new_n608_ = ~new_n605_ & new_n606_;
  assign new_n609_ = ~new_n607_ & ~new_n608_;
  assign new_n610_ = ~new_n470_ & new_n599_;
  assign new_n611_ = ~new_n600_ & ~new_n610_;
  assign new_n612_ = new_n609_ & new_n611_;
  assign new_n613_ = ~new_n600_ & ~new_n612_;
  assign new_n614_ = ~new_n468_ & ~new_n613_;
  assign new_n615_ = new_n468_ & new_n613_;
  assign new_n616_ = ~new_n614_ & ~new_n615_;
  assign new_n617_ = ~new_n603_ & ~new_n607_;
  assign new_n618_ = new_n616_ & ~new_n617_;
  assign new_n619_ = ~new_n616_ & new_n617_;
  assign new_n620_ = ~new_n618_ & ~new_n619_;
  assign new_n621_ = ~new_n609_ & ~new_n611_;
  assign new_n622_ = ~new_n612_ & ~new_n621_;
  assign new_n623_ = ~new_n595_ & ~new_n597_;
  assign new_n624_ = ~new_n598_ & ~new_n623_;
  assign new_n625_ = ~new_n565_ & ~new_n567_;
  assign new_n626_ = ~new_n568_ & ~new_n625_;
  assign new_n627_ = ~\p_input[0]  & ~\p_input[256] ;
  assign new_n628_ = \p_input[0]  & \p_input[256] ;
  assign new_n629_ = ~new_n627_ & ~new_n628_;
  assign new_n630_ = ~new_n626_ & new_n629_;
  assign new_n631_ = ~new_n624_ & new_n630_;
  assign new_n632_ = ~new_n622_ & new_n631_;
  assign new_n633_ = ~new_n620_ & new_n632_;
  assign new_n634_ = ~new_n614_ & ~new_n618_;
  assign new_n635_ = new_n633_ & new_n634_;
  assign new_n636_ = ~\p_input[47]  & ~\p_input[271] ;
  assign new_n637_ = \p_input[47]  & \p_input[271] ;
  assign new_n638_ = ~new_n636_ & ~new_n637_;
  assign new_n639_ = ~\p_input[46]  & ~\p_input[270] ;
  assign new_n640_ = \p_input[46]  & \p_input[270] ;
  assign new_n641_ = ~new_n639_ & ~new_n640_;
  assign new_n642_ = ~new_n638_ & ~new_n641_;
  assign new_n643_ = new_n638_ & new_n641_;
  assign new_n644_ = ~new_n642_ & ~new_n643_;
  assign new_n645_ = ~\p_input[48]  & ~\p_input[272] ;
  assign new_n646_ = \p_input[48]  & \p_input[272] ;
  assign new_n647_ = ~new_n645_ & ~new_n646_;
  assign new_n648_ = ~new_n644_ & ~new_n647_;
  assign new_n649_ = new_n644_ & new_n647_;
  assign new_n650_ = ~new_n648_ & ~new_n649_;
  assign new_n651_ = ~\p_input[42]  & ~\p_input[266] ;
  assign new_n652_ = \p_input[42]  & \p_input[266] ;
  assign new_n653_ = ~new_n651_ & ~new_n652_;
  assign new_n654_ = ~new_n650_ & ~new_n653_;
  assign new_n655_ = new_n650_ & new_n653_;
  assign new_n656_ = ~new_n654_ & ~new_n655_;
  assign new_n657_ = ~\p_input[44]  & ~\p_input[268] ;
  assign new_n658_ = \p_input[44]  & \p_input[268] ;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign new_n660_ = ~\p_input[43]  & ~\p_input[267] ;
  assign new_n661_ = \p_input[43]  & \p_input[267] ;
  assign new_n662_ = ~new_n660_ & ~new_n661_;
  assign new_n663_ = ~new_n659_ & ~new_n662_;
  assign new_n664_ = new_n659_ & new_n662_;
  assign new_n665_ = ~new_n663_ & ~new_n664_;
  assign new_n666_ = ~\p_input[45]  & ~\p_input[269] ;
  assign new_n667_ = \p_input[45]  & \p_input[269] ;
  assign new_n668_ = ~new_n666_ & ~new_n667_;
  assign new_n669_ = ~new_n665_ & ~new_n668_;
  assign new_n670_ = new_n665_ & new_n668_;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = new_n656_ & ~new_n671_;
  assign new_n673_ = ~new_n654_ & ~new_n672_;
  assign new_n674_ = ~new_n643_ & ~new_n649_;
  assign new_n675_ = ~new_n673_ & new_n674_;
  assign new_n676_ = new_n673_ & ~new_n674_;
  assign new_n677_ = ~new_n675_ & ~new_n676_;
  assign new_n678_ = ~new_n664_ & ~new_n670_;
  assign new_n679_ = new_n677_ & new_n678_;
  assign new_n680_ = ~new_n675_ & ~new_n679_;
  assign new_n681_ = ~new_n677_ & ~new_n678_;
  assign new_n682_ = ~new_n679_ & ~new_n681_;
  assign new_n683_ = ~new_n656_ & new_n671_;
  assign new_n684_ = ~new_n672_ & ~new_n683_;
  assign new_n685_ = ~\p_input[34]  & ~\p_input[258] ;
  assign new_n686_ = \p_input[34]  & \p_input[258] ;
  assign new_n687_ = ~new_n685_ & ~new_n686_;
  assign new_n688_ = new_n684_ & ~new_n687_;
  assign new_n689_ = ~\p_input[40]  & ~\p_input[264] ;
  assign new_n690_ = \p_input[40]  & \p_input[264] ;
  assign new_n691_ = ~new_n689_ & ~new_n690_;
  assign new_n692_ = ~\p_input[39]  & ~\p_input[263] ;
  assign new_n693_ = \p_input[39]  & \p_input[263] ;
  assign new_n694_ = ~new_n692_ & ~new_n693_;
  assign new_n695_ = ~new_n691_ & ~new_n694_;
  assign new_n696_ = new_n691_ & new_n694_;
  assign new_n697_ = ~new_n695_ & ~new_n696_;
  assign new_n698_ = ~\p_input[41]  & ~\p_input[265] ;
  assign new_n699_ = \p_input[41]  & \p_input[265] ;
  assign new_n700_ = ~new_n698_ & ~new_n699_;
  assign new_n701_ = ~new_n697_ & ~new_n700_;
  assign new_n702_ = new_n697_ & new_n700_;
  assign new_n703_ = ~new_n701_ & ~new_n702_;
  assign new_n704_ = ~\p_input[35]  & ~\p_input[259] ;
  assign new_n705_ = \p_input[35]  & \p_input[259] ;
  assign new_n706_ = ~new_n704_ & ~new_n705_;
  assign new_n707_ = ~new_n703_ & ~new_n706_;
  assign new_n708_ = new_n703_ & new_n706_;
  assign new_n709_ = ~new_n707_ & ~new_n708_;
  assign new_n710_ = ~\p_input[37]  & ~\p_input[261] ;
  assign new_n711_ = \p_input[37]  & \p_input[261] ;
  assign new_n712_ = ~new_n710_ & ~new_n711_;
  assign new_n713_ = ~\p_input[36]  & ~\p_input[260] ;
  assign new_n714_ = \p_input[36]  & \p_input[260] ;
  assign new_n715_ = ~new_n713_ & ~new_n714_;
  assign new_n716_ = ~new_n712_ & ~new_n715_;
  assign new_n717_ = new_n712_ & new_n715_;
  assign new_n718_ = ~new_n716_ & ~new_n717_;
  assign new_n719_ = ~\p_input[38]  & ~\p_input[262] ;
  assign new_n720_ = \p_input[38]  & \p_input[262] ;
  assign new_n721_ = ~new_n719_ & ~new_n720_;
  assign new_n722_ = ~new_n718_ & ~new_n721_;
  assign new_n723_ = new_n718_ & new_n721_;
  assign new_n724_ = ~new_n722_ & ~new_n723_;
  assign new_n725_ = new_n709_ & ~new_n724_;
  assign new_n726_ = ~new_n709_ & new_n724_;
  assign new_n727_ = ~new_n725_ & ~new_n726_;
  assign new_n728_ = ~new_n684_ & new_n687_;
  assign new_n729_ = ~new_n688_ & ~new_n728_;
  assign new_n730_ = new_n727_ & new_n729_;
  assign new_n731_ = ~new_n688_ & ~new_n730_;
  assign new_n732_ = new_n682_ & ~new_n731_;
  assign new_n733_ = ~new_n707_ & ~new_n725_;
  assign new_n734_ = ~new_n696_ & ~new_n702_;
  assign new_n735_ = ~new_n733_ & new_n734_;
  assign new_n736_ = new_n733_ & ~new_n734_;
  assign new_n737_ = ~new_n735_ & ~new_n736_;
  assign new_n738_ = ~new_n717_ & ~new_n723_;
  assign new_n739_ = new_n737_ & new_n738_;
  assign new_n740_ = ~new_n737_ & ~new_n738_;
  assign new_n741_ = ~new_n739_ & ~new_n740_;
  assign new_n742_ = ~new_n682_ & new_n731_;
  assign new_n743_ = ~new_n732_ & ~new_n742_;
  assign new_n744_ = new_n741_ & new_n743_;
  assign new_n745_ = ~new_n732_ & ~new_n744_;
  assign new_n746_ = ~new_n680_ & ~new_n745_;
  assign new_n747_ = new_n680_ & new_n745_;
  assign new_n748_ = ~new_n746_ & ~new_n747_;
  assign new_n749_ = ~new_n735_ & ~new_n739_;
  assign new_n750_ = new_n748_ & ~new_n749_;
  assign new_n751_ = ~new_n748_ & new_n749_;
  assign new_n752_ = ~new_n750_ & ~new_n751_;
  assign new_n753_ = ~\p_input[62]  & ~\p_input[286] ;
  assign new_n754_ = \p_input[62]  & \p_input[286] ;
  assign new_n755_ = ~new_n753_ & ~new_n754_;
  assign new_n756_ = ~\p_input[61]  & ~\p_input[285] ;
  assign new_n757_ = \p_input[61]  & \p_input[285] ;
  assign new_n758_ = ~new_n756_ & ~new_n757_;
  assign new_n759_ = new_n755_ & new_n758_;
  assign new_n760_ = ~new_n755_ & ~new_n758_;
  assign new_n761_ = ~new_n759_ & ~new_n760_;
  assign new_n762_ = ~\p_input[63]  & ~\p_input[287] ;
  assign new_n763_ = \p_input[63]  & \p_input[287] ;
  assign new_n764_ = ~new_n762_ & ~new_n763_;
  assign new_n765_ = ~new_n761_ & ~new_n764_;
  assign new_n766_ = new_n761_ & new_n764_;
  assign new_n767_ = ~new_n765_ & ~new_n766_;
  assign new_n768_ = ~\p_input[57]  & ~\p_input[281] ;
  assign new_n769_ = \p_input[57]  & \p_input[281] ;
  assign new_n770_ = ~new_n768_ & ~new_n769_;
  assign new_n771_ = ~new_n767_ & ~new_n770_;
  assign new_n772_ = new_n767_ & new_n770_;
  assign new_n773_ = ~new_n771_ & ~new_n772_;
  assign new_n774_ = ~\p_input[59]  & ~\p_input[283] ;
  assign new_n775_ = \p_input[59]  & \p_input[283] ;
  assign new_n776_ = ~new_n774_ & ~new_n775_;
  assign new_n777_ = ~\p_input[58]  & ~\p_input[282] ;
  assign new_n778_ = \p_input[58]  & \p_input[282] ;
  assign new_n779_ = ~new_n777_ & ~new_n778_;
  assign new_n780_ = ~new_n776_ & ~new_n779_;
  assign new_n781_ = new_n776_ & new_n779_;
  assign new_n782_ = ~new_n780_ & ~new_n781_;
  assign new_n783_ = ~\p_input[60]  & ~\p_input[284] ;
  assign new_n784_ = \p_input[60]  & \p_input[284] ;
  assign new_n785_ = ~new_n783_ & ~new_n784_;
  assign new_n786_ = ~new_n782_ & ~new_n785_;
  assign new_n787_ = new_n782_ & new_n785_;
  assign new_n788_ = ~new_n786_ & ~new_n787_;
  assign new_n789_ = new_n773_ & ~new_n788_;
  assign new_n790_ = ~new_n771_ & ~new_n789_;
  assign new_n791_ = ~new_n759_ & ~new_n766_;
  assign new_n792_ = ~new_n790_ & new_n791_;
  assign new_n793_ = new_n790_ & ~new_n791_;
  assign new_n794_ = ~new_n792_ & ~new_n793_;
  assign new_n795_ = ~new_n781_ & ~new_n787_;
  assign new_n796_ = new_n794_ & new_n795_;
  assign new_n797_ = ~new_n792_ & ~new_n796_;
  assign new_n798_ = ~new_n794_ & ~new_n795_;
  assign new_n799_ = ~new_n796_ & ~new_n798_;
  assign new_n800_ = ~new_n773_ & new_n788_;
  assign new_n801_ = ~new_n789_ & ~new_n800_;
  assign new_n802_ = ~\p_input[49]  & ~\p_input[273] ;
  assign new_n803_ = \p_input[49]  & \p_input[273] ;
  assign new_n804_ = ~new_n802_ & ~new_n803_;
  assign new_n805_ = new_n801_ & ~new_n804_;
  assign new_n806_ = ~\p_input[55]  & ~\p_input[279] ;
  assign new_n807_ = \p_input[55]  & \p_input[279] ;
  assign new_n808_ = ~new_n806_ & ~new_n807_;
  assign new_n809_ = ~\p_input[54]  & ~\p_input[278] ;
  assign new_n810_ = \p_input[54]  & \p_input[278] ;
  assign new_n811_ = ~new_n809_ & ~new_n810_;
  assign new_n812_ = ~new_n808_ & ~new_n811_;
  assign new_n813_ = new_n808_ & new_n811_;
  assign new_n814_ = ~new_n812_ & ~new_n813_;
  assign new_n815_ = ~\p_input[56]  & ~\p_input[280] ;
  assign new_n816_ = \p_input[56]  & \p_input[280] ;
  assign new_n817_ = ~new_n815_ & ~new_n816_;
  assign new_n818_ = ~new_n814_ & ~new_n817_;
  assign new_n819_ = new_n814_ & new_n817_;
  assign new_n820_ = ~new_n818_ & ~new_n819_;
  assign new_n821_ = ~\p_input[50]  & ~\p_input[274] ;
  assign new_n822_ = \p_input[50]  & \p_input[274] ;
  assign new_n823_ = ~new_n821_ & ~new_n822_;
  assign new_n824_ = ~new_n820_ & ~new_n823_;
  assign new_n825_ = new_n820_ & new_n823_;
  assign new_n826_ = ~new_n824_ & ~new_n825_;
  assign new_n827_ = ~\p_input[52]  & ~\p_input[276] ;
  assign new_n828_ = \p_input[52]  & \p_input[276] ;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = ~\p_input[51]  & ~\p_input[275] ;
  assign new_n831_ = \p_input[51]  & \p_input[275] ;
  assign new_n832_ = ~new_n830_ & ~new_n831_;
  assign new_n833_ = ~new_n829_ & ~new_n832_;
  assign new_n834_ = new_n829_ & new_n832_;
  assign new_n835_ = ~new_n833_ & ~new_n834_;
  assign new_n836_ = ~\p_input[53]  & ~\p_input[277] ;
  assign new_n837_ = \p_input[53]  & \p_input[277] ;
  assign new_n838_ = ~new_n836_ & ~new_n837_;
  assign new_n839_ = ~new_n835_ & ~new_n838_;
  assign new_n840_ = new_n835_ & new_n838_;
  assign new_n841_ = ~new_n839_ & ~new_n840_;
  assign new_n842_ = new_n826_ & ~new_n841_;
  assign new_n843_ = ~new_n826_ & new_n841_;
  assign new_n844_ = ~new_n842_ & ~new_n843_;
  assign new_n845_ = ~new_n801_ & new_n804_;
  assign new_n846_ = ~new_n805_ & ~new_n845_;
  assign new_n847_ = new_n844_ & new_n846_;
  assign new_n848_ = ~new_n805_ & ~new_n847_;
  assign new_n849_ = new_n799_ & ~new_n848_;
  assign new_n850_ = ~new_n824_ & ~new_n842_;
  assign new_n851_ = ~new_n813_ & ~new_n819_;
  assign new_n852_ = ~new_n850_ & new_n851_;
  assign new_n853_ = new_n850_ & ~new_n851_;
  assign new_n854_ = ~new_n852_ & ~new_n853_;
  assign new_n855_ = ~new_n834_ & ~new_n840_;
  assign new_n856_ = new_n854_ & new_n855_;
  assign new_n857_ = ~new_n854_ & ~new_n855_;
  assign new_n858_ = ~new_n856_ & ~new_n857_;
  assign new_n859_ = ~new_n799_ & new_n848_;
  assign new_n860_ = ~new_n849_ & ~new_n859_;
  assign new_n861_ = new_n858_ & new_n860_;
  assign new_n862_ = ~new_n849_ & ~new_n861_;
  assign new_n863_ = ~new_n797_ & ~new_n862_;
  assign new_n864_ = new_n797_ & new_n862_;
  assign new_n865_ = ~new_n863_ & ~new_n864_;
  assign new_n866_ = ~new_n852_ & ~new_n856_;
  assign new_n867_ = new_n865_ & ~new_n866_;
  assign new_n868_ = ~new_n865_ & new_n866_;
  assign new_n869_ = ~new_n867_ & ~new_n868_;
  assign new_n870_ = ~new_n858_ & ~new_n860_;
  assign new_n871_ = ~new_n861_ & ~new_n870_;
  assign new_n872_ = ~new_n844_ & ~new_n846_;
  assign new_n873_ = ~new_n847_ & ~new_n872_;
  assign new_n874_ = ~\p_input[33]  & ~\p_input[257] ;
  assign new_n875_ = \p_input[33]  & \p_input[257] ;
  assign new_n876_ = ~new_n874_ & ~new_n875_;
  assign new_n877_ = new_n873_ & ~new_n876_;
  assign new_n878_ = ~new_n727_ & ~new_n729_;
  assign new_n879_ = ~new_n730_ & ~new_n878_;
  assign new_n880_ = ~new_n873_ & new_n876_;
  assign new_n881_ = ~new_n877_ & ~new_n880_;
  assign new_n882_ = new_n879_ & new_n881_;
  assign new_n883_ = ~new_n877_ & ~new_n882_;
  assign new_n884_ = new_n871_ & ~new_n883_;
  assign new_n885_ = ~new_n741_ & ~new_n743_;
  assign new_n886_ = ~new_n744_ & ~new_n885_;
  assign new_n887_ = ~new_n871_ & new_n883_;
  assign new_n888_ = ~new_n884_ & ~new_n887_;
  assign new_n889_ = new_n886_ & new_n888_;
  assign new_n890_ = ~new_n884_ & ~new_n889_;
  assign new_n891_ = new_n869_ & ~new_n890_;
  assign new_n892_ = ~new_n869_ & new_n890_;
  assign new_n893_ = ~new_n891_ & ~new_n892_;
  assign new_n894_ = new_n752_ & new_n893_;
  assign new_n895_ = ~new_n752_ & ~new_n893_;
  assign new_n896_ = ~new_n894_ & ~new_n895_;
  assign new_n897_ = ~new_n886_ & ~new_n888_;
  assign new_n898_ = ~new_n889_ & ~new_n897_;
  assign new_n899_ = ~new_n879_ & ~new_n881_;
  assign new_n900_ = ~new_n882_ & ~new_n899_;
  assign new_n901_ = ~\p_input[32]  & ~\p_input[256] ;
  assign new_n902_ = \p_input[32]  & \p_input[256] ;
  assign new_n903_ = ~new_n901_ & ~new_n902_;
  assign new_n904_ = ~new_n900_ & new_n903_;
  assign new_n905_ = ~new_n898_ & new_n904_;
  assign new_n906_ = ~new_n896_ & new_n905_;
  assign new_n907_ = ~new_n863_ & ~new_n867_;
  assign new_n908_ = ~new_n891_ & ~new_n894_;
  assign new_n909_ = ~new_n907_ & ~new_n908_;
  assign new_n910_ = new_n907_ & new_n908_;
  assign new_n911_ = ~new_n909_ & ~new_n910_;
  assign new_n912_ = ~new_n746_ & ~new_n750_;
  assign new_n913_ = new_n911_ & ~new_n912_;
  assign new_n914_ = ~new_n911_ & new_n912_;
  assign new_n915_ = ~new_n913_ & ~new_n914_;
  assign new_n916_ = new_n906_ & ~new_n915_;
  assign new_n917_ = ~new_n909_ & ~new_n913_;
  assign new_n918_ = new_n916_ & new_n917_;
  assign new_n919_ = ~\p_input[79]  & ~\p_input[271] ;
  assign new_n920_ = \p_input[79]  & \p_input[271] ;
  assign new_n921_ = ~new_n919_ & ~new_n920_;
  assign new_n922_ = ~\p_input[78]  & ~\p_input[270] ;
  assign new_n923_ = \p_input[78]  & \p_input[270] ;
  assign new_n924_ = ~new_n922_ & ~new_n923_;
  assign new_n925_ = ~new_n921_ & ~new_n924_;
  assign new_n926_ = new_n921_ & new_n924_;
  assign new_n927_ = ~new_n925_ & ~new_n926_;
  assign new_n928_ = ~\p_input[80]  & ~\p_input[272] ;
  assign new_n929_ = \p_input[80]  & \p_input[272] ;
  assign new_n930_ = ~new_n928_ & ~new_n929_;
  assign new_n931_ = ~new_n927_ & ~new_n930_;
  assign new_n932_ = new_n927_ & new_n930_;
  assign new_n933_ = ~new_n931_ & ~new_n932_;
  assign new_n934_ = ~\p_input[74]  & ~\p_input[266] ;
  assign new_n935_ = \p_input[74]  & \p_input[266] ;
  assign new_n936_ = ~new_n934_ & ~new_n935_;
  assign new_n937_ = ~new_n933_ & ~new_n936_;
  assign new_n938_ = new_n933_ & new_n936_;
  assign new_n939_ = ~new_n937_ & ~new_n938_;
  assign new_n940_ = ~\p_input[76]  & ~\p_input[268] ;
  assign new_n941_ = \p_input[76]  & \p_input[268] ;
  assign new_n942_ = ~new_n940_ & ~new_n941_;
  assign new_n943_ = ~\p_input[75]  & ~\p_input[267] ;
  assign new_n944_ = \p_input[75]  & \p_input[267] ;
  assign new_n945_ = ~new_n943_ & ~new_n944_;
  assign new_n946_ = ~new_n942_ & ~new_n945_;
  assign new_n947_ = new_n942_ & new_n945_;
  assign new_n948_ = ~new_n946_ & ~new_n947_;
  assign new_n949_ = ~\p_input[77]  & ~\p_input[269] ;
  assign new_n950_ = \p_input[77]  & \p_input[269] ;
  assign new_n951_ = ~new_n949_ & ~new_n950_;
  assign new_n952_ = ~new_n948_ & ~new_n951_;
  assign new_n953_ = new_n948_ & new_n951_;
  assign new_n954_ = ~new_n952_ & ~new_n953_;
  assign new_n955_ = new_n939_ & ~new_n954_;
  assign new_n956_ = ~new_n937_ & ~new_n955_;
  assign new_n957_ = ~new_n926_ & ~new_n932_;
  assign new_n958_ = ~new_n956_ & new_n957_;
  assign new_n959_ = new_n956_ & ~new_n957_;
  assign new_n960_ = ~new_n958_ & ~new_n959_;
  assign new_n961_ = ~new_n947_ & ~new_n953_;
  assign new_n962_ = new_n960_ & new_n961_;
  assign new_n963_ = ~new_n958_ & ~new_n962_;
  assign new_n964_ = ~new_n960_ & ~new_n961_;
  assign new_n965_ = ~new_n962_ & ~new_n964_;
  assign new_n966_ = ~new_n939_ & new_n954_;
  assign new_n967_ = ~new_n955_ & ~new_n966_;
  assign new_n968_ = ~\p_input[66]  & ~\p_input[258] ;
  assign new_n969_ = \p_input[66]  & \p_input[258] ;
  assign new_n970_ = ~new_n968_ & ~new_n969_;
  assign new_n971_ = new_n967_ & ~new_n970_;
  assign new_n972_ = ~\p_input[72]  & ~\p_input[264] ;
  assign new_n973_ = \p_input[72]  & \p_input[264] ;
  assign new_n974_ = ~new_n972_ & ~new_n973_;
  assign new_n975_ = ~\p_input[71]  & ~\p_input[263] ;
  assign new_n976_ = \p_input[71]  & \p_input[263] ;
  assign new_n977_ = ~new_n975_ & ~new_n976_;
  assign new_n978_ = ~new_n974_ & ~new_n977_;
  assign new_n979_ = new_n974_ & new_n977_;
  assign new_n980_ = ~new_n978_ & ~new_n979_;
  assign new_n981_ = ~\p_input[73]  & ~\p_input[265] ;
  assign new_n982_ = \p_input[73]  & \p_input[265] ;
  assign new_n983_ = ~new_n981_ & ~new_n982_;
  assign new_n984_ = ~new_n980_ & ~new_n983_;
  assign new_n985_ = new_n980_ & new_n983_;
  assign new_n986_ = ~new_n984_ & ~new_n985_;
  assign new_n987_ = ~\p_input[67]  & ~\p_input[259] ;
  assign new_n988_ = \p_input[67]  & \p_input[259] ;
  assign new_n989_ = ~new_n987_ & ~new_n988_;
  assign new_n990_ = ~new_n986_ & ~new_n989_;
  assign new_n991_ = new_n986_ & new_n989_;
  assign new_n992_ = ~new_n990_ & ~new_n991_;
  assign new_n993_ = ~\p_input[69]  & ~\p_input[261] ;
  assign new_n994_ = \p_input[69]  & \p_input[261] ;
  assign new_n995_ = ~new_n993_ & ~new_n994_;
  assign new_n996_ = ~\p_input[68]  & ~\p_input[260] ;
  assign new_n997_ = \p_input[68]  & \p_input[260] ;
  assign new_n998_ = ~new_n996_ & ~new_n997_;
  assign new_n999_ = ~new_n995_ & ~new_n998_;
  assign new_n1000_ = new_n995_ & new_n998_;
  assign new_n1001_ = ~new_n999_ & ~new_n1000_;
  assign new_n1002_ = ~\p_input[70]  & ~\p_input[262] ;
  assign new_n1003_ = \p_input[70]  & \p_input[262] ;
  assign new_n1004_ = ~new_n1002_ & ~new_n1003_;
  assign new_n1005_ = ~new_n1001_ & ~new_n1004_;
  assign new_n1006_ = new_n1001_ & new_n1004_;
  assign new_n1007_ = ~new_n1005_ & ~new_n1006_;
  assign new_n1008_ = new_n992_ & ~new_n1007_;
  assign new_n1009_ = ~new_n992_ & new_n1007_;
  assign new_n1010_ = ~new_n1008_ & ~new_n1009_;
  assign new_n1011_ = ~new_n967_ & new_n970_;
  assign new_n1012_ = ~new_n971_ & ~new_n1011_;
  assign new_n1013_ = new_n1010_ & new_n1012_;
  assign new_n1014_ = ~new_n971_ & ~new_n1013_;
  assign new_n1015_ = new_n965_ & ~new_n1014_;
  assign new_n1016_ = ~new_n990_ & ~new_n1008_;
  assign new_n1017_ = ~new_n979_ & ~new_n985_;
  assign new_n1018_ = ~new_n1016_ & new_n1017_;
  assign new_n1019_ = new_n1016_ & ~new_n1017_;
  assign new_n1020_ = ~new_n1018_ & ~new_n1019_;
  assign new_n1021_ = ~new_n1000_ & ~new_n1006_;
  assign new_n1022_ = new_n1020_ & new_n1021_;
  assign new_n1023_ = ~new_n1020_ & ~new_n1021_;
  assign new_n1024_ = ~new_n1022_ & ~new_n1023_;
  assign new_n1025_ = ~new_n965_ & new_n1014_;
  assign new_n1026_ = ~new_n1015_ & ~new_n1025_;
  assign new_n1027_ = new_n1024_ & new_n1026_;
  assign new_n1028_ = ~new_n1015_ & ~new_n1027_;
  assign new_n1029_ = ~new_n963_ & ~new_n1028_;
  assign new_n1030_ = new_n963_ & new_n1028_;
  assign new_n1031_ = ~new_n1029_ & ~new_n1030_;
  assign new_n1032_ = ~new_n1018_ & ~new_n1022_;
  assign new_n1033_ = new_n1031_ & ~new_n1032_;
  assign new_n1034_ = ~new_n1031_ & new_n1032_;
  assign new_n1035_ = ~new_n1033_ & ~new_n1034_;
  assign new_n1036_ = ~\p_input[94]  & ~\p_input[286] ;
  assign new_n1037_ = \p_input[94]  & \p_input[286] ;
  assign new_n1038_ = ~new_n1036_ & ~new_n1037_;
  assign new_n1039_ = ~\p_input[93]  & ~\p_input[285] ;
  assign new_n1040_ = \p_input[93]  & \p_input[285] ;
  assign new_n1041_ = ~new_n1039_ & ~new_n1040_;
  assign new_n1042_ = new_n1038_ & new_n1041_;
  assign new_n1043_ = ~new_n1038_ & ~new_n1041_;
  assign new_n1044_ = ~new_n1042_ & ~new_n1043_;
  assign new_n1045_ = ~\p_input[95]  & ~\p_input[287] ;
  assign new_n1046_ = \p_input[95]  & \p_input[287] ;
  assign new_n1047_ = ~new_n1045_ & ~new_n1046_;
  assign new_n1048_ = ~new_n1044_ & ~new_n1047_;
  assign new_n1049_ = new_n1044_ & new_n1047_;
  assign new_n1050_ = ~new_n1048_ & ~new_n1049_;
  assign new_n1051_ = ~\p_input[89]  & ~\p_input[281] ;
  assign new_n1052_ = \p_input[89]  & \p_input[281] ;
  assign new_n1053_ = ~new_n1051_ & ~new_n1052_;
  assign new_n1054_ = ~new_n1050_ & ~new_n1053_;
  assign new_n1055_ = new_n1050_ & new_n1053_;
  assign new_n1056_ = ~new_n1054_ & ~new_n1055_;
  assign new_n1057_ = ~\p_input[91]  & ~\p_input[283] ;
  assign new_n1058_ = \p_input[91]  & \p_input[283] ;
  assign new_n1059_ = ~new_n1057_ & ~new_n1058_;
  assign new_n1060_ = ~\p_input[90]  & ~\p_input[282] ;
  assign new_n1061_ = \p_input[90]  & \p_input[282] ;
  assign new_n1062_ = ~new_n1060_ & ~new_n1061_;
  assign new_n1063_ = ~new_n1059_ & ~new_n1062_;
  assign new_n1064_ = new_n1059_ & new_n1062_;
  assign new_n1065_ = ~new_n1063_ & ~new_n1064_;
  assign new_n1066_ = ~\p_input[92]  & ~\p_input[284] ;
  assign new_n1067_ = \p_input[92]  & \p_input[284] ;
  assign new_n1068_ = ~new_n1066_ & ~new_n1067_;
  assign new_n1069_ = ~new_n1065_ & ~new_n1068_;
  assign new_n1070_ = new_n1065_ & new_n1068_;
  assign new_n1071_ = ~new_n1069_ & ~new_n1070_;
  assign new_n1072_ = new_n1056_ & ~new_n1071_;
  assign new_n1073_ = ~new_n1054_ & ~new_n1072_;
  assign new_n1074_ = ~new_n1042_ & ~new_n1049_;
  assign new_n1075_ = ~new_n1073_ & new_n1074_;
  assign new_n1076_ = new_n1073_ & ~new_n1074_;
  assign new_n1077_ = ~new_n1075_ & ~new_n1076_;
  assign new_n1078_ = ~new_n1064_ & ~new_n1070_;
  assign new_n1079_ = new_n1077_ & new_n1078_;
  assign new_n1080_ = ~new_n1075_ & ~new_n1079_;
  assign new_n1081_ = ~new_n1077_ & ~new_n1078_;
  assign new_n1082_ = ~new_n1079_ & ~new_n1081_;
  assign new_n1083_ = ~new_n1056_ & new_n1071_;
  assign new_n1084_ = ~new_n1072_ & ~new_n1083_;
  assign new_n1085_ = ~\p_input[81]  & ~\p_input[273] ;
  assign new_n1086_ = \p_input[81]  & \p_input[273] ;
  assign new_n1087_ = ~new_n1085_ & ~new_n1086_;
  assign new_n1088_ = new_n1084_ & ~new_n1087_;
  assign new_n1089_ = ~\p_input[87]  & ~\p_input[279] ;
  assign new_n1090_ = \p_input[87]  & \p_input[279] ;
  assign new_n1091_ = ~new_n1089_ & ~new_n1090_;
  assign new_n1092_ = ~\p_input[86]  & ~\p_input[278] ;
  assign new_n1093_ = \p_input[86]  & \p_input[278] ;
  assign new_n1094_ = ~new_n1092_ & ~new_n1093_;
  assign new_n1095_ = ~new_n1091_ & ~new_n1094_;
  assign new_n1096_ = new_n1091_ & new_n1094_;
  assign new_n1097_ = ~new_n1095_ & ~new_n1096_;
  assign new_n1098_ = ~\p_input[88]  & ~\p_input[280] ;
  assign new_n1099_ = \p_input[88]  & \p_input[280] ;
  assign new_n1100_ = ~new_n1098_ & ~new_n1099_;
  assign new_n1101_ = ~new_n1097_ & ~new_n1100_;
  assign new_n1102_ = new_n1097_ & new_n1100_;
  assign new_n1103_ = ~new_n1101_ & ~new_n1102_;
  assign new_n1104_ = ~\p_input[82]  & ~\p_input[274] ;
  assign new_n1105_ = \p_input[82]  & \p_input[274] ;
  assign new_n1106_ = ~new_n1104_ & ~new_n1105_;
  assign new_n1107_ = ~new_n1103_ & ~new_n1106_;
  assign new_n1108_ = new_n1103_ & new_n1106_;
  assign new_n1109_ = ~new_n1107_ & ~new_n1108_;
  assign new_n1110_ = ~\p_input[84]  & ~\p_input[276] ;
  assign new_n1111_ = \p_input[84]  & \p_input[276] ;
  assign new_n1112_ = ~new_n1110_ & ~new_n1111_;
  assign new_n1113_ = ~\p_input[83]  & ~\p_input[275] ;
  assign new_n1114_ = \p_input[83]  & \p_input[275] ;
  assign new_n1115_ = ~new_n1113_ & ~new_n1114_;
  assign new_n1116_ = ~new_n1112_ & ~new_n1115_;
  assign new_n1117_ = new_n1112_ & new_n1115_;
  assign new_n1118_ = ~new_n1116_ & ~new_n1117_;
  assign new_n1119_ = ~\p_input[85]  & ~\p_input[277] ;
  assign new_n1120_ = \p_input[85]  & \p_input[277] ;
  assign new_n1121_ = ~new_n1119_ & ~new_n1120_;
  assign new_n1122_ = ~new_n1118_ & ~new_n1121_;
  assign new_n1123_ = new_n1118_ & new_n1121_;
  assign new_n1124_ = ~new_n1122_ & ~new_n1123_;
  assign new_n1125_ = new_n1109_ & ~new_n1124_;
  assign new_n1126_ = ~new_n1109_ & new_n1124_;
  assign new_n1127_ = ~new_n1125_ & ~new_n1126_;
  assign new_n1128_ = ~new_n1084_ & new_n1087_;
  assign new_n1129_ = ~new_n1088_ & ~new_n1128_;
  assign new_n1130_ = new_n1127_ & new_n1129_;
  assign new_n1131_ = ~new_n1088_ & ~new_n1130_;
  assign new_n1132_ = new_n1082_ & ~new_n1131_;
  assign new_n1133_ = ~new_n1107_ & ~new_n1125_;
  assign new_n1134_ = ~new_n1096_ & ~new_n1102_;
  assign new_n1135_ = ~new_n1133_ & new_n1134_;
  assign new_n1136_ = new_n1133_ & ~new_n1134_;
  assign new_n1137_ = ~new_n1135_ & ~new_n1136_;
  assign new_n1138_ = ~new_n1117_ & ~new_n1123_;
  assign new_n1139_ = new_n1137_ & new_n1138_;
  assign new_n1140_ = ~new_n1137_ & ~new_n1138_;
  assign new_n1141_ = ~new_n1139_ & ~new_n1140_;
  assign new_n1142_ = ~new_n1082_ & new_n1131_;
  assign new_n1143_ = ~new_n1132_ & ~new_n1142_;
  assign new_n1144_ = new_n1141_ & new_n1143_;
  assign new_n1145_ = ~new_n1132_ & ~new_n1144_;
  assign new_n1146_ = ~new_n1080_ & ~new_n1145_;
  assign new_n1147_ = new_n1080_ & new_n1145_;
  assign new_n1148_ = ~new_n1146_ & ~new_n1147_;
  assign new_n1149_ = ~new_n1135_ & ~new_n1139_;
  assign new_n1150_ = new_n1148_ & ~new_n1149_;
  assign new_n1151_ = ~new_n1148_ & new_n1149_;
  assign new_n1152_ = ~new_n1150_ & ~new_n1151_;
  assign new_n1153_ = ~new_n1141_ & ~new_n1143_;
  assign new_n1154_ = ~new_n1144_ & ~new_n1153_;
  assign new_n1155_ = ~new_n1127_ & ~new_n1129_;
  assign new_n1156_ = ~new_n1130_ & ~new_n1155_;
  assign new_n1157_ = ~\p_input[65]  & ~\p_input[257] ;
  assign new_n1158_ = \p_input[65]  & \p_input[257] ;
  assign new_n1159_ = ~new_n1157_ & ~new_n1158_;
  assign new_n1160_ = new_n1156_ & ~new_n1159_;
  assign new_n1161_ = ~new_n1010_ & ~new_n1012_;
  assign new_n1162_ = ~new_n1013_ & ~new_n1161_;
  assign new_n1163_ = ~new_n1156_ & new_n1159_;
  assign new_n1164_ = ~new_n1160_ & ~new_n1163_;
  assign new_n1165_ = new_n1162_ & new_n1164_;
  assign new_n1166_ = ~new_n1160_ & ~new_n1165_;
  assign new_n1167_ = new_n1154_ & ~new_n1166_;
  assign new_n1168_ = ~new_n1024_ & ~new_n1026_;
  assign new_n1169_ = ~new_n1027_ & ~new_n1168_;
  assign new_n1170_ = ~new_n1154_ & new_n1166_;
  assign new_n1171_ = ~new_n1167_ & ~new_n1170_;
  assign new_n1172_ = new_n1169_ & new_n1171_;
  assign new_n1173_ = ~new_n1167_ & ~new_n1172_;
  assign new_n1174_ = new_n1152_ & ~new_n1173_;
  assign new_n1175_ = ~new_n1152_ & new_n1173_;
  assign new_n1176_ = ~new_n1174_ & ~new_n1175_;
  assign new_n1177_ = new_n1035_ & new_n1176_;
  assign new_n1178_ = ~new_n1035_ & ~new_n1176_;
  assign new_n1179_ = ~new_n1177_ & ~new_n1178_;
  assign new_n1180_ = ~new_n1169_ & ~new_n1171_;
  assign new_n1181_ = ~new_n1172_ & ~new_n1180_;
  assign new_n1182_ = ~new_n1162_ & ~new_n1164_;
  assign new_n1183_ = ~new_n1165_ & ~new_n1182_;
  assign new_n1184_ = ~\p_input[64]  & ~\p_input[256] ;
  assign new_n1185_ = \p_input[64]  & \p_input[256] ;
  assign new_n1186_ = ~new_n1184_ & ~new_n1185_;
  assign new_n1187_ = ~new_n1183_ & new_n1186_;
  assign new_n1188_ = ~new_n1181_ & new_n1187_;
  assign new_n1189_ = ~new_n1179_ & new_n1188_;
  assign new_n1190_ = ~new_n1146_ & ~new_n1150_;
  assign new_n1191_ = ~new_n1174_ & ~new_n1177_;
  assign new_n1192_ = ~new_n1190_ & ~new_n1191_;
  assign new_n1193_ = new_n1190_ & new_n1191_;
  assign new_n1194_ = ~new_n1192_ & ~new_n1193_;
  assign new_n1195_ = ~new_n1029_ & ~new_n1033_;
  assign new_n1196_ = new_n1194_ & ~new_n1195_;
  assign new_n1197_ = ~new_n1194_ & new_n1195_;
  assign new_n1198_ = ~new_n1196_ & ~new_n1197_;
  assign new_n1199_ = new_n1189_ & ~new_n1198_;
  assign new_n1200_ = ~new_n1192_ & ~new_n1196_;
  assign new_n1201_ = new_n1199_ & new_n1200_;
  assign new_n1202_ = ~\p_input[111]  & ~\p_input[271] ;
  assign new_n1203_ = \p_input[111]  & \p_input[271] ;
  assign new_n1204_ = ~new_n1202_ & ~new_n1203_;
  assign new_n1205_ = ~\p_input[110]  & ~\p_input[270] ;
  assign new_n1206_ = \p_input[110]  & \p_input[270] ;
  assign new_n1207_ = ~new_n1205_ & ~new_n1206_;
  assign new_n1208_ = ~new_n1204_ & ~new_n1207_;
  assign new_n1209_ = new_n1204_ & new_n1207_;
  assign new_n1210_ = ~new_n1208_ & ~new_n1209_;
  assign new_n1211_ = ~\p_input[112]  & ~\p_input[272] ;
  assign new_n1212_ = \p_input[112]  & \p_input[272] ;
  assign new_n1213_ = ~new_n1211_ & ~new_n1212_;
  assign new_n1214_ = ~new_n1210_ & ~new_n1213_;
  assign new_n1215_ = new_n1210_ & new_n1213_;
  assign new_n1216_ = ~new_n1214_ & ~new_n1215_;
  assign new_n1217_ = ~\p_input[106]  & ~\p_input[266] ;
  assign new_n1218_ = \p_input[106]  & \p_input[266] ;
  assign new_n1219_ = ~new_n1217_ & ~new_n1218_;
  assign new_n1220_ = ~new_n1216_ & ~new_n1219_;
  assign new_n1221_ = new_n1216_ & new_n1219_;
  assign new_n1222_ = ~new_n1220_ & ~new_n1221_;
  assign new_n1223_ = ~\p_input[108]  & ~\p_input[268] ;
  assign new_n1224_ = \p_input[108]  & \p_input[268] ;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = ~\p_input[107]  & ~\p_input[267] ;
  assign new_n1227_ = \p_input[107]  & \p_input[267] ;
  assign new_n1228_ = ~new_n1226_ & ~new_n1227_;
  assign new_n1229_ = ~new_n1225_ & ~new_n1228_;
  assign new_n1230_ = new_n1225_ & new_n1228_;
  assign new_n1231_ = ~new_n1229_ & ~new_n1230_;
  assign new_n1232_ = ~\p_input[109]  & ~\p_input[269] ;
  assign new_n1233_ = \p_input[109]  & \p_input[269] ;
  assign new_n1234_ = ~new_n1232_ & ~new_n1233_;
  assign new_n1235_ = ~new_n1231_ & ~new_n1234_;
  assign new_n1236_ = new_n1231_ & new_n1234_;
  assign new_n1237_ = ~new_n1235_ & ~new_n1236_;
  assign new_n1238_ = new_n1222_ & ~new_n1237_;
  assign new_n1239_ = ~new_n1220_ & ~new_n1238_;
  assign new_n1240_ = ~new_n1209_ & ~new_n1215_;
  assign new_n1241_ = ~new_n1239_ & new_n1240_;
  assign new_n1242_ = new_n1239_ & ~new_n1240_;
  assign new_n1243_ = ~new_n1241_ & ~new_n1242_;
  assign new_n1244_ = ~new_n1230_ & ~new_n1236_;
  assign new_n1245_ = new_n1243_ & new_n1244_;
  assign new_n1246_ = ~new_n1241_ & ~new_n1245_;
  assign new_n1247_ = ~new_n1243_ & ~new_n1244_;
  assign new_n1248_ = ~new_n1245_ & ~new_n1247_;
  assign new_n1249_ = ~new_n1222_ & new_n1237_;
  assign new_n1250_ = ~new_n1238_ & ~new_n1249_;
  assign new_n1251_ = ~\p_input[98]  & ~\p_input[258] ;
  assign new_n1252_ = \p_input[98]  & \p_input[258] ;
  assign new_n1253_ = ~new_n1251_ & ~new_n1252_;
  assign new_n1254_ = new_n1250_ & ~new_n1253_;
  assign new_n1255_ = ~\p_input[104]  & ~\p_input[264] ;
  assign new_n1256_ = \p_input[104]  & \p_input[264] ;
  assign new_n1257_ = ~new_n1255_ & ~new_n1256_;
  assign new_n1258_ = ~\p_input[103]  & ~\p_input[263] ;
  assign new_n1259_ = \p_input[103]  & \p_input[263] ;
  assign new_n1260_ = ~new_n1258_ & ~new_n1259_;
  assign new_n1261_ = ~new_n1257_ & ~new_n1260_;
  assign new_n1262_ = new_n1257_ & new_n1260_;
  assign new_n1263_ = ~new_n1261_ & ~new_n1262_;
  assign new_n1264_ = ~\p_input[105]  & ~\p_input[265] ;
  assign new_n1265_ = \p_input[105]  & \p_input[265] ;
  assign new_n1266_ = ~new_n1264_ & ~new_n1265_;
  assign new_n1267_ = ~new_n1263_ & ~new_n1266_;
  assign new_n1268_ = new_n1263_ & new_n1266_;
  assign new_n1269_ = ~new_n1267_ & ~new_n1268_;
  assign new_n1270_ = ~\p_input[99]  & ~\p_input[259] ;
  assign new_n1271_ = \p_input[99]  & \p_input[259] ;
  assign new_n1272_ = ~new_n1270_ & ~new_n1271_;
  assign new_n1273_ = ~new_n1269_ & ~new_n1272_;
  assign new_n1274_ = new_n1269_ & new_n1272_;
  assign new_n1275_ = ~new_n1273_ & ~new_n1274_;
  assign new_n1276_ = ~\p_input[101]  & ~\p_input[261] ;
  assign new_n1277_ = \p_input[101]  & \p_input[261] ;
  assign new_n1278_ = ~new_n1276_ & ~new_n1277_;
  assign new_n1279_ = ~\p_input[100]  & ~\p_input[260] ;
  assign new_n1280_ = \p_input[100]  & \p_input[260] ;
  assign new_n1281_ = ~new_n1279_ & ~new_n1280_;
  assign new_n1282_ = ~new_n1278_ & ~new_n1281_;
  assign new_n1283_ = new_n1278_ & new_n1281_;
  assign new_n1284_ = ~new_n1282_ & ~new_n1283_;
  assign new_n1285_ = ~\p_input[102]  & ~\p_input[262] ;
  assign new_n1286_ = \p_input[102]  & \p_input[262] ;
  assign new_n1287_ = ~new_n1285_ & ~new_n1286_;
  assign new_n1288_ = ~new_n1284_ & ~new_n1287_;
  assign new_n1289_ = new_n1284_ & new_n1287_;
  assign new_n1290_ = ~new_n1288_ & ~new_n1289_;
  assign new_n1291_ = new_n1275_ & ~new_n1290_;
  assign new_n1292_ = ~new_n1275_ & new_n1290_;
  assign new_n1293_ = ~new_n1291_ & ~new_n1292_;
  assign new_n1294_ = ~new_n1250_ & new_n1253_;
  assign new_n1295_ = ~new_n1254_ & ~new_n1294_;
  assign new_n1296_ = new_n1293_ & new_n1295_;
  assign new_n1297_ = ~new_n1254_ & ~new_n1296_;
  assign new_n1298_ = new_n1248_ & ~new_n1297_;
  assign new_n1299_ = ~new_n1273_ & ~new_n1291_;
  assign new_n1300_ = ~new_n1262_ & ~new_n1268_;
  assign new_n1301_ = ~new_n1299_ & new_n1300_;
  assign new_n1302_ = new_n1299_ & ~new_n1300_;
  assign new_n1303_ = ~new_n1301_ & ~new_n1302_;
  assign new_n1304_ = ~new_n1283_ & ~new_n1289_;
  assign new_n1305_ = new_n1303_ & new_n1304_;
  assign new_n1306_ = ~new_n1303_ & ~new_n1304_;
  assign new_n1307_ = ~new_n1305_ & ~new_n1306_;
  assign new_n1308_ = ~new_n1248_ & new_n1297_;
  assign new_n1309_ = ~new_n1298_ & ~new_n1308_;
  assign new_n1310_ = new_n1307_ & new_n1309_;
  assign new_n1311_ = ~new_n1298_ & ~new_n1310_;
  assign new_n1312_ = ~new_n1246_ & ~new_n1311_;
  assign new_n1313_ = new_n1246_ & new_n1311_;
  assign new_n1314_ = ~new_n1312_ & ~new_n1313_;
  assign new_n1315_ = ~new_n1301_ & ~new_n1305_;
  assign new_n1316_ = new_n1314_ & ~new_n1315_;
  assign new_n1317_ = ~new_n1314_ & new_n1315_;
  assign new_n1318_ = ~new_n1316_ & ~new_n1317_;
  assign new_n1319_ = ~\p_input[126]  & ~\p_input[286] ;
  assign new_n1320_ = \p_input[126]  & \p_input[286] ;
  assign new_n1321_ = ~new_n1319_ & ~new_n1320_;
  assign new_n1322_ = ~\p_input[125]  & ~\p_input[285] ;
  assign new_n1323_ = \p_input[125]  & \p_input[285] ;
  assign new_n1324_ = ~new_n1322_ & ~new_n1323_;
  assign new_n1325_ = new_n1321_ & new_n1324_;
  assign new_n1326_ = ~new_n1321_ & ~new_n1324_;
  assign new_n1327_ = ~new_n1325_ & ~new_n1326_;
  assign new_n1328_ = ~\p_input[127]  & ~\p_input[287] ;
  assign new_n1329_ = \p_input[127]  & \p_input[287] ;
  assign new_n1330_ = ~new_n1328_ & ~new_n1329_;
  assign new_n1331_ = ~new_n1327_ & ~new_n1330_;
  assign new_n1332_ = new_n1327_ & new_n1330_;
  assign new_n1333_ = ~new_n1331_ & ~new_n1332_;
  assign new_n1334_ = ~\p_input[121]  & ~\p_input[281] ;
  assign new_n1335_ = \p_input[121]  & \p_input[281] ;
  assign new_n1336_ = ~new_n1334_ & ~new_n1335_;
  assign new_n1337_ = ~new_n1333_ & ~new_n1336_;
  assign new_n1338_ = new_n1333_ & new_n1336_;
  assign new_n1339_ = ~new_n1337_ & ~new_n1338_;
  assign new_n1340_ = ~\p_input[123]  & ~\p_input[283] ;
  assign new_n1341_ = \p_input[123]  & \p_input[283] ;
  assign new_n1342_ = ~new_n1340_ & ~new_n1341_;
  assign new_n1343_ = ~\p_input[122]  & ~\p_input[282] ;
  assign new_n1344_ = \p_input[122]  & \p_input[282] ;
  assign new_n1345_ = ~new_n1343_ & ~new_n1344_;
  assign new_n1346_ = ~new_n1342_ & ~new_n1345_;
  assign new_n1347_ = new_n1342_ & new_n1345_;
  assign new_n1348_ = ~new_n1346_ & ~new_n1347_;
  assign new_n1349_ = ~\p_input[124]  & ~\p_input[284] ;
  assign new_n1350_ = \p_input[124]  & \p_input[284] ;
  assign new_n1351_ = ~new_n1349_ & ~new_n1350_;
  assign new_n1352_ = ~new_n1348_ & ~new_n1351_;
  assign new_n1353_ = new_n1348_ & new_n1351_;
  assign new_n1354_ = ~new_n1352_ & ~new_n1353_;
  assign new_n1355_ = new_n1339_ & ~new_n1354_;
  assign new_n1356_ = ~new_n1337_ & ~new_n1355_;
  assign new_n1357_ = ~new_n1325_ & ~new_n1332_;
  assign new_n1358_ = ~new_n1356_ & new_n1357_;
  assign new_n1359_ = new_n1356_ & ~new_n1357_;
  assign new_n1360_ = ~new_n1358_ & ~new_n1359_;
  assign new_n1361_ = ~new_n1347_ & ~new_n1353_;
  assign new_n1362_ = new_n1360_ & new_n1361_;
  assign new_n1363_ = ~new_n1358_ & ~new_n1362_;
  assign new_n1364_ = ~new_n1360_ & ~new_n1361_;
  assign new_n1365_ = ~new_n1362_ & ~new_n1364_;
  assign new_n1366_ = ~new_n1339_ & new_n1354_;
  assign new_n1367_ = ~new_n1355_ & ~new_n1366_;
  assign new_n1368_ = ~\p_input[113]  & ~\p_input[273] ;
  assign new_n1369_ = \p_input[113]  & \p_input[273] ;
  assign new_n1370_ = ~new_n1368_ & ~new_n1369_;
  assign new_n1371_ = new_n1367_ & ~new_n1370_;
  assign new_n1372_ = ~\p_input[119]  & ~\p_input[279] ;
  assign new_n1373_ = \p_input[119]  & \p_input[279] ;
  assign new_n1374_ = ~new_n1372_ & ~new_n1373_;
  assign new_n1375_ = ~\p_input[118]  & ~\p_input[278] ;
  assign new_n1376_ = \p_input[118]  & \p_input[278] ;
  assign new_n1377_ = ~new_n1375_ & ~new_n1376_;
  assign new_n1378_ = ~new_n1374_ & ~new_n1377_;
  assign new_n1379_ = new_n1374_ & new_n1377_;
  assign new_n1380_ = ~new_n1378_ & ~new_n1379_;
  assign new_n1381_ = ~\p_input[120]  & ~\p_input[280] ;
  assign new_n1382_ = \p_input[120]  & \p_input[280] ;
  assign new_n1383_ = ~new_n1381_ & ~new_n1382_;
  assign new_n1384_ = ~new_n1380_ & ~new_n1383_;
  assign new_n1385_ = new_n1380_ & new_n1383_;
  assign new_n1386_ = ~new_n1384_ & ~new_n1385_;
  assign new_n1387_ = ~\p_input[114]  & ~\p_input[274] ;
  assign new_n1388_ = \p_input[114]  & \p_input[274] ;
  assign new_n1389_ = ~new_n1387_ & ~new_n1388_;
  assign new_n1390_ = ~new_n1386_ & ~new_n1389_;
  assign new_n1391_ = new_n1386_ & new_n1389_;
  assign new_n1392_ = ~new_n1390_ & ~new_n1391_;
  assign new_n1393_ = ~\p_input[116]  & ~\p_input[276] ;
  assign new_n1394_ = \p_input[116]  & \p_input[276] ;
  assign new_n1395_ = ~new_n1393_ & ~new_n1394_;
  assign new_n1396_ = ~\p_input[115]  & ~\p_input[275] ;
  assign new_n1397_ = \p_input[115]  & \p_input[275] ;
  assign new_n1398_ = ~new_n1396_ & ~new_n1397_;
  assign new_n1399_ = ~new_n1395_ & ~new_n1398_;
  assign new_n1400_ = new_n1395_ & new_n1398_;
  assign new_n1401_ = ~new_n1399_ & ~new_n1400_;
  assign new_n1402_ = ~\p_input[117]  & ~\p_input[277] ;
  assign new_n1403_ = \p_input[117]  & \p_input[277] ;
  assign new_n1404_ = ~new_n1402_ & ~new_n1403_;
  assign new_n1405_ = ~new_n1401_ & ~new_n1404_;
  assign new_n1406_ = new_n1401_ & new_n1404_;
  assign new_n1407_ = ~new_n1405_ & ~new_n1406_;
  assign new_n1408_ = new_n1392_ & ~new_n1407_;
  assign new_n1409_ = ~new_n1392_ & new_n1407_;
  assign new_n1410_ = ~new_n1408_ & ~new_n1409_;
  assign new_n1411_ = ~new_n1367_ & new_n1370_;
  assign new_n1412_ = ~new_n1371_ & ~new_n1411_;
  assign new_n1413_ = new_n1410_ & new_n1412_;
  assign new_n1414_ = ~new_n1371_ & ~new_n1413_;
  assign new_n1415_ = new_n1365_ & ~new_n1414_;
  assign new_n1416_ = ~new_n1390_ & ~new_n1408_;
  assign new_n1417_ = ~new_n1379_ & ~new_n1385_;
  assign new_n1418_ = ~new_n1416_ & new_n1417_;
  assign new_n1419_ = new_n1416_ & ~new_n1417_;
  assign new_n1420_ = ~new_n1418_ & ~new_n1419_;
  assign new_n1421_ = ~new_n1400_ & ~new_n1406_;
  assign new_n1422_ = new_n1420_ & new_n1421_;
  assign new_n1423_ = ~new_n1420_ & ~new_n1421_;
  assign new_n1424_ = ~new_n1422_ & ~new_n1423_;
  assign new_n1425_ = ~new_n1365_ & new_n1414_;
  assign new_n1426_ = ~new_n1415_ & ~new_n1425_;
  assign new_n1427_ = new_n1424_ & new_n1426_;
  assign new_n1428_ = ~new_n1415_ & ~new_n1427_;
  assign new_n1429_ = ~new_n1363_ & ~new_n1428_;
  assign new_n1430_ = new_n1363_ & new_n1428_;
  assign new_n1431_ = ~new_n1429_ & ~new_n1430_;
  assign new_n1432_ = ~new_n1418_ & ~new_n1422_;
  assign new_n1433_ = new_n1431_ & ~new_n1432_;
  assign new_n1434_ = ~new_n1431_ & new_n1432_;
  assign new_n1435_ = ~new_n1433_ & ~new_n1434_;
  assign new_n1436_ = ~new_n1424_ & ~new_n1426_;
  assign new_n1437_ = ~new_n1427_ & ~new_n1436_;
  assign new_n1438_ = ~new_n1410_ & ~new_n1412_;
  assign new_n1439_ = ~new_n1413_ & ~new_n1438_;
  assign new_n1440_ = ~\p_input[97]  & ~\p_input[257] ;
  assign new_n1441_ = \p_input[97]  & \p_input[257] ;
  assign new_n1442_ = ~new_n1440_ & ~new_n1441_;
  assign new_n1443_ = new_n1439_ & ~new_n1442_;
  assign new_n1444_ = ~new_n1293_ & ~new_n1295_;
  assign new_n1445_ = ~new_n1296_ & ~new_n1444_;
  assign new_n1446_ = ~new_n1439_ & new_n1442_;
  assign new_n1447_ = ~new_n1443_ & ~new_n1446_;
  assign new_n1448_ = new_n1445_ & new_n1447_;
  assign new_n1449_ = ~new_n1443_ & ~new_n1448_;
  assign new_n1450_ = new_n1437_ & ~new_n1449_;
  assign new_n1451_ = ~new_n1307_ & ~new_n1309_;
  assign new_n1452_ = ~new_n1310_ & ~new_n1451_;
  assign new_n1453_ = ~new_n1437_ & new_n1449_;
  assign new_n1454_ = ~new_n1450_ & ~new_n1453_;
  assign new_n1455_ = new_n1452_ & new_n1454_;
  assign new_n1456_ = ~new_n1450_ & ~new_n1455_;
  assign new_n1457_ = new_n1435_ & ~new_n1456_;
  assign new_n1458_ = ~new_n1435_ & new_n1456_;
  assign new_n1459_ = ~new_n1457_ & ~new_n1458_;
  assign new_n1460_ = new_n1318_ & new_n1459_;
  assign new_n1461_ = ~new_n1318_ & ~new_n1459_;
  assign new_n1462_ = ~new_n1460_ & ~new_n1461_;
  assign new_n1463_ = ~new_n1452_ & ~new_n1454_;
  assign new_n1464_ = ~new_n1455_ & ~new_n1463_;
  assign new_n1465_ = ~new_n1445_ & ~new_n1447_;
  assign new_n1466_ = ~new_n1448_ & ~new_n1465_;
  assign new_n1467_ = ~\p_input[96]  & ~\p_input[256] ;
  assign new_n1468_ = \p_input[96]  & \p_input[256] ;
  assign new_n1469_ = ~new_n1467_ & ~new_n1468_;
  assign new_n1470_ = ~new_n1466_ & new_n1469_;
  assign new_n1471_ = ~new_n1464_ & new_n1470_;
  assign new_n1472_ = ~new_n1462_ & new_n1471_;
  assign new_n1473_ = ~new_n1429_ & ~new_n1433_;
  assign new_n1474_ = ~new_n1457_ & ~new_n1460_;
  assign new_n1475_ = ~new_n1473_ & ~new_n1474_;
  assign new_n1476_ = new_n1473_ & new_n1474_;
  assign new_n1477_ = ~new_n1475_ & ~new_n1476_;
  assign new_n1478_ = ~new_n1312_ & ~new_n1316_;
  assign new_n1479_ = new_n1477_ & ~new_n1478_;
  assign new_n1480_ = ~new_n1477_ & new_n1478_;
  assign new_n1481_ = ~new_n1479_ & ~new_n1480_;
  assign new_n1482_ = new_n1472_ & ~new_n1481_;
  assign new_n1483_ = ~new_n1475_ & ~new_n1479_;
  assign new_n1484_ = new_n1482_ & new_n1483_;
  assign new_n1485_ = ~\p_input[175]  & ~\p_input[271] ;
  assign new_n1486_ = \p_input[175]  & \p_input[271] ;
  assign new_n1487_ = ~new_n1485_ & ~new_n1486_;
  assign new_n1488_ = ~\p_input[174]  & ~\p_input[270] ;
  assign new_n1489_ = \p_input[174]  & \p_input[270] ;
  assign new_n1490_ = ~new_n1488_ & ~new_n1489_;
  assign new_n1491_ = ~new_n1487_ & ~new_n1490_;
  assign new_n1492_ = new_n1487_ & new_n1490_;
  assign new_n1493_ = ~new_n1491_ & ~new_n1492_;
  assign new_n1494_ = ~\p_input[176]  & ~\p_input[272] ;
  assign new_n1495_ = \p_input[176]  & \p_input[272] ;
  assign new_n1496_ = ~new_n1494_ & ~new_n1495_;
  assign new_n1497_ = ~new_n1493_ & ~new_n1496_;
  assign new_n1498_ = new_n1493_ & new_n1496_;
  assign new_n1499_ = ~new_n1497_ & ~new_n1498_;
  assign new_n1500_ = ~\p_input[170]  & ~\p_input[266] ;
  assign new_n1501_ = \p_input[170]  & \p_input[266] ;
  assign new_n1502_ = ~new_n1500_ & ~new_n1501_;
  assign new_n1503_ = ~new_n1499_ & ~new_n1502_;
  assign new_n1504_ = new_n1499_ & new_n1502_;
  assign new_n1505_ = ~new_n1503_ & ~new_n1504_;
  assign new_n1506_ = ~\p_input[172]  & ~\p_input[268] ;
  assign new_n1507_ = \p_input[172]  & \p_input[268] ;
  assign new_n1508_ = ~new_n1506_ & ~new_n1507_;
  assign new_n1509_ = ~\p_input[171]  & ~\p_input[267] ;
  assign new_n1510_ = \p_input[171]  & \p_input[267] ;
  assign new_n1511_ = ~new_n1509_ & ~new_n1510_;
  assign new_n1512_ = ~new_n1508_ & ~new_n1511_;
  assign new_n1513_ = new_n1508_ & new_n1511_;
  assign new_n1514_ = ~new_n1512_ & ~new_n1513_;
  assign new_n1515_ = ~\p_input[173]  & ~\p_input[269] ;
  assign new_n1516_ = \p_input[173]  & \p_input[269] ;
  assign new_n1517_ = ~new_n1515_ & ~new_n1516_;
  assign new_n1518_ = ~new_n1514_ & ~new_n1517_;
  assign new_n1519_ = new_n1514_ & new_n1517_;
  assign new_n1520_ = ~new_n1518_ & ~new_n1519_;
  assign new_n1521_ = new_n1505_ & ~new_n1520_;
  assign new_n1522_ = ~new_n1503_ & ~new_n1521_;
  assign new_n1523_ = ~new_n1492_ & ~new_n1498_;
  assign new_n1524_ = ~new_n1522_ & new_n1523_;
  assign new_n1525_ = new_n1522_ & ~new_n1523_;
  assign new_n1526_ = ~new_n1524_ & ~new_n1525_;
  assign new_n1527_ = ~new_n1513_ & ~new_n1519_;
  assign new_n1528_ = new_n1526_ & new_n1527_;
  assign new_n1529_ = ~new_n1524_ & ~new_n1528_;
  assign new_n1530_ = ~new_n1526_ & ~new_n1527_;
  assign new_n1531_ = ~new_n1528_ & ~new_n1530_;
  assign new_n1532_ = ~new_n1505_ & new_n1520_;
  assign new_n1533_ = ~new_n1521_ & ~new_n1532_;
  assign new_n1534_ = ~\p_input[162]  & ~\p_input[258] ;
  assign new_n1535_ = \p_input[162]  & \p_input[258] ;
  assign new_n1536_ = ~new_n1534_ & ~new_n1535_;
  assign new_n1537_ = new_n1533_ & ~new_n1536_;
  assign new_n1538_ = ~\p_input[168]  & ~\p_input[264] ;
  assign new_n1539_ = \p_input[168]  & \p_input[264] ;
  assign new_n1540_ = ~new_n1538_ & ~new_n1539_;
  assign new_n1541_ = ~\p_input[167]  & ~\p_input[263] ;
  assign new_n1542_ = \p_input[167]  & \p_input[263] ;
  assign new_n1543_ = ~new_n1541_ & ~new_n1542_;
  assign new_n1544_ = ~new_n1540_ & ~new_n1543_;
  assign new_n1545_ = new_n1540_ & new_n1543_;
  assign new_n1546_ = ~new_n1544_ & ~new_n1545_;
  assign new_n1547_ = ~\p_input[169]  & ~\p_input[265] ;
  assign new_n1548_ = \p_input[169]  & \p_input[265] ;
  assign new_n1549_ = ~new_n1547_ & ~new_n1548_;
  assign new_n1550_ = ~new_n1546_ & ~new_n1549_;
  assign new_n1551_ = new_n1546_ & new_n1549_;
  assign new_n1552_ = ~new_n1550_ & ~new_n1551_;
  assign new_n1553_ = ~\p_input[163]  & ~\p_input[259] ;
  assign new_n1554_ = \p_input[163]  & \p_input[259] ;
  assign new_n1555_ = ~new_n1553_ & ~new_n1554_;
  assign new_n1556_ = ~new_n1552_ & ~new_n1555_;
  assign new_n1557_ = new_n1552_ & new_n1555_;
  assign new_n1558_ = ~new_n1556_ & ~new_n1557_;
  assign new_n1559_ = ~\p_input[165]  & ~\p_input[261] ;
  assign new_n1560_ = \p_input[165]  & \p_input[261] ;
  assign new_n1561_ = ~new_n1559_ & ~new_n1560_;
  assign new_n1562_ = ~\p_input[164]  & ~\p_input[260] ;
  assign new_n1563_ = \p_input[164]  & \p_input[260] ;
  assign new_n1564_ = ~new_n1562_ & ~new_n1563_;
  assign new_n1565_ = ~new_n1561_ & ~new_n1564_;
  assign new_n1566_ = new_n1561_ & new_n1564_;
  assign new_n1567_ = ~new_n1565_ & ~new_n1566_;
  assign new_n1568_ = ~\p_input[166]  & ~\p_input[262] ;
  assign new_n1569_ = \p_input[166]  & \p_input[262] ;
  assign new_n1570_ = ~new_n1568_ & ~new_n1569_;
  assign new_n1571_ = ~new_n1567_ & ~new_n1570_;
  assign new_n1572_ = new_n1567_ & new_n1570_;
  assign new_n1573_ = ~new_n1571_ & ~new_n1572_;
  assign new_n1574_ = new_n1558_ & ~new_n1573_;
  assign new_n1575_ = ~new_n1558_ & new_n1573_;
  assign new_n1576_ = ~new_n1574_ & ~new_n1575_;
  assign new_n1577_ = ~new_n1533_ & new_n1536_;
  assign new_n1578_ = ~new_n1537_ & ~new_n1577_;
  assign new_n1579_ = new_n1576_ & new_n1578_;
  assign new_n1580_ = ~new_n1537_ & ~new_n1579_;
  assign new_n1581_ = new_n1531_ & ~new_n1580_;
  assign new_n1582_ = ~new_n1556_ & ~new_n1574_;
  assign new_n1583_ = ~new_n1545_ & ~new_n1551_;
  assign new_n1584_ = ~new_n1582_ & new_n1583_;
  assign new_n1585_ = new_n1582_ & ~new_n1583_;
  assign new_n1586_ = ~new_n1584_ & ~new_n1585_;
  assign new_n1587_ = ~new_n1566_ & ~new_n1572_;
  assign new_n1588_ = new_n1586_ & new_n1587_;
  assign new_n1589_ = ~new_n1586_ & ~new_n1587_;
  assign new_n1590_ = ~new_n1588_ & ~new_n1589_;
  assign new_n1591_ = ~new_n1531_ & new_n1580_;
  assign new_n1592_ = ~new_n1581_ & ~new_n1591_;
  assign new_n1593_ = new_n1590_ & new_n1592_;
  assign new_n1594_ = ~new_n1581_ & ~new_n1593_;
  assign new_n1595_ = ~new_n1529_ & ~new_n1594_;
  assign new_n1596_ = new_n1529_ & new_n1594_;
  assign new_n1597_ = ~new_n1595_ & ~new_n1596_;
  assign new_n1598_ = ~new_n1584_ & ~new_n1588_;
  assign new_n1599_ = new_n1597_ & ~new_n1598_;
  assign new_n1600_ = ~new_n1597_ & new_n1598_;
  assign new_n1601_ = ~new_n1599_ & ~new_n1600_;
  assign new_n1602_ = ~\p_input[190]  & ~\p_input[286] ;
  assign new_n1603_ = \p_input[190]  & \p_input[286] ;
  assign new_n1604_ = ~new_n1602_ & ~new_n1603_;
  assign new_n1605_ = ~\p_input[189]  & ~\p_input[285] ;
  assign new_n1606_ = \p_input[189]  & \p_input[285] ;
  assign new_n1607_ = ~new_n1605_ & ~new_n1606_;
  assign new_n1608_ = new_n1604_ & new_n1607_;
  assign new_n1609_ = ~new_n1604_ & ~new_n1607_;
  assign new_n1610_ = ~new_n1608_ & ~new_n1609_;
  assign new_n1611_ = ~\p_input[191]  & ~\p_input[287] ;
  assign new_n1612_ = \p_input[191]  & \p_input[287] ;
  assign new_n1613_ = ~new_n1611_ & ~new_n1612_;
  assign new_n1614_ = ~new_n1610_ & ~new_n1613_;
  assign new_n1615_ = new_n1610_ & new_n1613_;
  assign new_n1616_ = ~new_n1614_ & ~new_n1615_;
  assign new_n1617_ = ~\p_input[185]  & ~\p_input[281] ;
  assign new_n1618_ = \p_input[185]  & \p_input[281] ;
  assign new_n1619_ = ~new_n1617_ & ~new_n1618_;
  assign new_n1620_ = ~new_n1616_ & ~new_n1619_;
  assign new_n1621_ = new_n1616_ & new_n1619_;
  assign new_n1622_ = ~new_n1620_ & ~new_n1621_;
  assign new_n1623_ = ~\p_input[187]  & ~\p_input[283] ;
  assign new_n1624_ = \p_input[187]  & \p_input[283] ;
  assign new_n1625_ = ~new_n1623_ & ~new_n1624_;
  assign new_n1626_ = ~\p_input[186]  & ~\p_input[282] ;
  assign new_n1627_ = \p_input[186]  & \p_input[282] ;
  assign new_n1628_ = ~new_n1626_ & ~new_n1627_;
  assign new_n1629_ = ~new_n1625_ & ~new_n1628_;
  assign new_n1630_ = new_n1625_ & new_n1628_;
  assign new_n1631_ = ~new_n1629_ & ~new_n1630_;
  assign new_n1632_ = ~\p_input[188]  & ~\p_input[284] ;
  assign new_n1633_ = \p_input[188]  & \p_input[284] ;
  assign new_n1634_ = ~new_n1632_ & ~new_n1633_;
  assign new_n1635_ = ~new_n1631_ & ~new_n1634_;
  assign new_n1636_ = new_n1631_ & new_n1634_;
  assign new_n1637_ = ~new_n1635_ & ~new_n1636_;
  assign new_n1638_ = new_n1622_ & ~new_n1637_;
  assign new_n1639_ = ~new_n1620_ & ~new_n1638_;
  assign new_n1640_ = ~new_n1608_ & ~new_n1615_;
  assign new_n1641_ = ~new_n1639_ & new_n1640_;
  assign new_n1642_ = new_n1639_ & ~new_n1640_;
  assign new_n1643_ = ~new_n1641_ & ~new_n1642_;
  assign new_n1644_ = ~new_n1630_ & ~new_n1636_;
  assign new_n1645_ = new_n1643_ & new_n1644_;
  assign new_n1646_ = ~new_n1641_ & ~new_n1645_;
  assign new_n1647_ = ~new_n1643_ & ~new_n1644_;
  assign new_n1648_ = ~new_n1645_ & ~new_n1647_;
  assign new_n1649_ = ~new_n1622_ & new_n1637_;
  assign new_n1650_ = ~new_n1638_ & ~new_n1649_;
  assign new_n1651_ = ~\p_input[177]  & ~\p_input[273] ;
  assign new_n1652_ = \p_input[177]  & \p_input[273] ;
  assign new_n1653_ = ~new_n1651_ & ~new_n1652_;
  assign new_n1654_ = new_n1650_ & ~new_n1653_;
  assign new_n1655_ = ~\p_input[183]  & ~\p_input[279] ;
  assign new_n1656_ = \p_input[183]  & \p_input[279] ;
  assign new_n1657_ = ~new_n1655_ & ~new_n1656_;
  assign new_n1658_ = ~\p_input[182]  & ~\p_input[278] ;
  assign new_n1659_ = \p_input[182]  & \p_input[278] ;
  assign new_n1660_ = ~new_n1658_ & ~new_n1659_;
  assign new_n1661_ = ~new_n1657_ & ~new_n1660_;
  assign new_n1662_ = new_n1657_ & new_n1660_;
  assign new_n1663_ = ~new_n1661_ & ~new_n1662_;
  assign new_n1664_ = ~\p_input[184]  & ~\p_input[280] ;
  assign new_n1665_ = \p_input[184]  & \p_input[280] ;
  assign new_n1666_ = ~new_n1664_ & ~new_n1665_;
  assign new_n1667_ = ~new_n1663_ & ~new_n1666_;
  assign new_n1668_ = new_n1663_ & new_n1666_;
  assign new_n1669_ = ~new_n1667_ & ~new_n1668_;
  assign new_n1670_ = ~\p_input[178]  & ~\p_input[274] ;
  assign new_n1671_ = \p_input[178]  & \p_input[274] ;
  assign new_n1672_ = ~new_n1670_ & ~new_n1671_;
  assign new_n1673_ = ~new_n1669_ & ~new_n1672_;
  assign new_n1674_ = new_n1669_ & new_n1672_;
  assign new_n1675_ = ~new_n1673_ & ~new_n1674_;
  assign new_n1676_ = ~\p_input[180]  & ~\p_input[276] ;
  assign new_n1677_ = \p_input[180]  & \p_input[276] ;
  assign new_n1678_ = ~new_n1676_ & ~new_n1677_;
  assign new_n1679_ = ~\p_input[179]  & ~\p_input[275] ;
  assign new_n1680_ = \p_input[179]  & \p_input[275] ;
  assign new_n1681_ = ~new_n1679_ & ~new_n1680_;
  assign new_n1682_ = ~new_n1678_ & ~new_n1681_;
  assign new_n1683_ = new_n1678_ & new_n1681_;
  assign new_n1684_ = ~new_n1682_ & ~new_n1683_;
  assign new_n1685_ = ~\p_input[181]  & ~\p_input[277] ;
  assign new_n1686_ = \p_input[181]  & \p_input[277] ;
  assign new_n1687_ = ~new_n1685_ & ~new_n1686_;
  assign new_n1688_ = ~new_n1684_ & ~new_n1687_;
  assign new_n1689_ = new_n1684_ & new_n1687_;
  assign new_n1690_ = ~new_n1688_ & ~new_n1689_;
  assign new_n1691_ = new_n1675_ & ~new_n1690_;
  assign new_n1692_ = ~new_n1675_ & new_n1690_;
  assign new_n1693_ = ~new_n1691_ & ~new_n1692_;
  assign new_n1694_ = ~new_n1650_ & new_n1653_;
  assign new_n1695_ = ~new_n1654_ & ~new_n1694_;
  assign new_n1696_ = new_n1693_ & new_n1695_;
  assign new_n1697_ = ~new_n1654_ & ~new_n1696_;
  assign new_n1698_ = new_n1648_ & ~new_n1697_;
  assign new_n1699_ = ~new_n1673_ & ~new_n1691_;
  assign new_n1700_ = ~new_n1662_ & ~new_n1668_;
  assign new_n1701_ = ~new_n1699_ & new_n1700_;
  assign new_n1702_ = new_n1699_ & ~new_n1700_;
  assign new_n1703_ = ~new_n1701_ & ~new_n1702_;
  assign new_n1704_ = ~new_n1683_ & ~new_n1689_;
  assign new_n1705_ = new_n1703_ & new_n1704_;
  assign new_n1706_ = ~new_n1703_ & ~new_n1704_;
  assign new_n1707_ = ~new_n1705_ & ~new_n1706_;
  assign new_n1708_ = ~new_n1648_ & new_n1697_;
  assign new_n1709_ = ~new_n1698_ & ~new_n1708_;
  assign new_n1710_ = new_n1707_ & new_n1709_;
  assign new_n1711_ = ~new_n1698_ & ~new_n1710_;
  assign new_n1712_ = ~new_n1646_ & ~new_n1711_;
  assign new_n1713_ = new_n1646_ & new_n1711_;
  assign new_n1714_ = ~new_n1712_ & ~new_n1713_;
  assign new_n1715_ = ~new_n1701_ & ~new_n1705_;
  assign new_n1716_ = new_n1714_ & ~new_n1715_;
  assign new_n1717_ = ~new_n1714_ & new_n1715_;
  assign new_n1718_ = ~new_n1716_ & ~new_n1717_;
  assign new_n1719_ = ~new_n1707_ & ~new_n1709_;
  assign new_n1720_ = ~new_n1710_ & ~new_n1719_;
  assign new_n1721_ = ~new_n1693_ & ~new_n1695_;
  assign new_n1722_ = ~new_n1696_ & ~new_n1721_;
  assign new_n1723_ = ~\p_input[161]  & ~\p_input[257] ;
  assign new_n1724_ = \p_input[161]  & \p_input[257] ;
  assign new_n1725_ = ~new_n1723_ & ~new_n1724_;
  assign new_n1726_ = new_n1722_ & ~new_n1725_;
  assign new_n1727_ = ~new_n1576_ & ~new_n1578_;
  assign new_n1728_ = ~new_n1579_ & ~new_n1727_;
  assign new_n1729_ = ~new_n1722_ & new_n1725_;
  assign new_n1730_ = ~new_n1726_ & ~new_n1729_;
  assign new_n1731_ = new_n1728_ & new_n1730_;
  assign new_n1732_ = ~new_n1726_ & ~new_n1731_;
  assign new_n1733_ = new_n1720_ & ~new_n1732_;
  assign new_n1734_ = ~new_n1590_ & ~new_n1592_;
  assign new_n1735_ = ~new_n1593_ & ~new_n1734_;
  assign new_n1736_ = ~new_n1720_ & new_n1732_;
  assign new_n1737_ = ~new_n1733_ & ~new_n1736_;
  assign new_n1738_ = new_n1735_ & new_n1737_;
  assign new_n1739_ = ~new_n1733_ & ~new_n1738_;
  assign new_n1740_ = new_n1718_ & ~new_n1739_;
  assign new_n1741_ = ~new_n1718_ & new_n1739_;
  assign new_n1742_ = ~new_n1740_ & ~new_n1741_;
  assign new_n1743_ = new_n1601_ & new_n1742_;
  assign new_n1744_ = ~new_n1601_ & ~new_n1742_;
  assign new_n1745_ = ~new_n1743_ & ~new_n1744_;
  assign new_n1746_ = ~new_n1735_ & ~new_n1737_;
  assign new_n1747_ = ~new_n1738_ & ~new_n1746_;
  assign new_n1748_ = ~new_n1728_ & ~new_n1730_;
  assign new_n1749_ = ~new_n1731_ & ~new_n1748_;
  assign new_n1750_ = ~\p_input[160]  & ~\p_input[256] ;
  assign new_n1751_ = \p_input[160]  & \p_input[256] ;
  assign new_n1752_ = ~new_n1750_ & ~new_n1751_;
  assign new_n1753_ = ~new_n1749_ & new_n1752_;
  assign new_n1754_ = ~new_n1747_ & new_n1753_;
  assign new_n1755_ = ~new_n1745_ & new_n1754_;
  assign new_n1756_ = ~new_n1712_ & ~new_n1716_;
  assign new_n1757_ = ~new_n1740_ & ~new_n1743_;
  assign new_n1758_ = ~new_n1756_ & ~new_n1757_;
  assign new_n1759_ = new_n1756_ & new_n1757_;
  assign new_n1760_ = ~new_n1758_ & ~new_n1759_;
  assign new_n1761_ = ~new_n1595_ & ~new_n1599_;
  assign new_n1762_ = new_n1760_ & ~new_n1761_;
  assign new_n1763_ = ~new_n1760_ & new_n1761_;
  assign new_n1764_ = ~new_n1762_ & ~new_n1763_;
  assign new_n1765_ = new_n1755_ & ~new_n1764_;
  assign new_n1766_ = ~new_n1758_ & ~new_n1762_;
  assign new_n1767_ = new_n1765_ & new_n1766_;
  assign new_n1768_ = ~\p_input[254]  & ~\p_input[286] ;
  assign new_n1769_ = \p_input[254]  & \p_input[286] ;
  assign new_n1770_ = ~new_n1768_ & ~new_n1769_;
  assign new_n1771_ = ~\p_input[253]  & ~\p_input[285] ;
  assign new_n1772_ = \p_input[253]  & \p_input[285] ;
  assign new_n1773_ = ~new_n1771_ & ~new_n1772_;
  assign new_n1774_ = new_n1770_ & new_n1773_;
  assign new_n1775_ = ~new_n1770_ & ~new_n1773_;
  assign new_n1776_ = ~new_n1774_ & ~new_n1775_;
  assign new_n1777_ = ~\p_input[255]  & ~\p_input[287] ;
  assign new_n1778_ = \p_input[255]  & \p_input[287] ;
  assign new_n1779_ = ~new_n1777_ & ~new_n1778_;
  assign new_n1780_ = new_n1776_ & new_n1779_;
  assign new_n1781_ = ~new_n1774_ & ~new_n1780_;
  assign new_n1782_ = ~new_n1776_ & ~new_n1779_;
  assign new_n1783_ = ~new_n1780_ & ~new_n1782_;
  assign new_n1784_ = ~\p_input[249]  & ~\p_input[281] ;
  assign new_n1785_ = \p_input[249]  & \p_input[281] ;
  assign new_n1786_ = ~new_n1784_ & ~new_n1785_;
  assign new_n1787_ = new_n1783_ & new_n1786_;
  assign new_n1788_ = ~new_n1783_ & ~new_n1786_;
  assign new_n1789_ = ~\p_input[251]  & ~\p_input[283] ;
  assign new_n1790_ = \p_input[251]  & \p_input[283] ;
  assign new_n1791_ = ~new_n1789_ & ~new_n1790_;
  assign new_n1792_ = ~\p_input[250]  & ~\p_input[282] ;
  assign new_n1793_ = \p_input[250]  & \p_input[282] ;
  assign new_n1794_ = ~new_n1792_ & ~new_n1793_;
  assign new_n1795_ = ~new_n1791_ & ~new_n1794_;
  assign new_n1796_ = new_n1791_ & new_n1794_;
  assign new_n1797_ = ~new_n1795_ & ~new_n1796_;
  assign new_n1798_ = ~\p_input[252]  & ~\p_input[284] ;
  assign new_n1799_ = \p_input[252]  & \p_input[284] ;
  assign new_n1800_ = ~new_n1798_ & ~new_n1799_;
  assign new_n1801_ = ~new_n1797_ & ~new_n1800_;
  assign new_n1802_ = new_n1797_ & new_n1800_;
  assign new_n1803_ = ~new_n1801_ & ~new_n1802_;
  assign new_n1804_ = ~new_n1788_ & new_n1803_;
  assign new_n1805_ = ~new_n1787_ & ~new_n1804_;
  assign new_n1806_ = new_n1781_ & new_n1805_;
  assign new_n1807_ = ~new_n1781_ & ~new_n1805_;
  assign new_n1808_ = ~new_n1806_ & ~new_n1807_;
  assign new_n1809_ = ~new_n1796_ & ~new_n1802_;
  assign new_n1810_ = new_n1808_ & new_n1809_;
  assign new_n1811_ = ~new_n1806_ & ~new_n1810_;
  assign new_n1812_ = ~new_n1808_ & ~new_n1809_;
  assign new_n1813_ = ~new_n1810_ & ~new_n1812_;
  assign new_n1814_ = ~new_n1787_ & ~new_n1788_;
  assign new_n1815_ = ~new_n1803_ & new_n1814_;
  assign new_n1816_ = new_n1803_ & ~new_n1814_;
  assign new_n1817_ = ~new_n1815_ & ~new_n1816_;
  assign new_n1818_ = ~\p_input[241]  & ~\p_input[273] ;
  assign new_n1819_ = \p_input[241]  & \p_input[273] ;
  assign new_n1820_ = ~new_n1818_ & ~new_n1819_;
  assign new_n1821_ = ~new_n1817_ & new_n1820_;
  assign new_n1822_ = new_n1817_ & ~new_n1820_;
  assign new_n1823_ = ~\p_input[247]  & ~\p_input[279] ;
  assign new_n1824_ = \p_input[247]  & \p_input[279] ;
  assign new_n1825_ = ~new_n1823_ & ~new_n1824_;
  assign new_n1826_ = ~\p_input[246]  & ~\p_input[278] ;
  assign new_n1827_ = \p_input[246]  & \p_input[278] ;
  assign new_n1828_ = ~new_n1826_ & ~new_n1827_;
  assign new_n1829_ = ~new_n1825_ & ~new_n1828_;
  assign new_n1830_ = new_n1825_ & new_n1828_;
  assign new_n1831_ = ~new_n1829_ & ~new_n1830_;
  assign new_n1832_ = ~\p_input[248]  & ~\p_input[280] ;
  assign new_n1833_ = \p_input[248]  & \p_input[280] ;
  assign new_n1834_ = ~new_n1832_ & ~new_n1833_;
  assign new_n1835_ = ~new_n1831_ & ~new_n1834_;
  assign new_n1836_ = new_n1831_ & new_n1834_;
  assign new_n1837_ = ~new_n1835_ & ~new_n1836_;
  assign new_n1838_ = ~\p_input[242]  & ~\p_input[274] ;
  assign new_n1839_ = \p_input[242]  & \p_input[274] ;
  assign new_n1840_ = ~new_n1838_ & ~new_n1839_;
  assign new_n1841_ = ~new_n1837_ & ~new_n1840_;
  assign new_n1842_ = new_n1837_ & new_n1840_;
  assign new_n1843_ = ~new_n1841_ & ~new_n1842_;
  assign new_n1844_ = ~\p_input[244]  & ~\p_input[276] ;
  assign new_n1845_ = \p_input[244]  & \p_input[276] ;
  assign new_n1846_ = ~new_n1844_ & ~new_n1845_;
  assign new_n1847_ = ~\p_input[243]  & ~\p_input[275] ;
  assign new_n1848_ = \p_input[243]  & \p_input[275] ;
  assign new_n1849_ = ~new_n1847_ & ~new_n1848_;
  assign new_n1850_ = ~new_n1846_ & ~new_n1849_;
  assign new_n1851_ = new_n1846_ & new_n1849_;
  assign new_n1852_ = ~new_n1850_ & ~new_n1851_;
  assign new_n1853_ = ~\p_input[245]  & ~\p_input[277] ;
  assign new_n1854_ = \p_input[245]  & \p_input[277] ;
  assign new_n1855_ = ~new_n1853_ & ~new_n1854_;
  assign new_n1856_ = ~new_n1852_ & ~new_n1855_;
  assign new_n1857_ = new_n1852_ & new_n1855_;
  assign new_n1858_ = ~new_n1856_ & ~new_n1857_;
  assign new_n1859_ = new_n1843_ & ~new_n1858_;
  assign new_n1860_ = ~new_n1843_ & new_n1858_;
  assign new_n1861_ = ~new_n1859_ & ~new_n1860_;
  assign new_n1862_ = ~new_n1822_ & ~new_n1861_;
  assign new_n1863_ = ~new_n1821_ & ~new_n1862_;
  assign new_n1864_ = new_n1813_ & new_n1863_;
  assign new_n1865_ = ~new_n1813_ & ~new_n1863_;
  assign new_n1866_ = ~new_n1841_ & ~new_n1859_;
  assign new_n1867_ = ~new_n1830_ & ~new_n1836_;
  assign new_n1868_ = ~new_n1866_ & new_n1867_;
  assign new_n1869_ = new_n1866_ & ~new_n1867_;
  assign new_n1870_ = ~new_n1868_ & ~new_n1869_;
  assign new_n1871_ = ~new_n1851_ & ~new_n1857_;
  assign new_n1872_ = new_n1870_ & new_n1871_;
  assign new_n1873_ = ~new_n1870_ & ~new_n1871_;
  assign new_n1874_ = ~new_n1872_ & ~new_n1873_;
  assign new_n1875_ = ~new_n1865_ & new_n1874_;
  assign new_n1876_ = ~new_n1864_ & ~new_n1875_;
  assign new_n1877_ = ~new_n1811_ & ~new_n1876_;
  assign new_n1878_ = new_n1811_ & new_n1876_;
  assign new_n1879_ = ~new_n1877_ & ~new_n1878_;
  assign new_n1880_ = ~new_n1868_ & ~new_n1872_;
  assign new_n1881_ = new_n1879_ & ~new_n1880_;
  assign new_n1882_ = ~new_n1877_ & ~new_n1881_;
  assign new_n1883_ = ~new_n1879_ & new_n1880_;
  assign new_n1884_ = ~new_n1881_ & ~new_n1883_;
  assign new_n1885_ = ~\p_input[225]  & ~\p_input[257] ;
  assign new_n1886_ = \p_input[225]  & \p_input[257] ;
  assign new_n1887_ = ~new_n1885_ & ~new_n1886_;
  assign new_n1888_ = ~new_n1821_ & ~new_n1822_;
  assign new_n1889_ = ~new_n1861_ & new_n1888_;
  assign new_n1890_ = new_n1861_ & ~new_n1888_;
  assign new_n1891_ = ~new_n1889_ & ~new_n1890_;
  assign new_n1892_ = ~new_n1887_ & ~new_n1891_;
  assign new_n1893_ = new_n1887_ & new_n1891_;
  assign new_n1894_ = ~\p_input[232]  & ~\p_input[264] ;
  assign new_n1895_ = \p_input[232]  & \p_input[264] ;
  assign new_n1896_ = ~new_n1894_ & ~new_n1895_;
  assign new_n1897_ = ~\p_input[231]  & ~\p_input[263] ;
  assign new_n1898_ = \p_input[231]  & \p_input[263] ;
  assign new_n1899_ = ~new_n1897_ & ~new_n1898_;
  assign new_n1900_ = ~new_n1896_ & ~new_n1899_;
  assign new_n1901_ = new_n1896_ & new_n1899_;
  assign new_n1902_ = ~new_n1900_ & ~new_n1901_;
  assign new_n1903_ = ~\p_input[233]  & ~\p_input[265] ;
  assign new_n1904_ = \p_input[233]  & \p_input[265] ;
  assign new_n1905_ = ~new_n1903_ & ~new_n1904_;
  assign new_n1906_ = ~new_n1902_ & ~new_n1905_;
  assign new_n1907_ = new_n1902_ & new_n1905_;
  assign new_n1908_ = ~new_n1906_ & ~new_n1907_;
  assign new_n1909_ = ~\p_input[227]  & ~\p_input[259] ;
  assign new_n1910_ = \p_input[227]  & \p_input[259] ;
  assign new_n1911_ = ~new_n1909_ & ~new_n1910_;
  assign new_n1912_ = ~new_n1908_ & ~new_n1911_;
  assign new_n1913_ = new_n1908_ & new_n1911_;
  assign new_n1914_ = ~new_n1912_ & ~new_n1913_;
  assign new_n1915_ = ~\p_input[229]  & ~\p_input[261] ;
  assign new_n1916_ = \p_input[229]  & \p_input[261] ;
  assign new_n1917_ = ~new_n1915_ & ~new_n1916_;
  assign new_n1918_ = ~\p_input[228]  & ~\p_input[260] ;
  assign new_n1919_ = \p_input[228]  & \p_input[260] ;
  assign new_n1920_ = ~new_n1918_ & ~new_n1919_;
  assign new_n1921_ = ~new_n1917_ & ~new_n1920_;
  assign new_n1922_ = new_n1917_ & new_n1920_;
  assign new_n1923_ = ~new_n1921_ & ~new_n1922_;
  assign new_n1924_ = ~\p_input[230]  & ~\p_input[262] ;
  assign new_n1925_ = \p_input[230]  & \p_input[262] ;
  assign new_n1926_ = ~new_n1924_ & ~new_n1925_;
  assign new_n1927_ = ~new_n1923_ & ~new_n1926_;
  assign new_n1928_ = new_n1923_ & new_n1926_;
  assign new_n1929_ = ~new_n1927_ & ~new_n1928_;
  assign new_n1930_ = new_n1914_ & ~new_n1929_;
  assign new_n1931_ = ~new_n1914_ & new_n1929_;
  assign new_n1932_ = ~new_n1930_ & ~new_n1931_;
  assign new_n1933_ = ~\p_input[239]  & ~\p_input[271] ;
  assign new_n1934_ = \p_input[239]  & \p_input[271] ;
  assign new_n1935_ = ~new_n1933_ & ~new_n1934_;
  assign new_n1936_ = ~\p_input[238]  & ~\p_input[270] ;
  assign new_n1937_ = \p_input[238]  & \p_input[270] ;
  assign new_n1938_ = ~new_n1936_ & ~new_n1937_;
  assign new_n1939_ = ~new_n1935_ & ~new_n1938_;
  assign new_n1940_ = new_n1935_ & new_n1938_;
  assign new_n1941_ = ~new_n1939_ & ~new_n1940_;
  assign new_n1942_ = ~\p_input[240]  & ~\p_input[272] ;
  assign new_n1943_ = \p_input[240]  & \p_input[272] ;
  assign new_n1944_ = ~new_n1942_ & ~new_n1943_;
  assign new_n1945_ = ~new_n1941_ & ~new_n1944_;
  assign new_n1946_ = new_n1941_ & new_n1944_;
  assign new_n1947_ = ~new_n1945_ & ~new_n1946_;
  assign new_n1948_ = ~\p_input[234]  & ~\p_input[266] ;
  assign new_n1949_ = \p_input[234]  & \p_input[266] ;
  assign new_n1950_ = ~new_n1948_ & ~new_n1949_;
  assign new_n1951_ = ~new_n1947_ & ~new_n1950_;
  assign new_n1952_ = new_n1947_ & new_n1950_;
  assign new_n1953_ = ~new_n1951_ & ~new_n1952_;
  assign new_n1954_ = ~\p_input[236]  & ~\p_input[268] ;
  assign new_n1955_ = \p_input[236]  & \p_input[268] ;
  assign new_n1956_ = ~new_n1954_ & ~new_n1955_;
  assign new_n1957_ = ~\p_input[235]  & ~\p_input[267] ;
  assign new_n1958_ = \p_input[235]  & \p_input[267] ;
  assign new_n1959_ = ~new_n1957_ & ~new_n1958_;
  assign new_n1960_ = ~new_n1956_ & ~new_n1959_;
  assign new_n1961_ = new_n1956_ & new_n1959_;
  assign new_n1962_ = ~new_n1960_ & ~new_n1961_;
  assign new_n1963_ = ~\p_input[237]  & ~\p_input[269] ;
  assign new_n1964_ = \p_input[237]  & \p_input[269] ;
  assign new_n1965_ = ~new_n1963_ & ~new_n1964_;
  assign new_n1966_ = ~new_n1962_ & ~new_n1965_;
  assign new_n1967_ = new_n1962_ & new_n1965_;
  assign new_n1968_ = ~new_n1966_ & ~new_n1967_;
  assign new_n1969_ = new_n1953_ & ~new_n1968_;
  assign new_n1970_ = ~new_n1953_ & new_n1968_;
  assign new_n1971_ = ~new_n1969_ & ~new_n1970_;
  assign new_n1972_ = ~\p_input[226]  & ~\p_input[258] ;
  assign new_n1973_ = \p_input[226]  & \p_input[258] ;
  assign new_n1974_ = ~new_n1972_ & ~new_n1973_;
  assign new_n1975_ = new_n1971_ & ~new_n1974_;
  assign new_n1976_ = ~new_n1971_ & new_n1974_;
  assign new_n1977_ = ~new_n1975_ & ~new_n1976_;
  assign new_n1978_ = new_n1932_ & new_n1977_;
  assign new_n1979_ = ~new_n1932_ & ~new_n1977_;
  assign new_n1980_ = ~new_n1978_ & ~new_n1979_;
  assign new_n1981_ = ~new_n1893_ & new_n1980_;
  assign new_n1982_ = ~new_n1892_ & ~new_n1981_;
  assign new_n1983_ = ~new_n1864_ & ~new_n1865_;
  assign new_n1984_ = ~new_n1874_ & new_n1983_;
  assign new_n1985_ = new_n1874_ & ~new_n1983_;
  assign new_n1986_ = ~new_n1984_ & ~new_n1985_;
  assign new_n1987_ = new_n1982_ & new_n1986_;
  assign new_n1988_ = ~new_n1982_ & ~new_n1986_;
  assign new_n1989_ = ~new_n1912_ & ~new_n1930_;
  assign new_n1990_ = ~new_n1901_ & ~new_n1907_;
  assign new_n1991_ = ~new_n1989_ & new_n1990_;
  assign new_n1992_ = new_n1989_ & ~new_n1990_;
  assign new_n1993_ = ~new_n1991_ & ~new_n1992_;
  assign new_n1994_ = ~new_n1922_ & ~new_n1928_;
  assign new_n1995_ = new_n1993_ & new_n1994_;
  assign new_n1996_ = ~new_n1993_ & ~new_n1994_;
  assign new_n1997_ = ~new_n1995_ & ~new_n1996_;
  assign new_n1998_ = ~new_n1951_ & ~new_n1969_;
  assign new_n1999_ = ~new_n1940_ & ~new_n1946_;
  assign new_n2000_ = ~new_n1998_ & new_n1999_;
  assign new_n2001_ = new_n1998_ & ~new_n1999_;
  assign new_n2002_ = ~new_n2000_ & ~new_n2001_;
  assign new_n2003_ = ~new_n1961_ & ~new_n1967_;
  assign new_n2004_ = new_n2002_ & new_n2003_;
  assign new_n2005_ = ~new_n2002_ & ~new_n2003_;
  assign new_n2006_ = ~new_n2004_ & ~new_n2005_;
  assign new_n2007_ = ~new_n1975_ & ~new_n1978_;
  assign new_n2008_ = new_n2006_ & ~new_n2007_;
  assign new_n2009_ = ~new_n2006_ & new_n2007_;
  assign new_n2010_ = ~new_n2008_ & ~new_n2009_;
  assign new_n2011_ = new_n1997_ & new_n2010_;
  assign new_n2012_ = ~new_n1997_ & ~new_n2010_;
  assign new_n2013_ = ~new_n2011_ & ~new_n2012_;
  assign new_n2014_ = ~new_n1988_ & ~new_n2013_;
  assign new_n2015_ = ~new_n1987_ & ~new_n2014_;
  assign new_n2016_ = ~new_n1884_ & ~new_n2015_;
  assign new_n2017_ = new_n1884_ & new_n2015_;
  assign new_n2018_ = ~new_n1997_ & ~new_n2008_;
  assign new_n2019_ = ~new_n2009_ & ~new_n2018_;
  assign new_n2020_ = ~new_n2000_ & ~new_n2004_;
  assign new_n2021_ = new_n2019_ & ~new_n2020_;
  assign new_n2022_ = ~new_n2019_ & new_n2020_;
  assign new_n2023_ = ~new_n2021_ & ~new_n2022_;
  assign new_n2024_ = ~new_n1991_ & ~new_n1995_;
  assign new_n2025_ = new_n2023_ & ~new_n2024_;
  assign new_n2026_ = ~new_n2023_ & new_n2024_;
  assign new_n2027_ = ~new_n2025_ & ~new_n2026_;
  assign new_n2028_ = ~new_n2017_ & ~new_n2027_;
  assign new_n2029_ = ~new_n2016_ & ~new_n2028_;
  assign new_n2030_ = ~new_n1882_ & new_n2029_;
  assign new_n2031_ = new_n1882_ & ~new_n2029_;
  assign new_n2032_ = ~new_n2030_ & ~new_n2031_;
  assign new_n2033_ = ~new_n2021_ & ~new_n2025_;
  assign new_n2034_ = new_n2032_ & ~new_n2033_;
  assign new_n2035_ = ~new_n2032_ & new_n2033_;
  assign new_n2036_ = ~new_n2034_ & ~new_n2035_;
  assign new_n2037_ = ~\p_input[224]  & ~\p_input[256] ;
  assign new_n2038_ = \p_input[224]  & \p_input[256] ;
  assign new_n2039_ = ~new_n2037_ & ~new_n2038_;
  assign new_n2040_ = ~new_n1892_ & ~new_n1893_;
  assign new_n2041_ = new_n1980_ & new_n2040_;
  assign new_n2042_ = ~new_n1980_ & ~new_n2040_;
  assign new_n2043_ = ~new_n2041_ & ~new_n2042_;
  assign new_n2044_ = new_n2039_ & ~new_n2043_;
  assign new_n2045_ = ~new_n1987_ & ~new_n1988_;
  assign new_n2046_ = ~new_n2013_ & new_n2045_;
  assign new_n2047_ = new_n2013_ & ~new_n2045_;
  assign new_n2048_ = ~new_n2046_ & ~new_n2047_;
  assign new_n2049_ = new_n2044_ & new_n2048_;
  assign new_n2050_ = ~new_n2016_ & ~new_n2017_;
  assign new_n2051_ = ~new_n2027_ & new_n2050_;
  assign new_n2052_ = new_n2027_ & ~new_n2050_;
  assign new_n2053_ = ~new_n2051_ & ~new_n2052_;
  assign new_n2054_ = new_n2049_ & new_n2053_;
  assign new_n2055_ = ~new_n2036_ & new_n2054_;
  assign new_n2056_ = ~new_n2030_ & ~new_n2034_;
  assign new_n2057_ = new_n2055_ & new_n2056_;
  assign new_n2058_ = ~\p_input[222]  & ~\p_input[286] ;
  assign new_n2059_ = \p_input[222]  & \p_input[286] ;
  assign new_n2060_ = ~new_n2058_ & ~new_n2059_;
  assign new_n2061_ = ~\p_input[221]  & ~\p_input[285] ;
  assign new_n2062_ = \p_input[221]  & \p_input[285] ;
  assign new_n2063_ = ~new_n2061_ & ~new_n2062_;
  assign new_n2064_ = new_n2060_ & new_n2063_;
  assign new_n2065_ = ~new_n2060_ & ~new_n2063_;
  assign new_n2066_ = ~new_n2064_ & ~new_n2065_;
  assign new_n2067_ = ~\p_input[223]  & ~\p_input[287] ;
  assign new_n2068_ = \p_input[223]  & \p_input[287] ;
  assign new_n2069_ = ~new_n2067_ & ~new_n2068_;
  assign new_n2070_ = new_n2066_ & new_n2069_;
  assign new_n2071_ = ~new_n2064_ & ~new_n2070_;
  assign new_n2072_ = ~new_n2066_ & ~new_n2069_;
  assign new_n2073_ = ~new_n2070_ & ~new_n2072_;
  assign new_n2074_ = ~\p_input[217]  & ~\p_input[281] ;
  assign new_n2075_ = \p_input[217]  & \p_input[281] ;
  assign new_n2076_ = ~new_n2074_ & ~new_n2075_;
  assign new_n2077_ = new_n2073_ & new_n2076_;
  assign new_n2078_ = ~new_n2073_ & ~new_n2076_;
  assign new_n2079_ = ~\p_input[219]  & ~\p_input[283] ;
  assign new_n2080_ = \p_input[219]  & \p_input[283] ;
  assign new_n2081_ = ~new_n2079_ & ~new_n2080_;
  assign new_n2082_ = ~\p_input[218]  & ~\p_input[282] ;
  assign new_n2083_ = \p_input[218]  & \p_input[282] ;
  assign new_n2084_ = ~new_n2082_ & ~new_n2083_;
  assign new_n2085_ = ~new_n2081_ & ~new_n2084_;
  assign new_n2086_ = new_n2081_ & new_n2084_;
  assign new_n2087_ = ~new_n2085_ & ~new_n2086_;
  assign new_n2088_ = ~\p_input[220]  & ~\p_input[284] ;
  assign new_n2089_ = \p_input[220]  & \p_input[284] ;
  assign new_n2090_ = ~new_n2088_ & ~new_n2089_;
  assign new_n2091_ = ~new_n2087_ & ~new_n2090_;
  assign new_n2092_ = new_n2087_ & new_n2090_;
  assign new_n2093_ = ~new_n2091_ & ~new_n2092_;
  assign new_n2094_ = ~new_n2078_ & new_n2093_;
  assign new_n2095_ = ~new_n2077_ & ~new_n2094_;
  assign new_n2096_ = new_n2071_ & new_n2095_;
  assign new_n2097_ = ~new_n2071_ & ~new_n2095_;
  assign new_n2098_ = ~new_n2096_ & ~new_n2097_;
  assign new_n2099_ = ~new_n2086_ & ~new_n2092_;
  assign new_n2100_ = new_n2098_ & new_n2099_;
  assign new_n2101_ = ~new_n2096_ & ~new_n2100_;
  assign new_n2102_ = ~new_n2098_ & ~new_n2099_;
  assign new_n2103_ = ~new_n2100_ & ~new_n2102_;
  assign new_n2104_ = ~new_n2077_ & ~new_n2078_;
  assign new_n2105_ = ~new_n2093_ & new_n2104_;
  assign new_n2106_ = new_n2093_ & ~new_n2104_;
  assign new_n2107_ = ~new_n2105_ & ~new_n2106_;
  assign new_n2108_ = ~\p_input[209]  & ~\p_input[273] ;
  assign new_n2109_ = \p_input[209]  & \p_input[273] ;
  assign new_n2110_ = ~new_n2108_ & ~new_n2109_;
  assign new_n2111_ = ~new_n2107_ & new_n2110_;
  assign new_n2112_ = new_n2107_ & ~new_n2110_;
  assign new_n2113_ = ~\p_input[215]  & ~\p_input[279] ;
  assign new_n2114_ = \p_input[215]  & \p_input[279] ;
  assign new_n2115_ = ~new_n2113_ & ~new_n2114_;
  assign new_n2116_ = ~\p_input[214]  & ~\p_input[278] ;
  assign new_n2117_ = \p_input[214]  & \p_input[278] ;
  assign new_n2118_ = ~new_n2116_ & ~new_n2117_;
  assign new_n2119_ = ~new_n2115_ & ~new_n2118_;
  assign new_n2120_ = new_n2115_ & new_n2118_;
  assign new_n2121_ = ~new_n2119_ & ~new_n2120_;
  assign new_n2122_ = ~\p_input[216]  & ~\p_input[280] ;
  assign new_n2123_ = \p_input[216]  & \p_input[280] ;
  assign new_n2124_ = ~new_n2122_ & ~new_n2123_;
  assign new_n2125_ = ~new_n2121_ & ~new_n2124_;
  assign new_n2126_ = new_n2121_ & new_n2124_;
  assign new_n2127_ = ~new_n2125_ & ~new_n2126_;
  assign new_n2128_ = ~\p_input[210]  & ~\p_input[274] ;
  assign new_n2129_ = \p_input[210]  & \p_input[274] ;
  assign new_n2130_ = ~new_n2128_ & ~new_n2129_;
  assign new_n2131_ = ~new_n2127_ & ~new_n2130_;
  assign new_n2132_ = new_n2127_ & new_n2130_;
  assign new_n2133_ = ~new_n2131_ & ~new_n2132_;
  assign new_n2134_ = ~\p_input[212]  & ~\p_input[276] ;
  assign new_n2135_ = \p_input[212]  & \p_input[276] ;
  assign new_n2136_ = ~new_n2134_ & ~new_n2135_;
  assign new_n2137_ = ~\p_input[211]  & ~\p_input[275] ;
  assign new_n2138_ = \p_input[211]  & \p_input[275] ;
  assign new_n2139_ = ~new_n2137_ & ~new_n2138_;
  assign new_n2140_ = ~new_n2136_ & ~new_n2139_;
  assign new_n2141_ = new_n2136_ & new_n2139_;
  assign new_n2142_ = ~new_n2140_ & ~new_n2141_;
  assign new_n2143_ = ~\p_input[213]  & ~\p_input[277] ;
  assign new_n2144_ = \p_input[213]  & \p_input[277] ;
  assign new_n2145_ = ~new_n2143_ & ~new_n2144_;
  assign new_n2146_ = ~new_n2142_ & ~new_n2145_;
  assign new_n2147_ = new_n2142_ & new_n2145_;
  assign new_n2148_ = ~new_n2146_ & ~new_n2147_;
  assign new_n2149_ = new_n2133_ & ~new_n2148_;
  assign new_n2150_ = ~new_n2133_ & new_n2148_;
  assign new_n2151_ = ~new_n2149_ & ~new_n2150_;
  assign new_n2152_ = ~new_n2112_ & ~new_n2151_;
  assign new_n2153_ = ~new_n2111_ & ~new_n2152_;
  assign new_n2154_ = new_n2103_ & new_n2153_;
  assign new_n2155_ = ~new_n2103_ & ~new_n2153_;
  assign new_n2156_ = ~new_n2131_ & ~new_n2149_;
  assign new_n2157_ = ~new_n2120_ & ~new_n2126_;
  assign new_n2158_ = ~new_n2156_ & new_n2157_;
  assign new_n2159_ = new_n2156_ & ~new_n2157_;
  assign new_n2160_ = ~new_n2158_ & ~new_n2159_;
  assign new_n2161_ = ~new_n2141_ & ~new_n2147_;
  assign new_n2162_ = new_n2160_ & new_n2161_;
  assign new_n2163_ = ~new_n2160_ & ~new_n2161_;
  assign new_n2164_ = ~new_n2162_ & ~new_n2163_;
  assign new_n2165_ = ~new_n2155_ & new_n2164_;
  assign new_n2166_ = ~new_n2154_ & ~new_n2165_;
  assign new_n2167_ = ~new_n2101_ & ~new_n2166_;
  assign new_n2168_ = new_n2101_ & new_n2166_;
  assign new_n2169_ = ~new_n2167_ & ~new_n2168_;
  assign new_n2170_ = ~new_n2158_ & ~new_n2162_;
  assign new_n2171_ = new_n2169_ & ~new_n2170_;
  assign new_n2172_ = ~new_n2167_ & ~new_n2171_;
  assign new_n2173_ = ~new_n2169_ & new_n2170_;
  assign new_n2174_ = ~new_n2171_ & ~new_n2173_;
  assign new_n2175_ = ~\p_input[193]  & ~\p_input[257] ;
  assign new_n2176_ = \p_input[193]  & \p_input[257] ;
  assign new_n2177_ = ~new_n2175_ & ~new_n2176_;
  assign new_n2178_ = ~new_n2111_ & ~new_n2112_;
  assign new_n2179_ = ~new_n2151_ & new_n2178_;
  assign new_n2180_ = new_n2151_ & ~new_n2178_;
  assign new_n2181_ = ~new_n2179_ & ~new_n2180_;
  assign new_n2182_ = ~new_n2177_ & ~new_n2181_;
  assign new_n2183_ = new_n2177_ & new_n2181_;
  assign new_n2184_ = ~\p_input[200]  & ~\p_input[264] ;
  assign new_n2185_ = \p_input[200]  & \p_input[264] ;
  assign new_n2186_ = ~new_n2184_ & ~new_n2185_;
  assign new_n2187_ = ~\p_input[199]  & ~\p_input[263] ;
  assign new_n2188_ = \p_input[199]  & \p_input[263] ;
  assign new_n2189_ = ~new_n2187_ & ~new_n2188_;
  assign new_n2190_ = ~new_n2186_ & ~new_n2189_;
  assign new_n2191_ = new_n2186_ & new_n2189_;
  assign new_n2192_ = ~new_n2190_ & ~new_n2191_;
  assign new_n2193_ = ~\p_input[201]  & ~\p_input[265] ;
  assign new_n2194_ = \p_input[201]  & \p_input[265] ;
  assign new_n2195_ = ~new_n2193_ & ~new_n2194_;
  assign new_n2196_ = ~new_n2192_ & ~new_n2195_;
  assign new_n2197_ = new_n2192_ & new_n2195_;
  assign new_n2198_ = ~new_n2196_ & ~new_n2197_;
  assign new_n2199_ = ~\p_input[195]  & ~\p_input[259] ;
  assign new_n2200_ = \p_input[195]  & \p_input[259] ;
  assign new_n2201_ = ~new_n2199_ & ~new_n2200_;
  assign new_n2202_ = ~new_n2198_ & ~new_n2201_;
  assign new_n2203_ = new_n2198_ & new_n2201_;
  assign new_n2204_ = ~new_n2202_ & ~new_n2203_;
  assign new_n2205_ = ~\p_input[197]  & ~\p_input[261] ;
  assign new_n2206_ = \p_input[197]  & \p_input[261] ;
  assign new_n2207_ = ~new_n2205_ & ~new_n2206_;
  assign new_n2208_ = ~\p_input[196]  & ~\p_input[260] ;
  assign new_n2209_ = \p_input[196]  & \p_input[260] ;
  assign new_n2210_ = ~new_n2208_ & ~new_n2209_;
  assign new_n2211_ = ~new_n2207_ & ~new_n2210_;
  assign new_n2212_ = new_n2207_ & new_n2210_;
  assign new_n2213_ = ~new_n2211_ & ~new_n2212_;
  assign new_n2214_ = ~\p_input[198]  & ~\p_input[262] ;
  assign new_n2215_ = \p_input[198]  & \p_input[262] ;
  assign new_n2216_ = ~new_n2214_ & ~new_n2215_;
  assign new_n2217_ = ~new_n2213_ & ~new_n2216_;
  assign new_n2218_ = new_n2213_ & new_n2216_;
  assign new_n2219_ = ~new_n2217_ & ~new_n2218_;
  assign new_n2220_ = new_n2204_ & ~new_n2219_;
  assign new_n2221_ = ~new_n2204_ & new_n2219_;
  assign new_n2222_ = ~new_n2220_ & ~new_n2221_;
  assign new_n2223_ = ~\p_input[207]  & ~\p_input[271] ;
  assign new_n2224_ = \p_input[207]  & \p_input[271] ;
  assign new_n2225_ = ~new_n2223_ & ~new_n2224_;
  assign new_n2226_ = ~\p_input[206]  & ~\p_input[270] ;
  assign new_n2227_ = \p_input[206]  & \p_input[270] ;
  assign new_n2228_ = ~new_n2226_ & ~new_n2227_;
  assign new_n2229_ = ~new_n2225_ & ~new_n2228_;
  assign new_n2230_ = new_n2225_ & new_n2228_;
  assign new_n2231_ = ~new_n2229_ & ~new_n2230_;
  assign new_n2232_ = ~\p_input[208]  & ~\p_input[272] ;
  assign new_n2233_ = \p_input[208]  & \p_input[272] ;
  assign new_n2234_ = ~new_n2232_ & ~new_n2233_;
  assign new_n2235_ = ~new_n2231_ & ~new_n2234_;
  assign new_n2236_ = new_n2231_ & new_n2234_;
  assign new_n2237_ = ~new_n2235_ & ~new_n2236_;
  assign new_n2238_ = ~\p_input[202]  & ~\p_input[266] ;
  assign new_n2239_ = \p_input[202]  & \p_input[266] ;
  assign new_n2240_ = ~new_n2238_ & ~new_n2239_;
  assign new_n2241_ = ~new_n2237_ & ~new_n2240_;
  assign new_n2242_ = new_n2237_ & new_n2240_;
  assign new_n2243_ = ~new_n2241_ & ~new_n2242_;
  assign new_n2244_ = ~\p_input[204]  & ~\p_input[268] ;
  assign new_n2245_ = \p_input[204]  & \p_input[268] ;
  assign new_n2246_ = ~new_n2244_ & ~new_n2245_;
  assign new_n2247_ = ~\p_input[203]  & ~\p_input[267] ;
  assign new_n2248_ = \p_input[203]  & \p_input[267] ;
  assign new_n2249_ = ~new_n2247_ & ~new_n2248_;
  assign new_n2250_ = ~new_n2246_ & ~new_n2249_;
  assign new_n2251_ = new_n2246_ & new_n2249_;
  assign new_n2252_ = ~new_n2250_ & ~new_n2251_;
  assign new_n2253_ = ~\p_input[205]  & ~\p_input[269] ;
  assign new_n2254_ = \p_input[205]  & \p_input[269] ;
  assign new_n2255_ = ~new_n2253_ & ~new_n2254_;
  assign new_n2256_ = ~new_n2252_ & ~new_n2255_;
  assign new_n2257_ = new_n2252_ & new_n2255_;
  assign new_n2258_ = ~new_n2256_ & ~new_n2257_;
  assign new_n2259_ = new_n2243_ & ~new_n2258_;
  assign new_n2260_ = ~new_n2243_ & new_n2258_;
  assign new_n2261_ = ~new_n2259_ & ~new_n2260_;
  assign new_n2262_ = ~\p_input[194]  & ~\p_input[258] ;
  assign new_n2263_ = \p_input[194]  & \p_input[258] ;
  assign new_n2264_ = ~new_n2262_ & ~new_n2263_;
  assign new_n2265_ = new_n2261_ & ~new_n2264_;
  assign new_n2266_ = ~new_n2261_ & new_n2264_;
  assign new_n2267_ = ~new_n2265_ & ~new_n2266_;
  assign new_n2268_ = new_n2222_ & new_n2267_;
  assign new_n2269_ = ~new_n2222_ & ~new_n2267_;
  assign new_n2270_ = ~new_n2268_ & ~new_n2269_;
  assign new_n2271_ = ~new_n2183_ & new_n2270_;
  assign new_n2272_ = ~new_n2182_ & ~new_n2271_;
  assign new_n2273_ = ~new_n2154_ & ~new_n2155_;
  assign new_n2274_ = ~new_n2164_ & new_n2273_;
  assign new_n2275_ = new_n2164_ & ~new_n2273_;
  assign new_n2276_ = ~new_n2274_ & ~new_n2275_;
  assign new_n2277_ = new_n2272_ & new_n2276_;
  assign new_n2278_ = ~new_n2272_ & ~new_n2276_;
  assign new_n2279_ = ~new_n2202_ & ~new_n2220_;
  assign new_n2280_ = ~new_n2191_ & ~new_n2197_;
  assign new_n2281_ = ~new_n2279_ & new_n2280_;
  assign new_n2282_ = new_n2279_ & ~new_n2280_;
  assign new_n2283_ = ~new_n2281_ & ~new_n2282_;
  assign new_n2284_ = ~new_n2212_ & ~new_n2218_;
  assign new_n2285_ = new_n2283_ & new_n2284_;
  assign new_n2286_ = ~new_n2283_ & ~new_n2284_;
  assign new_n2287_ = ~new_n2285_ & ~new_n2286_;
  assign new_n2288_ = ~new_n2241_ & ~new_n2259_;
  assign new_n2289_ = ~new_n2230_ & ~new_n2236_;
  assign new_n2290_ = ~new_n2288_ & new_n2289_;
  assign new_n2291_ = new_n2288_ & ~new_n2289_;
  assign new_n2292_ = ~new_n2290_ & ~new_n2291_;
  assign new_n2293_ = ~new_n2251_ & ~new_n2257_;
  assign new_n2294_ = new_n2292_ & new_n2293_;
  assign new_n2295_ = ~new_n2292_ & ~new_n2293_;
  assign new_n2296_ = ~new_n2294_ & ~new_n2295_;
  assign new_n2297_ = ~new_n2265_ & ~new_n2268_;
  assign new_n2298_ = new_n2296_ & ~new_n2297_;
  assign new_n2299_ = ~new_n2296_ & new_n2297_;
  assign new_n2300_ = ~new_n2298_ & ~new_n2299_;
  assign new_n2301_ = new_n2287_ & new_n2300_;
  assign new_n2302_ = ~new_n2287_ & ~new_n2300_;
  assign new_n2303_ = ~new_n2301_ & ~new_n2302_;
  assign new_n2304_ = ~new_n2278_ & ~new_n2303_;
  assign new_n2305_ = ~new_n2277_ & ~new_n2304_;
  assign new_n2306_ = ~new_n2174_ & ~new_n2305_;
  assign new_n2307_ = new_n2174_ & new_n2305_;
  assign new_n2308_ = ~new_n2287_ & ~new_n2298_;
  assign new_n2309_ = ~new_n2299_ & ~new_n2308_;
  assign new_n2310_ = ~new_n2290_ & ~new_n2294_;
  assign new_n2311_ = new_n2309_ & ~new_n2310_;
  assign new_n2312_ = ~new_n2309_ & new_n2310_;
  assign new_n2313_ = ~new_n2311_ & ~new_n2312_;
  assign new_n2314_ = ~new_n2281_ & ~new_n2285_;
  assign new_n2315_ = new_n2313_ & ~new_n2314_;
  assign new_n2316_ = ~new_n2313_ & new_n2314_;
  assign new_n2317_ = ~new_n2315_ & ~new_n2316_;
  assign new_n2318_ = ~new_n2307_ & ~new_n2317_;
  assign new_n2319_ = ~new_n2306_ & ~new_n2318_;
  assign new_n2320_ = ~new_n2172_ & new_n2319_;
  assign new_n2321_ = new_n2172_ & ~new_n2319_;
  assign new_n2322_ = ~new_n2320_ & ~new_n2321_;
  assign new_n2323_ = ~new_n2311_ & ~new_n2315_;
  assign new_n2324_ = new_n2322_ & ~new_n2323_;
  assign new_n2325_ = ~new_n2322_ & new_n2323_;
  assign new_n2326_ = ~new_n2324_ & ~new_n2325_;
  assign new_n2327_ = ~\p_input[192]  & ~\p_input[256] ;
  assign new_n2328_ = \p_input[192]  & \p_input[256] ;
  assign new_n2329_ = ~new_n2327_ & ~new_n2328_;
  assign new_n2330_ = ~new_n2182_ & ~new_n2183_;
  assign new_n2331_ = new_n2270_ & new_n2330_;
  assign new_n2332_ = ~new_n2270_ & ~new_n2330_;
  assign new_n2333_ = ~new_n2331_ & ~new_n2332_;
  assign new_n2334_ = new_n2329_ & ~new_n2333_;
  assign new_n2335_ = ~new_n2277_ & ~new_n2278_;
  assign new_n2336_ = ~new_n2303_ & new_n2335_;
  assign new_n2337_ = new_n2303_ & ~new_n2335_;
  assign new_n2338_ = ~new_n2336_ & ~new_n2337_;
  assign new_n2339_ = new_n2334_ & new_n2338_;
  assign new_n2340_ = ~new_n2306_ & ~new_n2307_;
  assign new_n2341_ = ~new_n2317_ & new_n2340_;
  assign new_n2342_ = new_n2317_ & ~new_n2340_;
  assign new_n2343_ = ~new_n2341_ & ~new_n2342_;
  assign new_n2344_ = new_n2339_ & new_n2343_;
  assign new_n2345_ = ~new_n2326_ & new_n2344_;
  assign new_n2346_ = ~new_n2320_ & ~new_n2324_;
  assign new_n2347_ = new_n2345_ & new_n2346_;
  assign new_n2348_ = ~new_n2057_ & ~new_n2347_;
  assign new_n2349_ = new_n1767_ & ~new_n2348_;
  assign new_n2350_ = new_n2057_ & new_n2347_;
  assign new_n2351_ = ~new_n1767_ & new_n2350_;
  assign new_n2352_ = ~new_n2349_ & ~new_n2351_;
  assign new_n2353_ = ~\p_input[136]  & ~\p_input[264] ;
  assign new_n2354_ = \p_input[136]  & \p_input[264] ;
  assign new_n2355_ = ~new_n2353_ & ~new_n2354_;
  assign new_n2356_ = ~\p_input[135]  & ~\p_input[263] ;
  assign new_n2357_ = \p_input[135]  & \p_input[263] ;
  assign new_n2358_ = ~new_n2356_ & ~new_n2357_;
  assign new_n2359_ = ~new_n2355_ & ~new_n2358_;
  assign new_n2360_ = new_n2355_ & new_n2358_;
  assign new_n2361_ = ~new_n2359_ & ~new_n2360_;
  assign new_n2362_ = ~\p_input[137]  & ~\p_input[265] ;
  assign new_n2363_ = \p_input[137]  & \p_input[265] ;
  assign new_n2364_ = ~new_n2362_ & ~new_n2363_;
  assign new_n2365_ = ~new_n2361_ & ~new_n2364_;
  assign new_n2366_ = new_n2361_ & new_n2364_;
  assign new_n2367_ = ~new_n2365_ & ~new_n2366_;
  assign new_n2368_ = ~\p_input[131]  & ~\p_input[259] ;
  assign new_n2369_ = \p_input[131]  & \p_input[259] ;
  assign new_n2370_ = ~new_n2368_ & ~new_n2369_;
  assign new_n2371_ = ~new_n2367_ & ~new_n2370_;
  assign new_n2372_ = new_n2367_ & new_n2370_;
  assign new_n2373_ = ~new_n2371_ & ~new_n2372_;
  assign new_n2374_ = ~\p_input[133]  & ~\p_input[261] ;
  assign new_n2375_ = \p_input[133]  & \p_input[261] ;
  assign new_n2376_ = ~new_n2374_ & ~new_n2375_;
  assign new_n2377_ = ~\p_input[132]  & ~\p_input[260] ;
  assign new_n2378_ = \p_input[132]  & \p_input[260] ;
  assign new_n2379_ = ~new_n2377_ & ~new_n2378_;
  assign new_n2380_ = ~new_n2376_ & ~new_n2379_;
  assign new_n2381_ = new_n2376_ & new_n2379_;
  assign new_n2382_ = ~new_n2380_ & ~new_n2381_;
  assign new_n2383_ = ~\p_input[134]  & ~\p_input[262] ;
  assign new_n2384_ = \p_input[134]  & \p_input[262] ;
  assign new_n2385_ = ~new_n2383_ & ~new_n2384_;
  assign new_n2386_ = ~new_n2382_ & ~new_n2385_;
  assign new_n2387_ = new_n2382_ & new_n2385_;
  assign new_n2388_ = ~new_n2386_ & ~new_n2387_;
  assign new_n2389_ = new_n2373_ & ~new_n2388_;
  assign new_n2390_ = ~new_n2371_ & ~new_n2389_;
  assign new_n2391_ = ~new_n2360_ & ~new_n2366_;
  assign new_n2392_ = ~new_n2390_ & new_n2391_;
  assign new_n2393_ = new_n2390_ & ~new_n2391_;
  assign new_n2394_ = ~new_n2392_ & ~new_n2393_;
  assign new_n2395_ = ~new_n2381_ & ~new_n2387_;
  assign new_n2396_ = new_n2394_ & new_n2395_;
  assign new_n2397_ = ~new_n2394_ & ~new_n2395_;
  assign new_n2398_ = ~new_n2396_ & ~new_n2397_;
  assign new_n2399_ = ~\p_input[143]  & ~\p_input[271] ;
  assign new_n2400_ = \p_input[143]  & \p_input[271] ;
  assign new_n2401_ = ~new_n2399_ & ~new_n2400_;
  assign new_n2402_ = ~\p_input[142]  & ~\p_input[270] ;
  assign new_n2403_ = \p_input[142]  & \p_input[270] ;
  assign new_n2404_ = ~new_n2402_ & ~new_n2403_;
  assign new_n2405_ = ~new_n2401_ & ~new_n2404_;
  assign new_n2406_ = new_n2401_ & new_n2404_;
  assign new_n2407_ = ~new_n2405_ & ~new_n2406_;
  assign new_n2408_ = ~\p_input[144]  & ~\p_input[272] ;
  assign new_n2409_ = \p_input[144]  & \p_input[272] ;
  assign new_n2410_ = ~new_n2408_ & ~new_n2409_;
  assign new_n2411_ = ~new_n2407_ & ~new_n2410_;
  assign new_n2412_ = new_n2407_ & new_n2410_;
  assign new_n2413_ = ~new_n2411_ & ~new_n2412_;
  assign new_n2414_ = ~\p_input[138]  & ~\p_input[266] ;
  assign new_n2415_ = \p_input[138]  & \p_input[266] ;
  assign new_n2416_ = ~new_n2414_ & ~new_n2415_;
  assign new_n2417_ = ~new_n2413_ & ~new_n2416_;
  assign new_n2418_ = new_n2413_ & new_n2416_;
  assign new_n2419_ = ~new_n2417_ & ~new_n2418_;
  assign new_n2420_ = ~\p_input[140]  & ~\p_input[268] ;
  assign new_n2421_ = \p_input[140]  & \p_input[268] ;
  assign new_n2422_ = ~new_n2420_ & ~new_n2421_;
  assign new_n2423_ = ~\p_input[139]  & ~\p_input[267] ;
  assign new_n2424_ = \p_input[139]  & \p_input[267] ;
  assign new_n2425_ = ~new_n2423_ & ~new_n2424_;
  assign new_n2426_ = ~new_n2422_ & ~new_n2425_;
  assign new_n2427_ = new_n2422_ & new_n2425_;
  assign new_n2428_ = ~new_n2426_ & ~new_n2427_;
  assign new_n2429_ = ~\p_input[141]  & ~\p_input[269] ;
  assign new_n2430_ = \p_input[141]  & \p_input[269] ;
  assign new_n2431_ = ~new_n2429_ & ~new_n2430_;
  assign new_n2432_ = ~new_n2428_ & ~new_n2431_;
  assign new_n2433_ = new_n2428_ & new_n2431_;
  assign new_n2434_ = ~new_n2432_ & ~new_n2433_;
  assign new_n2435_ = new_n2419_ & ~new_n2434_;
  assign new_n2436_ = ~new_n2417_ & ~new_n2435_;
  assign new_n2437_ = ~new_n2406_ & ~new_n2412_;
  assign new_n2438_ = ~new_n2436_ & new_n2437_;
  assign new_n2439_ = new_n2436_ & ~new_n2437_;
  assign new_n2440_ = ~new_n2438_ & ~new_n2439_;
  assign new_n2441_ = ~new_n2427_ & ~new_n2433_;
  assign new_n2442_ = new_n2440_ & new_n2441_;
  assign new_n2443_ = ~new_n2440_ & ~new_n2441_;
  assign new_n2444_ = ~new_n2442_ & ~new_n2443_;
  assign new_n2445_ = ~new_n2419_ & new_n2434_;
  assign new_n2446_ = ~new_n2435_ & ~new_n2445_;
  assign new_n2447_ = ~\p_input[130]  & ~\p_input[258] ;
  assign new_n2448_ = \p_input[130]  & \p_input[258] ;
  assign new_n2449_ = ~new_n2447_ & ~new_n2448_;
  assign new_n2450_ = new_n2446_ & ~new_n2449_;
  assign new_n2451_ = ~new_n2373_ & new_n2388_;
  assign new_n2452_ = ~new_n2389_ & ~new_n2451_;
  assign new_n2453_ = ~new_n2446_ & new_n2449_;
  assign new_n2454_ = ~new_n2450_ & ~new_n2453_;
  assign new_n2455_ = new_n2452_ & new_n2454_;
  assign new_n2456_ = ~new_n2450_ & ~new_n2455_;
  assign new_n2457_ = new_n2444_ & ~new_n2456_;
  assign new_n2458_ = ~new_n2444_ & new_n2456_;
  assign new_n2459_ = ~new_n2457_ & ~new_n2458_;
  assign new_n2460_ = new_n2398_ & new_n2459_;
  assign new_n2461_ = ~new_n2398_ & ~new_n2459_;
  assign new_n2462_ = ~new_n2460_ & ~new_n2461_;
  assign new_n2463_ = ~\p_input[151]  & ~\p_input[279] ;
  assign new_n2464_ = \p_input[151]  & \p_input[279] ;
  assign new_n2465_ = ~new_n2463_ & ~new_n2464_;
  assign new_n2466_ = ~\p_input[150]  & ~\p_input[278] ;
  assign new_n2467_ = \p_input[150]  & \p_input[278] ;
  assign new_n2468_ = ~new_n2466_ & ~new_n2467_;
  assign new_n2469_ = ~new_n2465_ & ~new_n2468_;
  assign new_n2470_ = new_n2465_ & new_n2468_;
  assign new_n2471_ = ~new_n2469_ & ~new_n2470_;
  assign new_n2472_ = ~\p_input[152]  & ~\p_input[280] ;
  assign new_n2473_ = \p_input[152]  & \p_input[280] ;
  assign new_n2474_ = ~new_n2472_ & ~new_n2473_;
  assign new_n2475_ = ~new_n2471_ & ~new_n2474_;
  assign new_n2476_ = new_n2471_ & new_n2474_;
  assign new_n2477_ = ~new_n2475_ & ~new_n2476_;
  assign new_n2478_ = ~\p_input[146]  & ~\p_input[274] ;
  assign new_n2479_ = \p_input[146]  & \p_input[274] ;
  assign new_n2480_ = ~new_n2478_ & ~new_n2479_;
  assign new_n2481_ = ~new_n2477_ & ~new_n2480_;
  assign new_n2482_ = new_n2477_ & new_n2480_;
  assign new_n2483_ = ~new_n2481_ & ~new_n2482_;
  assign new_n2484_ = ~\p_input[148]  & ~\p_input[276] ;
  assign new_n2485_ = \p_input[148]  & \p_input[276] ;
  assign new_n2486_ = ~new_n2484_ & ~new_n2485_;
  assign new_n2487_ = ~\p_input[147]  & ~\p_input[275] ;
  assign new_n2488_ = \p_input[147]  & \p_input[275] ;
  assign new_n2489_ = ~new_n2487_ & ~new_n2488_;
  assign new_n2490_ = ~new_n2486_ & ~new_n2489_;
  assign new_n2491_ = new_n2486_ & new_n2489_;
  assign new_n2492_ = ~new_n2490_ & ~new_n2491_;
  assign new_n2493_ = ~\p_input[149]  & ~\p_input[277] ;
  assign new_n2494_ = \p_input[149]  & \p_input[277] ;
  assign new_n2495_ = ~new_n2493_ & ~new_n2494_;
  assign new_n2496_ = ~new_n2492_ & ~new_n2495_;
  assign new_n2497_ = new_n2492_ & new_n2495_;
  assign new_n2498_ = ~new_n2496_ & ~new_n2497_;
  assign new_n2499_ = new_n2483_ & ~new_n2498_;
  assign new_n2500_ = ~new_n2481_ & ~new_n2499_;
  assign new_n2501_ = ~new_n2470_ & ~new_n2476_;
  assign new_n2502_ = ~new_n2500_ & new_n2501_;
  assign new_n2503_ = new_n2500_ & ~new_n2501_;
  assign new_n2504_ = ~new_n2502_ & ~new_n2503_;
  assign new_n2505_ = ~new_n2491_ & ~new_n2497_;
  assign new_n2506_ = new_n2504_ & new_n2505_;
  assign new_n2507_ = ~new_n2504_ & ~new_n2505_;
  assign new_n2508_ = ~new_n2506_ & ~new_n2507_;
  assign new_n2509_ = ~\p_input[158]  & ~\p_input[286] ;
  assign new_n2510_ = \p_input[158]  & \p_input[286] ;
  assign new_n2511_ = ~new_n2509_ & ~new_n2510_;
  assign new_n2512_ = ~\p_input[157]  & ~\p_input[285] ;
  assign new_n2513_ = \p_input[157]  & \p_input[285] ;
  assign new_n2514_ = ~new_n2512_ & ~new_n2513_;
  assign new_n2515_ = new_n2511_ & new_n2514_;
  assign new_n2516_ = ~new_n2511_ & ~new_n2514_;
  assign new_n2517_ = ~new_n2515_ & ~new_n2516_;
  assign new_n2518_ = ~\p_input[159]  & ~\p_input[287] ;
  assign new_n2519_ = \p_input[159]  & \p_input[287] ;
  assign new_n2520_ = ~new_n2518_ & ~new_n2519_;
  assign new_n2521_ = ~new_n2517_ & ~new_n2520_;
  assign new_n2522_ = new_n2517_ & new_n2520_;
  assign new_n2523_ = ~new_n2521_ & ~new_n2522_;
  assign new_n2524_ = ~\p_input[153]  & ~\p_input[281] ;
  assign new_n2525_ = \p_input[153]  & \p_input[281] ;
  assign new_n2526_ = ~new_n2524_ & ~new_n2525_;
  assign new_n2527_ = ~new_n2523_ & ~new_n2526_;
  assign new_n2528_ = new_n2523_ & new_n2526_;
  assign new_n2529_ = ~new_n2527_ & ~new_n2528_;
  assign new_n2530_ = ~\p_input[155]  & ~\p_input[283] ;
  assign new_n2531_ = \p_input[155]  & \p_input[283] ;
  assign new_n2532_ = ~new_n2530_ & ~new_n2531_;
  assign new_n2533_ = ~\p_input[154]  & ~\p_input[282] ;
  assign new_n2534_ = \p_input[154]  & \p_input[282] ;
  assign new_n2535_ = ~new_n2533_ & ~new_n2534_;
  assign new_n2536_ = ~new_n2532_ & ~new_n2535_;
  assign new_n2537_ = new_n2532_ & new_n2535_;
  assign new_n2538_ = ~new_n2536_ & ~new_n2537_;
  assign new_n2539_ = ~\p_input[156]  & ~\p_input[284] ;
  assign new_n2540_ = \p_input[156]  & \p_input[284] ;
  assign new_n2541_ = ~new_n2539_ & ~new_n2540_;
  assign new_n2542_ = ~new_n2538_ & ~new_n2541_;
  assign new_n2543_ = new_n2538_ & new_n2541_;
  assign new_n2544_ = ~new_n2542_ & ~new_n2543_;
  assign new_n2545_ = new_n2529_ & ~new_n2544_;
  assign new_n2546_ = ~new_n2527_ & ~new_n2545_;
  assign new_n2547_ = ~new_n2515_ & ~new_n2522_;
  assign new_n2548_ = ~new_n2546_ & new_n2547_;
  assign new_n2549_ = new_n2546_ & ~new_n2547_;
  assign new_n2550_ = ~new_n2548_ & ~new_n2549_;
  assign new_n2551_ = ~new_n2537_ & ~new_n2543_;
  assign new_n2552_ = new_n2550_ & new_n2551_;
  assign new_n2553_ = ~new_n2550_ & ~new_n2551_;
  assign new_n2554_ = ~new_n2552_ & ~new_n2553_;
  assign new_n2555_ = ~new_n2529_ & new_n2544_;
  assign new_n2556_ = ~new_n2545_ & ~new_n2555_;
  assign new_n2557_ = ~\p_input[145]  & ~\p_input[273] ;
  assign new_n2558_ = \p_input[145]  & \p_input[273] ;
  assign new_n2559_ = ~new_n2557_ & ~new_n2558_;
  assign new_n2560_ = new_n2556_ & ~new_n2559_;
  assign new_n2561_ = ~new_n2483_ & new_n2498_;
  assign new_n2562_ = ~new_n2499_ & ~new_n2561_;
  assign new_n2563_ = ~new_n2556_ & new_n2559_;
  assign new_n2564_ = ~new_n2560_ & ~new_n2563_;
  assign new_n2565_ = new_n2562_ & new_n2564_;
  assign new_n2566_ = ~new_n2560_ & ~new_n2565_;
  assign new_n2567_ = new_n2554_ & ~new_n2566_;
  assign new_n2568_ = ~new_n2554_ & new_n2566_;
  assign new_n2569_ = ~new_n2567_ & ~new_n2568_;
  assign new_n2570_ = new_n2508_ & new_n2569_;
  assign new_n2571_ = ~new_n2508_ & ~new_n2569_;
  assign new_n2572_ = ~new_n2570_ & ~new_n2571_;
  assign new_n2573_ = ~new_n2562_ & ~new_n2564_;
  assign new_n2574_ = ~new_n2565_ & ~new_n2573_;
  assign new_n2575_ = ~\p_input[129]  & ~\p_input[257] ;
  assign new_n2576_ = \p_input[129]  & \p_input[257] ;
  assign new_n2577_ = ~new_n2575_ & ~new_n2576_;
  assign new_n2578_ = new_n2574_ & ~new_n2577_;
  assign new_n2579_ = ~new_n2452_ & ~new_n2454_;
  assign new_n2580_ = ~new_n2455_ & ~new_n2579_;
  assign new_n2581_ = ~new_n2574_ & new_n2577_;
  assign new_n2582_ = ~new_n2578_ & ~new_n2581_;
  assign new_n2583_ = new_n2580_ & new_n2582_;
  assign new_n2584_ = ~new_n2578_ & ~new_n2583_;
  assign new_n2585_ = new_n2572_ & ~new_n2584_;
  assign new_n2586_ = ~new_n2572_ & new_n2584_;
  assign new_n2587_ = ~new_n2585_ & ~new_n2586_;
  assign new_n2588_ = new_n2462_ & new_n2587_;
  assign new_n2589_ = ~new_n2462_ & ~new_n2587_;
  assign new_n2590_ = ~new_n2588_ & ~new_n2589_;
  assign new_n2591_ = ~new_n2580_ & ~new_n2582_;
  assign new_n2592_ = ~new_n2583_ & ~new_n2591_;
  assign new_n2593_ = ~\p_input[128]  & ~\p_input[256] ;
  assign new_n2594_ = \p_input[128]  & \p_input[256] ;
  assign new_n2595_ = ~new_n2593_ & ~new_n2594_;
  assign new_n2596_ = ~new_n2592_ & new_n2595_;
  assign new_n2597_ = ~new_n2590_ & new_n2596_;
  assign new_n2598_ = ~new_n2438_ & ~new_n2442_;
  assign new_n2599_ = ~new_n2457_ & ~new_n2460_;
  assign new_n2600_ = ~new_n2598_ & ~new_n2599_;
  assign new_n2601_ = new_n2598_ & new_n2599_;
  assign new_n2602_ = ~new_n2600_ & ~new_n2601_;
  assign new_n2603_ = ~new_n2392_ & ~new_n2396_;
  assign new_n2604_ = new_n2602_ & ~new_n2603_;
  assign new_n2605_ = ~new_n2602_ & new_n2603_;
  assign new_n2606_ = ~new_n2604_ & ~new_n2605_;
  assign new_n2607_ = ~new_n2548_ & ~new_n2552_;
  assign new_n2608_ = ~new_n2567_ & ~new_n2570_;
  assign new_n2609_ = ~new_n2607_ & ~new_n2608_;
  assign new_n2610_ = new_n2607_ & new_n2608_;
  assign new_n2611_ = ~new_n2609_ & ~new_n2610_;
  assign new_n2612_ = ~new_n2502_ & ~new_n2506_;
  assign new_n2613_ = new_n2611_ & ~new_n2612_;
  assign new_n2614_ = ~new_n2611_ & new_n2612_;
  assign new_n2615_ = ~new_n2613_ & ~new_n2614_;
  assign new_n2616_ = ~new_n2585_ & ~new_n2588_;
  assign new_n2617_ = new_n2615_ & ~new_n2616_;
  assign new_n2618_ = ~new_n2615_ & new_n2616_;
  assign new_n2619_ = ~new_n2617_ & ~new_n2618_;
  assign new_n2620_ = new_n2606_ & new_n2619_;
  assign new_n2621_ = ~new_n2606_ & ~new_n2619_;
  assign new_n2622_ = ~new_n2620_ & ~new_n2621_;
  assign new_n2623_ = new_n2597_ & ~new_n2622_;
  assign new_n2624_ = ~new_n2609_ & ~new_n2613_;
  assign new_n2625_ = ~new_n2617_ & ~new_n2620_;
  assign new_n2626_ = ~new_n2624_ & ~new_n2625_;
  assign new_n2627_ = new_n2624_ & new_n2625_;
  assign new_n2628_ = ~new_n2626_ & ~new_n2627_;
  assign new_n2629_ = ~new_n2600_ & ~new_n2604_;
  assign new_n2630_ = new_n2628_ & ~new_n2629_;
  assign new_n2631_ = ~new_n2628_ & new_n2629_;
  assign new_n2632_ = ~new_n2630_ & ~new_n2631_;
  assign new_n2633_ = new_n2623_ & ~new_n2632_;
  assign new_n2634_ = ~new_n2626_ & ~new_n2630_;
  assign new_n2635_ = new_n2633_ & new_n2634_;
  assign new_n2636_ = ~new_n2352_ & new_n2635_;
  assign new_n2637_ = new_n1767_ & new_n2350_;
  assign new_n2638_ = ~new_n2635_ & new_n2637_;
  assign new_n2639_ = ~new_n2636_ & ~new_n2638_;
  assign new_n2640_ = new_n1484_ & ~new_n2639_;
  assign new_n2641_ = new_n2635_ & new_n2637_;
  assign new_n2642_ = ~new_n2640_ & ~new_n2641_;
  assign new_n2643_ = new_n1201_ & ~new_n2642_;
  assign new_n2644_ = new_n2640_ & new_n2641_;
  assign new_n2645_ = ~new_n1201_ & new_n2644_;
  assign new_n2646_ = ~new_n2643_ & ~new_n2645_;
  assign new_n2647_ = new_n918_ & ~new_n2646_;
  assign new_n2648_ = new_n1201_ & new_n2644_;
  assign new_n2649_ = ~new_n918_ & new_n2648_;
  assign new_n2650_ = ~new_n2647_ & ~new_n2649_;
  assign new_n2651_ = new_n635_ & ~new_n2650_;
  assign new_n2652_ = new_n918_ & new_n2648_;
  assign new_n2653_ = ~new_n2651_ & new_n2652_;
  assign new_n2654_ = new_n2326_ & ~new_n2344_;
  assign new_n2655_ = ~new_n2345_ & ~new_n2654_;
  assign new_n2656_ = new_n2036_ & ~new_n2054_;
  assign new_n2657_ = ~new_n2055_ & ~new_n2656_;
  assign new_n2658_ = new_n2655_ & ~new_n2657_;
  assign new_n2659_ = new_n2057_ & ~new_n2347_;
  assign new_n2660_ = ~new_n2055_ & ~new_n2056_;
  assign new_n2661_ = ~new_n2057_ & ~new_n2660_;
  assign new_n2662_ = ~new_n2345_ & ~new_n2346_;
  assign new_n2663_ = ~new_n2347_ & ~new_n2662_;
  assign new_n2664_ = new_n2661_ & ~new_n2663_;
  assign new_n2665_ = ~new_n2655_ & new_n2657_;
  assign new_n2666_ = ~new_n2049_ & ~new_n2053_;
  assign new_n2667_ = ~new_n2054_ & ~new_n2666_;
  assign new_n2668_ = ~new_n2339_ & ~new_n2343_;
  assign new_n2669_ = ~new_n2344_ & ~new_n2668_;
  assign new_n2670_ = ~new_n2667_ & new_n2669_;
  assign new_n2671_ = new_n2667_ & ~new_n2669_;
  assign new_n2672_ = ~new_n2334_ & ~new_n2338_;
  assign new_n2673_ = ~new_n2339_ & ~new_n2672_;
  assign new_n2674_ = ~new_n2044_ & ~new_n2048_;
  assign new_n2675_ = ~new_n2049_ & ~new_n2674_;
  assign new_n2676_ = new_n2673_ & ~new_n2675_;
  assign new_n2677_ = ~new_n2329_ & new_n2333_;
  assign new_n2678_ = ~new_n2334_ & ~new_n2677_;
  assign new_n2679_ = ~new_n2338_ & new_n2675_;
  assign new_n2680_ = ~new_n2039_ & new_n2043_;
  assign new_n2681_ = ~new_n2044_ & ~new_n2680_;
  assign new_n2682_ = new_n2678_ & ~new_n2681_;
  assign new_n2683_ = ~new_n2679_ & new_n2682_;
  assign new_n2684_ = ~new_n2676_ & ~new_n2683_;
  assign new_n2685_ = ~new_n2671_ & ~new_n2684_;
  assign new_n2686_ = ~new_n2670_ & ~new_n2685_;
  assign new_n2687_ = ~new_n2658_ & new_n2686_;
  assign new_n2688_ = ~new_n2664_ & ~new_n2665_;
  assign new_n2689_ = ~new_n2687_ & new_n2688_;
  assign new_n2690_ = ~new_n2661_ & new_n2663_;
  assign new_n2691_ = ~new_n2057_ & new_n2347_;
  assign new_n2692_ = ~new_n2690_ & ~new_n2691_;
  assign new_n2693_ = ~new_n2689_ & new_n2692_;
  assign new_n2694_ = ~new_n2659_ & ~new_n2693_;
  assign new_n2695_ = new_n2658_ & ~new_n2694_;
  assign new_n2696_ = ~new_n2658_ & ~new_n2665_;
  assign new_n2697_ = ~new_n2694_ & ~new_n2696_;
  assign new_n2698_ = new_n2657_ & ~new_n2697_;
  assign new_n2699_ = ~new_n2695_ & ~new_n2698_;
  assign new_n2700_ = ~new_n1755_ & new_n1764_;
  assign new_n2701_ = ~new_n1765_ & ~new_n2700_;
  assign new_n2702_ = new_n1747_ & ~new_n1753_;
  assign new_n2703_ = ~new_n1754_ & ~new_n2702_;
  assign new_n2704_ = ~new_n2675_ & ~new_n2694_;
  assign new_n2705_ = ~new_n2673_ & new_n2694_;
  assign new_n2706_ = ~new_n2704_ & ~new_n2705_;
  assign new_n2707_ = new_n2703_ & ~new_n2706_;
  assign new_n2708_ = new_n1749_ & ~new_n1752_;
  assign new_n2709_ = ~new_n1753_ & ~new_n2708_;
  assign new_n2710_ = ~new_n2681_ & ~new_n2694_;
  assign new_n2711_ = ~new_n2678_ & new_n2694_;
  assign new_n2712_ = ~new_n2710_ & ~new_n2711_;
  assign new_n2713_ = new_n2709_ & ~new_n2712_;
  assign new_n2714_ = ~new_n2707_ & ~new_n2713_;
  assign new_n2715_ = new_n1747_ & new_n2706_;
  assign new_n2716_ = new_n1745_ & ~new_n1754_;
  assign new_n2717_ = ~new_n1755_ & ~new_n2716_;
  assign new_n2718_ = ~new_n2667_ & ~new_n2694_;
  assign new_n2719_ = ~new_n2669_ & new_n2694_;
  assign new_n2720_ = ~new_n2718_ & ~new_n2719_;
  assign new_n2721_ = ~new_n2717_ & new_n2720_;
  assign new_n2722_ = ~new_n2715_ & ~new_n2721_;
  assign new_n2723_ = ~new_n2714_ & new_n2722_;
  assign new_n2724_ = ~new_n2655_ & ~new_n2697_;
  assign new_n2725_ = ~new_n2695_ & ~new_n2724_;
  assign new_n2726_ = new_n2701_ & ~new_n2725_;
  assign new_n2727_ = new_n2717_ & ~new_n2720_;
  assign new_n2728_ = ~new_n2726_ & ~new_n2727_;
  assign new_n2729_ = ~new_n2723_ & new_n2728_;
  assign new_n2730_ = ~new_n1765_ & ~new_n1766_;
  assign new_n2731_ = ~new_n1767_ & ~new_n2730_;
  assign new_n2732_ = ~new_n2664_ & ~new_n2690_;
  assign new_n2733_ = ~new_n2694_ & ~new_n2732_;
  assign new_n2734_ = ~new_n2663_ & ~new_n2733_;
  assign new_n2735_ = new_n2659_ & ~new_n2662_;
  assign new_n2736_ = ~new_n2734_ & ~new_n2735_;
  assign new_n2737_ = ~new_n2731_ & new_n2736_;
  assign new_n2738_ = ~new_n2701_ & new_n2725_;
  assign new_n2739_ = ~new_n1767_ & ~new_n2348_;
  assign new_n2740_ = ~new_n2737_ & ~new_n2739_;
  assign new_n2741_ = ~new_n2738_ & new_n2740_;
  assign new_n2742_ = ~new_n2729_ & new_n2741_;
  assign new_n2743_ = ~new_n1767_ & new_n2736_;
  assign new_n2744_ = new_n2348_ & ~new_n2730_;
  assign new_n2745_ = ~new_n2743_ & new_n2744_;
  assign new_n2746_ = ~new_n2742_ & ~new_n2745_;
  assign new_n2747_ = new_n2701_ & new_n2746_;
  assign new_n2748_ = new_n2725_ & ~new_n2746_;
  assign new_n2749_ = ~new_n2747_ & ~new_n2748_;
  assign new_n2750_ = new_n2699_ & ~new_n2749_;
  assign new_n2751_ = new_n2349_ & ~new_n2350_;
  assign new_n2752_ = new_n2706_ & ~new_n2746_;
  assign new_n2753_ = new_n2703_ & new_n2746_;
  assign new_n2754_ = ~new_n2752_ & ~new_n2753_;
  assign new_n2755_ = new_n2673_ & ~new_n2694_;
  assign new_n2756_ = new_n2675_ & new_n2694_;
  assign new_n2757_ = ~new_n2755_ & ~new_n2756_;
  assign new_n2758_ = new_n2754_ & ~new_n2757_;
  assign new_n2759_ = ~new_n2709_ & new_n2746_;
  assign new_n2760_ = ~new_n2712_ & ~new_n2746_;
  assign new_n2761_ = ~new_n2759_ & ~new_n2760_;
  assign new_n2762_ = new_n2678_ & ~new_n2694_;
  assign new_n2763_ = new_n2681_ & new_n2694_;
  assign new_n2764_ = ~new_n2762_ & ~new_n2763_;
  assign new_n2765_ = new_n2761_ & new_n2764_;
  assign new_n2766_ = ~new_n2758_ & new_n2765_;
  assign new_n2767_ = ~new_n2754_ & new_n2757_;
  assign new_n2768_ = new_n2669_ & ~new_n2694_;
  assign new_n2769_ = new_n2667_ & new_n2694_;
  assign new_n2770_ = ~new_n2768_ & ~new_n2769_;
  assign new_n2771_ = new_n2717_ & new_n2746_;
  assign new_n2772_ = new_n2720_ & ~new_n2746_;
  assign new_n2773_ = ~new_n2771_ & ~new_n2772_;
  assign new_n2774_ = new_n2770_ & ~new_n2773_;
  assign new_n2775_ = ~new_n2767_ & ~new_n2774_;
  assign new_n2776_ = ~new_n2766_ & new_n2775_;
  assign new_n2777_ = ~new_n2699_ & new_n2749_;
  assign new_n2778_ = ~new_n2770_ & new_n2773_;
  assign new_n2779_ = ~new_n2777_ & ~new_n2778_;
  assign new_n2780_ = ~new_n2776_ & new_n2779_;
  assign new_n2781_ = new_n2661_ & ~new_n2733_;
  assign new_n2782_ = ~new_n2735_ & ~new_n2781_;
  assign new_n2783_ = new_n2731_ & new_n2746_;
  assign new_n2784_ = new_n2736_ & ~new_n2746_;
  assign new_n2785_ = ~new_n2783_ & ~new_n2784_;
  assign new_n2786_ = new_n2782_ & ~new_n2785_;
  assign new_n2787_ = ~new_n2750_ & ~new_n2786_;
  assign new_n2788_ = ~new_n2780_ & new_n2787_;
  assign new_n2789_ = ~new_n2782_ & new_n2785_;
  assign new_n2790_ = ~new_n2351_ & ~new_n2789_;
  assign new_n2791_ = ~new_n2788_ & new_n2790_;
  assign new_n2792_ = ~new_n2751_ & ~new_n2791_;
  assign new_n2793_ = new_n2750_ & new_n2792_;
  assign new_n2794_ = ~new_n2750_ & ~new_n2777_;
  assign new_n2795_ = new_n2792_ & ~new_n2794_;
  assign new_n2796_ = ~new_n2699_ & ~new_n2795_;
  assign new_n2797_ = ~new_n2793_ & ~new_n2796_;
  assign new_n2798_ = ~new_n2623_ & new_n2632_;
  assign new_n2799_ = ~new_n2633_ & ~new_n2798_;
  assign new_n2800_ = new_n2592_ & ~new_n2595_;
  assign new_n2801_ = ~new_n2596_ & ~new_n2800_;
  assign new_n2802_ = ~new_n2764_ & new_n2792_;
  assign new_n2803_ = new_n2761_ & ~new_n2792_;
  assign new_n2804_ = ~new_n2802_ & ~new_n2803_;
  assign new_n2805_ = new_n2801_ & new_n2804_;
  assign new_n2806_ = ~new_n2590_ & new_n2805_;
  assign new_n2807_ = ~new_n2757_ & new_n2792_;
  assign new_n2808_ = ~new_n2754_ & ~new_n2792_;
  assign new_n2809_ = ~new_n2807_ & ~new_n2808_;
  assign new_n2810_ = ~new_n2806_ & ~new_n2809_;
  assign new_n2811_ = new_n2590_ & ~new_n2596_;
  assign new_n2812_ = ~new_n2597_ & ~new_n2811_;
  assign new_n2813_ = ~new_n2805_ & ~new_n2812_;
  assign new_n2814_ = ~new_n2597_ & new_n2622_;
  assign new_n2815_ = ~new_n2623_ & ~new_n2814_;
  assign new_n2816_ = ~new_n2770_ & new_n2792_;
  assign new_n2817_ = ~new_n2773_ & ~new_n2792_;
  assign new_n2818_ = ~new_n2816_ & ~new_n2817_;
  assign new_n2819_ = ~new_n2815_ & ~new_n2818_;
  assign new_n2820_ = ~new_n2813_ & ~new_n2819_;
  assign new_n2821_ = ~new_n2810_ & new_n2820_;
  assign new_n2822_ = new_n2815_ & new_n2818_;
  assign new_n2823_ = new_n2749_ & ~new_n2795_;
  assign new_n2824_ = ~new_n2793_ & ~new_n2823_;
  assign new_n2825_ = new_n2799_ & ~new_n2824_;
  assign new_n2826_ = ~new_n2822_ & ~new_n2825_;
  assign new_n2827_ = ~new_n2821_ & new_n2826_;
  assign new_n2828_ = ~new_n2799_ & new_n2824_;
  assign new_n2829_ = ~new_n2633_ & ~new_n2634_;
  assign new_n2830_ = ~new_n2635_ & ~new_n2829_;
  assign new_n2831_ = new_n2786_ & new_n2792_;
  assign new_n2832_ = ~new_n2786_ & ~new_n2789_;
  assign new_n2833_ = new_n2792_ & ~new_n2832_;
  assign new_n2834_ = new_n2785_ & ~new_n2833_;
  assign new_n2835_ = ~new_n2831_ & ~new_n2834_;
  assign new_n2836_ = ~new_n2830_ & new_n2835_;
  assign new_n2837_ = ~new_n2352_ & ~new_n2635_;
  assign new_n2838_ = ~new_n2828_ & ~new_n2837_;
  assign new_n2839_ = ~new_n2836_ & new_n2838_;
  assign new_n2840_ = ~new_n2827_ & new_n2839_;
  assign new_n2841_ = ~new_n2635_ & new_n2835_;
  assign new_n2842_ = new_n2352_ & ~new_n2829_;
  assign new_n2843_ = ~new_n2841_ & new_n2842_;
  assign new_n2844_ = ~new_n2840_ & ~new_n2843_;
  assign new_n2845_ = new_n2799_ & new_n2844_;
  assign new_n2846_ = new_n2824_ & ~new_n2844_;
  assign new_n2847_ = ~new_n2845_ & ~new_n2846_;
  assign new_n2848_ = new_n2797_ & ~new_n2847_;
  assign new_n2849_ = new_n2636_ & ~new_n2637_;
  assign new_n2850_ = ~new_n2754_ & new_n2792_;
  assign new_n2851_ = ~new_n2757_ & ~new_n2792_;
  assign new_n2852_ = ~new_n2850_ & ~new_n2851_;
  assign new_n2853_ = ~new_n2809_ & ~new_n2844_;
  assign new_n2854_ = new_n2812_ & new_n2844_;
  assign new_n2855_ = ~new_n2853_ & ~new_n2854_;
  assign new_n2856_ = ~new_n2852_ & new_n2855_;
  assign new_n2857_ = ~new_n2761_ & new_n2792_;
  assign new_n2858_ = new_n2764_ & ~new_n2792_;
  assign new_n2859_ = ~new_n2857_ & ~new_n2858_;
  assign new_n2860_ = ~new_n2801_ & new_n2844_;
  assign new_n2861_ = new_n2804_ & ~new_n2844_;
  assign new_n2862_ = ~new_n2860_ & ~new_n2861_;
  assign new_n2863_ = ~new_n2859_ & new_n2862_;
  assign new_n2864_ = ~new_n2856_ & new_n2863_;
  assign new_n2865_ = new_n2852_ & ~new_n2855_;
  assign new_n2866_ = new_n2770_ & ~new_n2792_;
  assign new_n2867_ = new_n2773_ & new_n2792_;
  assign new_n2868_ = ~new_n2866_ & ~new_n2867_;
  assign new_n2869_ = ~new_n2818_ & ~new_n2844_;
  assign new_n2870_ = new_n2815_ & new_n2844_;
  assign new_n2871_ = ~new_n2869_ & ~new_n2870_;
  assign new_n2872_ = ~new_n2868_ & ~new_n2871_;
  assign new_n2873_ = ~new_n2865_ & ~new_n2872_;
  assign new_n2874_ = ~new_n2864_ & new_n2873_;
  assign new_n2875_ = ~new_n2797_ & new_n2847_;
  assign new_n2876_ = new_n2868_ & new_n2871_;
  assign new_n2877_ = ~new_n2875_ & ~new_n2876_;
  assign new_n2878_ = ~new_n2874_ & new_n2877_;
  assign new_n2879_ = ~new_n2782_ & ~new_n2833_;
  assign new_n2880_ = ~new_n2831_ & ~new_n2879_;
  assign new_n2881_ = new_n2830_ & new_n2844_;
  assign new_n2882_ = new_n2835_ & ~new_n2844_;
  assign new_n2883_ = ~new_n2881_ & ~new_n2882_;
  assign new_n2884_ = new_n2880_ & ~new_n2883_;
  assign new_n2885_ = ~new_n2848_ & ~new_n2884_;
  assign new_n2886_ = ~new_n2878_ & new_n2885_;
  assign new_n2887_ = ~new_n2880_ & new_n2883_;
  assign new_n2888_ = ~new_n2638_ & ~new_n2887_;
  assign new_n2889_ = ~new_n2886_ & new_n2888_;
  assign new_n2890_ = ~new_n2849_ & ~new_n2889_;
  assign new_n2891_ = new_n2848_ & new_n2890_;
  assign new_n2892_ = ~new_n2848_ & ~new_n2875_;
  assign new_n2893_ = new_n2890_ & ~new_n2892_;
  assign new_n2894_ = ~new_n2797_ & ~new_n2893_;
  assign new_n2895_ = ~new_n2891_ & ~new_n2894_;
  assign new_n2896_ = ~new_n1472_ & new_n1481_;
  assign new_n2897_ = ~new_n1482_ & ~new_n2896_;
  assign new_n2898_ = new_n1464_ & ~new_n1470_;
  assign new_n2899_ = ~new_n1471_ & ~new_n2898_;
  assign new_n2900_ = ~new_n2855_ & ~new_n2890_;
  assign new_n2901_ = ~new_n2852_ & new_n2890_;
  assign new_n2902_ = ~new_n2900_ & ~new_n2901_;
  assign new_n2903_ = new_n2899_ & new_n2902_;
  assign new_n2904_ = new_n1466_ & ~new_n1469_;
  assign new_n2905_ = ~new_n1470_ & ~new_n2904_;
  assign new_n2906_ = ~new_n2859_ & new_n2890_;
  assign new_n2907_ = ~new_n2862_ & ~new_n2890_;
  assign new_n2908_ = ~new_n2906_ & ~new_n2907_;
  assign new_n2909_ = new_n2905_ & ~new_n2908_;
  assign new_n2910_ = ~new_n2903_ & ~new_n2909_;
  assign new_n2911_ = new_n1464_ & ~new_n2902_;
  assign new_n2912_ = new_n1462_ & ~new_n1471_;
  assign new_n2913_ = ~new_n1472_ & ~new_n2912_;
  assign new_n2914_ = ~new_n2868_ & new_n2890_;
  assign new_n2915_ = new_n2871_ & ~new_n2890_;
  assign new_n2916_ = ~new_n2914_ & ~new_n2915_;
  assign new_n2917_ = ~new_n2913_ & new_n2916_;
  assign new_n2918_ = ~new_n2911_ & ~new_n2917_;
  assign new_n2919_ = ~new_n2910_ & new_n2918_;
  assign new_n2920_ = new_n2847_ & ~new_n2893_;
  assign new_n2921_ = ~new_n2891_ & ~new_n2920_;
  assign new_n2922_ = new_n2897_ & ~new_n2921_;
  assign new_n2923_ = new_n2913_ & ~new_n2916_;
  assign new_n2924_ = ~new_n2922_ & ~new_n2923_;
  assign new_n2925_ = ~new_n2919_ & new_n2924_;
  assign new_n2926_ = ~new_n1482_ & ~new_n1483_;
  assign new_n2927_ = ~new_n1484_ & ~new_n2926_;
  assign new_n2928_ = new_n2884_ & new_n2890_;
  assign new_n2929_ = ~new_n2884_ & ~new_n2887_;
  assign new_n2930_ = new_n2890_ & ~new_n2929_;
  assign new_n2931_ = new_n2883_ & ~new_n2930_;
  assign new_n2932_ = ~new_n2928_ & ~new_n2931_;
  assign new_n2933_ = ~new_n2927_ & new_n2932_;
  assign new_n2934_ = ~new_n2897_ & new_n2921_;
  assign new_n2935_ = ~new_n1484_ & ~new_n2639_;
  assign new_n2936_ = ~new_n2933_ & ~new_n2935_;
  assign new_n2937_ = ~new_n2934_ & new_n2936_;
  assign new_n2938_ = ~new_n2925_ & new_n2937_;
  assign new_n2939_ = ~new_n1484_ & new_n2932_;
  assign new_n2940_ = new_n2639_ & ~new_n2926_;
  assign new_n2941_ = ~new_n2939_ & new_n2940_;
  assign new_n2942_ = ~new_n2938_ & ~new_n2941_;
  assign new_n2943_ = new_n2897_ & new_n2942_;
  assign new_n2944_ = new_n2921_ & ~new_n2942_;
  assign new_n2945_ = ~new_n2943_ & ~new_n2944_;
  assign new_n2946_ = new_n2895_ & ~new_n2945_;
  assign new_n2947_ = new_n2640_ & ~new_n2641_;
  assign new_n2948_ = ~new_n2902_ & ~new_n2942_;
  assign new_n2949_ = new_n2899_ & new_n2942_;
  assign new_n2950_ = ~new_n2948_ & ~new_n2949_;
  assign new_n2951_ = new_n2852_ & ~new_n2890_;
  assign new_n2952_ = new_n2855_ & new_n2890_;
  assign new_n2953_ = ~new_n2951_ & ~new_n2952_;
  assign new_n2954_ = new_n2950_ & new_n2953_;
  assign new_n2955_ = new_n2859_ & ~new_n2890_;
  assign new_n2956_ = new_n2862_ & new_n2890_;
  assign new_n2957_ = ~new_n2955_ & ~new_n2956_;
  assign new_n2958_ = ~new_n2905_ & new_n2942_;
  assign new_n2959_ = ~new_n2908_ & ~new_n2942_;
  assign new_n2960_ = ~new_n2958_ & ~new_n2959_;
  assign new_n2961_ = new_n2957_ & new_n2960_;
  assign new_n2962_ = ~new_n2954_ & new_n2961_;
  assign new_n2963_ = ~new_n2950_ & ~new_n2953_;
  assign new_n2964_ = ~new_n2871_ & new_n2890_;
  assign new_n2965_ = new_n2868_ & ~new_n2890_;
  assign new_n2966_ = ~new_n2964_ & ~new_n2965_;
  assign new_n2967_ = new_n2913_ & new_n2942_;
  assign new_n2968_ = new_n2916_ & ~new_n2942_;
  assign new_n2969_ = ~new_n2967_ & ~new_n2968_;
  assign new_n2970_ = new_n2966_ & ~new_n2969_;
  assign new_n2971_ = ~new_n2963_ & ~new_n2970_;
  assign new_n2972_ = ~new_n2962_ & new_n2971_;
  assign new_n2973_ = ~new_n2895_ & new_n2945_;
  assign new_n2974_ = ~new_n2966_ & new_n2969_;
  assign new_n2975_ = ~new_n2973_ & ~new_n2974_;
  assign new_n2976_ = ~new_n2972_ & new_n2975_;
  assign new_n2977_ = ~new_n2880_ & ~new_n2930_;
  assign new_n2978_ = ~new_n2928_ & ~new_n2977_;
  assign new_n2979_ = new_n2927_ & new_n2942_;
  assign new_n2980_ = new_n2932_ & ~new_n2942_;
  assign new_n2981_ = ~new_n2979_ & ~new_n2980_;
  assign new_n2982_ = new_n2978_ & ~new_n2981_;
  assign new_n2983_ = ~new_n2946_ & ~new_n2982_;
  assign new_n2984_ = ~new_n2976_ & new_n2983_;
  assign new_n2985_ = ~new_n2978_ & new_n2981_;
  assign new_n2986_ = ~new_n2640_ & new_n2641_;
  assign new_n2987_ = ~new_n2985_ & ~new_n2986_;
  assign new_n2988_ = ~new_n2984_ & new_n2987_;
  assign new_n2989_ = ~new_n2947_ & ~new_n2988_;
  assign new_n2990_ = new_n2946_ & new_n2989_;
  assign new_n2991_ = ~new_n2946_ & ~new_n2973_;
  assign new_n2992_ = new_n2989_ & ~new_n2991_;
  assign new_n2993_ = ~new_n2895_ & ~new_n2992_;
  assign new_n2994_ = ~new_n2990_ & ~new_n2993_;
  assign new_n2995_ = ~new_n1189_ & new_n1198_;
  assign new_n2996_ = ~new_n1199_ & ~new_n2995_;
  assign new_n2997_ = new_n1181_ & ~new_n1187_;
  assign new_n2998_ = ~new_n1188_ & ~new_n2997_;
  assign new_n2999_ = ~new_n2953_ & new_n2989_;
  assign new_n3000_ = new_n2950_ & ~new_n2989_;
  assign new_n3001_ = ~new_n2999_ & ~new_n3000_;
  assign new_n3002_ = new_n2998_ & ~new_n3001_;
  assign new_n3003_ = new_n1183_ & ~new_n1186_;
  assign new_n3004_ = ~new_n1187_ & ~new_n3003_;
  assign new_n3005_ = ~new_n2957_ & new_n2989_;
  assign new_n3006_ = new_n2960_ & ~new_n2989_;
  assign new_n3007_ = ~new_n3005_ & ~new_n3006_;
  assign new_n3008_ = new_n3004_ & new_n3007_;
  assign new_n3009_ = ~new_n3002_ & ~new_n3008_;
  assign new_n3010_ = new_n1181_ & new_n3001_;
  assign new_n3011_ = new_n1179_ & ~new_n1188_;
  assign new_n3012_ = ~new_n1189_ & ~new_n3011_;
  assign new_n3013_ = ~new_n2966_ & new_n2989_;
  assign new_n3014_ = ~new_n2969_ & ~new_n2989_;
  assign new_n3015_ = ~new_n3013_ & ~new_n3014_;
  assign new_n3016_ = ~new_n3012_ & ~new_n3015_;
  assign new_n3017_ = ~new_n3010_ & ~new_n3016_;
  assign new_n3018_ = ~new_n3009_ & new_n3017_;
  assign new_n3019_ = new_n2945_ & ~new_n2992_;
  assign new_n3020_ = ~new_n2990_ & ~new_n3019_;
  assign new_n3021_ = new_n2996_ & ~new_n3020_;
  assign new_n3022_ = new_n3012_ & new_n3015_;
  assign new_n3023_ = ~new_n3021_ & ~new_n3022_;
  assign new_n3024_ = ~new_n3018_ & new_n3023_;
  assign new_n3025_ = ~new_n1199_ & ~new_n1200_;
  assign new_n3026_ = ~new_n1201_ & ~new_n3025_;
  assign new_n3027_ = new_n2982_ & new_n2989_;
  assign new_n3028_ = ~new_n2982_ & ~new_n2985_;
  assign new_n3029_ = new_n2989_ & ~new_n3028_;
  assign new_n3030_ = new_n2981_ & ~new_n3029_;
  assign new_n3031_ = ~new_n3027_ & ~new_n3030_;
  assign new_n3032_ = ~new_n3026_ & new_n3031_;
  assign new_n3033_ = ~new_n2996_ & new_n3020_;
  assign new_n3034_ = ~new_n1201_ & ~new_n2642_;
  assign new_n3035_ = ~new_n3032_ & ~new_n3034_;
  assign new_n3036_ = ~new_n3033_ & new_n3035_;
  assign new_n3037_ = ~new_n3024_ & new_n3036_;
  assign new_n3038_ = ~new_n1201_ & new_n3031_;
  assign new_n3039_ = new_n2642_ & ~new_n3025_;
  assign new_n3040_ = ~new_n3038_ & new_n3039_;
  assign new_n3041_ = ~new_n3037_ & ~new_n3040_;
  assign new_n3042_ = new_n2996_ & new_n3041_;
  assign new_n3043_ = new_n3020_ & ~new_n3041_;
  assign new_n3044_ = ~new_n3042_ & ~new_n3043_;
  assign new_n3045_ = new_n2994_ & ~new_n3044_;
  assign new_n3046_ = new_n2643_ & ~new_n2644_;
  assign new_n3047_ = new_n3001_ & ~new_n3041_;
  assign new_n3048_ = new_n2998_ & new_n3041_;
  assign new_n3049_ = ~new_n3047_ & ~new_n3048_;
  assign new_n3050_ = ~new_n2953_ & ~new_n2989_;
  assign new_n3051_ = new_n2950_ & new_n2989_;
  assign new_n3052_ = ~new_n3050_ & ~new_n3051_;
  assign new_n3053_ = new_n3049_ & new_n3052_;
  assign new_n3054_ = new_n2957_ & ~new_n2989_;
  assign new_n3055_ = ~new_n2960_ & new_n2989_;
  assign new_n3056_ = ~new_n3054_ & ~new_n3055_;
  assign new_n3057_ = ~new_n3004_ & new_n3041_;
  assign new_n3058_ = new_n3007_ & ~new_n3041_;
  assign new_n3059_ = ~new_n3057_ & ~new_n3058_;
  assign new_n3060_ = ~new_n3056_ & new_n3059_;
  assign new_n3061_ = ~new_n3053_ & new_n3060_;
  assign new_n3062_ = ~new_n3049_ & ~new_n3052_;
  assign new_n3063_ = new_n2966_ & ~new_n2989_;
  assign new_n3064_ = new_n2969_ & new_n2989_;
  assign new_n3065_ = ~new_n3063_ & ~new_n3064_;
  assign new_n3066_ = ~new_n3015_ & ~new_n3041_;
  assign new_n3067_ = new_n3012_ & new_n3041_;
  assign new_n3068_ = ~new_n3066_ & ~new_n3067_;
  assign new_n3069_ = ~new_n3065_ & ~new_n3068_;
  assign new_n3070_ = ~new_n3062_ & ~new_n3069_;
  assign new_n3071_ = ~new_n3061_ & new_n3070_;
  assign new_n3072_ = ~new_n2994_ & new_n3044_;
  assign new_n3073_ = new_n3065_ & new_n3068_;
  assign new_n3074_ = ~new_n3072_ & ~new_n3073_;
  assign new_n3075_ = ~new_n3071_ & new_n3074_;
  assign new_n3076_ = ~new_n2978_ & ~new_n3029_;
  assign new_n3077_ = ~new_n3027_ & ~new_n3076_;
  assign new_n3078_ = new_n3026_ & new_n3041_;
  assign new_n3079_ = new_n3031_ & ~new_n3041_;
  assign new_n3080_ = ~new_n3078_ & ~new_n3079_;
  assign new_n3081_ = new_n3077_ & ~new_n3080_;
  assign new_n3082_ = ~new_n3045_ & ~new_n3081_;
  assign new_n3083_ = ~new_n3075_ & new_n3082_;
  assign new_n3084_ = ~new_n3077_ & new_n3080_;
  assign new_n3085_ = ~new_n2645_ & ~new_n3084_;
  assign new_n3086_ = ~new_n3083_ & new_n3085_;
  assign new_n3087_ = ~new_n3046_ & ~new_n3086_;
  assign new_n3088_ = new_n3045_ & new_n3087_;
  assign new_n3089_ = ~new_n3045_ & ~new_n3072_;
  assign new_n3090_ = new_n3087_ & ~new_n3089_;
  assign new_n3091_ = ~new_n2994_ & ~new_n3090_;
  assign new_n3092_ = ~new_n3088_ & ~new_n3091_;
  assign new_n3093_ = ~new_n906_ & new_n915_;
  assign new_n3094_ = ~new_n916_ & ~new_n3093_;
  assign new_n3095_ = new_n898_ & ~new_n904_;
  assign new_n3096_ = ~new_n905_ & ~new_n3095_;
  assign new_n3097_ = ~new_n3052_ & new_n3087_;
  assign new_n3098_ = new_n3049_ & ~new_n3087_;
  assign new_n3099_ = ~new_n3097_ & ~new_n3098_;
  assign new_n3100_ = new_n3096_ & ~new_n3099_;
  assign new_n3101_ = new_n900_ & ~new_n903_;
  assign new_n3102_ = ~new_n904_ & ~new_n3101_;
  assign new_n3103_ = new_n3059_ & ~new_n3087_;
  assign new_n3104_ = new_n3056_ & new_n3087_;
  assign new_n3105_ = ~new_n3103_ & ~new_n3104_;
  assign new_n3106_ = new_n3102_ & new_n3105_;
  assign new_n3107_ = ~new_n3100_ & ~new_n3106_;
  assign new_n3108_ = new_n898_ & new_n3099_;
  assign new_n3109_ = new_n896_ & ~new_n905_;
  assign new_n3110_ = ~new_n906_ & ~new_n3109_;
  assign new_n3111_ = ~new_n3065_ & new_n3087_;
  assign new_n3112_ = new_n3068_ & ~new_n3087_;
  assign new_n3113_ = ~new_n3111_ & ~new_n3112_;
  assign new_n3114_ = ~new_n3110_ & new_n3113_;
  assign new_n3115_ = ~new_n3108_ & ~new_n3114_;
  assign new_n3116_ = ~new_n3107_ & new_n3115_;
  assign new_n3117_ = new_n3044_ & ~new_n3090_;
  assign new_n3118_ = ~new_n3088_ & ~new_n3117_;
  assign new_n3119_ = new_n3094_ & ~new_n3118_;
  assign new_n3120_ = new_n3110_ & ~new_n3113_;
  assign new_n3121_ = ~new_n3119_ & ~new_n3120_;
  assign new_n3122_ = ~new_n3116_ & new_n3121_;
  assign new_n3123_ = ~new_n916_ & ~new_n917_;
  assign new_n3124_ = ~new_n918_ & ~new_n3123_;
  assign new_n3125_ = new_n3081_ & new_n3087_;
  assign new_n3126_ = ~new_n3081_ & ~new_n3084_;
  assign new_n3127_ = new_n3087_ & ~new_n3126_;
  assign new_n3128_ = new_n3080_ & ~new_n3127_;
  assign new_n3129_ = ~new_n3125_ & ~new_n3128_;
  assign new_n3130_ = ~new_n3124_ & new_n3129_;
  assign new_n3131_ = ~new_n3094_ & new_n3118_;
  assign new_n3132_ = ~new_n918_ & ~new_n2646_;
  assign new_n3133_ = ~new_n3130_ & ~new_n3132_;
  assign new_n3134_ = ~new_n3131_ & new_n3133_;
  assign new_n3135_ = ~new_n3122_ & new_n3134_;
  assign new_n3136_ = ~new_n918_ & new_n3129_;
  assign new_n3137_ = new_n2646_ & ~new_n3123_;
  assign new_n3138_ = ~new_n3136_ & new_n3137_;
  assign new_n3139_ = ~new_n3135_ & ~new_n3138_;
  assign new_n3140_ = new_n3094_ & new_n3139_;
  assign new_n3141_ = new_n3118_ & ~new_n3139_;
  assign new_n3142_ = ~new_n3140_ & ~new_n3141_;
  assign new_n3143_ = new_n3092_ & ~new_n3142_;
  assign new_n3144_ = new_n2647_ & ~new_n2648_;
  assign new_n3145_ = new_n3099_ & ~new_n3139_;
  assign new_n3146_ = new_n3096_ & new_n3139_;
  assign new_n3147_ = ~new_n3145_ & ~new_n3146_;
  assign new_n3148_ = ~new_n3052_ & ~new_n3087_;
  assign new_n3149_ = new_n3049_ & new_n3087_;
  assign new_n3150_ = ~new_n3148_ & ~new_n3149_;
  assign new_n3151_ = new_n3147_ & new_n3150_;
  assign new_n3152_ = ~new_n3102_ & new_n3139_;
  assign new_n3153_ = new_n3105_ & ~new_n3139_;
  assign new_n3154_ = ~new_n3152_ & ~new_n3153_;
  assign new_n3155_ = ~new_n3056_ & ~new_n3087_;
  assign new_n3156_ = ~new_n3059_ & new_n3087_;
  assign new_n3157_ = ~new_n3155_ & ~new_n3156_;
  assign new_n3158_ = new_n3154_ & ~new_n3157_;
  assign new_n3159_ = ~new_n3151_ & new_n3158_;
  assign new_n3160_ = ~new_n3147_ & ~new_n3150_;
  assign new_n3161_ = ~new_n3068_ & new_n3087_;
  assign new_n3162_ = new_n3065_ & ~new_n3087_;
  assign new_n3163_ = ~new_n3161_ & ~new_n3162_;
  assign new_n3164_ = new_n3110_ & new_n3139_;
  assign new_n3165_ = new_n3113_ & ~new_n3139_;
  assign new_n3166_ = ~new_n3164_ & ~new_n3165_;
  assign new_n3167_ = new_n3163_ & ~new_n3166_;
  assign new_n3168_ = ~new_n3160_ & ~new_n3167_;
  assign new_n3169_ = ~new_n3159_ & new_n3168_;
  assign new_n3170_ = ~new_n3092_ & new_n3142_;
  assign new_n3171_ = ~new_n3163_ & new_n3166_;
  assign new_n3172_ = ~new_n3170_ & ~new_n3171_;
  assign new_n3173_ = ~new_n3169_ & new_n3172_;
  assign new_n3174_ = ~new_n3077_ & ~new_n3127_;
  assign new_n3175_ = ~new_n3125_ & ~new_n3174_;
  assign new_n3176_ = new_n3124_ & new_n3139_;
  assign new_n3177_ = new_n3129_ & ~new_n3139_;
  assign new_n3178_ = ~new_n3176_ & ~new_n3177_;
  assign new_n3179_ = new_n3175_ & ~new_n3178_;
  assign new_n3180_ = ~new_n3143_ & ~new_n3179_;
  assign new_n3181_ = ~new_n3173_ & new_n3180_;
  assign new_n3182_ = ~new_n3175_ & new_n3178_;
  assign new_n3183_ = ~new_n2649_ & ~new_n3182_;
  assign new_n3184_ = ~new_n3181_ & new_n3183_;
  assign new_n3185_ = ~new_n3144_ & ~new_n3184_;
  assign new_n3186_ = new_n3143_ & new_n3185_;
  assign new_n3187_ = ~new_n3143_ & ~new_n3170_;
  assign new_n3188_ = new_n3185_ & ~new_n3187_;
  assign new_n3189_ = ~new_n3092_ & ~new_n3188_;
  assign new_n3190_ = ~new_n3186_ & ~new_n3189_;
  assign new_n3191_ = new_n3142_ & ~new_n3188_;
  assign new_n3192_ = ~new_n3186_ & ~new_n3191_;
  assign new_n3193_ = new_n624_ & ~new_n630_;
  assign new_n3194_ = ~new_n631_ & ~new_n3193_;
  assign new_n3195_ = ~new_n3150_ & new_n3185_;
  assign new_n3196_ = new_n3147_ & ~new_n3185_;
  assign new_n3197_ = ~new_n3195_ & ~new_n3196_;
  assign new_n3198_ = new_n3194_ & ~new_n3197_;
  assign new_n3199_ = new_n626_ & ~new_n629_;
  assign new_n3200_ = ~new_n630_ & ~new_n3199_;
  assign new_n3201_ = ~new_n3157_ & new_n3185_;
  assign new_n3202_ = ~new_n3154_ & ~new_n3185_;
  assign new_n3203_ = ~new_n3201_ & ~new_n3202_;
  assign new_n3204_ = new_n3200_ & ~new_n3203_;
  assign new_n3205_ = ~new_n3198_ & ~new_n3204_;
  assign new_n3206_ = new_n624_ & new_n3197_;
  assign new_n3207_ = new_n622_ & ~new_n631_;
  assign new_n3208_ = ~new_n632_ & ~new_n3207_;
  assign new_n3209_ = ~new_n3163_ & new_n3185_;
  assign new_n3210_ = ~new_n3166_ & ~new_n3185_;
  assign new_n3211_ = ~new_n3209_ & ~new_n3210_;
  assign new_n3212_ = ~new_n3208_ & ~new_n3211_;
  assign new_n3213_ = ~new_n3206_ & ~new_n3212_;
  assign new_n3214_ = ~new_n3205_ & new_n3213_;
  assign new_n3215_ = new_n620_ & ~new_n632_;
  assign new_n3216_ = ~new_n633_ & ~new_n3215_;
  assign new_n3217_ = ~new_n3192_ & new_n3216_;
  assign new_n3218_ = new_n3208_ & new_n3211_;
  assign new_n3219_ = ~new_n3217_ & ~new_n3218_;
  assign new_n3220_ = ~new_n3214_ & new_n3219_;
  assign new_n3221_ = new_n3179_ & new_n3185_;
  assign new_n3222_ = ~new_n3179_ & ~new_n3182_;
  assign new_n3223_ = new_n3185_ & ~new_n3222_;
  assign new_n3224_ = new_n3178_ & ~new_n3223_;
  assign new_n3225_ = ~new_n3221_ & ~new_n3224_;
  assign new_n3226_ = ~new_n633_ & ~new_n634_;
  assign new_n3227_ = ~new_n635_ & ~new_n3226_;
  assign new_n3228_ = new_n3225_ & ~new_n3227_;
  assign new_n3229_ = new_n3192_ & ~new_n3216_;
  assign new_n3230_ = ~new_n635_ & ~new_n2650_;
  assign new_n3231_ = ~new_n3228_ & ~new_n3230_;
  assign new_n3232_ = ~new_n3229_ & new_n3231_;
  assign new_n3233_ = ~new_n3220_ & new_n3232_;
  assign new_n3234_ = ~new_n635_ & new_n3225_;
  assign new_n3235_ = new_n2650_ & ~new_n3226_;
  assign new_n3236_ = ~new_n3234_ & new_n3235_;
  assign new_n3237_ = ~new_n3233_ & ~new_n3236_;
  assign new_n3238_ = ~new_n3192_ & ~new_n3237_;
  assign new_n3239_ = ~new_n3216_ & new_n3237_;
  assign new_n3240_ = ~new_n3238_ & ~new_n3239_;
  assign new_n3241_ = new_n3190_ & new_n3240_;
  assign new_n3242_ = ~new_n3166_ & new_n3185_;
  assign new_n3243_ = ~new_n3163_ & ~new_n3185_;
  assign new_n3244_ = ~new_n3242_ & ~new_n3243_;
  assign new_n3245_ = ~new_n3211_ & ~new_n3237_;
  assign new_n3246_ = new_n3208_ & new_n3237_;
  assign new_n3247_ = ~new_n3245_ & ~new_n3246_;
  assign new_n3248_ = new_n3244_ & ~new_n3247_;
  assign new_n3249_ = ~new_n3147_ & new_n3185_;
  assign new_n3250_ = new_n3150_ & ~new_n3185_;
  assign new_n3251_ = ~new_n3249_ & ~new_n3250_;
  assign new_n3252_ = ~new_n3200_ & new_n3237_;
  assign new_n3253_ = ~new_n3203_ & ~new_n3237_;
  assign new_n3254_ = new_n3154_ & new_n3185_;
  assign new_n3255_ = new_n3157_ & ~new_n3185_;
  assign new_n3256_ = ~new_n3254_ & ~new_n3255_;
  assign new_n3257_ = ~new_n3252_ & new_n3256_;
  assign new_n3258_ = ~new_n3253_ & new_n3257_;
  assign new_n3259_ = ~new_n3194_ & new_n3237_;
  assign new_n3260_ = ~new_n3197_ & ~new_n3237_;
  assign new_n3261_ = ~new_n3259_ & ~new_n3260_;
  assign new_n3262_ = new_n3258_ & new_n3261_;
  assign new_n3263_ = ~new_n3251_ & ~new_n3262_;
  assign new_n3264_ = ~new_n3244_ & new_n3247_;
  assign new_n3265_ = ~new_n3258_ & ~new_n3261_;
  assign new_n3266_ = ~new_n3264_ & ~new_n3265_;
  assign new_n3267_ = ~new_n3263_ & new_n3266_;
  assign new_n3268_ = ~new_n3241_ & ~new_n3248_;
  assign new_n3269_ = ~new_n3267_ & new_n3268_;
  assign new_n3270_ = ~new_n3175_ & ~new_n3223_;
  assign new_n3271_ = ~new_n3221_ & ~new_n3270_;
  assign new_n3272_ = new_n3225_ & ~new_n3237_;
  assign new_n3273_ = new_n3227_ & new_n3237_;
  assign new_n3274_ = ~new_n3272_ & ~new_n3273_;
  assign new_n3275_ = ~new_n3271_ & new_n3274_;
  assign new_n3276_ = ~new_n3190_ & ~new_n3240_;
  assign new_n3277_ = ~new_n3275_ & ~new_n3276_;
  assign new_n3278_ = ~new_n3269_ & new_n3277_;
  assign new_n3279_ = new_n2651_ & ~new_n2652_;
  assign new_n3280_ = new_n3271_ & ~new_n3274_;
  assign new_n3281_ = ~new_n3279_ & ~new_n3280_;
  assign new_n3282_ = ~new_n3278_ & new_n3281_;
  assign new_n3283_ = ~new_n2653_ & ~new_n3282_;
  assign new_n3284_ = \p_input[192]  & ~new_n2694_;
  assign new_n3285_ = \p_input[224]  & new_n2694_;
  assign new_n3286_ = ~new_n3284_ & ~new_n3285_;
  assign new_n3287_ = ~new_n2792_ & ~new_n3286_;
  assign new_n3288_ = ~\p_input[224]  & ~new_n2694_;
  assign new_n3289_ = ~\p_input[192]  & new_n2694_;
  assign new_n3290_ = ~new_n3288_ & ~new_n3289_;
  assign new_n3291_ = ~new_n2746_ & ~new_n3290_;
  assign new_n3292_ = ~\p_input[160]  & new_n2746_;
  assign new_n3293_ = ~new_n3291_ & ~new_n3292_;
  assign new_n3294_ = new_n2792_ & new_n3293_;
  assign new_n3295_ = ~new_n3287_ & ~new_n3294_;
  assign new_n3296_ = ~new_n2890_ & ~new_n3295_;
  assign new_n3297_ = new_n2792_ & ~new_n3286_;
  assign new_n3298_ = ~new_n2792_ & new_n3293_;
  assign new_n3299_ = ~new_n3297_ & ~new_n3298_;
  assign new_n3300_ = ~new_n2844_ & ~new_n3299_;
  assign new_n3301_ = \p_input[128]  & new_n2844_;
  assign new_n3302_ = ~new_n3300_ & ~new_n3301_;
  assign new_n3303_ = new_n2890_ & ~new_n3302_;
  assign new_n3304_ = ~new_n3296_ & ~new_n3303_;
  assign new_n3305_ = ~new_n2989_ & ~new_n3304_;
  assign new_n3306_ = new_n2890_ & ~new_n3295_;
  assign new_n3307_ = ~new_n2890_ & ~new_n3302_;
  assign new_n3308_ = ~new_n3306_ & ~new_n3307_;
  assign new_n3309_ = ~new_n2942_ & ~new_n3308_;
  assign new_n3310_ = \p_input[96]  & new_n2942_;
  assign new_n3311_ = ~new_n3309_ & ~new_n3310_;
  assign new_n3312_ = new_n2989_ & ~new_n3311_;
  assign new_n3313_ = ~new_n3305_ & ~new_n3312_;
  assign new_n3314_ = ~new_n3087_ & ~new_n3313_;
  assign new_n3315_ = new_n2989_ & ~new_n3304_;
  assign new_n3316_ = ~new_n2989_ & ~new_n3311_;
  assign new_n3317_ = ~new_n3315_ & ~new_n3316_;
  assign new_n3318_ = ~new_n3041_ & ~new_n3317_;
  assign new_n3319_ = \p_input[64]  & new_n3041_;
  assign new_n3320_ = ~new_n3318_ & ~new_n3319_;
  assign new_n3321_ = new_n3087_ & ~new_n3320_;
  assign new_n3322_ = ~new_n3314_ & ~new_n3321_;
  assign new_n3323_ = ~new_n3185_ & ~new_n3322_;
  assign new_n3324_ = new_n3087_ & ~new_n3313_;
  assign new_n3325_ = ~new_n3087_ & ~new_n3320_;
  assign new_n3326_ = ~new_n3324_ & ~new_n3325_;
  assign new_n3327_ = ~new_n3139_ & ~new_n3326_;
  assign new_n3328_ = \p_input[32]  & new_n3139_;
  assign new_n3329_ = ~new_n3327_ & ~new_n3328_;
  assign new_n3330_ = new_n3185_ & ~new_n3329_;
  assign new_n3331_ = ~new_n3323_ & ~new_n3330_;
  assign new_n3332_ = new_n3283_ & ~new_n3331_;
  assign new_n3333_ = new_n3185_ & ~new_n3322_;
  assign new_n3334_ = ~new_n3185_ & ~new_n3329_;
  assign new_n3335_ = ~new_n3333_ & ~new_n3334_;
  assign new_n3336_ = ~new_n3237_ & ~new_n3335_;
  assign new_n3337_ = \p_input[0]  & new_n3237_;
  assign new_n3338_ = ~new_n3336_ & ~new_n3337_;
  assign new_n3339_ = ~new_n3283_ & ~new_n3338_;
  assign \o[0]  = new_n3332_ | new_n3339_;
  assign new_n3341_ = \p_input[193]  & ~new_n2694_;
  assign new_n3342_ = \p_input[225]  & new_n2694_;
  assign new_n3343_ = ~new_n3341_ & ~new_n3342_;
  assign new_n3344_ = ~new_n2792_ & ~new_n3343_;
  assign new_n3345_ = ~\p_input[225]  & ~new_n2694_;
  assign new_n3346_ = ~\p_input[193]  & new_n2694_;
  assign new_n3347_ = ~new_n3345_ & ~new_n3346_;
  assign new_n3348_ = ~new_n2746_ & ~new_n3347_;
  assign new_n3349_ = ~\p_input[161]  & new_n2746_;
  assign new_n3350_ = ~new_n3348_ & ~new_n3349_;
  assign new_n3351_ = new_n2792_ & new_n3350_;
  assign new_n3352_ = ~new_n3344_ & ~new_n3351_;
  assign new_n3353_ = ~new_n2890_ & ~new_n3352_;
  assign new_n3354_ = new_n2792_ & ~new_n3343_;
  assign new_n3355_ = ~new_n2792_ & new_n3350_;
  assign new_n3356_ = ~new_n3354_ & ~new_n3355_;
  assign new_n3357_ = ~new_n2844_ & ~new_n3356_;
  assign new_n3358_ = \p_input[129]  & new_n2844_;
  assign new_n3359_ = ~new_n3357_ & ~new_n3358_;
  assign new_n3360_ = new_n2890_ & ~new_n3359_;
  assign new_n3361_ = ~new_n3353_ & ~new_n3360_;
  assign new_n3362_ = ~new_n2989_ & ~new_n3361_;
  assign new_n3363_ = new_n2890_ & ~new_n3352_;
  assign new_n3364_ = ~new_n2890_ & ~new_n3359_;
  assign new_n3365_ = ~new_n3363_ & ~new_n3364_;
  assign new_n3366_ = ~new_n2942_ & ~new_n3365_;
  assign new_n3367_ = \p_input[97]  & new_n2942_;
  assign new_n3368_ = ~new_n3366_ & ~new_n3367_;
  assign new_n3369_ = new_n2989_ & ~new_n3368_;
  assign new_n3370_ = ~new_n3362_ & ~new_n3369_;
  assign new_n3371_ = ~new_n3087_ & ~new_n3370_;
  assign new_n3372_ = new_n2989_ & ~new_n3361_;
  assign new_n3373_ = ~new_n2989_ & ~new_n3368_;
  assign new_n3374_ = ~new_n3372_ & ~new_n3373_;
  assign new_n3375_ = ~new_n3041_ & ~new_n3374_;
  assign new_n3376_ = \p_input[65]  & new_n3041_;
  assign new_n3377_ = ~new_n3375_ & ~new_n3376_;
  assign new_n3378_ = new_n3087_ & ~new_n3377_;
  assign new_n3379_ = ~new_n3371_ & ~new_n3378_;
  assign new_n3380_ = ~new_n3185_ & ~new_n3379_;
  assign new_n3381_ = new_n3087_ & ~new_n3370_;
  assign new_n3382_ = ~new_n3087_ & ~new_n3377_;
  assign new_n3383_ = ~new_n3381_ & ~new_n3382_;
  assign new_n3384_ = ~new_n3139_ & ~new_n3383_;
  assign new_n3385_ = \p_input[33]  & new_n3139_;
  assign new_n3386_ = ~new_n3384_ & ~new_n3385_;
  assign new_n3387_ = new_n3185_ & ~new_n3386_;
  assign new_n3388_ = ~new_n3380_ & ~new_n3387_;
  assign new_n3389_ = new_n3283_ & ~new_n3388_;
  assign new_n3390_ = new_n3185_ & ~new_n3379_;
  assign new_n3391_ = ~new_n3185_ & ~new_n3386_;
  assign new_n3392_ = ~new_n3390_ & ~new_n3391_;
  assign new_n3393_ = ~new_n3237_ & ~new_n3392_;
  assign new_n3394_ = \p_input[1]  & new_n3237_;
  assign new_n3395_ = ~new_n3393_ & ~new_n3394_;
  assign new_n3396_ = ~new_n3283_ & ~new_n3395_;
  assign \o[1]  = new_n3389_ | new_n3396_;
  assign new_n3398_ = \p_input[194]  & ~new_n2694_;
  assign new_n3399_ = \p_input[226]  & new_n2694_;
  assign new_n3400_ = ~new_n3398_ & ~new_n3399_;
  assign new_n3401_ = ~new_n2792_ & ~new_n3400_;
  assign new_n3402_ = ~\p_input[226]  & ~new_n2694_;
  assign new_n3403_ = ~\p_input[194]  & new_n2694_;
  assign new_n3404_ = ~new_n3402_ & ~new_n3403_;
  assign new_n3405_ = ~new_n2746_ & ~new_n3404_;
  assign new_n3406_ = ~\p_input[162]  & new_n2746_;
  assign new_n3407_ = ~new_n3405_ & ~new_n3406_;
  assign new_n3408_ = new_n2792_ & new_n3407_;
  assign new_n3409_ = ~new_n3401_ & ~new_n3408_;
  assign new_n3410_ = ~new_n2890_ & ~new_n3409_;
  assign new_n3411_ = new_n2792_ & ~new_n3400_;
  assign new_n3412_ = ~new_n2792_ & new_n3407_;
  assign new_n3413_ = ~new_n3411_ & ~new_n3412_;
  assign new_n3414_ = ~new_n2844_ & ~new_n3413_;
  assign new_n3415_ = \p_input[130]  & new_n2844_;
  assign new_n3416_ = ~new_n3414_ & ~new_n3415_;
  assign new_n3417_ = new_n2890_ & ~new_n3416_;
  assign new_n3418_ = ~new_n3410_ & ~new_n3417_;
  assign new_n3419_ = ~new_n2989_ & ~new_n3418_;
  assign new_n3420_ = new_n2890_ & ~new_n3409_;
  assign new_n3421_ = ~new_n2890_ & ~new_n3416_;
  assign new_n3422_ = ~new_n3420_ & ~new_n3421_;
  assign new_n3423_ = ~new_n2942_ & ~new_n3422_;
  assign new_n3424_ = \p_input[98]  & new_n2942_;
  assign new_n3425_ = ~new_n3423_ & ~new_n3424_;
  assign new_n3426_ = new_n2989_ & ~new_n3425_;
  assign new_n3427_ = ~new_n3419_ & ~new_n3426_;
  assign new_n3428_ = ~new_n3087_ & ~new_n3427_;
  assign new_n3429_ = new_n2989_ & ~new_n3418_;
  assign new_n3430_ = ~new_n2989_ & ~new_n3425_;
  assign new_n3431_ = ~new_n3429_ & ~new_n3430_;
  assign new_n3432_ = ~new_n3041_ & ~new_n3431_;
  assign new_n3433_ = \p_input[66]  & new_n3041_;
  assign new_n3434_ = ~new_n3432_ & ~new_n3433_;
  assign new_n3435_ = new_n3087_ & ~new_n3434_;
  assign new_n3436_ = ~new_n3428_ & ~new_n3435_;
  assign new_n3437_ = ~new_n3185_ & ~new_n3436_;
  assign new_n3438_ = new_n3087_ & ~new_n3427_;
  assign new_n3439_ = ~new_n3087_ & ~new_n3434_;
  assign new_n3440_ = ~new_n3438_ & ~new_n3439_;
  assign new_n3441_ = ~new_n3139_ & ~new_n3440_;
  assign new_n3442_ = \p_input[34]  & new_n3139_;
  assign new_n3443_ = ~new_n3441_ & ~new_n3442_;
  assign new_n3444_ = new_n3185_ & ~new_n3443_;
  assign new_n3445_ = ~new_n3437_ & ~new_n3444_;
  assign new_n3446_ = new_n3283_ & ~new_n3445_;
  assign new_n3447_ = new_n3185_ & ~new_n3436_;
  assign new_n3448_ = ~new_n3185_ & ~new_n3443_;
  assign new_n3449_ = ~new_n3447_ & ~new_n3448_;
  assign new_n3450_ = ~new_n3237_ & ~new_n3449_;
  assign new_n3451_ = \p_input[2]  & new_n3237_;
  assign new_n3452_ = ~new_n3450_ & ~new_n3451_;
  assign new_n3453_ = ~new_n3283_ & ~new_n3452_;
  assign \o[2]  = new_n3446_ | new_n3453_;
  assign new_n3455_ = \p_input[195]  & ~new_n2694_;
  assign new_n3456_ = \p_input[227]  & new_n2694_;
  assign new_n3457_ = ~new_n3455_ & ~new_n3456_;
  assign new_n3458_ = ~new_n2792_ & ~new_n3457_;
  assign new_n3459_ = ~\p_input[227]  & ~new_n2694_;
  assign new_n3460_ = ~\p_input[195]  & new_n2694_;
  assign new_n3461_ = ~new_n3459_ & ~new_n3460_;
  assign new_n3462_ = ~new_n2746_ & ~new_n3461_;
  assign new_n3463_ = ~\p_input[163]  & new_n2746_;
  assign new_n3464_ = ~new_n3462_ & ~new_n3463_;
  assign new_n3465_ = new_n2792_ & new_n3464_;
  assign new_n3466_ = ~new_n3458_ & ~new_n3465_;
  assign new_n3467_ = ~new_n2890_ & ~new_n3466_;
  assign new_n3468_ = new_n2792_ & ~new_n3457_;
  assign new_n3469_ = ~new_n2792_ & new_n3464_;
  assign new_n3470_ = ~new_n3468_ & ~new_n3469_;
  assign new_n3471_ = ~new_n2844_ & ~new_n3470_;
  assign new_n3472_ = \p_input[131]  & new_n2844_;
  assign new_n3473_ = ~new_n3471_ & ~new_n3472_;
  assign new_n3474_ = new_n2890_ & ~new_n3473_;
  assign new_n3475_ = ~new_n3467_ & ~new_n3474_;
  assign new_n3476_ = ~new_n2989_ & ~new_n3475_;
  assign new_n3477_ = new_n2890_ & ~new_n3466_;
  assign new_n3478_ = ~new_n2890_ & ~new_n3473_;
  assign new_n3479_ = ~new_n3477_ & ~new_n3478_;
  assign new_n3480_ = ~new_n2942_ & ~new_n3479_;
  assign new_n3481_ = \p_input[99]  & new_n2942_;
  assign new_n3482_ = ~new_n3480_ & ~new_n3481_;
  assign new_n3483_ = new_n2989_ & ~new_n3482_;
  assign new_n3484_ = ~new_n3476_ & ~new_n3483_;
  assign new_n3485_ = ~new_n3087_ & ~new_n3484_;
  assign new_n3486_ = new_n2989_ & ~new_n3475_;
  assign new_n3487_ = ~new_n2989_ & ~new_n3482_;
  assign new_n3488_ = ~new_n3486_ & ~new_n3487_;
  assign new_n3489_ = ~new_n3041_ & ~new_n3488_;
  assign new_n3490_ = \p_input[67]  & new_n3041_;
  assign new_n3491_ = ~new_n3489_ & ~new_n3490_;
  assign new_n3492_ = new_n3087_ & ~new_n3491_;
  assign new_n3493_ = ~new_n3485_ & ~new_n3492_;
  assign new_n3494_ = ~new_n3185_ & ~new_n3493_;
  assign new_n3495_ = new_n3087_ & ~new_n3484_;
  assign new_n3496_ = ~new_n3087_ & ~new_n3491_;
  assign new_n3497_ = ~new_n3495_ & ~new_n3496_;
  assign new_n3498_ = ~new_n3139_ & ~new_n3497_;
  assign new_n3499_ = \p_input[35]  & new_n3139_;
  assign new_n3500_ = ~new_n3498_ & ~new_n3499_;
  assign new_n3501_ = new_n3185_ & ~new_n3500_;
  assign new_n3502_ = ~new_n3494_ & ~new_n3501_;
  assign new_n3503_ = new_n3283_ & ~new_n3502_;
  assign new_n3504_ = new_n3185_ & ~new_n3493_;
  assign new_n3505_ = ~new_n3185_ & ~new_n3500_;
  assign new_n3506_ = ~new_n3504_ & ~new_n3505_;
  assign new_n3507_ = ~new_n3237_ & ~new_n3506_;
  assign new_n3508_ = \p_input[3]  & new_n3237_;
  assign new_n3509_ = ~new_n3507_ & ~new_n3508_;
  assign new_n3510_ = ~new_n3283_ & ~new_n3509_;
  assign \o[3]  = new_n3503_ | new_n3510_;
  assign new_n3512_ = \p_input[196]  & ~new_n2694_;
  assign new_n3513_ = \p_input[228]  & new_n2694_;
  assign new_n3514_ = ~new_n3512_ & ~new_n3513_;
  assign new_n3515_ = ~new_n2792_ & ~new_n3514_;
  assign new_n3516_ = ~\p_input[228]  & ~new_n2694_;
  assign new_n3517_ = ~\p_input[196]  & new_n2694_;
  assign new_n3518_ = ~new_n3516_ & ~new_n3517_;
  assign new_n3519_ = ~new_n2746_ & ~new_n3518_;
  assign new_n3520_ = ~\p_input[164]  & new_n2746_;
  assign new_n3521_ = ~new_n3519_ & ~new_n3520_;
  assign new_n3522_ = new_n2792_ & new_n3521_;
  assign new_n3523_ = ~new_n3515_ & ~new_n3522_;
  assign new_n3524_ = ~new_n2890_ & ~new_n3523_;
  assign new_n3525_ = new_n2792_ & ~new_n3514_;
  assign new_n3526_ = ~new_n2792_ & new_n3521_;
  assign new_n3527_ = ~new_n3525_ & ~new_n3526_;
  assign new_n3528_ = ~new_n2844_ & ~new_n3527_;
  assign new_n3529_ = \p_input[132]  & new_n2844_;
  assign new_n3530_ = ~new_n3528_ & ~new_n3529_;
  assign new_n3531_ = new_n2890_ & ~new_n3530_;
  assign new_n3532_ = ~new_n3524_ & ~new_n3531_;
  assign new_n3533_ = ~new_n2989_ & ~new_n3532_;
  assign new_n3534_ = new_n2890_ & ~new_n3523_;
  assign new_n3535_ = ~new_n2890_ & ~new_n3530_;
  assign new_n3536_ = ~new_n3534_ & ~new_n3535_;
  assign new_n3537_ = ~new_n2942_ & ~new_n3536_;
  assign new_n3538_ = \p_input[100]  & new_n2942_;
  assign new_n3539_ = ~new_n3537_ & ~new_n3538_;
  assign new_n3540_ = new_n2989_ & ~new_n3539_;
  assign new_n3541_ = ~new_n3533_ & ~new_n3540_;
  assign new_n3542_ = ~new_n3087_ & ~new_n3541_;
  assign new_n3543_ = new_n2989_ & ~new_n3532_;
  assign new_n3544_ = ~new_n2989_ & ~new_n3539_;
  assign new_n3545_ = ~new_n3543_ & ~new_n3544_;
  assign new_n3546_ = ~new_n3041_ & ~new_n3545_;
  assign new_n3547_ = \p_input[68]  & new_n3041_;
  assign new_n3548_ = ~new_n3546_ & ~new_n3547_;
  assign new_n3549_ = new_n3087_ & ~new_n3548_;
  assign new_n3550_ = ~new_n3542_ & ~new_n3549_;
  assign new_n3551_ = ~new_n3185_ & ~new_n3550_;
  assign new_n3552_ = new_n3087_ & ~new_n3541_;
  assign new_n3553_ = ~new_n3087_ & ~new_n3548_;
  assign new_n3554_ = ~new_n3552_ & ~new_n3553_;
  assign new_n3555_ = ~new_n3139_ & ~new_n3554_;
  assign new_n3556_ = \p_input[36]  & new_n3139_;
  assign new_n3557_ = ~new_n3555_ & ~new_n3556_;
  assign new_n3558_ = new_n3185_ & ~new_n3557_;
  assign new_n3559_ = ~new_n3551_ & ~new_n3558_;
  assign new_n3560_ = new_n3283_ & ~new_n3559_;
  assign new_n3561_ = new_n3185_ & ~new_n3550_;
  assign new_n3562_ = ~new_n3185_ & ~new_n3557_;
  assign new_n3563_ = ~new_n3561_ & ~new_n3562_;
  assign new_n3564_ = ~new_n3237_ & ~new_n3563_;
  assign new_n3565_ = \p_input[4]  & new_n3237_;
  assign new_n3566_ = ~new_n3564_ & ~new_n3565_;
  assign new_n3567_ = ~new_n3283_ & ~new_n3566_;
  assign \o[4]  = new_n3560_ | new_n3567_;
  assign new_n3569_ = \p_input[197]  & ~new_n2694_;
  assign new_n3570_ = \p_input[229]  & new_n2694_;
  assign new_n3571_ = ~new_n3569_ & ~new_n3570_;
  assign new_n3572_ = ~new_n2792_ & ~new_n3571_;
  assign new_n3573_ = ~\p_input[229]  & ~new_n2694_;
  assign new_n3574_ = ~\p_input[197]  & new_n2694_;
  assign new_n3575_ = ~new_n3573_ & ~new_n3574_;
  assign new_n3576_ = ~new_n2746_ & ~new_n3575_;
  assign new_n3577_ = ~\p_input[165]  & new_n2746_;
  assign new_n3578_ = ~new_n3576_ & ~new_n3577_;
  assign new_n3579_ = new_n2792_ & new_n3578_;
  assign new_n3580_ = ~new_n3572_ & ~new_n3579_;
  assign new_n3581_ = ~new_n2890_ & ~new_n3580_;
  assign new_n3582_ = new_n2792_ & ~new_n3571_;
  assign new_n3583_ = ~new_n2792_ & new_n3578_;
  assign new_n3584_ = ~new_n3582_ & ~new_n3583_;
  assign new_n3585_ = ~new_n2844_ & ~new_n3584_;
  assign new_n3586_ = \p_input[133]  & new_n2844_;
  assign new_n3587_ = ~new_n3585_ & ~new_n3586_;
  assign new_n3588_ = new_n2890_ & ~new_n3587_;
  assign new_n3589_ = ~new_n3581_ & ~new_n3588_;
  assign new_n3590_ = ~new_n2989_ & ~new_n3589_;
  assign new_n3591_ = new_n2890_ & ~new_n3580_;
  assign new_n3592_ = ~new_n2890_ & ~new_n3587_;
  assign new_n3593_ = ~new_n3591_ & ~new_n3592_;
  assign new_n3594_ = ~new_n2942_ & ~new_n3593_;
  assign new_n3595_ = \p_input[101]  & new_n2942_;
  assign new_n3596_ = ~new_n3594_ & ~new_n3595_;
  assign new_n3597_ = new_n2989_ & ~new_n3596_;
  assign new_n3598_ = ~new_n3590_ & ~new_n3597_;
  assign new_n3599_ = ~new_n3087_ & ~new_n3598_;
  assign new_n3600_ = new_n2989_ & ~new_n3589_;
  assign new_n3601_ = ~new_n2989_ & ~new_n3596_;
  assign new_n3602_ = ~new_n3600_ & ~new_n3601_;
  assign new_n3603_ = ~new_n3041_ & ~new_n3602_;
  assign new_n3604_ = \p_input[69]  & new_n3041_;
  assign new_n3605_ = ~new_n3603_ & ~new_n3604_;
  assign new_n3606_ = new_n3087_ & ~new_n3605_;
  assign new_n3607_ = ~new_n3599_ & ~new_n3606_;
  assign new_n3608_ = ~new_n3185_ & ~new_n3607_;
  assign new_n3609_ = new_n3087_ & ~new_n3598_;
  assign new_n3610_ = ~new_n3087_ & ~new_n3605_;
  assign new_n3611_ = ~new_n3609_ & ~new_n3610_;
  assign new_n3612_ = ~new_n3139_ & ~new_n3611_;
  assign new_n3613_ = \p_input[37]  & new_n3139_;
  assign new_n3614_ = ~new_n3612_ & ~new_n3613_;
  assign new_n3615_ = new_n3185_ & ~new_n3614_;
  assign new_n3616_ = ~new_n3608_ & ~new_n3615_;
  assign new_n3617_ = new_n3283_ & ~new_n3616_;
  assign new_n3618_ = new_n3185_ & ~new_n3607_;
  assign new_n3619_ = ~new_n3185_ & ~new_n3614_;
  assign new_n3620_ = ~new_n3618_ & ~new_n3619_;
  assign new_n3621_ = ~new_n3237_ & ~new_n3620_;
  assign new_n3622_ = \p_input[5]  & new_n3237_;
  assign new_n3623_ = ~new_n3621_ & ~new_n3622_;
  assign new_n3624_ = ~new_n3283_ & ~new_n3623_;
  assign \o[5]  = new_n3617_ | new_n3624_;
  assign new_n3626_ = \p_input[198]  & ~new_n2694_;
  assign new_n3627_ = \p_input[230]  & new_n2694_;
  assign new_n3628_ = ~new_n3626_ & ~new_n3627_;
  assign new_n3629_ = ~new_n2792_ & ~new_n3628_;
  assign new_n3630_ = ~\p_input[230]  & ~new_n2694_;
  assign new_n3631_ = ~\p_input[198]  & new_n2694_;
  assign new_n3632_ = ~new_n3630_ & ~new_n3631_;
  assign new_n3633_ = ~new_n2746_ & ~new_n3632_;
  assign new_n3634_ = ~\p_input[166]  & new_n2746_;
  assign new_n3635_ = ~new_n3633_ & ~new_n3634_;
  assign new_n3636_ = new_n2792_ & new_n3635_;
  assign new_n3637_ = ~new_n3629_ & ~new_n3636_;
  assign new_n3638_ = ~new_n2890_ & ~new_n3637_;
  assign new_n3639_ = new_n2792_ & ~new_n3628_;
  assign new_n3640_ = ~new_n2792_ & new_n3635_;
  assign new_n3641_ = ~new_n3639_ & ~new_n3640_;
  assign new_n3642_ = ~new_n2844_ & ~new_n3641_;
  assign new_n3643_ = \p_input[134]  & new_n2844_;
  assign new_n3644_ = ~new_n3642_ & ~new_n3643_;
  assign new_n3645_ = new_n2890_ & ~new_n3644_;
  assign new_n3646_ = ~new_n3638_ & ~new_n3645_;
  assign new_n3647_ = ~new_n2989_ & ~new_n3646_;
  assign new_n3648_ = new_n2890_ & ~new_n3637_;
  assign new_n3649_ = ~new_n2890_ & ~new_n3644_;
  assign new_n3650_ = ~new_n3648_ & ~new_n3649_;
  assign new_n3651_ = ~new_n2942_ & ~new_n3650_;
  assign new_n3652_ = \p_input[102]  & new_n2942_;
  assign new_n3653_ = ~new_n3651_ & ~new_n3652_;
  assign new_n3654_ = new_n2989_ & ~new_n3653_;
  assign new_n3655_ = ~new_n3647_ & ~new_n3654_;
  assign new_n3656_ = ~new_n3087_ & ~new_n3655_;
  assign new_n3657_ = new_n2989_ & ~new_n3646_;
  assign new_n3658_ = ~new_n2989_ & ~new_n3653_;
  assign new_n3659_ = ~new_n3657_ & ~new_n3658_;
  assign new_n3660_ = ~new_n3041_ & ~new_n3659_;
  assign new_n3661_ = \p_input[70]  & new_n3041_;
  assign new_n3662_ = ~new_n3660_ & ~new_n3661_;
  assign new_n3663_ = new_n3087_ & ~new_n3662_;
  assign new_n3664_ = ~new_n3656_ & ~new_n3663_;
  assign new_n3665_ = ~new_n3185_ & ~new_n3664_;
  assign new_n3666_ = new_n3087_ & ~new_n3655_;
  assign new_n3667_ = ~new_n3087_ & ~new_n3662_;
  assign new_n3668_ = ~new_n3666_ & ~new_n3667_;
  assign new_n3669_ = ~new_n3139_ & ~new_n3668_;
  assign new_n3670_ = \p_input[38]  & new_n3139_;
  assign new_n3671_ = ~new_n3669_ & ~new_n3670_;
  assign new_n3672_ = new_n3185_ & ~new_n3671_;
  assign new_n3673_ = ~new_n3665_ & ~new_n3672_;
  assign new_n3674_ = new_n3283_ & ~new_n3673_;
  assign new_n3675_ = new_n3185_ & ~new_n3664_;
  assign new_n3676_ = ~new_n3185_ & ~new_n3671_;
  assign new_n3677_ = ~new_n3675_ & ~new_n3676_;
  assign new_n3678_ = ~new_n3237_ & ~new_n3677_;
  assign new_n3679_ = \p_input[6]  & new_n3237_;
  assign new_n3680_ = ~new_n3678_ & ~new_n3679_;
  assign new_n3681_ = ~new_n3283_ & ~new_n3680_;
  assign \o[6]  = new_n3674_ | new_n3681_;
  assign new_n3683_ = \p_input[199]  & ~new_n2694_;
  assign new_n3684_ = \p_input[231]  & new_n2694_;
  assign new_n3685_ = ~new_n3683_ & ~new_n3684_;
  assign new_n3686_ = ~new_n2792_ & ~new_n3685_;
  assign new_n3687_ = ~\p_input[231]  & ~new_n2694_;
  assign new_n3688_ = ~\p_input[199]  & new_n2694_;
  assign new_n3689_ = ~new_n3687_ & ~new_n3688_;
  assign new_n3690_ = ~new_n2746_ & ~new_n3689_;
  assign new_n3691_ = ~\p_input[167]  & new_n2746_;
  assign new_n3692_ = ~new_n3690_ & ~new_n3691_;
  assign new_n3693_ = new_n2792_ & new_n3692_;
  assign new_n3694_ = ~new_n3686_ & ~new_n3693_;
  assign new_n3695_ = ~new_n2890_ & ~new_n3694_;
  assign new_n3696_ = new_n2792_ & ~new_n3685_;
  assign new_n3697_ = ~new_n2792_ & new_n3692_;
  assign new_n3698_ = ~new_n3696_ & ~new_n3697_;
  assign new_n3699_ = ~new_n2844_ & ~new_n3698_;
  assign new_n3700_ = \p_input[135]  & new_n2844_;
  assign new_n3701_ = ~new_n3699_ & ~new_n3700_;
  assign new_n3702_ = new_n2890_ & ~new_n3701_;
  assign new_n3703_ = ~new_n3695_ & ~new_n3702_;
  assign new_n3704_ = ~new_n2989_ & ~new_n3703_;
  assign new_n3705_ = new_n2890_ & ~new_n3694_;
  assign new_n3706_ = ~new_n2890_ & ~new_n3701_;
  assign new_n3707_ = ~new_n3705_ & ~new_n3706_;
  assign new_n3708_ = ~new_n2942_ & ~new_n3707_;
  assign new_n3709_ = \p_input[103]  & new_n2942_;
  assign new_n3710_ = ~new_n3708_ & ~new_n3709_;
  assign new_n3711_ = new_n2989_ & ~new_n3710_;
  assign new_n3712_ = ~new_n3704_ & ~new_n3711_;
  assign new_n3713_ = ~new_n3087_ & ~new_n3712_;
  assign new_n3714_ = new_n2989_ & ~new_n3703_;
  assign new_n3715_ = ~new_n2989_ & ~new_n3710_;
  assign new_n3716_ = ~new_n3714_ & ~new_n3715_;
  assign new_n3717_ = ~new_n3041_ & ~new_n3716_;
  assign new_n3718_ = \p_input[71]  & new_n3041_;
  assign new_n3719_ = ~new_n3717_ & ~new_n3718_;
  assign new_n3720_ = new_n3087_ & ~new_n3719_;
  assign new_n3721_ = ~new_n3713_ & ~new_n3720_;
  assign new_n3722_ = ~new_n3185_ & ~new_n3721_;
  assign new_n3723_ = new_n3087_ & ~new_n3712_;
  assign new_n3724_ = ~new_n3087_ & ~new_n3719_;
  assign new_n3725_ = ~new_n3723_ & ~new_n3724_;
  assign new_n3726_ = ~new_n3139_ & ~new_n3725_;
  assign new_n3727_ = \p_input[39]  & new_n3139_;
  assign new_n3728_ = ~new_n3726_ & ~new_n3727_;
  assign new_n3729_ = new_n3185_ & ~new_n3728_;
  assign new_n3730_ = ~new_n3722_ & ~new_n3729_;
  assign new_n3731_ = new_n3283_ & ~new_n3730_;
  assign new_n3732_ = new_n3185_ & ~new_n3721_;
  assign new_n3733_ = ~new_n3185_ & ~new_n3728_;
  assign new_n3734_ = ~new_n3732_ & ~new_n3733_;
  assign new_n3735_ = ~new_n3237_ & ~new_n3734_;
  assign new_n3736_ = \p_input[7]  & new_n3237_;
  assign new_n3737_ = ~new_n3735_ & ~new_n3736_;
  assign new_n3738_ = ~new_n3283_ & ~new_n3737_;
  assign \o[7]  = new_n3731_ | new_n3738_;
  assign new_n3740_ = \p_input[200]  & ~new_n2694_;
  assign new_n3741_ = \p_input[232]  & new_n2694_;
  assign new_n3742_ = ~new_n3740_ & ~new_n3741_;
  assign new_n3743_ = ~new_n2792_ & ~new_n3742_;
  assign new_n3744_ = ~\p_input[232]  & ~new_n2694_;
  assign new_n3745_ = ~\p_input[200]  & new_n2694_;
  assign new_n3746_ = ~new_n3744_ & ~new_n3745_;
  assign new_n3747_ = ~new_n2746_ & ~new_n3746_;
  assign new_n3748_ = ~\p_input[168]  & new_n2746_;
  assign new_n3749_ = ~new_n3747_ & ~new_n3748_;
  assign new_n3750_ = new_n2792_ & new_n3749_;
  assign new_n3751_ = ~new_n3743_ & ~new_n3750_;
  assign new_n3752_ = ~new_n2890_ & ~new_n3751_;
  assign new_n3753_ = new_n2792_ & ~new_n3742_;
  assign new_n3754_ = ~new_n2792_ & new_n3749_;
  assign new_n3755_ = ~new_n3753_ & ~new_n3754_;
  assign new_n3756_ = ~new_n2844_ & ~new_n3755_;
  assign new_n3757_ = \p_input[136]  & new_n2844_;
  assign new_n3758_ = ~new_n3756_ & ~new_n3757_;
  assign new_n3759_ = new_n2890_ & ~new_n3758_;
  assign new_n3760_ = ~new_n3752_ & ~new_n3759_;
  assign new_n3761_ = ~new_n2989_ & ~new_n3760_;
  assign new_n3762_ = new_n2890_ & ~new_n3751_;
  assign new_n3763_ = ~new_n2890_ & ~new_n3758_;
  assign new_n3764_ = ~new_n3762_ & ~new_n3763_;
  assign new_n3765_ = ~new_n2942_ & ~new_n3764_;
  assign new_n3766_ = \p_input[104]  & new_n2942_;
  assign new_n3767_ = ~new_n3765_ & ~new_n3766_;
  assign new_n3768_ = new_n2989_ & ~new_n3767_;
  assign new_n3769_ = ~new_n3761_ & ~new_n3768_;
  assign new_n3770_ = ~new_n3087_ & ~new_n3769_;
  assign new_n3771_ = new_n2989_ & ~new_n3760_;
  assign new_n3772_ = ~new_n2989_ & ~new_n3767_;
  assign new_n3773_ = ~new_n3771_ & ~new_n3772_;
  assign new_n3774_ = ~new_n3041_ & ~new_n3773_;
  assign new_n3775_ = \p_input[72]  & new_n3041_;
  assign new_n3776_ = ~new_n3774_ & ~new_n3775_;
  assign new_n3777_ = new_n3087_ & ~new_n3776_;
  assign new_n3778_ = ~new_n3770_ & ~new_n3777_;
  assign new_n3779_ = ~new_n3185_ & ~new_n3778_;
  assign new_n3780_ = new_n3087_ & ~new_n3769_;
  assign new_n3781_ = ~new_n3087_ & ~new_n3776_;
  assign new_n3782_ = ~new_n3780_ & ~new_n3781_;
  assign new_n3783_ = ~new_n3139_ & ~new_n3782_;
  assign new_n3784_ = \p_input[40]  & new_n3139_;
  assign new_n3785_ = ~new_n3783_ & ~new_n3784_;
  assign new_n3786_ = new_n3185_ & ~new_n3785_;
  assign new_n3787_ = ~new_n3779_ & ~new_n3786_;
  assign new_n3788_ = new_n3283_ & ~new_n3787_;
  assign new_n3789_ = new_n3185_ & ~new_n3778_;
  assign new_n3790_ = ~new_n3185_ & ~new_n3785_;
  assign new_n3791_ = ~new_n3789_ & ~new_n3790_;
  assign new_n3792_ = ~new_n3237_ & ~new_n3791_;
  assign new_n3793_ = \p_input[8]  & new_n3237_;
  assign new_n3794_ = ~new_n3792_ & ~new_n3793_;
  assign new_n3795_ = ~new_n3283_ & ~new_n3794_;
  assign \o[8]  = new_n3788_ | new_n3795_;
  assign new_n3797_ = \p_input[201]  & ~new_n2694_;
  assign new_n3798_ = \p_input[233]  & new_n2694_;
  assign new_n3799_ = ~new_n3797_ & ~new_n3798_;
  assign new_n3800_ = ~new_n2792_ & ~new_n3799_;
  assign new_n3801_ = ~\p_input[233]  & ~new_n2694_;
  assign new_n3802_ = ~\p_input[201]  & new_n2694_;
  assign new_n3803_ = ~new_n3801_ & ~new_n3802_;
  assign new_n3804_ = ~new_n2746_ & ~new_n3803_;
  assign new_n3805_ = ~\p_input[169]  & new_n2746_;
  assign new_n3806_ = ~new_n3804_ & ~new_n3805_;
  assign new_n3807_ = new_n2792_ & new_n3806_;
  assign new_n3808_ = ~new_n3800_ & ~new_n3807_;
  assign new_n3809_ = ~new_n2890_ & ~new_n3808_;
  assign new_n3810_ = new_n2792_ & ~new_n3799_;
  assign new_n3811_ = ~new_n2792_ & new_n3806_;
  assign new_n3812_ = ~new_n3810_ & ~new_n3811_;
  assign new_n3813_ = ~new_n2844_ & ~new_n3812_;
  assign new_n3814_ = \p_input[137]  & new_n2844_;
  assign new_n3815_ = ~new_n3813_ & ~new_n3814_;
  assign new_n3816_ = new_n2890_ & ~new_n3815_;
  assign new_n3817_ = ~new_n3809_ & ~new_n3816_;
  assign new_n3818_ = ~new_n2989_ & ~new_n3817_;
  assign new_n3819_ = new_n2890_ & ~new_n3808_;
  assign new_n3820_ = ~new_n2890_ & ~new_n3815_;
  assign new_n3821_ = ~new_n3819_ & ~new_n3820_;
  assign new_n3822_ = ~new_n2942_ & ~new_n3821_;
  assign new_n3823_ = \p_input[105]  & new_n2942_;
  assign new_n3824_ = ~new_n3822_ & ~new_n3823_;
  assign new_n3825_ = new_n2989_ & ~new_n3824_;
  assign new_n3826_ = ~new_n3818_ & ~new_n3825_;
  assign new_n3827_ = ~new_n3087_ & ~new_n3826_;
  assign new_n3828_ = new_n2989_ & ~new_n3817_;
  assign new_n3829_ = ~new_n2989_ & ~new_n3824_;
  assign new_n3830_ = ~new_n3828_ & ~new_n3829_;
  assign new_n3831_ = ~new_n3041_ & ~new_n3830_;
  assign new_n3832_ = \p_input[73]  & new_n3041_;
  assign new_n3833_ = ~new_n3831_ & ~new_n3832_;
  assign new_n3834_ = new_n3087_ & ~new_n3833_;
  assign new_n3835_ = ~new_n3827_ & ~new_n3834_;
  assign new_n3836_ = ~new_n3185_ & ~new_n3835_;
  assign new_n3837_ = new_n3087_ & ~new_n3826_;
  assign new_n3838_ = ~new_n3087_ & ~new_n3833_;
  assign new_n3839_ = ~new_n3837_ & ~new_n3838_;
  assign new_n3840_ = ~new_n3139_ & ~new_n3839_;
  assign new_n3841_ = \p_input[41]  & new_n3139_;
  assign new_n3842_ = ~new_n3840_ & ~new_n3841_;
  assign new_n3843_ = new_n3185_ & ~new_n3842_;
  assign new_n3844_ = ~new_n3836_ & ~new_n3843_;
  assign new_n3845_ = new_n3283_ & ~new_n3844_;
  assign new_n3846_ = new_n3185_ & ~new_n3835_;
  assign new_n3847_ = ~new_n3185_ & ~new_n3842_;
  assign new_n3848_ = ~new_n3846_ & ~new_n3847_;
  assign new_n3849_ = ~new_n3237_ & ~new_n3848_;
  assign new_n3850_ = \p_input[9]  & new_n3237_;
  assign new_n3851_ = ~new_n3849_ & ~new_n3850_;
  assign new_n3852_ = ~new_n3283_ & ~new_n3851_;
  assign \o[9]  = new_n3845_ | new_n3852_;
  assign new_n3854_ = \p_input[202]  & ~new_n2694_;
  assign new_n3855_ = \p_input[234]  & new_n2694_;
  assign new_n3856_ = ~new_n3854_ & ~new_n3855_;
  assign new_n3857_ = ~new_n2792_ & ~new_n3856_;
  assign new_n3858_ = ~\p_input[234]  & ~new_n2694_;
  assign new_n3859_ = ~\p_input[202]  & new_n2694_;
  assign new_n3860_ = ~new_n3858_ & ~new_n3859_;
  assign new_n3861_ = ~new_n2746_ & ~new_n3860_;
  assign new_n3862_ = ~\p_input[170]  & new_n2746_;
  assign new_n3863_ = ~new_n3861_ & ~new_n3862_;
  assign new_n3864_ = new_n2792_ & new_n3863_;
  assign new_n3865_ = ~new_n3857_ & ~new_n3864_;
  assign new_n3866_ = ~new_n2890_ & ~new_n3865_;
  assign new_n3867_ = new_n2792_ & ~new_n3856_;
  assign new_n3868_ = ~new_n2792_ & new_n3863_;
  assign new_n3869_ = ~new_n3867_ & ~new_n3868_;
  assign new_n3870_ = ~new_n2844_ & ~new_n3869_;
  assign new_n3871_ = \p_input[138]  & new_n2844_;
  assign new_n3872_ = ~new_n3870_ & ~new_n3871_;
  assign new_n3873_ = new_n2890_ & ~new_n3872_;
  assign new_n3874_ = ~new_n3866_ & ~new_n3873_;
  assign new_n3875_ = ~new_n2989_ & ~new_n3874_;
  assign new_n3876_ = new_n2890_ & ~new_n3865_;
  assign new_n3877_ = ~new_n2890_ & ~new_n3872_;
  assign new_n3878_ = ~new_n3876_ & ~new_n3877_;
  assign new_n3879_ = ~new_n2942_ & ~new_n3878_;
  assign new_n3880_ = \p_input[106]  & new_n2942_;
  assign new_n3881_ = ~new_n3879_ & ~new_n3880_;
  assign new_n3882_ = new_n2989_ & ~new_n3881_;
  assign new_n3883_ = ~new_n3875_ & ~new_n3882_;
  assign new_n3884_ = ~new_n3087_ & ~new_n3883_;
  assign new_n3885_ = new_n2989_ & ~new_n3874_;
  assign new_n3886_ = ~new_n2989_ & ~new_n3881_;
  assign new_n3887_ = ~new_n3885_ & ~new_n3886_;
  assign new_n3888_ = ~new_n3041_ & ~new_n3887_;
  assign new_n3889_ = \p_input[74]  & new_n3041_;
  assign new_n3890_ = ~new_n3888_ & ~new_n3889_;
  assign new_n3891_ = new_n3087_ & ~new_n3890_;
  assign new_n3892_ = ~new_n3884_ & ~new_n3891_;
  assign new_n3893_ = ~new_n3185_ & ~new_n3892_;
  assign new_n3894_ = new_n3087_ & ~new_n3883_;
  assign new_n3895_ = ~new_n3087_ & ~new_n3890_;
  assign new_n3896_ = ~new_n3894_ & ~new_n3895_;
  assign new_n3897_ = ~new_n3139_ & ~new_n3896_;
  assign new_n3898_ = \p_input[42]  & new_n3139_;
  assign new_n3899_ = ~new_n3897_ & ~new_n3898_;
  assign new_n3900_ = new_n3185_ & ~new_n3899_;
  assign new_n3901_ = ~new_n3893_ & ~new_n3900_;
  assign new_n3902_ = new_n3283_ & ~new_n3901_;
  assign new_n3903_ = new_n3185_ & ~new_n3892_;
  assign new_n3904_ = ~new_n3185_ & ~new_n3899_;
  assign new_n3905_ = ~new_n3903_ & ~new_n3904_;
  assign new_n3906_ = ~new_n3237_ & ~new_n3905_;
  assign new_n3907_ = \p_input[10]  & new_n3237_;
  assign new_n3908_ = ~new_n3906_ & ~new_n3907_;
  assign new_n3909_ = ~new_n3283_ & ~new_n3908_;
  assign \o[10]  = new_n3902_ | new_n3909_;
  assign new_n3911_ = \p_input[203]  & ~new_n2694_;
  assign new_n3912_ = \p_input[235]  & new_n2694_;
  assign new_n3913_ = ~new_n3911_ & ~new_n3912_;
  assign new_n3914_ = ~new_n2792_ & ~new_n3913_;
  assign new_n3915_ = ~\p_input[235]  & ~new_n2694_;
  assign new_n3916_ = ~\p_input[203]  & new_n2694_;
  assign new_n3917_ = ~new_n3915_ & ~new_n3916_;
  assign new_n3918_ = ~new_n2746_ & ~new_n3917_;
  assign new_n3919_ = ~\p_input[171]  & new_n2746_;
  assign new_n3920_ = ~new_n3918_ & ~new_n3919_;
  assign new_n3921_ = new_n2792_ & new_n3920_;
  assign new_n3922_ = ~new_n3914_ & ~new_n3921_;
  assign new_n3923_ = ~new_n2890_ & ~new_n3922_;
  assign new_n3924_ = new_n2792_ & ~new_n3913_;
  assign new_n3925_ = ~new_n2792_ & new_n3920_;
  assign new_n3926_ = ~new_n3924_ & ~new_n3925_;
  assign new_n3927_ = ~new_n2844_ & ~new_n3926_;
  assign new_n3928_ = \p_input[139]  & new_n2844_;
  assign new_n3929_ = ~new_n3927_ & ~new_n3928_;
  assign new_n3930_ = new_n2890_ & ~new_n3929_;
  assign new_n3931_ = ~new_n3923_ & ~new_n3930_;
  assign new_n3932_ = ~new_n2989_ & ~new_n3931_;
  assign new_n3933_ = new_n2890_ & ~new_n3922_;
  assign new_n3934_ = ~new_n2890_ & ~new_n3929_;
  assign new_n3935_ = ~new_n3933_ & ~new_n3934_;
  assign new_n3936_ = ~new_n2942_ & ~new_n3935_;
  assign new_n3937_ = \p_input[107]  & new_n2942_;
  assign new_n3938_ = ~new_n3936_ & ~new_n3937_;
  assign new_n3939_ = new_n2989_ & ~new_n3938_;
  assign new_n3940_ = ~new_n3932_ & ~new_n3939_;
  assign new_n3941_ = ~new_n3087_ & ~new_n3940_;
  assign new_n3942_ = new_n2989_ & ~new_n3931_;
  assign new_n3943_ = ~new_n2989_ & ~new_n3938_;
  assign new_n3944_ = ~new_n3942_ & ~new_n3943_;
  assign new_n3945_ = ~new_n3041_ & ~new_n3944_;
  assign new_n3946_ = \p_input[75]  & new_n3041_;
  assign new_n3947_ = ~new_n3945_ & ~new_n3946_;
  assign new_n3948_ = new_n3087_ & ~new_n3947_;
  assign new_n3949_ = ~new_n3941_ & ~new_n3948_;
  assign new_n3950_ = ~new_n3185_ & ~new_n3949_;
  assign new_n3951_ = new_n3087_ & ~new_n3940_;
  assign new_n3952_ = ~new_n3087_ & ~new_n3947_;
  assign new_n3953_ = ~new_n3951_ & ~new_n3952_;
  assign new_n3954_ = ~new_n3139_ & ~new_n3953_;
  assign new_n3955_ = \p_input[43]  & new_n3139_;
  assign new_n3956_ = ~new_n3954_ & ~new_n3955_;
  assign new_n3957_ = new_n3185_ & ~new_n3956_;
  assign new_n3958_ = ~new_n3950_ & ~new_n3957_;
  assign new_n3959_ = new_n3283_ & ~new_n3958_;
  assign new_n3960_ = new_n3185_ & ~new_n3949_;
  assign new_n3961_ = ~new_n3185_ & ~new_n3956_;
  assign new_n3962_ = ~new_n3960_ & ~new_n3961_;
  assign new_n3963_ = ~new_n3237_ & ~new_n3962_;
  assign new_n3964_ = \p_input[11]  & new_n3237_;
  assign new_n3965_ = ~new_n3963_ & ~new_n3964_;
  assign new_n3966_ = ~new_n3283_ & ~new_n3965_;
  assign \o[11]  = new_n3959_ | new_n3966_;
  assign new_n3968_ = \p_input[204]  & ~new_n2694_;
  assign new_n3969_ = \p_input[236]  & new_n2694_;
  assign new_n3970_ = ~new_n3968_ & ~new_n3969_;
  assign new_n3971_ = ~new_n2792_ & ~new_n3970_;
  assign new_n3972_ = ~\p_input[236]  & ~new_n2694_;
  assign new_n3973_ = ~\p_input[204]  & new_n2694_;
  assign new_n3974_ = ~new_n3972_ & ~new_n3973_;
  assign new_n3975_ = ~new_n2746_ & ~new_n3974_;
  assign new_n3976_ = ~\p_input[172]  & new_n2746_;
  assign new_n3977_ = ~new_n3975_ & ~new_n3976_;
  assign new_n3978_ = new_n2792_ & new_n3977_;
  assign new_n3979_ = ~new_n3971_ & ~new_n3978_;
  assign new_n3980_ = ~new_n2890_ & ~new_n3979_;
  assign new_n3981_ = new_n2792_ & ~new_n3970_;
  assign new_n3982_ = ~new_n2792_ & new_n3977_;
  assign new_n3983_ = ~new_n3981_ & ~new_n3982_;
  assign new_n3984_ = ~new_n2844_ & ~new_n3983_;
  assign new_n3985_ = \p_input[140]  & new_n2844_;
  assign new_n3986_ = ~new_n3984_ & ~new_n3985_;
  assign new_n3987_ = new_n2890_ & ~new_n3986_;
  assign new_n3988_ = ~new_n3980_ & ~new_n3987_;
  assign new_n3989_ = ~new_n2989_ & ~new_n3988_;
  assign new_n3990_ = new_n2890_ & ~new_n3979_;
  assign new_n3991_ = ~new_n2890_ & ~new_n3986_;
  assign new_n3992_ = ~new_n3990_ & ~new_n3991_;
  assign new_n3993_ = ~new_n2942_ & ~new_n3992_;
  assign new_n3994_ = \p_input[108]  & new_n2942_;
  assign new_n3995_ = ~new_n3993_ & ~new_n3994_;
  assign new_n3996_ = new_n2989_ & ~new_n3995_;
  assign new_n3997_ = ~new_n3989_ & ~new_n3996_;
  assign new_n3998_ = ~new_n3087_ & ~new_n3997_;
  assign new_n3999_ = new_n2989_ & ~new_n3988_;
  assign new_n4000_ = ~new_n2989_ & ~new_n3995_;
  assign new_n4001_ = ~new_n3999_ & ~new_n4000_;
  assign new_n4002_ = ~new_n3041_ & ~new_n4001_;
  assign new_n4003_ = \p_input[76]  & new_n3041_;
  assign new_n4004_ = ~new_n4002_ & ~new_n4003_;
  assign new_n4005_ = new_n3087_ & ~new_n4004_;
  assign new_n4006_ = ~new_n3998_ & ~new_n4005_;
  assign new_n4007_ = ~new_n3185_ & ~new_n4006_;
  assign new_n4008_ = new_n3087_ & ~new_n3997_;
  assign new_n4009_ = ~new_n3087_ & ~new_n4004_;
  assign new_n4010_ = ~new_n4008_ & ~new_n4009_;
  assign new_n4011_ = ~new_n3139_ & ~new_n4010_;
  assign new_n4012_ = \p_input[44]  & new_n3139_;
  assign new_n4013_ = ~new_n4011_ & ~new_n4012_;
  assign new_n4014_ = new_n3185_ & ~new_n4013_;
  assign new_n4015_ = ~new_n4007_ & ~new_n4014_;
  assign new_n4016_ = new_n3283_ & ~new_n4015_;
  assign new_n4017_ = new_n3185_ & ~new_n4006_;
  assign new_n4018_ = ~new_n3185_ & ~new_n4013_;
  assign new_n4019_ = ~new_n4017_ & ~new_n4018_;
  assign new_n4020_ = ~new_n3237_ & ~new_n4019_;
  assign new_n4021_ = \p_input[12]  & new_n3237_;
  assign new_n4022_ = ~new_n4020_ & ~new_n4021_;
  assign new_n4023_ = ~new_n3283_ & ~new_n4022_;
  assign \o[12]  = new_n4016_ | new_n4023_;
  assign new_n4025_ = \p_input[205]  & ~new_n2694_;
  assign new_n4026_ = \p_input[237]  & new_n2694_;
  assign new_n4027_ = ~new_n4025_ & ~new_n4026_;
  assign new_n4028_ = ~new_n2792_ & ~new_n4027_;
  assign new_n4029_ = ~\p_input[237]  & ~new_n2694_;
  assign new_n4030_ = ~\p_input[205]  & new_n2694_;
  assign new_n4031_ = ~new_n4029_ & ~new_n4030_;
  assign new_n4032_ = ~new_n2746_ & ~new_n4031_;
  assign new_n4033_ = ~\p_input[173]  & new_n2746_;
  assign new_n4034_ = ~new_n4032_ & ~new_n4033_;
  assign new_n4035_ = new_n2792_ & new_n4034_;
  assign new_n4036_ = ~new_n4028_ & ~new_n4035_;
  assign new_n4037_ = ~new_n2890_ & ~new_n4036_;
  assign new_n4038_ = new_n2792_ & ~new_n4027_;
  assign new_n4039_ = ~new_n2792_ & new_n4034_;
  assign new_n4040_ = ~new_n4038_ & ~new_n4039_;
  assign new_n4041_ = ~new_n2844_ & ~new_n4040_;
  assign new_n4042_ = \p_input[141]  & new_n2844_;
  assign new_n4043_ = ~new_n4041_ & ~new_n4042_;
  assign new_n4044_ = new_n2890_ & ~new_n4043_;
  assign new_n4045_ = ~new_n4037_ & ~new_n4044_;
  assign new_n4046_ = ~new_n2989_ & ~new_n4045_;
  assign new_n4047_ = new_n2890_ & ~new_n4036_;
  assign new_n4048_ = ~new_n2890_ & ~new_n4043_;
  assign new_n4049_ = ~new_n4047_ & ~new_n4048_;
  assign new_n4050_ = ~new_n2942_ & ~new_n4049_;
  assign new_n4051_ = \p_input[109]  & new_n2942_;
  assign new_n4052_ = ~new_n4050_ & ~new_n4051_;
  assign new_n4053_ = new_n2989_ & ~new_n4052_;
  assign new_n4054_ = ~new_n4046_ & ~new_n4053_;
  assign new_n4055_ = ~new_n3087_ & ~new_n4054_;
  assign new_n4056_ = new_n2989_ & ~new_n4045_;
  assign new_n4057_ = ~new_n2989_ & ~new_n4052_;
  assign new_n4058_ = ~new_n4056_ & ~new_n4057_;
  assign new_n4059_ = ~new_n3041_ & ~new_n4058_;
  assign new_n4060_ = \p_input[77]  & new_n3041_;
  assign new_n4061_ = ~new_n4059_ & ~new_n4060_;
  assign new_n4062_ = new_n3087_ & ~new_n4061_;
  assign new_n4063_ = ~new_n4055_ & ~new_n4062_;
  assign new_n4064_ = ~new_n3185_ & ~new_n4063_;
  assign new_n4065_ = new_n3087_ & ~new_n4054_;
  assign new_n4066_ = ~new_n3087_ & ~new_n4061_;
  assign new_n4067_ = ~new_n4065_ & ~new_n4066_;
  assign new_n4068_ = ~new_n3139_ & ~new_n4067_;
  assign new_n4069_ = \p_input[45]  & new_n3139_;
  assign new_n4070_ = ~new_n4068_ & ~new_n4069_;
  assign new_n4071_ = new_n3185_ & ~new_n4070_;
  assign new_n4072_ = ~new_n4064_ & ~new_n4071_;
  assign new_n4073_ = new_n3283_ & ~new_n4072_;
  assign new_n4074_ = new_n3185_ & ~new_n4063_;
  assign new_n4075_ = ~new_n3185_ & ~new_n4070_;
  assign new_n4076_ = ~new_n4074_ & ~new_n4075_;
  assign new_n4077_ = ~new_n3237_ & ~new_n4076_;
  assign new_n4078_ = \p_input[13]  & new_n3237_;
  assign new_n4079_ = ~new_n4077_ & ~new_n4078_;
  assign new_n4080_ = ~new_n3283_ & ~new_n4079_;
  assign \o[13]  = new_n4073_ | new_n4080_;
  assign new_n4082_ = \p_input[206]  & ~new_n2694_;
  assign new_n4083_ = \p_input[238]  & new_n2694_;
  assign new_n4084_ = ~new_n4082_ & ~new_n4083_;
  assign new_n4085_ = ~new_n2792_ & ~new_n4084_;
  assign new_n4086_ = ~\p_input[238]  & ~new_n2694_;
  assign new_n4087_ = ~\p_input[206]  & new_n2694_;
  assign new_n4088_ = ~new_n4086_ & ~new_n4087_;
  assign new_n4089_ = ~new_n2746_ & ~new_n4088_;
  assign new_n4090_ = ~\p_input[174]  & new_n2746_;
  assign new_n4091_ = ~new_n4089_ & ~new_n4090_;
  assign new_n4092_ = new_n2792_ & new_n4091_;
  assign new_n4093_ = ~new_n4085_ & ~new_n4092_;
  assign new_n4094_ = ~new_n2890_ & ~new_n4093_;
  assign new_n4095_ = new_n2792_ & ~new_n4084_;
  assign new_n4096_ = ~new_n2792_ & new_n4091_;
  assign new_n4097_ = ~new_n4095_ & ~new_n4096_;
  assign new_n4098_ = ~new_n2844_ & ~new_n4097_;
  assign new_n4099_ = \p_input[142]  & new_n2844_;
  assign new_n4100_ = ~new_n4098_ & ~new_n4099_;
  assign new_n4101_ = new_n2890_ & ~new_n4100_;
  assign new_n4102_ = ~new_n4094_ & ~new_n4101_;
  assign new_n4103_ = ~new_n2989_ & ~new_n4102_;
  assign new_n4104_ = new_n2890_ & ~new_n4093_;
  assign new_n4105_ = ~new_n2890_ & ~new_n4100_;
  assign new_n4106_ = ~new_n4104_ & ~new_n4105_;
  assign new_n4107_ = ~new_n2942_ & ~new_n4106_;
  assign new_n4108_ = \p_input[110]  & new_n2942_;
  assign new_n4109_ = ~new_n4107_ & ~new_n4108_;
  assign new_n4110_ = new_n2989_ & ~new_n4109_;
  assign new_n4111_ = ~new_n4103_ & ~new_n4110_;
  assign new_n4112_ = ~new_n3087_ & ~new_n4111_;
  assign new_n4113_ = new_n2989_ & ~new_n4102_;
  assign new_n4114_ = ~new_n2989_ & ~new_n4109_;
  assign new_n4115_ = ~new_n4113_ & ~new_n4114_;
  assign new_n4116_ = ~new_n3041_ & ~new_n4115_;
  assign new_n4117_ = \p_input[78]  & new_n3041_;
  assign new_n4118_ = ~new_n4116_ & ~new_n4117_;
  assign new_n4119_ = new_n3087_ & ~new_n4118_;
  assign new_n4120_ = ~new_n4112_ & ~new_n4119_;
  assign new_n4121_ = ~new_n3185_ & ~new_n4120_;
  assign new_n4122_ = new_n3087_ & ~new_n4111_;
  assign new_n4123_ = ~new_n3087_ & ~new_n4118_;
  assign new_n4124_ = ~new_n4122_ & ~new_n4123_;
  assign new_n4125_ = ~new_n3139_ & ~new_n4124_;
  assign new_n4126_ = \p_input[46]  & new_n3139_;
  assign new_n4127_ = ~new_n4125_ & ~new_n4126_;
  assign new_n4128_ = new_n3185_ & ~new_n4127_;
  assign new_n4129_ = ~new_n4121_ & ~new_n4128_;
  assign new_n4130_ = new_n3283_ & ~new_n4129_;
  assign new_n4131_ = new_n3185_ & ~new_n4120_;
  assign new_n4132_ = ~new_n3185_ & ~new_n4127_;
  assign new_n4133_ = ~new_n4131_ & ~new_n4132_;
  assign new_n4134_ = ~new_n3237_ & ~new_n4133_;
  assign new_n4135_ = \p_input[14]  & new_n3237_;
  assign new_n4136_ = ~new_n4134_ & ~new_n4135_;
  assign new_n4137_ = ~new_n3283_ & ~new_n4136_;
  assign \o[14]  = new_n4130_ | new_n4137_;
  assign new_n4139_ = \p_input[207]  & ~new_n2694_;
  assign new_n4140_ = \p_input[239]  & new_n2694_;
  assign new_n4141_ = ~new_n4139_ & ~new_n4140_;
  assign new_n4142_ = ~new_n2792_ & ~new_n4141_;
  assign new_n4143_ = ~\p_input[239]  & ~new_n2694_;
  assign new_n4144_ = ~\p_input[207]  & new_n2694_;
  assign new_n4145_ = ~new_n4143_ & ~new_n4144_;
  assign new_n4146_ = ~new_n2746_ & ~new_n4145_;
  assign new_n4147_ = ~\p_input[175]  & new_n2746_;
  assign new_n4148_ = ~new_n4146_ & ~new_n4147_;
  assign new_n4149_ = new_n2792_ & new_n4148_;
  assign new_n4150_ = ~new_n4142_ & ~new_n4149_;
  assign new_n4151_ = ~new_n2890_ & ~new_n4150_;
  assign new_n4152_ = new_n2792_ & ~new_n4141_;
  assign new_n4153_ = ~new_n2792_ & new_n4148_;
  assign new_n4154_ = ~new_n4152_ & ~new_n4153_;
  assign new_n4155_ = ~new_n2844_ & ~new_n4154_;
  assign new_n4156_ = \p_input[143]  & new_n2844_;
  assign new_n4157_ = ~new_n4155_ & ~new_n4156_;
  assign new_n4158_ = new_n2890_ & ~new_n4157_;
  assign new_n4159_ = ~new_n4151_ & ~new_n4158_;
  assign new_n4160_ = ~new_n2989_ & ~new_n4159_;
  assign new_n4161_ = new_n2890_ & ~new_n4150_;
  assign new_n4162_ = ~new_n2890_ & ~new_n4157_;
  assign new_n4163_ = ~new_n4161_ & ~new_n4162_;
  assign new_n4164_ = ~new_n2942_ & ~new_n4163_;
  assign new_n4165_ = \p_input[111]  & new_n2942_;
  assign new_n4166_ = ~new_n4164_ & ~new_n4165_;
  assign new_n4167_ = new_n2989_ & ~new_n4166_;
  assign new_n4168_ = ~new_n4160_ & ~new_n4167_;
  assign new_n4169_ = ~new_n3087_ & ~new_n4168_;
  assign new_n4170_ = new_n2989_ & ~new_n4159_;
  assign new_n4171_ = ~new_n2989_ & ~new_n4166_;
  assign new_n4172_ = ~new_n4170_ & ~new_n4171_;
  assign new_n4173_ = ~new_n3041_ & ~new_n4172_;
  assign new_n4174_ = \p_input[79]  & new_n3041_;
  assign new_n4175_ = ~new_n4173_ & ~new_n4174_;
  assign new_n4176_ = new_n3087_ & ~new_n4175_;
  assign new_n4177_ = ~new_n4169_ & ~new_n4176_;
  assign new_n4178_ = ~new_n3185_ & ~new_n4177_;
  assign new_n4179_ = new_n3087_ & ~new_n4168_;
  assign new_n4180_ = ~new_n3087_ & ~new_n4175_;
  assign new_n4181_ = ~new_n4179_ & ~new_n4180_;
  assign new_n4182_ = ~new_n3139_ & ~new_n4181_;
  assign new_n4183_ = \p_input[47]  & new_n3139_;
  assign new_n4184_ = ~new_n4182_ & ~new_n4183_;
  assign new_n4185_ = new_n3185_ & ~new_n4184_;
  assign new_n4186_ = ~new_n4178_ & ~new_n4185_;
  assign new_n4187_ = new_n3283_ & ~new_n4186_;
  assign new_n4188_ = new_n3185_ & ~new_n4177_;
  assign new_n4189_ = ~new_n3185_ & ~new_n4184_;
  assign new_n4190_ = ~new_n4188_ & ~new_n4189_;
  assign new_n4191_ = ~new_n3237_ & ~new_n4190_;
  assign new_n4192_ = \p_input[15]  & new_n3237_;
  assign new_n4193_ = ~new_n4191_ & ~new_n4192_;
  assign new_n4194_ = ~new_n3283_ & ~new_n4193_;
  assign \o[15]  = new_n4187_ | new_n4194_;
  assign new_n4196_ = \p_input[208]  & ~new_n2694_;
  assign new_n4197_ = \p_input[240]  & new_n2694_;
  assign new_n4198_ = ~new_n4196_ & ~new_n4197_;
  assign new_n4199_ = ~new_n2792_ & ~new_n4198_;
  assign new_n4200_ = ~\p_input[240]  & ~new_n2694_;
  assign new_n4201_ = ~\p_input[208]  & new_n2694_;
  assign new_n4202_ = ~new_n4200_ & ~new_n4201_;
  assign new_n4203_ = ~new_n2746_ & ~new_n4202_;
  assign new_n4204_ = ~\p_input[176]  & new_n2746_;
  assign new_n4205_ = ~new_n4203_ & ~new_n4204_;
  assign new_n4206_ = new_n2792_ & new_n4205_;
  assign new_n4207_ = ~new_n4199_ & ~new_n4206_;
  assign new_n4208_ = ~new_n2890_ & ~new_n4207_;
  assign new_n4209_ = new_n2792_ & ~new_n4198_;
  assign new_n4210_ = ~new_n2792_ & new_n4205_;
  assign new_n4211_ = ~new_n4209_ & ~new_n4210_;
  assign new_n4212_ = ~new_n2844_ & ~new_n4211_;
  assign new_n4213_ = \p_input[144]  & new_n2844_;
  assign new_n4214_ = ~new_n4212_ & ~new_n4213_;
  assign new_n4215_ = new_n2890_ & ~new_n4214_;
  assign new_n4216_ = ~new_n4208_ & ~new_n4215_;
  assign new_n4217_ = ~new_n2989_ & ~new_n4216_;
  assign new_n4218_ = new_n2890_ & ~new_n4207_;
  assign new_n4219_ = ~new_n2890_ & ~new_n4214_;
  assign new_n4220_ = ~new_n4218_ & ~new_n4219_;
  assign new_n4221_ = ~new_n2942_ & ~new_n4220_;
  assign new_n4222_ = \p_input[112]  & new_n2942_;
  assign new_n4223_ = ~new_n4221_ & ~new_n4222_;
  assign new_n4224_ = new_n2989_ & ~new_n4223_;
  assign new_n4225_ = ~new_n4217_ & ~new_n4224_;
  assign new_n4226_ = ~new_n3087_ & ~new_n4225_;
  assign new_n4227_ = new_n2989_ & ~new_n4216_;
  assign new_n4228_ = ~new_n2989_ & ~new_n4223_;
  assign new_n4229_ = ~new_n4227_ & ~new_n4228_;
  assign new_n4230_ = ~new_n3041_ & ~new_n4229_;
  assign new_n4231_ = \p_input[80]  & new_n3041_;
  assign new_n4232_ = ~new_n4230_ & ~new_n4231_;
  assign new_n4233_ = new_n3087_ & ~new_n4232_;
  assign new_n4234_ = ~new_n4226_ & ~new_n4233_;
  assign new_n4235_ = ~new_n3185_ & ~new_n4234_;
  assign new_n4236_ = new_n3087_ & ~new_n4225_;
  assign new_n4237_ = ~new_n3087_ & ~new_n4232_;
  assign new_n4238_ = ~new_n4236_ & ~new_n4237_;
  assign new_n4239_ = ~new_n3139_ & ~new_n4238_;
  assign new_n4240_ = \p_input[48]  & new_n3139_;
  assign new_n4241_ = ~new_n4239_ & ~new_n4240_;
  assign new_n4242_ = new_n3185_ & ~new_n4241_;
  assign new_n4243_ = ~new_n4235_ & ~new_n4242_;
  assign new_n4244_ = new_n3283_ & ~new_n4243_;
  assign new_n4245_ = new_n3185_ & ~new_n4234_;
  assign new_n4246_ = ~new_n3185_ & ~new_n4241_;
  assign new_n4247_ = ~new_n4245_ & ~new_n4246_;
  assign new_n4248_ = ~new_n3237_ & ~new_n4247_;
  assign new_n4249_ = \p_input[16]  & new_n3237_;
  assign new_n4250_ = ~new_n4248_ & ~new_n4249_;
  assign new_n4251_ = ~new_n3283_ & ~new_n4250_;
  assign \o[16]  = new_n4244_ | new_n4251_;
  assign new_n4253_ = \p_input[209]  & ~new_n2694_;
  assign new_n4254_ = \p_input[241]  & new_n2694_;
  assign new_n4255_ = ~new_n4253_ & ~new_n4254_;
  assign new_n4256_ = ~new_n2792_ & ~new_n4255_;
  assign new_n4257_ = ~\p_input[241]  & ~new_n2694_;
  assign new_n4258_ = ~\p_input[209]  & new_n2694_;
  assign new_n4259_ = ~new_n4257_ & ~new_n4258_;
  assign new_n4260_ = ~new_n2746_ & ~new_n4259_;
  assign new_n4261_ = ~\p_input[177]  & new_n2746_;
  assign new_n4262_ = ~new_n4260_ & ~new_n4261_;
  assign new_n4263_ = new_n2792_ & new_n4262_;
  assign new_n4264_ = ~new_n4256_ & ~new_n4263_;
  assign new_n4265_ = ~new_n2890_ & ~new_n4264_;
  assign new_n4266_ = new_n2792_ & ~new_n4255_;
  assign new_n4267_ = ~new_n2792_ & new_n4262_;
  assign new_n4268_ = ~new_n4266_ & ~new_n4267_;
  assign new_n4269_ = ~new_n2844_ & ~new_n4268_;
  assign new_n4270_ = \p_input[145]  & new_n2844_;
  assign new_n4271_ = ~new_n4269_ & ~new_n4270_;
  assign new_n4272_ = new_n2890_ & ~new_n4271_;
  assign new_n4273_ = ~new_n4265_ & ~new_n4272_;
  assign new_n4274_ = ~new_n2989_ & ~new_n4273_;
  assign new_n4275_ = new_n2890_ & ~new_n4264_;
  assign new_n4276_ = ~new_n2890_ & ~new_n4271_;
  assign new_n4277_ = ~new_n4275_ & ~new_n4276_;
  assign new_n4278_ = ~new_n2942_ & ~new_n4277_;
  assign new_n4279_ = \p_input[113]  & new_n2942_;
  assign new_n4280_ = ~new_n4278_ & ~new_n4279_;
  assign new_n4281_ = new_n2989_ & ~new_n4280_;
  assign new_n4282_ = ~new_n4274_ & ~new_n4281_;
  assign new_n4283_ = ~new_n3087_ & ~new_n4282_;
  assign new_n4284_ = new_n2989_ & ~new_n4273_;
  assign new_n4285_ = ~new_n2989_ & ~new_n4280_;
  assign new_n4286_ = ~new_n4284_ & ~new_n4285_;
  assign new_n4287_ = ~new_n3041_ & ~new_n4286_;
  assign new_n4288_ = \p_input[81]  & new_n3041_;
  assign new_n4289_ = ~new_n4287_ & ~new_n4288_;
  assign new_n4290_ = new_n3087_ & ~new_n4289_;
  assign new_n4291_ = ~new_n4283_ & ~new_n4290_;
  assign new_n4292_ = ~new_n3185_ & ~new_n4291_;
  assign new_n4293_ = new_n3087_ & ~new_n4282_;
  assign new_n4294_ = ~new_n3087_ & ~new_n4289_;
  assign new_n4295_ = ~new_n4293_ & ~new_n4294_;
  assign new_n4296_ = ~new_n3139_ & ~new_n4295_;
  assign new_n4297_ = \p_input[49]  & new_n3139_;
  assign new_n4298_ = ~new_n4296_ & ~new_n4297_;
  assign new_n4299_ = new_n3185_ & ~new_n4298_;
  assign new_n4300_ = ~new_n4292_ & ~new_n4299_;
  assign new_n4301_ = new_n3283_ & ~new_n4300_;
  assign new_n4302_ = new_n3185_ & ~new_n4291_;
  assign new_n4303_ = ~new_n3185_ & ~new_n4298_;
  assign new_n4304_ = ~new_n4302_ & ~new_n4303_;
  assign new_n4305_ = ~new_n3237_ & ~new_n4304_;
  assign new_n4306_ = \p_input[17]  & new_n3237_;
  assign new_n4307_ = ~new_n4305_ & ~new_n4306_;
  assign new_n4308_ = ~new_n3283_ & ~new_n4307_;
  assign \o[17]  = new_n4301_ | new_n4308_;
  assign new_n4310_ = \p_input[210]  & ~new_n2694_;
  assign new_n4311_ = \p_input[242]  & new_n2694_;
  assign new_n4312_ = ~new_n4310_ & ~new_n4311_;
  assign new_n4313_ = ~new_n2792_ & ~new_n4312_;
  assign new_n4314_ = ~\p_input[242]  & ~new_n2694_;
  assign new_n4315_ = ~\p_input[210]  & new_n2694_;
  assign new_n4316_ = ~new_n4314_ & ~new_n4315_;
  assign new_n4317_ = ~new_n2746_ & ~new_n4316_;
  assign new_n4318_ = ~\p_input[178]  & new_n2746_;
  assign new_n4319_ = ~new_n4317_ & ~new_n4318_;
  assign new_n4320_ = new_n2792_ & new_n4319_;
  assign new_n4321_ = ~new_n4313_ & ~new_n4320_;
  assign new_n4322_ = ~new_n2890_ & ~new_n4321_;
  assign new_n4323_ = new_n2792_ & ~new_n4312_;
  assign new_n4324_ = ~new_n2792_ & new_n4319_;
  assign new_n4325_ = ~new_n4323_ & ~new_n4324_;
  assign new_n4326_ = ~new_n2844_ & ~new_n4325_;
  assign new_n4327_ = \p_input[146]  & new_n2844_;
  assign new_n4328_ = ~new_n4326_ & ~new_n4327_;
  assign new_n4329_ = new_n2890_ & ~new_n4328_;
  assign new_n4330_ = ~new_n4322_ & ~new_n4329_;
  assign new_n4331_ = ~new_n2989_ & ~new_n4330_;
  assign new_n4332_ = new_n2890_ & ~new_n4321_;
  assign new_n4333_ = ~new_n2890_ & ~new_n4328_;
  assign new_n4334_ = ~new_n4332_ & ~new_n4333_;
  assign new_n4335_ = ~new_n2942_ & ~new_n4334_;
  assign new_n4336_ = \p_input[114]  & new_n2942_;
  assign new_n4337_ = ~new_n4335_ & ~new_n4336_;
  assign new_n4338_ = new_n2989_ & ~new_n4337_;
  assign new_n4339_ = ~new_n4331_ & ~new_n4338_;
  assign new_n4340_ = ~new_n3087_ & ~new_n4339_;
  assign new_n4341_ = new_n2989_ & ~new_n4330_;
  assign new_n4342_ = ~new_n2989_ & ~new_n4337_;
  assign new_n4343_ = ~new_n4341_ & ~new_n4342_;
  assign new_n4344_ = ~new_n3041_ & ~new_n4343_;
  assign new_n4345_ = \p_input[82]  & new_n3041_;
  assign new_n4346_ = ~new_n4344_ & ~new_n4345_;
  assign new_n4347_ = new_n3087_ & ~new_n4346_;
  assign new_n4348_ = ~new_n4340_ & ~new_n4347_;
  assign new_n4349_ = ~new_n3185_ & ~new_n4348_;
  assign new_n4350_ = new_n3087_ & ~new_n4339_;
  assign new_n4351_ = ~new_n3087_ & ~new_n4346_;
  assign new_n4352_ = ~new_n4350_ & ~new_n4351_;
  assign new_n4353_ = ~new_n3139_ & ~new_n4352_;
  assign new_n4354_ = \p_input[50]  & new_n3139_;
  assign new_n4355_ = ~new_n4353_ & ~new_n4354_;
  assign new_n4356_ = new_n3185_ & ~new_n4355_;
  assign new_n4357_ = ~new_n4349_ & ~new_n4356_;
  assign new_n4358_ = new_n3283_ & ~new_n4357_;
  assign new_n4359_ = new_n3185_ & ~new_n4348_;
  assign new_n4360_ = ~new_n3185_ & ~new_n4355_;
  assign new_n4361_ = ~new_n4359_ & ~new_n4360_;
  assign new_n4362_ = ~new_n3237_ & ~new_n4361_;
  assign new_n4363_ = \p_input[18]  & new_n3237_;
  assign new_n4364_ = ~new_n4362_ & ~new_n4363_;
  assign new_n4365_ = ~new_n3283_ & ~new_n4364_;
  assign \o[18]  = new_n4358_ | new_n4365_;
  assign new_n4367_ = \p_input[211]  & ~new_n2694_;
  assign new_n4368_ = \p_input[243]  & new_n2694_;
  assign new_n4369_ = ~new_n4367_ & ~new_n4368_;
  assign new_n4370_ = ~new_n2792_ & ~new_n4369_;
  assign new_n4371_ = ~\p_input[243]  & ~new_n2694_;
  assign new_n4372_ = ~\p_input[211]  & new_n2694_;
  assign new_n4373_ = ~new_n4371_ & ~new_n4372_;
  assign new_n4374_ = ~new_n2746_ & ~new_n4373_;
  assign new_n4375_ = ~\p_input[179]  & new_n2746_;
  assign new_n4376_ = ~new_n4374_ & ~new_n4375_;
  assign new_n4377_ = new_n2792_ & new_n4376_;
  assign new_n4378_ = ~new_n4370_ & ~new_n4377_;
  assign new_n4379_ = ~new_n2890_ & ~new_n4378_;
  assign new_n4380_ = new_n2792_ & ~new_n4369_;
  assign new_n4381_ = ~new_n2792_ & new_n4376_;
  assign new_n4382_ = ~new_n4380_ & ~new_n4381_;
  assign new_n4383_ = ~new_n2844_ & ~new_n4382_;
  assign new_n4384_ = \p_input[147]  & new_n2844_;
  assign new_n4385_ = ~new_n4383_ & ~new_n4384_;
  assign new_n4386_ = new_n2890_ & ~new_n4385_;
  assign new_n4387_ = ~new_n4379_ & ~new_n4386_;
  assign new_n4388_ = ~new_n2989_ & ~new_n4387_;
  assign new_n4389_ = new_n2890_ & ~new_n4378_;
  assign new_n4390_ = ~new_n2890_ & ~new_n4385_;
  assign new_n4391_ = ~new_n4389_ & ~new_n4390_;
  assign new_n4392_ = ~new_n2942_ & ~new_n4391_;
  assign new_n4393_ = \p_input[115]  & new_n2942_;
  assign new_n4394_ = ~new_n4392_ & ~new_n4393_;
  assign new_n4395_ = new_n2989_ & ~new_n4394_;
  assign new_n4396_ = ~new_n4388_ & ~new_n4395_;
  assign new_n4397_ = ~new_n3087_ & ~new_n4396_;
  assign new_n4398_ = new_n2989_ & ~new_n4387_;
  assign new_n4399_ = ~new_n2989_ & ~new_n4394_;
  assign new_n4400_ = ~new_n4398_ & ~new_n4399_;
  assign new_n4401_ = ~new_n3041_ & ~new_n4400_;
  assign new_n4402_ = \p_input[83]  & new_n3041_;
  assign new_n4403_ = ~new_n4401_ & ~new_n4402_;
  assign new_n4404_ = new_n3087_ & ~new_n4403_;
  assign new_n4405_ = ~new_n4397_ & ~new_n4404_;
  assign new_n4406_ = ~new_n3185_ & ~new_n4405_;
  assign new_n4407_ = new_n3087_ & ~new_n4396_;
  assign new_n4408_ = ~new_n3087_ & ~new_n4403_;
  assign new_n4409_ = ~new_n4407_ & ~new_n4408_;
  assign new_n4410_ = ~new_n3139_ & ~new_n4409_;
  assign new_n4411_ = \p_input[51]  & new_n3139_;
  assign new_n4412_ = ~new_n4410_ & ~new_n4411_;
  assign new_n4413_ = new_n3185_ & ~new_n4412_;
  assign new_n4414_ = ~new_n4406_ & ~new_n4413_;
  assign new_n4415_ = new_n3283_ & ~new_n4414_;
  assign new_n4416_ = new_n3185_ & ~new_n4405_;
  assign new_n4417_ = ~new_n3185_ & ~new_n4412_;
  assign new_n4418_ = ~new_n4416_ & ~new_n4417_;
  assign new_n4419_ = ~new_n3237_ & ~new_n4418_;
  assign new_n4420_ = \p_input[19]  & new_n3237_;
  assign new_n4421_ = ~new_n4419_ & ~new_n4420_;
  assign new_n4422_ = ~new_n3283_ & ~new_n4421_;
  assign \o[19]  = new_n4415_ | new_n4422_;
  assign new_n4424_ = \p_input[212]  & ~new_n2694_;
  assign new_n4425_ = \p_input[244]  & new_n2694_;
  assign new_n4426_ = ~new_n4424_ & ~new_n4425_;
  assign new_n4427_ = ~new_n2792_ & ~new_n4426_;
  assign new_n4428_ = ~\p_input[244]  & ~new_n2694_;
  assign new_n4429_ = ~\p_input[212]  & new_n2694_;
  assign new_n4430_ = ~new_n4428_ & ~new_n4429_;
  assign new_n4431_ = ~new_n2746_ & ~new_n4430_;
  assign new_n4432_ = ~\p_input[180]  & new_n2746_;
  assign new_n4433_ = ~new_n4431_ & ~new_n4432_;
  assign new_n4434_ = new_n2792_ & new_n4433_;
  assign new_n4435_ = ~new_n4427_ & ~new_n4434_;
  assign new_n4436_ = ~new_n2890_ & ~new_n4435_;
  assign new_n4437_ = new_n2792_ & ~new_n4426_;
  assign new_n4438_ = ~new_n2792_ & new_n4433_;
  assign new_n4439_ = ~new_n4437_ & ~new_n4438_;
  assign new_n4440_ = ~new_n2844_ & ~new_n4439_;
  assign new_n4441_ = \p_input[148]  & new_n2844_;
  assign new_n4442_ = ~new_n4440_ & ~new_n4441_;
  assign new_n4443_ = new_n2890_ & ~new_n4442_;
  assign new_n4444_ = ~new_n4436_ & ~new_n4443_;
  assign new_n4445_ = ~new_n2989_ & ~new_n4444_;
  assign new_n4446_ = new_n2890_ & ~new_n4435_;
  assign new_n4447_ = ~new_n2890_ & ~new_n4442_;
  assign new_n4448_ = ~new_n4446_ & ~new_n4447_;
  assign new_n4449_ = ~new_n2942_ & ~new_n4448_;
  assign new_n4450_ = \p_input[116]  & new_n2942_;
  assign new_n4451_ = ~new_n4449_ & ~new_n4450_;
  assign new_n4452_ = new_n2989_ & ~new_n4451_;
  assign new_n4453_ = ~new_n4445_ & ~new_n4452_;
  assign new_n4454_ = ~new_n3087_ & ~new_n4453_;
  assign new_n4455_ = new_n2989_ & ~new_n4444_;
  assign new_n4456_ = ~new_n2989_ & ~new_n4451_;
  assign new_n4457_ = ~new_n4455_ & ~new_n4456_;
  assign new_n4458_ = ~new_n3041_ & ~new_n4457_;
  assign new_n4459_ = \p_input[84]  & new_n3041_;
  assign new_n4460_ = ~new_n4458_ & ~new_n4459_;
  assign new_n4461_ = new_n3087_ & ~new_n4460_;
  assign new_n4462_ = ~new_n4454_ & ~new_n4461_;
  assign new_n4463_ = ~new_n3185_ & ~new_n4462_;
  assign new_n4464_ = new_n3087_ & ~new_n4453_;
  assign new_n4465_ = ~new_n3087_ & ~new_n4460_;
  assign new_n4466_ = ~new_n4464_ & ~new_n4465_;
  assign new_n4467_ = ~new_n3139_ & ~new_n4466_;
  assign new_n4468_ = \p_input[52]  & new_n3139_;
  assign new_n4469_ = ~new_n4467_ & ~new_n4468_;
  assign new_n4470_ = new_n3185_ & ~new_n4469_;
  assign new_n4471_ = ~new_n4463_ & ~new_n4470_;
  assign new_n4472_ = new_n3283_ & ~new_n4471_;
  assign new_n4473_ = new_n3185_ & ~new_n4462_;
  assign new_n4474_ = ~new_n3185_ & ~new_n4469_;
  assign new_n4475_ = ~new_n4473_ & ~new_n4474_;
  assign new_n4476_ = ~new_n3237_ & ~new_n4475_;
  assign new_n4477_ = \p_input[20]  & new_n3237_;
  assign new_n4478_ = ~new_n4476_ & ~new_n4477_;
  assign new_n4479_ = ~new_n3283_ & ~new_n4478_;
  assign \o[20]  = new_n4472_ | new_n4479_;
  assign new_n4481_ = \p_input[213]  & ~new_n2694_;
  assign new_n4482_ = \p_input[245]  & new_n2694_;
  assign new_n4483_ = ~new_n4481_ & ~new_n4482_;
  assign new_n4484_ = ~new_n2792_ & ~new_n4483_;
  assign new_n4485_ = ~\p_input[245]  & ~new_n2694_;
  assign new_n4486_ = ~\p_input[213]  & new_n2694_;
  assign new_n4487_ = ~new_n4485_ & ~new_n4486_;
  assign new_n4488_ = ~new_n2746_ & ~new_n4487_;
  assign new_n4489_ = ~\p_input[181]  & new_n2746_;
  assign new_n4490_ = ~new_n4488_ & ~new_n4489_;
  assign new_n4491_ = new_n2792_ & new_n4490_;
  assign new_n4492_ = ~new_n4484_ & ~new_n4491_;
  assign new_n4493_ = ~new_n2890_ & ~new_n4492_;
  assign new_n4494_ = new_n2792_ & ~new_n4483_;
  assign new_n4495_ = ~new_n2792_ & new_n4490_;
  assign new_n4496_ = ~new_n4494_ & ~new_n4495_;
  assign new_n4497_ = ~new_n2844_ & ~new_n4496_;
  assign new_n4498_ = \p_input[149]  & new_n2844_;
  assign new_n4499_ = ~new_n4497_ & ~new_n4498_;
  assign new_n4500_ = new_n2890_ & ~new_n4499_;
  assign new_n4501_ = ~new_n4493_ & ~new_n4500_;
  assign new_n4502_ = ~new_n2989_ & ~new_n4501_;
  assign new_n4503_ = new_n2890_ & ~new_n4492_;
  assign new_n4504_ = ~new_n2890_ & ~new_n4499_;
  assign new_n4505_ = ~new_n4503_ & ~new_n4504_;
  assign new_n4506_ = ~new_n2942_ & ~new_n4505_;
  assign new_n4507_ = \p_input[117]  & new_n2942_;
  assign new_n4508_ = ~new_n4506_ & ~new_n4507_;
  assign new_n4509_ = new_n2989_ & ~new_n4508_;
  assign new_n4510_ = ~new_n4502_ & ~new_n4509_;
  assign new_n4511_ = ~new_n3087_ & ~new_n4510_;
  assign new_n4512_ = new_n2989_ & ~new_n4501_;
  assign new_n4513_ = ~new_n2989_ & ~new_n4508_;
  assign new_n4514_ = ~new_n4512_ & ~new_n4513_;
  assign new_n4515_ = ~new_n3041_ & ~new_n4514_;
  assign new_n4516_ = \p_input[85]  & new_n3041_;
  assign new_n4517_ = ~new_n4515_ & ~new_n4516_;
  assign new_n4518_ = new_n3087_ & ~new_n4517_;
  assign new_n4519_ = ~new_n4511_ & ~new_n4518_;
  assign new_n4520_ = ~new_n3185_ & ~new_n4519_;
  assign new_n4521_ = new_n3087_ & ~new_n4510_;
  assign new_n4522_ = ~new_n3087_ & ~new_n4517_;
  assign new_n4523_ = ~new_n4521_ & ~new_n4522_;
  assign new_n4524_ = ~new_n3139_ & ~new_n4523_;
  assign new_n4525_ = \p_input[53]  & new_n3139_;
  assign new_n4526_ = ~new_n4524_ & ~new_n4525_;
  assign new_n4527_ = new_n3185_ & ~new_n4526_;
  assign new_n4528_ = ~new_n4520_ & ~new_n4527_;
  assign new_n4529_ = new_n3283_ & ~new_n4528_;
  assign new_n4530_ = new_n3185_ & ~new_n4519_;
  assign new_n4531_ = ~new_n3185_ & ~new_n4526_;
  assign new_n4532_ = ~new_n4530_ & ~new_n4531_;
  assign new_n4533_ = ~new_n3237_ & ~new_n4532_;
  assign new_n4534_ = \p_input[21]  & new_n3237_;
  assign new_n4535_ = ~new_n4533_ & ~new_n4534_;
  assign new_n4536_ = ~new_n3283_ & ~new_n4535_;
  assign \o[21]  = new_n4529_ | new_n4536_;
  assign new_n4538_ = \p_input[214]  & ~new_n2694_;
  assign new_n4539_ = \p_input[246]  & new_n2694_;
  assign new_n4540_ = ~new_n4538_ & ~new_n4539_;
  assign new_n4541_ = ~new_n2792_ & ~new_n4540_;
  assign new_n4542_ = ~\p_input[246]  & ~new_n2694_;
  assign new_n4543_ = ~\p_input[214]  & new_n2694_;
  assign new_n4544_ = ~new_n4542_ & ~new_n4543_;
  assign new_n4545_ = ~new_n2746_ & ~new_n4544_;
  assign new_n4546_ = ~\p_input[182]  & new_n2746_;
  assign new_n4547_ = ~new_n4545_ & ~new_n4546_;
  assign new_n4548_ = new_n2792_ & new_n4547_;
  assign new_n4549_ = ~new_n4541_ & ~new_n4548_;
  assign new_n4550_ = ~new_n2890_ & ~new_n4549_;
  assign new_n4551_ = new_n2792_ & ~new_n4540_;
  assign new_n4552_ = ~new_n2792_ & new_n4547_;
  assign new_n4553_ = ~new_n4551_ & ~new_n4552_;
  assign new_n4554_ = ~new_n2844_ & ~new_n4553_;
  assign new_n4555_ = \p_input[150]  & new_n2844_;
  assign new_n4556_ = ~new_n4554_ & ~new_n4555_;
  assign new_n4557_ = new_n2890_ & ~new_n4556_;
  assign new_n4558_ = ~new_n4550_ & ~new_n4557_;
  assign new_n4559_ = ~new_n2989_ & ~new_n4558_;
  assign new_n4560_ = new_n2890_ & ~new_n4549_;
  assign new_n4561_ = ~new_n2890_ & ~new_n4556_;
  assign new_n4562_ = ~new_n4560_ & ~new_n4561_;
  assign new_n4563_ = ~new_n2942_ & ~new_n4562_;
  assign new_n4564_ = \p_input[118]  & new_n2942_;
  assign new_n4565_ = ~new_n4563_ & ~new_n4564_;
  assign new_n4566_ = new_n2989_ & ~new_n4565_;
  assign new_n4567_ = ~new_n4559_ & ~new_n4566_;
  assign new_n4568_ = ~new_n3087_ & ~new_n4567_;
  assign new_n4569_ = new_n2989_ & ~new_n4558_;
  assign new_n4570_ = ~new_n2989_ & ~new_n4565_;
  assign new_n4571_ = ~new_n4569_ & ~new_n4570_;
  assign new_n4572_ = ~new_n3041_ & ~new_n4571_;
  assign new_n4573_ = \p_input[86]  & new_n3041_;
  assign new_n4574_ = ~new_n4572_ & ~new_n4573_;
  assign new_n4575_ = new_n3087_ & ~new_n4574_;
  assign new_n4576_ = ~new_n4568_ & ~new_n4575_;
  assign new_n4577_ = ~new_n3185_ & ~new_n4576_;
  assign new_n4578_ = new_n3087_ & ~new_n4567_;
  assign new_n4579_ = ~new_n3087_ & ~new_n4574_;
  assign new_n4580_ = ~new_n4578_ & ~new_n4579_;
  assign new_n4581_ = ~new_n3139_ & ~new_n4580_;
  assign new_n4582_ = \p_input[54]  & new_n3139_;
  assign new_n4583_ = ~new_n4581_ & ~new_n4582_;
  assign new_n4584_ = new_n3185_ & ~new_n4583_;
  assign new_n4585_ = ~new_n4577_ & ~new_n4584_;
  assign new_n4586_ = new_n3283_ & ~new_n4585_;
  assign new_n4587_ = new_n3185_ & ~new_n4576_;
  assign new_n4588_ = ~new_n3185_ & ~new_n4583_;
  assign new_n4589_ = ~new_n4587_ & ~new_n4588_;
  assign new_n4590_ = ~new_n3237_ & ~new_n4589_;
  assign new_n4591_ = \p_input[22]  & new_n3237_;
  assign new_n4592_ = ~new_n4590_ & ~new_n4591_;
  assign new_n4593_ = ~new_n3283_ & ~new_n4592_;
  assign \o[22]  = new_n4586_ | new_n4593_;
  assign new_n4595_ = \p_input[215]  & ~new_n2694_;
  assign new_n4596_ = \p_input[247]  & new_n2694_;
  assign new_n4597_ = ~new_n4595_ & ~new_n4596_;
  assign new_n4598_ = ~new_n2792_ & ~new_n4597_;
  assign new_n4599_ = ~\p_input[247]  & ~new_n2694_;
  assign new_n4600_ = ~\p_input[215]  & new_n2694_;
  assign new_n4601_ = ~new_n4599_ & ~new_n4600_;
  assign new_n4602_ = ~new_n2746_ & ~new_n4601_;
  assign new_n4603_ = ~\p_input[183]  & new_n2746_;
  assign new_n4604_ = ~new_n4602_ & ~new_n4603_;
  assign new_n4605_ = new_n2792_ & new_n4604_;
  assign new_n4606_ = ~new_n4598_ & ~new_n4605_;
  assign new_n4607_ = ~new_n2890_ & ~new_n4606_;
  assign new_n4608_ = new_n2792_ & ~new_n4597_;
  assign new_n4609_ = ~new_n2792_ & new_n4604_;
  assign new_n4610_ = ~new_n4608_ & ~new_n4609_;
  assign new_n4611_ = ~new_n2844_ & ~new_n4610_;
  assign new_n4612_ = \p_input[151]  & new_n2844_;
  assign new_n4613_ = ~new_n4611_ & ~new_n4612_;
  assign new_n4614_ = new_n2890_ & ~new_n4613_;
  assign new_n4615_ = ~new_n4607_ & ~new_n4614_;
  assign new_n4616_ = ~new_n2989_ & ~new_n4615_;
  assign new_n4617_ = new_n2890_ & ~new_n4606_;
  assign new_n4618_ = ~new_n2890_ & ~new_n4613_;
  assign new_n4619_ = ~new_n4617_ & ~new_n4618_;
  assign new_n4620_ = ~new_n2942_ & ~new_n4619_;
  assign new_n4621_ = \p_input[119]  & new_n2942_;
  assign new_n4622_ = ~new_n4620_ & ~new_n4621_;
  assign new_n4623_ = new_n2989_ & ~new_n4622_;
  assign new_n4624_ = ~new_n4616_ & ~new_n4623_;
  assign new_n4625_ = ~new_n3087_ & ~new_n4624_;
  assign new_n4626_ = new_n2989_ & ~new_n4615_;
  assign new_n4627_ = ~new_n2989_ & ~new_n4622_;
  assign new_n4628_ = ~new_n4626_ & ~new_n4627_;
  assign new_n4629_ = ~new_n3041_ & ~new_n4628_;
  assign new_n4630_ = \p_input[87]  & new_n3041_;
  assign new_n4631_ = ~new_n4629_ & ~new_n4630_;
  assign new_n4632_ = new_n3087_ & ~new_n4631_;
  assign new_n4633_ = ~new_n4625_ & ~new_n4632_;
  assign new_n4634_ = ~new_n3185_ & ~new_n4633_;
  assign new_n4635_ = new_n3087_ & ~new_n4624_;
  assign new_n4636_ = ~new_n3087_ & ~new_n4631_;
  assign new_n4637_ = ~new_n4635_ & ~new_n4636_;
  assign new_n4638_ = ~new_n3139_ & ~new_n4637_;
  assign new_n4639_ = \p_input[55]  & new_n3139_;
  assign new_n4640_ = ~new_n4638_ & ~new_n4639_;
  assign new_n4641_ = new_n3185_ & ~new_n4640_;
  assign new_n4642_ = ~new_n4634_ & ~new_n4641_;
  assign new_n4643_ = new_n3283_ & ~new_n4642_;
  assign new_n4644_ = new_n3185_ & ~new_n4633_;
  assign new_n4645_ = ~new_n3185_ & ~new_n4640_;
  assign new_n4646_ = ~new_n4644_ & ~new_n4645_;
  assign new_n4647_ = ~new_n3237_ & ~new_n4646_;
  assign new_n4648_ = \p_input[23]  & new_n3237_;
  assign new_n4649_ = ~new_n4647_ & ~new_n4648_;
  assign new_n4650_ = ~new_n3283_ & ~new_n4649_;
  assign \o[23]  = new_n4643_ | new_n4650_;
  assign new_n4652_ = \p_input[216]  & ~new_n2694_;
  assign new_n4653_ = \p_input[248]  & new_n2694_;
  assign new_n4654_ = ~new_n4652_ & ~new_n4653_;
  assign new_n4655_ = ~new_n2792_ & ~new_n4654_;
  assign new_n4656_ = ~\p_input[248]  & ~new_n2694_;
  assign new_n4657_ = ~\p_input[216]  & new_n2694_;
  assign new_n4658_ = ~new_n4656_ & ~new_n4657_;
  assign new_n4659_ = ~new_n2746_ & ~new_n4658_;
  assign new_n4660_ = ~\p_input[184]  & new_n2746_;
  assign new_n4661_ = ~new_n4659_ & ~new_n4660_;
  assign new_n4662_ = new_n2792_ & new_n4661_;
  assign new_n4663_ = ~new_n4655_ & ~new_n4662_;
  assign new_n4664_ = ~new_n2890_ & ~new_n4663_;
  assign new_n4665_ = new_n2792_ & ~new_n4654_;
  assign new_n4666_ = ~new_n2792_ & new_n4661_;
  assign new_n4667_ = ~new_n4665_ & ~new_n4666_;
  assign new_n4668_ = ~new_n2844_ & ~new_n4667_;
  assign new_n4669_ = \p_input[152]  & new_n2844_;
  assign new_n4670_ = ~new_n4668_ & ~new_n4669_;
  assign new_n4671_ = new_n2890_ & ~new_n4670_;
  assign new_n4672_ = ~new_n4664_ & ~new_n4671_;
  assign new_n4673_ = ~new_n2989_ & ~new_n4672_;
  assign new_n4674_ = new_n2890_ & ~new_n4663_;
  assign new_n4675_ = ~new_n2890_ & ~new_n4670_;
  assign new_n4676_ = ~new_n4674_ & ~new_n4675_;
  assign new_n4677_ = ~new_n2942_ & ~new_n4676_;
  assign new_n4678_ = \p_input[120]  & new_n2942_;
  assign new_n4679_ = ~new_n4677_ & ~new_n4678_;
  assign new_n4680_ = new_n2989_ & ~new_n4679_;
  assign new_n4681_ = ~new_n4673_ & ~new_n4680_;
  assign new_n4682_ = ~new_n3087_ & ~new_n4681_;
  assign new_n4683_ = new_n2989_ & ~new_n4672_;
  assign new_n4684_ = ~new_n2989_ & ~new_n4679_;
  assign new_n4685_ = ~new_n4683_ & ~new_n4684_;
  assign new_n4686_ = ~new_n3041_ & ~new_n4685_;
  assign new_n4687_ = \p_input[88]  & new_n3041_;
  assign new_n4688_ = ~new_n4686_ & ~new_n4687_;
  assign new_n4689_ = new_n3087_ & ~new_n4688_;
  assign new_n4690_ = ~new_n4682_ & ~new_n4689_;
  assign new_n4691_ = ~new_n3185_ & ~new_n4690_;
  assign new_n4692_ = new_n3087_ & ~new_n4681_;
  assign new_n4693_ = ~new_n3087_ & ~new_n4688_;
  assign new_n4694_ = ~new_n4692_ & ~new_n4693_;
  assign new_n4695_ = ~new_n3139_ & ~new_n4694_;
  assign new_n4696_ = \p_input[56]  & new_n3139_;
  assign new_n4697_ = ~new_n4695_ & ~new_n4696_;
  assign new_n4698_ = new_n3185_ & ~new_n4697_;
  assign new_n4699_ = ~new_n4691_ & ~new_n4698_;
  assign new_n4700_ = new_n3283_ & ~new_n4699_;
  assign new_n4701_ = new_n3185_ & ~new_n4690_;
  assign new_n4702_ = ~new_n3185_ & ~new_n4697_;
  assign new_n4703_ = ~new_n4701_ & ~new_n4702_;
  assign new_n4704_ = ~new_n3237_ & ~new_n4703_;
  assign new_n4705_ = \p_input[24]  & new_n3237_;
  assign new_n4706_ = ~new_n4704_ & ~new_n4705_;
  assign new_n4707_ = ~new_n3283_ & ~new_n4706_;
  assign \o[24]  = new_n4700_ | new_n4707_;
  assign new_n4709_ = \p_input[217]  & ~new_n2694_;
  assign new_n4710_ = \p_input[249]  & new_n2694_;
  assign new_n4711_ = ~new_n4709_ & ~new_n4710_;
  assign new_n4712_ = ~new_n2792_ & ~new_n4711_;
  assign new_n4713_ = ~\p_input[249]  & ~new_n2694_;
  assign new_n4714_ = ~\p_input[217]  & new_n2694_;
  assign new_n4715_ = ~new_n4713_ & ~new_n4714_;
  assign new_n4716_ = ~new_n2746_ & ~new_n4715_;
  assign new_n4717_ = ~\p_input[185]  & new_n2746_;
  assign new_n4718_ = ~new_n4716_ & ~new_n4717_;
  assign new_n4719_ = new_n2792_ & new_n4718_;
  assign new_n4720_ = ~new_n4712_ & ~new_n4719_;
  assign new_n4721_ = ~new_n2890_ & ~new_n4720_;
  assign new_n4722_ = new_n2792_ & ~new_n4711_;
  assign new_n4723_ = ~new_n2792_ & new_n4718_;
  assign new_n4724_ = ~new_n4722_ & ~new_n4723_;
  assign new_n4725_ = ~new_n2844_ & ~new_n4724_;
  assign new_n4726_ = \p_input[153]  & new_n2844_;
  assign new_n4727_ = ~new_n4725_ & ~new_n4726_;
  assign new_n4728_ = new_n2890_ & ~new_n4727_;
  assign new_n4729_ = ~new_n4721_ & ~new_n4728_;
  assign new_n4730_ = ~new_n2989_ & ~new_n4729_;
  assign new_n4731_ = new_n2890_ & ~new_n4720_;
  assign new_n4732_ = ~new_n2890_ & ~new_n4727_;
  assign new_n4733_ = ~new_n4731_ & ~new_n4732_;
  assign new_n4734_ = ~new_n2942_ & ~new_n4733_;
  assign new_n4735_ = \p_input[121]  & new_n2942_;
  assign new_n4736_ = ~new_n4734_ & ~new_n4735_;
  assign new_n4737_ = new_n2989_ & ~new_n4736_;
  assign new_n4738_ = ~new_n4730_ & ~new_n4737_;
  assign new_n4739_ = ~new_n3087_ & ~new_n4738_;
  assign new_n4740_ = new_n2989_ & ~new_n4729_;
  assign new_n4741_ = ~new_n2989_ & ~new_n4736_;
  assign new_n4742_ = ~new_n4740_ & ~new_n4741_;
  assign new_n4743_ = ~new_n3041_ & ~new_n4742_;
  assign new_n4744_ = \p_input[89]  & new_n3041_;
  assign new_n4745_ = ~new_n4743_ & ~new_n4744_;
  assign new_n4746_ = new_n3087_ & ~new_n4745_;
  assign new_n4747_ = ~new_n4739_ & ~new_n4746_;
  assign new_n4748_ = ~new_n3185_ & ~new_n4747_;
  assign new_n4749_ = new_n3087_ & ~new_n4738_;
  assign new_n4750_ = ~new_n3087_ & ~new_n4745_;
  assign new_n4751_ = ~new_n4749_ & ~new_n4750_;
  assign new_n4752_ = ~new_n3139_ & ~new_n4751_;
  assign new_n4753_ = \p_input[57]  & new_n3139_;
  assign new_n4754_ = ~new_n4752_ & ~new_n4753_;
  assign new_n4755_ = new_n3185_ & ~new_n4754_;
  assign new_n4756_ = ~new_n4748_ & ~new_n4755_;
  assign new_n4757_ = new_n3283_ & ~new_n4756_;
  assign new_n4758_ = new_n3185_ & ~new_n4747_;
  assign new_n4759_ = ~new_n3185_ & ~new_n4754_;
  assign new_n4760_ = ~new_n4758_ & ~new_n4759_;
  assign new_n4761_ = ~new_n3237_ & ~new_n4760_;
  assign new_n4762_ = \p_input[25]  & new_n3237_;
  assign new_n4763_ = ~new_n4761_ & ~new_n4762_;
  assign new_n4764_ = ~new_n3283_ & ~new_n4763_;
  assign \o[25]  = new_n4757_ | new_n4764_;
  assign new_n4766_ = \p_input[218]  & ~new_n2694_;
  assign new_n4767_ = \p_input[250]  & new_n2694_;
  assign new_n4768_ = ~new_n4766_ & ~new_n4767_;
  assign new_n4769_ = ~new_n2792_ & ~new_n4768_;
  assign new_n4770_ = ~\p_input[250]  & ~new_n2694_;
  assign new_n4771_ = ~\p_input[218]  & new_n2694_;
  assign new_n4772_ = ~new_n4770_ & ~new_n4771_;
  assign new_n4773_ = ~new_n2746_ & ~new_n4772_;
  assign new_n4774_ = ~\p_input[186]  & new_n2746_;
  assign new_n4775_ = ~new_n4773_ & ~new_n4774_;
  assign new_n4776_ = new_n2792_ & new_n4775_;
  assign new_n4777_ = ~new_n4769_ & ~new_n4776_;
  assign new_n4778_ = ~new_n2890_ & ~new_n4777_;
  assign new_n4779_ = new_n2792_ & ~new_n4768_;
  assign new_n4780_ = ~new_n2792_ & new_n4775_;
  assign new_n4781_ = ~new_n4779_ & ~new_n4780_;
  assign new_n4782_ = ~new_n2844_ & ~new_n4781_;
  assign new_n4783_ = \p_input[154]  & new_n2844_;
  assign new_n4784_ = ~new_n4782_ & ~new_n4783_;
  assign new_n4785_ = new_n2890_ & ~new_n4784_;
  assign new_n4786_ = ~new_n4778_ & ~new_n4785_;
  assign new_n4787_ = ~new_n2989_ & ~new_n4786_;
  assign new_n4788_ = new_n2890_ & ~new_n4777_;
  assign new_n4789_ = ~new_n2890_ & ~new_n4784_;
  assign new_n4790_ = ~new_n4788_ & ~new_n4789_;
  assign new_n4791_ = ~new_n2942_ & ~new_n4790_;
  assign new_n4792_ = \p_input[122]  & new_n2942_;
  assign new_n4793_ = ~new_n4791_ & ~new_n4792_;
  assign new_n4794_ = new_n2989_ & ~new_n4793_;
  assign new_n4795_ = ~new_n4787_ & ~new_n4794_;
  assign new_n4796_ = ~new_n3087_ & ~new_n4795_;
  assign new_n4797_ = new_n2989_ & ~new_n4786_;
  assign new_n4798_ = ~new_n2989_ & ~new_n4793_;
  assign new_n4799_ = ~new_n4797_ & ~new_n4798_;
  assign new_n4800_ = ~new_n3041_ & ~new_n4799_;
  assign new_n4801_ = \p_input[90]  & new_n3041_;
  assign new_n4802_ = ~new_n4800_ & ~new_n4801_;
  assign new_n4803_ = new_n3087_ & ~new_n4802_;
  assign new_n4804_ = ~new_n4796_ & ~new_n4803_;
  assign new_n4805_ = ~new_n3185_ & ~new_n4804_;
  assign new_n4806_ = new_n3087_ & ~new_n4795_;
  assign new_n4807_ = ~new_n3087_ & ~new_n4802_;
  assign new_n4808_ = ~new_n4806_ & ~new_n4807_;
  assign new_n4809_ = ~new_n3139_ & ~new_n4808_;
  assign new_n4810_ = \p_input[58]  & new_n3139_;
  assign new_n4811_ = ~new_n4809_ & ~new_n4810_;
  assign new_n4812_ = new_n3185_ & ~new_n4811_;
  assign new_n4813_ = ~new_n4805_ & ~new_n4812_;
  assign new_n4814_ = new_n3283_ & ~new_n4813_;
  assign new_n4815_ = new_n3185_ & ~new_n4804_;
  assign new_n4816_ = ~new_n3185_ & ~new_n4811_;
  assign new_n4817_ = ~new_n4815_ & ~new_n4816_;
  assign new_n4818_ = ~new_n3237_ & ~new_n4817_;
  assign new_n4819_ = \p_input[26]  & new_n3237_;
  assign new_n4820_ = ~new_n4818_ & ~new_n4819_;
  assign new_n4821_ = ~new_n3283_ & ~new_n4820_;
  assign \o[26]  = new_n4814_ | new_n4821_;
  assign new_n4823_ = \p_input[219]  & ~new_n2694_;
  assign new_n4824_ = \p_input[251]  & new_n2694_;
  assign new_n4825_ = ~new_n4823_ & ~new_n4824_;
  assign new_n4826_ = ~new_n2792_ & ~new_n4825_;
  assign new_n4827_ = ~\p_input[251]  & ~new_n2694_;
  assign new_n4828_ = ~\p_input[219]  & new_n2694_;
  assign new_n4829_ = ~new_n4827_ & ~new_n4828_;
  assign new_n4830_ = ~new_n2746_ & ~new_n4829_;
  assign new_n4831_ = ~\p_input[187]  & new_n2746_;
  assign new_n4832_ = ~new_n4830_ & ~new_n4831_;
  assign new_n4833_ = new_n2792_ & new_n4832_;
  assign new_n4834_ = ~new_n4826_ & ~new_n4833_;
  assign new_n4835_ = ~new_n2890_ & ~new_n4834_;
  assign new_n4836_ = new_n2792_ & ~new_n4825_;
  assign new_n4837_ = ~new_n2792_ & new_n4832_;
  assign new_n4838_ = ~new_n4836_ & ~new_n4837_;
  assign new_n4839_ = ~new_n2844_ & ~new_n4838_;
  assign new_n4840_ = \p_input[155]  & new_n2844_;
  assign new_n4841_ = ~new_n4839_ & ~new_n4840_;
  assign new_n4842_ = new_n2890_ & ~new_n4841_;
  assign new_n4843_ = ~new_n4835_ & ~new_n4842_;
  assign new_n4844_ = ~new_n2989_ & ~new_n4843_;
  assign new_n4845_ = new_n2890_ & ~new_n4834_;
  assign new_n4846_ = ~new_n2890_ & ~new_n4841_;
  assign new_n4847_ = ~new_n4845_ & ~new_n4846_;
  assign new_n4848_ = ~new_n2942_ & ~new_n4847_;
  assign new_n4849_ = \p_input[123]  & new_n2942_;
  assign new_n4850_ = ~new_n4848_ & ~new_n4849_;
  assign new_n4851_ = new_n2989_ & ~new_n4850_;
  assign new_n4852_ = ~new_n4844_ & ~new_n4851_;
  assign new_n4853_ = ~new_n3087_ & ~new_n4852_;
  assign new_n4854_ = new_n2989_ & ~new_n4843_;
  assign new_n4855_ = ~new_n2989_ & ~new_n4850_;
  assign new_n4856_ = ~new_n4854_ & ~new_n4855_;
  assign new_n4857_ = ~new_n3041_ & ~new_n4856_;
  assign new_n4858_ = \p_input[91]  & new_n3041_;
  assign new_n4859_ = ~new_n4857_ & ~new_n4858_;
  assign new_n4860_ = new_n3087_ & ~new_n4859_;
  assign new_n4861_ = ~new_n4853_ & ~new_n4860_;
  assign new_n4862_ = ~new_n3185_ & ~new_n4861_;
  assign new_n4863_ = new_n3087_ & ~new_n4852_;
  assign new_n4864_ = ~new_n3087_ & ~new_n4859_;
  assign new_n4865_ = ~new_n4863_ & ~new_n4864_;
  assign new_n4866_ = ~new_n3139_ & ~new_n4865_;
  assign new_n4867_ = \p_input[59]  & new_n3139_;
  assign new_n4868_ = ~new_n4866_ & ~new_n4867_;
  assign new_n4869_ = new_n3185_ & ~new_n4868_;
  assign new_n4870_ = ~new_n4862_ & ~new_n4869_;
  assign new_n4871_ = new_n3283_ & ~new_n4870_;
  assign new_n4872_ = new_n3185_ & ~new_n4861_;
  assign new_n4873_ = ~new_n3185_ & ~new_n4868_;
  assign new_n4874_ = ~new_n4872_ & ~new_n4873_;
  assign new_n4875_ = ~new_n3237_ & ~new_n4874_;
  assign new_n4876_ = \p_input[27]  & new_n3237_;
  assign new_n4877_ = ~new_n4875_ & ~new_n4876_;
  assign new_n4878_ = ~new_n3283_ & ~new_n4877_;
  assign \o[27]  = new_n4871_ | new_n4878_;
  assign new_n4880_ = \p_input[220]  & ~new_n2694_;
  assign new_n4881_ = \p_input[252]  & new_n2694_;
  assign new_n4882_ = ~new_n4880_ & ~new_n4881_;
  assign new_n4883_ = ~new_n2792_ & ~new_n4882_;
  assign new_n4884_ = ~\p_input[252]  & ~new_n2694_;
  assign new_n4885_ = ~\p_input[220]  & new_n2694_;
  assign new_n4886_ = ~new_n4884_ & ~new_n4885_;
  assign new_n4887_ = ~new_n2746_ & ~new_n4886_;
  assign new_n4888_ = ~\p_input[188]  & new_n2746_;
  assign new_n4889_ = ~new_n4887_ & ~new_n4888_;
  assign new_n4890_ = new_n2792_ & new_n4889_;
  assign new_n4891_ = ~new_n4883_ & ~new_n4890_;
  assign new_n4892_ = ~new_n2890_ & ~new_n4891_;
  assign new_n4893_ = new_n2792_ & ~new_n4882_;
  assign new_n4894_ = ~new_n2792_ & new_n4889_;
  assign new_n4895_ = ~new_n4893_ & ~new_n4894_;
  assign new_n4896_ = ~new_n2844_ & ~new_n4895_;
  assign new_n4897_ = \p_input[156]  & new_n2844_;
  assign new_n4898_ = ~new_n4896_ & ~new_n4897_;
  assign new_n4899_ = new_n2890_ & ~new_n4898_;
  assign new_n4900_ = ~new_n4892_ & ~new_n4899_;
  assign new_n4901_ = ~new_n2989_ & ~new_n4900_;
  assign new_n4902_ = new_n2890_ & ~new_n4891_;
  assign new_n4903_ = ~new_n2890_ & ~new_n4898_;
  assign new_n4904_ = ~new_n4902_ & ~new_n4903_;
  assign new_n4905_ = ~new_n2942_ & ~new_n4904_;
  assign new_n4906_ = \p_input[124]  & new_n2942_;
  assign new_n4907_ = ~new_n4905_ & ~new_n4906_;
  assign new_n4908_ = new_n2989_ & ~new_n4907_;
  assign new_n4909_ = ~new_n4901_ & ~new_n4908_;
  assign new_n4910_ = ~new_n3087_ & ~new_n4909_;
  assign new_n4911_ = new_n2989_ & ~new_n4900_;
  assign new_n4912_ = ~new_n2989_ & ~new_n4907_;
  assign new_n4913_ = ~new_n4911_ & ~new_n4912_;
  assign new_n4914_ = ~new_n3041_ & ~new_n4913_;
  assign new_n4915_ = \p_input[92]  & new_n3041_;
  assign new_n4916_ = ~new_n4914_ & ~new_n4915_;
  assign new_n4917_ = new_n3087_ & ~new_n4916_;
  assign new_n4918_ = ~new_n4910_ & ~new_n4917_;
  assign new_n4919_ = ~new_n3185_ & ~new_n4918_;
  assign new_n4920_ = new_n3087_ & ~new_n4909_;
  assign new_n4921_ = ~new_n3087_ & ~new_n4916_;
  assign new_n4922_ = ~new_n4920_ & ~new_n4921_;
  assign new_n4923_ = ~new_n3139_ & ~new_n4922_;
  assign new_n4924_ = \p_input[60]  & new_n3139_;
  assign new_n4925_ = ~new_n4923_ & ~new_n4924_;
  assign new_n4926_ = new_n3185_ & ~new_n4925_;
  assign new_n4927_ = ~new_n4919_ & ~new_n4926_;
  assign new_n4928_ = new_n3283_ & ~new_n4927_;
  assign new_n4929_ = new_n3185_ & ~new_n4918_;
  assign new_n4930_ = ~new_n3185_ & ~new_n4925_;
  assign new_n4931_ = ~new_n4929_ & ~new_n4930_;
  assign new_n4932_ = ~new_n3237_ & ~new_n4931_;
  assign new_n4933_ = \p_input[28]  & new_n3237_;
  assign new_n4934_ = ~new_n4932_ & ~new_n4933_;
  assign new_n4935_ = ~new_n3283_ & ~new_n4934_;
  assign \o[28]  = new_n4928_ | new_n4935_;
  assign new_n4937_ = \p_input[221]  & ~new_n2694_;
  assign new_n4938_ = \p_input[253]  & new_n2694_;
  assign new_n4939_ = ~new_n4937_ & ~new_n4938_;
  assign new_n4940_ = ~new_n2792_ & ~new_n4939_;
  assign new_n4941_ = ~\p_input[253]  & ~new_n2694_;
  assign new_n4942_ = ~\p_input[221]  & new_n2694_;
  assign new_n4943_ = ~new_n4941_ & ~new_n4942_;
  assign new_n4944_ = ~new_n2746_ & ~new_n4943_;
  assign new_n4945_ = ~\p_input[189]  & new_n2746_;
  assign new_n4946_ = ~new_n4944_ & ~new_n4945_;
  assign new_n4947_ = new_n2792_ & new_n4946_;
  assign new_n4948_ = ~new_n4940_ & ~new_n4947_;
  assign new_n4949_ = ~new_n2890_ & ~new_n4948_;
  assign new_n4950_ = new_n2792_ & ~new_n4939_;
  assign new_n4951_ = ~new_n2792_ & new_n4946_;
  assign new_n4952_ = ~new_n4950_ & ~new_n4951_;
  assign new_n4953_ = ~new_n2844_ & ~new_n4952_;
  assign new_n4954_ = \p_input[157]  & new_n2844_;
  assign new_n4955_ = ~new_n4953_ & ~new_n4954_;
  assign new_n4956_ = new_n2890_ & ~new_n4955_;
  assign new_n4957_ = ~new_n4949_ & ~new_n4956_;
  assign new_n4958_ = ~new_n2989_ & ~new_n4957_;
  assign new_n4959_ = new_n2890_ & ~new_n4948_;
  assign new_n4960_ = ~new_n2890_ & ~new_n4955_;
  assign new_n4961_ = ~new_n4959_ & ~new_n4960_;
  assign new_n4962_ = ~new_n2942_ & ~new_n4961_;
  assign new_n4963_ = \p_input[125]  & new_n2942_;
  assign new_n4964_ = ~new_n4962_ & ~new_n4963_;
  assign new_n4965_ = new_n2989_ & ~new_n4964_;
  assign new_n4966_ = ~new_n4958_ & ~new_n4965_;
  assign new_n4967_ = ~new_n3087_ & ~new_n4966_;
  assign new_n4968_ = new_n2989_ & ~new_n4957_;
  assign new_n4969_ = ~new_n2989_ & ~new_n4964_;
  assign new_n4970_ = ~new_n4968_ & ~new_n4969_;
  assign new_n4971_ = ~new_n3041_ & ~new_n4970_;
  assign new_n4972_ = \p_input[93]  & new_n3041_;
  assign new_n4973_ = ~new_n4971_ & ~new_n4972_;
  assign new_n4974_ = new_n3087_ & ~new_n4973_;
  assign new_n4975_ = ~new_n4967_ & ~new_n4974_;
  assign new_n4976_ = ~new_n3185_ & ~new_n4975_;
  assign new_n4977_ = new_n3087_ & ~new_n4966_;
  assign new_n4978_ = ~new_n3087_ & ~new_n4973_;
  assign new_n4979_ = ~new_n4977_ & ~new_n4978_;
  assign new_n4980_ = ~new_n3139_ & ~new_n4979_;
  assign new_n4981_ = \p_input[61]  & new_n3139_;
  assign new_n4982_ = ~new_n4980_ & ~new_n4981_;
  assign new_n4983_ = new_n3185_ & ~new_n4982_;
  assign new_n4984_ = ~new_n4976_ & ~new_n4983_;
  assign new_n4985_ = new_n3283_ & ~new_n4984_;
  assign new_n4986_ = new_n3185_ & ~new_n4975_;
  assign new_n4987_ = ~new_n3185_ & ~new_n4982_;
  assign new_n4988_ = ~new_n4986_ & ~new_n4987_;
  assign new_n4989_ = ~new_n3237_ & ~new_n4988_;
  assign new_n4990_ = \p_input[29]  & new_n3237_;
  assign new_n4991_ = ~new_n4989_ & ~new_n4990_;
  assign new_n4992_ = ~new_n3283_ & ~new_n4991_;
  assign \o[29]  = new_n4985_ | new_n4992_;
  assign new_n4994_ = \p_input[222]  & ~new_n2694_;
  assign new_n4995_ = \p_input[254]  & new_n2694_;
  assign new_n4996_ = ~new_n4994_ & ~new_n4995_;
  assign new_n4997_ = ~new_n2792_ & ~new_n4996_;
  assign new_n4998_ = ~\p_input[254]  & ~new_n2694_;
  assign new_n4999_ = ~\p_input[222]  & new_n2694_;
  assign new_n5000_ = ~new_n4998_ & ~new_n4999_;
  assign new_n5001_ = ~new_n2746_ & ~new_n5000_;
  assign new_n5002_ = ~\p_input[190]  & new_n2746_;
  assign new_n5003_ = ~new_n5001_ & ~new_n5002_;
  assign new_n5004_ = new_n2792_ & new_n5003_;
  assign new_n5005_ = ~new_n4997_ & ~new_n5004_;
  assign new_n5006_ = ~new_n2890_ & ~new_n5005_;
  assign new_n5007_ = new_n2792_ & ~new_n4996_;
  assign new_n5008_ = ~new_n2792_ & new_n5003_;
  assign new_n5009_ = ~new_n5007_ & ~new_n5008_;
  assign new_n5010_ = ~new_n2844_ & ~new_n5009_;
  assign new_n5011_ = \p_input[158]  & new_n2844_;
  assign new_n5012_ = ~new_n5010_ & ~new_n5011_;
  assign new_n5013_ = new_n2890_ & ~new_n5012_;
  assign new_n5014_ = ~new_n5006_ & ~new_n5013_;
  assign new_n5015_ = ~new_n2989_ & ~new_n5014_;
  assign new_n5016_ = new_n2890_ & ~new_n5005_;
  assign new_n5017_ = ~new_n2890_ & ~new_n5012_;
  assign new_n5018_ = ~new_n5016_ & ~new_n5017_;
  assign new_n5019_ = ~new_n2942_ & ~new_n5018_;
  assign new_n5020_ = \p_input[126]  & new_n2942_;
  assign new_n5021_ = ~new_n5019_ & ~new_n5020_;
  assign new_n5022_ = new_n2989_ & ~new_n5021_;
  assign new_n5023_ = ~new_n5015_ & ~new_n5022_;
  assign new_n5024_ = ~new_n3087_ & ~new_n5023_;
  assign new_n5025_ = new_n2989_ & ~new_n5014_;
  assign new_n5026_ = ~new_n2989_ & ~new_n5021_;
  assign new_n5027_ = ~new_n5025_ & ~new_n5026_;
  assign new_n5028_ = ~new_n3041_ & ~new_n5027_;
  assign new_n5029_ = \p_input[94]  & new_n3041_;
  assign new_n5030_ = ~new_n5028_ & ~new_n5029_;
  assign new_n5031_ = new_n3087_ & ~new_n5030_;
  assign new_n5032_ = ~new_n5024_ & ~new_n5031_;
  assign new_n5033_ = ~new_n3185_ & ~new_n5032_;
  assign new_n5034_ = new_n3087_ & ~new_n5023_;
  assign new_n5035_ = ~new_n3087_ & ~new_n5030_;
  assign new_n5036_ = ~new_n5034_ & ~new_n5035_;
  assign new_n5037_ = ~new_n3139_ & ~new_n5036_;
  assign new_n5038_ = \p_input[62]  & new_n3139_;
  assign new_n5039_ = ~new_n5037_ & ~new_n5038_;
  assign new_n5040_ = new_n3185_ & ~new_n5039_;
  assign new_n5041_ = ~new_n5033_ & ~new_n5040_;
  assign new_n5042_ = new_n3283_ & ~new_n5041_;
  assign new_n5043_ = new_n3185_ & ~new_n5032_;
  assign new_n5044_ = ~new_n3185_ & ~new_n5039_;
  assign new_n5045_ = ~new_n5043_ & ~new_n5044_;
  assign new_n5046_ = ~new_n3237_ & ~new_n5045_;
  assign new_n5047_ = \p_input[30]  & new_n3237_;
  assign new_n5048_ = ~new_n5046_ & ~new_n5047_;
  assign new_n5049_ = ~new_n3283_ & ~new_n5048_;
  assign \o[30]  = new_n5042_ | new_n5049_;
  assign new_n5051_ = \p_input[223]  & ~new_n2694_;
  assign new_n5052_ = \p_input[255]  & new_n2694_;
  assign new_n5053_ = ~new_n5051_ & ~new_n5052_;
  assign new_n5054_ = ~new_n2792_ & ~new_n5053_;
  assign new_n5055_ = ~\p_input[255]  & ~new_n2694_;
  assign new_n5056_ = ~\p_input[223]  & new_n2694_;
  assign new_n5057_ = ~new_n5055_ & ~new_n5056_;
  assign new_n5058_ = ~new_n2746_ & ~new_n5057_;
  assign new_n5059_ = ~\p_input[191]  & new_n2746_;
  assign new_n5060_ = ~new_n5058_ & ~new_n5059_;
  assign new_n5061_ = new_n2792_ & new_n5060_;
  assign new_n5062_ = ~new_n5054_ & ~new_n5061_;
  assign new_n5063_ = ~new_n2890_ & ~new_n5062_;
  assign new_n5064_ = new_n2792_ & ~new_n5053_;
  assign new_n5065_ = ~new_n2792_ & new_n5060_;
  assign new_n5066_ = ~new_n5064_ & ~new_n5065_;
  assign new_n5067_ = ~new_n2844_ & ~new_n5066_;
  assign new_n5068_ = \p_input[159]  & new_n2844_;
  assign new_n5069_ = ~new_n5067_ & ~new_n5068_;
  assign new_n5070_ = new_n2890_ & ~new_n5069_;
  assign new_n5071_ = ~new_n5063_ & ~new_n5070_;
  assign new_n5072_ = ~new_n2989_ & ~new_n5071_;
  assign new_n5073_ = new_n2890_ & ~new_n5062_;
  assign new_n5074_ = ~new_n2890_ & ~new_n5069_;
  assign new_n5075_ = ~new_n5073_ & ~new_n5074_;
  assign new_n5076_ = ~new_n2942_ & ~new_n5075_;
  assign new_n5077_ = \p_input[127]  & new_n2942_;
  assign new_n5078_ = ~new_n5076_ & ~new_n5077_;
  assign new_n5079_ = new_n2989_ & ~new_n5078_;
  assign new_n5080_ = ~new_n5072_ & ~new_n5079_;
  assign new_n5081_ = ~new_n3087_ & ~new_n5080_;
  assign new_n5082_ = new_n2989_ & ~new_n5071_;
  assign new_n5083_ = ~new_n2989_ & ~new_n5078_;
  assign new_n5084_ = ~new_n5082_ & ~new_n5083_;
  assign new_n5085_ = ~new_n3041_ & ~new_n5084_;
  assign new_n5086_ = \p_input[95]  & new_n3041_;
  assign new_n5087_ = ~new_n5085_ & ~new_n5086_;
  assign new_n5088_ = new_n3087_ & ~new_n5087_;
  assign new_n5089_ = ~new_n5081_ & ~new_n5088_;
  assign new_n5090_ = ~new_n3185_ & ~new_n5089_;
  assign new_n5091_ = new_n3087_ & ~new_n5080_;
  assign new_n5092_ = ~new_n3087_ & ~new_n5087_;
  assign new_n5093_ = ~new_n5091_ & ~new_n5092_;
  assign new_n5094_ = ~new_n3139_ & ~new_n5093_;
  assign new_n5095_ = \p_input[63]  & new_n3139_;
  assign new_n5096_ = ~new_n5094_ & ~new_n5095_;
  assign new_n5097_ = new_n3185_ & ~new_n5096_;
  assign new_n5098_ = ~new_n5090_ & ~new_n5097_;
  assign new_n5099_ = new_n3283_ & ~new_n5098_;
  assign new_n5100_ = new_n3185_ & ~new_n5089_;
  assign new_n5101_ = ~new_n3185_ & ~new_n5096_;
  assign new_n5102_ = ~new_n5100_ & ~new_n5101_;
  assign new_n5103_ = ~new_n3237_ & ~new_n5102_;
  assign new_n5104_ = \p_input[31]  & new_n3237_;
  assign new_n5105_ = ~new_n5103_ & ~new_n5104_;
  assign new_n5106_ = ~new_n3283_ & ~new_n5105_;
  assign \o[31]  = new_n5099_ | new_n5106_;
  assign new_n5108_ = ~new_n3283_ & ~new_n3331_;
  assign new_n5109_ = new_n3283_ & ~new_n3338_;
  assign \o[32]  = new_n5108_ | new_n5109_;
  assign new_n5111_ = ~new_n3283_ & ~new_n3388_;
  assign new_n5112_ = new_n3283_ & ~new_n3395_;
  assign \o[33]  = new_n5111_ | new_n5112_;
  assign new_n5114_ = ~new_n3283_ & ~new_n3445_;
  assign new_n5115_ = new_n3283_ & ~new_n3452_;
  assign \o[34]  = new_n5114_ | new_n5115_;
  assign new_n5117_ = ~new_n3283_ & ~new_n3502_;
  assign new_n5118_ = new_n3283_ & ~new_n3509_;
  assign \o[35]  = new_n5117_ | new_n5118_;
  assign new_n5120_ = ~new_n3283_ & ~new_n3559_;
  assign new_n5121_ = new_n3283_ & ~new_n3566_;
  assign \o[36]  = new_n5120_ | new_n5121_;
  assign new_n5123_ = ~new_n3283_ & ~new_n3616_;
  assign new_n5124_ = new_n3283_ & ~new_n3623_;
  assign \o[37]  = new_n5123_ | new_n5124_;
  assign new_n5126_ = ~new_n3283_ & ~new_n3673_;
  assign new_n5127_ = new_n3283_ & ~new_n3680_;
  assign \o[38]  = new_n5126_ | new_n5127_;
  assign new_n5129_ = ~new_n3283_ & ~new_n3730_;
  assign new_n5130_ = new_n3283_ & ~new_n3737_;
  assign \o[39]  = new_n5129_ | new_n5130_;
  assign new_n5132_ = ~new_n3283_ & ~new_n3787_;
  assign new_n5133_ = new_n3283_ & ~new_n3794_;
  assign \o[40]  = new_n5132_ | new_n5133_;
  assign new_n5135_ = ~new_n3283_ & ~new_n3844_;
  assign new_n5136_ = new_n3283_ & ~new_n3851_;
  assign \o[41]  = new_n5135_ | new_n5136_;
  assign new_n5138_ = ~new_n3283_ & ~new_n3901_;
  assign new_n5139_ = new_n3283_ & ~new_n3908_;
  assign \o[42]  = new_n5138_ | new_n5139_;
  assign new_n5141_ = ~new_n3283_ & ~new_n3958_;
  assign new_n5142_ = new_n3283_ & ~new_n3965_;
  assign \o[43]  = new_n5141_ | new_n5142_;
  assign new_n5144_ = ~new_n3283_ & ~new_n4015_;
  assign new_n5145_ = new_n3283_ & ~new_n4022_;
  assign \o[44]  = new_n5144_ | new_n5145_;
  assign new_n5147_ = ~new_n3283_ & ~new_n4072_;
  assign new_n5148_ = new_n3283_ & ~new_n4079_;
  assign \o[45]  = new_n5147_ | new_n5148_;
  assign new_n5150_ = ~new_n3283_ & ~new_n4129_;
  assign new_n5151_ = new_n3283_ & ~new_n4136_;
  assign \o[46]  = new_n5150_ | new_n5151_;
  assign new_n5153_ = ~new_n3283_ & ~new_n4186_;
  assign new_n5154_ = new_n3283_ & ~new_n4193_;
  assign \o[47]  = new_n5153_ | new_n5154_;
  assign new_n5156_ = ~new_n3283_ & ~new_n4243_;
  assign new_n5157_ = new_n3283_ & ~new_n4250_;
  assign \o[48]  = new_n5156_ | new_n5157_;
  assign new_n5159_ = ~new_n3283_ & ~new_n4300_;
  assign new_n5160_ = new_n3283_ & ~new_n4307_;
  assign \o[49]  = new_n5159_ | new_n5160_;
  assign new_n5162_ = ~new_n3283_ & ~new_n4357_;
  assign new_n5163_ = new_n3283_ & ~new_n4364_;
  assign \o[50]  = new_n5162_ | new_n5163_;
  assign new_n5165_ = ~new_n3283_ & ~new_n4414_;
  assign new_n5166_ = new_n3283_ & ~new_n4421_;
  assign \o[51]  = new_n5165_ | new_n5166_;
  assign new_n5168_ = ~new_n3283_ & ~new_n4471_;
  assign new_n5169_ = new_n3283_ & ~new_n4478_;
  assign \o[52]  = new_n5168_ | new_n5169_;
  assign new_n5171_ = ~new_n3283_ & ~new_n4528_;
  assign new_n5172_ = new_n3283_ & ~new_n4535_;
  assign \o[53]  = new_n5171_ | new_n5172_;
  assign new_n5174_ = ~new_n3283_ & ~new_n4585_;
  assign new_n5175_ = new_n3283_ & ~new_n4592_;
  assign \o[54]  = new_n5174_ | new_n5175_;
  assign new_n5177_ = ~new_n3283_ & ~new_n4642_;
  assign new_n5178_ = new_n3283_ & ~new_n4649_;
  assign \o[55]  = new_n5177_ | new_n5178_;
  assign new_n5180_ = ~new_n3283_ & ~new_n4699_;
  assign new_n5181_ = new_n3283_ & ~new_n4706_;
  assign \o[56]  = new_n5180_ | new_n5181_;
  assign new_n5183_ = ~new_n3283_ & ~new_n4756_;
  assign new_n5184_ = new_n3283_ & ~new_n4763_;
  assign \o[57]  = new_n5183_ | new_n5184_;
  assign new_n5186_ = ~new_n3283_ & ~new_n4813_;
  assign new_n5187_ = new_n3283_ & ~new_n4820_;
  assign \o[58]  = new_n5186_ | new_n5187_;
  assign new_n5189_ = ~new_n3283_ & ~new_n4870_;
  assign new_n5190_ = new_n3283_ & ~new_n4877_;
  assign \o[59]  = new_n5189_ | new_n5190_;
  assign new_n5192_ = ~new_n3283_ & ~new_n4927_;
  assign new_n5193_ = new_n3283_ & ~new_n4934_;
  assign \o[60]  = new_n5192_ | new_n5193_;
  assign new_n5195_ = ~new_n3283_ & ~new_n4984_;
  assign new_n5196_ = new_n3283_ & ~new_n4991_;
  assign \o[61]  = new_n5195_ | new_n5196_;
  assign new_n5198_ = ~new_n3283_ & ~new_n5041_;
  assign new_n5199_ = new_n3283_ & ~new_n5048_;
  assign \o[62]  = new_n5198_ | new_n5199_;
  assign new_n5201_ = ~new_n3283_ & ~new_n5098_;
  assign new_n5202_ = new_n3283_ & ~new_n5105_;
  assign \o[63]  = new_n5201_ | new_n5202_;
endmodule


