module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 ;
  wire n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 ;
  assign n1568 = x270 ^ x14 ;
  assign n1567 = x271 ^ x15 ;
  assign n1569 = n1568 ^ n1567 ;
  assign n1566 = x272 ^ x16 ;
  assign n1597 = n1568 ^ n1566 ;
  assign n1598 = n1569 & ~n1597 ;
  assign n1599 = n1598 ^ n1567 ;
  assign n1571 = x266 ^ x10 ;
  assign n1570 = n1569 ^ n1566 ;
  assign n1572 = n1571 ^ n1570 ;
  assign n1564 = x269 ^ x13 ;
  assign n1562 = x267 ^ x11 ;
  assign n1561 = x268 ^ x12 ;
  assign n1563 = n1562 ^ n1561 ;
  assign n1565 = n1564 ^ n1563 ;
  assign n1594 = n1571 ^ n1565 ;
  assign n1595 = n1572 & ~n1594 ;
  assign n1596 = n1595 ^ n1570 ;
  assign n1600 = n1599 ^ n1596 ;
  assign n1591 = n1564 ^ n1562 ;
  assign n1592 = n1563 & ~n1591 ;
  assign n1593 = n1592 ^ n1561 ;
  assign n1617 = n1599 ^ n1593 ;
  assign n1618 = n1600 & ~n1617 ;
  assign n1619 = n1618 ^ n1596 ;
  assign n1573 = n1572 ^ n1565 ;
  assign n1560 = x258 ^ x2 ;
  assign n1574 = n1573 ^ n1560 ;
  assign n1557 = x259 ^ x3 ;
  assign n1555 = x265 ^ x9 ;
  assign n1553 = x263 ^ x7 ;
  assign n1552 = x264 ^ x8 ;
  assign n1554 = n1553 ^ n1552 ;
  assign n1556 = n1555 ^ n1554 ;
  assign n1558 = n1557 ^ n1556 ;
  assign n1550 = x262 ^ x6 ;
  assign n1548 = x260 ^ x4 ;
  assign n1547 = x261 ^ x5 ;
  assign n1549 = n1548 ^ n1547 ;
  assign n1551 = n1550 ^ n1549 ;
  assign n1559 = n1558 ^ n1551 ;
  assign n1602 = n1573 ^ n1559 ;
  assign n1603 = n1574 & ~n1602 ;
  assign n1604 = n1603 ^ n1560 ;
  assign n1601 = n1600 ^ n1593 ;
  assign n1605 = n1604 ^ n1601 ;
  assign n1587 = n1550 ^ n1548 ;
  assign n1588 = n1549 & ~n1587 ;
  assign n1589 = n1588 ^ n1547 ;
  assign n1583 = n1556 ^ n1551 ;
  assign n1584 = ~n1558 & n1583 ;
  assign n1585 = n1584 ^ n1551 ;
  assign n1580 = n1555 ^ n1553 ;
  assign n1581 = n1554 & ~n1580 ;
  assign n1582 = n1581 ^ n1552 ;
  assign n1586 = n1585 ^ n1582 ;
  assign n1590 = n1589 ^ n1586 ;
  assign n1614 = n1601 ^ n1590 ;
  assign n1615 = n1605 & ~n1614 ;
  assign n1616 = n1615 ^ n1604 ;
  assign n1620 = n1619 ^ n1616 ;
  assign n1611 = n1589 ^ n1585 ;
  assign n1612 = n1586 & ~n1611 ;
  assign n1613 = n1612 ^ n1582 ;
  assign n1626 = n1619 ^ n1613 ;
  assign n1627 = n1620 & ~n1626 ;
  assign n1628 = n1627 ^ n1616 ;
  assign n1545 = x257 ^ x1 ;
  assign n1514 = x277 ^ x21 ;
  assign n1512 = x275 ^ x19 ;
  assign n1511 = x276 ^ x20 ;
  assign n1513 = n1512 ^ n1511 ;
  assign n1515 = n1514 ^ n1513 ;
  assign n1509 = x274 ^ x18 ;
  assign n1507 = x280 ^ x24 ;
  assign n1505 = x278 ^ x22 ;
  assign n1504 = x279 ^ x23 ;
  assign n1506 = n1505 ^ n1504 ;
  assign n1508 = n1507 ^ n1506 ;
  assign n1510 = n1509 ^ n1508 ;
  assign n1516 = n1515 ^ n1510 ;
  assign n1502 = x273 ^ x17 ;
  assign n1488 = x284 ^ x28 ;
  assign n1486 = x282 ^ x26 ;
  assign n1485 = x283 ^ x27 ;
  assign n1487 = n1486 ^ n1485 ;
  assign n1489 = n1488 ^ n1487 ;
  assign n1478 = x287 ^ x31 ;
  assign n1476 = x286 ^ x30 ;
  assign n1475 = x285 ^ x29 ;
  assign n1477 = n1476 ^ n1475 ;
  assign n1483 = n1478 ^ n1477 ;
  assign n1482 = x281 ^ x25 ;
  assign n1484 = n1483 ^ n1482 ;
  assign n1501 = n1489 ^ n1484 ;
  assign n1503 = n1502 ^ n1501 ;
  assign n1544 = n1516 ^ n1503 ;
  assign n1546 = n1545 ^ n1544 ;
  assign n1575 = n1574 ^ n1559 ;
  assign n1576 = n1575 ^ n1545 ;
  assign n1577 = n1546 & ~n1576 ;
  assign n1578 = n1577 ^ n1544 ;
  assign n1528 = n1514 ^ n1512 ;
  assign n1529 = n1513 & ~n1528 ;
  assign n1530 = n1529 ^ n1511 ;
  assign n1524 = n1507 ^ n1505 ;
  assign n1525 = n1506 & ~n1524 ;
  assign n1526 = n1525 ^ n1504 ;
  assign n1521 = n1515 ^ n1509 ;
  assign n1522 = n1510 & ~n1521 ;
  assign n1523 = n1522 ^ n1508 ;
  assign n1527 = n1526 ^ n1523 ;
  assign n1531 = n1530 ^ n1527 ;
  assign n1517 = n1516 ^ n1502 ;
  assign n1518 = n1503 & ~n1517 ;
  assign n1519 = n1518 ^ n1501 ;
  assign n1494 = n1488 ^ n1486 ;
  assign n1495 = n1487 & ~n1494 ;
  assign n1496 = n1495 ^ n1485 ;
  assign n1490 = n1489 ^ n1483 ;
  assign n1491 = n1484 & ~n1490 ;
  assign n1492 = n1491 ^ n1482 ;
  assign n1479 = n1478 ^ n1476 ;
  assign n1480 = n1477 & ~n1479 ;
  assign n1481 = n1480 ^ n1475 ;
  assign n1493 = n1492 ^ n1481 ;
  assign n1500 = n1496 ^ n1493 ;
  assign n1520 = n1519 ^ n1500 ;
  assign n1543 = n1531 ^ n1520 ;
  assign n1579 = n1578 ^ n1543 ;
  assign n1606 = n1605 ^ n1590 ;
  assign n1607 = n1606 ^ n1543 ;
  assign n1608 = n1579 & ~n1607 ;
  assign n1609 = n1608 ^ n1578 ;
  assign n1536 = n1530 ^ n1526 ;
  assign n1537 = n1527 & ~n1536 ;
  assign n1538 = n1537 ^ n1523 ;
  assign n1532 = n1531 ^ n1500 ;
  assign n1533 = n1520 & ~n1532 ;
  assign n1534 = n1533 ^ n1519 ;
  assign n1497 = n1496 ^ n1492 ;
  assign n1498 = n1493 & ~n1497 ;
  assign n1499 = n1498 ^ n1481 ;
  assign n1535 = n1534 ^ n1499 ;
  assign n1542 = n1538 ^ n1535 ;
  assign n1610 = n1609 ^ n1542 ;
  assign n1621 = n1620 ^ n1613 ;
  assign n1622 = n1621 ^ n1609 ;
  assign n1623 = n1610 & ~n1622 ;
  assign n1624 = n1623 ^ n1542 ;
  assign n1539 = n1538 ^ n1534 ;
  assign n1540 = n1535 & ~n1539 ;
  assign n1541 = n1540 ^ n1499 ;
  assign n1625 = n1624 ^ n1541 ;
  assign n1629 = n1628 ^ n1625 ;
  assign n1630 = n1606 ^ n1579 ;
  assign n1631 = n1575 ^ n1546 ;
  assign n1632 = x256 ^ x0 ;
  assign n1633 = n1631 & n1632 ;
  assign n1634 = n1630 & n1633 ;
  assign n1635 = n1621 ^ n1610 ;
  assign n1636 = n1634 & n1635 ;
  assign n1637 = n1629 & n1636 ;
  assign n1638 = n1628 ^ n1541 ;
  assign n1639 = ~n1625 & n1638 ;
  assign n1640 = n1639 ^ n1628 ;
  assign n1641 = n1637 & n1640 ;
  assign n387 = x258 ^ x34 ;
  assign n384 = x266 ^ x42 ;
  assign n382 = x272 ^ x48 ;
  assign n380 = x270 ^ x46 ;
  assign n379 = x271 ^ x47 ;
  assign n381 = n380 ^ n379 ;
  assign n383 = n382 ^ n381 ;
  assign n385 = n384 ^ n383 ;
  assign n377 = x269 ^ x45 ;
  assign n375 = x267 ^ x43 ;
  assign n374 = x268 ^ x44 ;
  assign n376 = n375 ^ n374 ;
  assign n378 = n377 ^ n376 ;
  assign n386 = n385 ^ n378 ;
  assign n388 = n387 ^ n386 ;
  assign n371 = x259 ^ x35 ;
  assign n369 = x265 ^ x41 ;
  assign n367 = x263 ^ x39 ;
  assign n366 = x264 ^ x40 ;
  assign n368 = n367 ^ n366 ;
  assign n370 = n369 ^ n368 ;
  assign n372 = n371 ^ n370 ;
  assign n364 = x262 ^ x38 ;
  assign n362 = x260 ^ x36 ;
  assign n361 = x261 ^ x37 ;
  assign n363 = n362 ^ n361 ;
  assign n365 = n364 ^ n363 ;
  assign n373 = n372 ^ n365 ;
  assign n416 = n387 ^ n373 ;
  assign n417 = n388 & ~n416 ;
  assign n418 = n417 ^ n386 ;
  assign n412 = n377 ^ n375 ;
  assign n413 = n376 & ~n412 ;
  assign n414 = n413 ^ n374 ;
  assign n408 = n382 ^ n380 ;
  assign n409 = n381 & ~n408 ;
  assign n410 = n409 ^ n379 ;
  assign n405 = n383 ^ n378 ;
  assign n406 = ~n385 & n405 ;
  assign n407 = n406 ^ n378 ;
  assign n411 = n410 ^ n407 ;
  assign n415 = n414 ^ n411 ;
  assign n419 = n418 ^ n415 ;
  assign n401 = n364 ^ n362 ;
  assign n402 = n363 & ~n401 ;
  assign n403 = n402 ^ n361 ;
  assign n397 = n370 ^ n365 ;
  assign n398 = ~n372 & n397 ;
  assign n399 = n398 ^ n365 ;
  assign n394 = n369 ^ n367 ;
  assign n395 = n368 & ~n394 ;
  assign n396 = n395 ^ n366 ;
  assign n400 = n399 ^ n396 ;
  assign n404 = n403 ^ n400 ;
  assign n431 = n418 ^ n404 ;
  assign n432 = n419 & ~n431 ;
  assign n433 = n432 ^ n415 ;
  assign n428 = n414 ^ n410 ;
  assign n429 = n411 & ~n428 ;
  assign n430 = n429 ^ n407 ;
  assign n434 = n433 ^ n430 ;
  assign n425 = n403 ^ n399 ;
  assign n426 = n400 & ~n425 ;
  assign n427 = n426 ^ n396 ;
  assign n440 = n430 ^ n427 ;
  assign n441 = ~n434 & n440 ;
  assign n442 = n441 ^ n427 ;
  assign n359 = x257 ^ x33 ;
  assign n325 = x277 ^ x53 ;
  assign n323 = x275 ^ x51 ;
  assign n322 = x276 ^ x52 ;
  assign n324 = n323 ^ n322 ;
  assign n326 = n325 ^ n324 ;
  assign n320 = x274 ^ x50 ;
  assign n318 = x280 ^ x56 ;
  assign n316 = x278 ^ x54 ;
  assign n315 = x279 ^ x55 ;
  assign n317 = n316 ^ n315 ;
  assign n319 = n318 ^ n317 ;
  assign n321 = n320 ^ n319 ;
  assign n327 = n326 ^ n321 ;
  assign n298 = x282 ^ x58 ;
  assign n297 = x283 ^ x59 ;
  assign n299 = n298 ^ n297 ;
  assign n296 = x284 ^ x60 ;
  assign n300 = n299 ^ n296 ;
  assign n294 = x281 ^ x57 ;
  assign n291 = x285 ^ x61 ;
  assign n290 = x286 ^ x62 ;
  assign n292 = n291 ^ n290 ;
  assign n289 = x287 ^ x63 ;
  assign n293 = n292 ^ n289 ;
  assign n295 = n294 ^ n293 ;
  assign n313 = n300 ^ n295 ;
  assign n312 = x273 ^ x49 ;
  assign n314 = n313 ^ n312 ;
  assign n358 = n327 ^ n314 ;
  assign n360 = n359 ^ n358 ;
  assign n389 = n388 ^ n373 ;
  assign n390 = n389 ^ n359 ;
  assign n391 = n360 & ~n390 ;
  assign n392 = n391 ^ n358 ;
  assign n339 = n325 ^ n323 ;
  assign n340 = n324 & ~n339 ;
  assign n341 = n340 ^ n322 ;
  assign n335 = n318 ^ n316 ;
  assign n336 = n317 & ~n335 ;
  assign n337 = n336 ^ n315 ;
  assign n332 = n326 ^ n320 ;
  assign n333 = n321 & ~n332 ;
  assign n334 = n333 ^ n319 ;
  assign n338 = n337 ^ n334 ;
  assign n342 = n341 ^ n338 ;
  assign n328 = n327 ^ n313 ;
  assign n329 = n314 & ~n328 ;
  assign n330 = n329 ^ n312 ;
  assign n308 = n297 ^ n296 ;
  assign n309 = ~n299 & n308 ;
  assign n310 = n309 ^ n296 ;
  assign n304 = n290 ^ n289 ;
  assign n305 = ~n292 & n304 ;
  assign n306 = n305 ^ n289 ;
  assign n301 = n300 ^ n294 ;
  assign n302 = n295 & ~n301 ;
  assign n303 = n302 ^ n293 ;
  assign n307 = n306 ^ n303 ;
  assign n311 = n310 ^ n307 ;
  assign n331 = n330 ^ n311 ;
  assign n357 = n342 ^ n331 ;
  assign n393 = n392 ^ n357 ;
  assign n420 = n419 ^ n404 ;
  assign n421 = n420 ^ n357 ;
  assign n422 = n393 & ~n421 ;
  assign n423 = n422 ^ n392 ;
  assign n350 = n341 ^ n337 ;
  assign n351 = n338 & ~n350 ;
  assign n352 = n351 ^ n334 ;
  assign n346 = n310 ^ n306 ;
  assign n347 = n307 & ~n346 ;
  assign n348 = n347 ^ n303 ;
  assign n343 = n342 ^ n330 ;
  assign n344 = n331 & ~n343 ;
  assign n345 = n344 ^ n311 ;
  assign n349 = n348 ^ n345 ;
  assign n356 = n352 ^ n349 ;
  assign n424 = n423 ^ n356 ;
  assign n435 = n434 ^ n427 ;
  assign n436 = n435 ^ n423 ;
  assign n437 = n424 & ~n436 ;
  assign n438 = n437 ^ n356 ;
  assign n353 = n352 ^ n348 ;
  assign n354 = n349 & ~n353 ;
  assign n355 = n354 ^ n345 ;
  assign n439 = n438 ^ n355 ;
  assign n443 = n442 ^ n439 ;
  assign n444 = n389 ^ n360 ;
  assign n445 = x256 ^ x32 ;
  assign n446 = n444 & n445 ;
  assign n447 = n420 ^ n393 ;
  assign n448 = n446 & n447 ;
  assign n449 = n435 ^ n424 ;
  assign n450 = n448 & n449 ;
  assign n451 = n443 & n450 ;
  assign n452 = n442 ^ n438 ;
  assign n453 = n439 & ~n452 ;
  assign n454 = n453 ^ n355 ;
  assign n455 = n451 & n454 ;
  assign n554 = x258 ^ x66 ;
  assign n551 = x266 ^ x74 ;
  assign n549 = x272 ^ x80 ;
  assign n547 = x270 ^ x78 ;
  assign n546 = x271 ^ x79 ;
  assign n548 = n547 ^ n546 ;
  assign n550 = n549 ^ n548 ;
  assign n552 = n551 ^ n550 ;
  assign n544 = x269 ^ x77 ;
  assign n542 = x267 ^ x75 ;
  assign n541 = x268 ^ x76 ;
  assign n543 = n542 ^ n541 ;
  assign n545 = n544 ^ n543 ;
  assign n553 = n552 ^ n545 ;
  assign n555 = n554 ^ n553 ;
  assign n538 = x259 ^ x67 ;
  assign n536 = x265 ^ x73 ;
  assign n534 = x263 ^ x71 ;
  assign n533 = x264 ^ x72 ;
  assign n535 = n534 ^ n533 ;
  assign n537 = n536 ^ n535 ;
  assign n539 = n538 ^ n537 ;
  assign n531 = x262 ^ x70 ;
  assign n529 = x260 ^ x68 ;
  assign n528 = x261 ^ x69 ;
  assign n530 = n529 ^ n528 ;
  assign n532 = n531 ^ n530 ;
  assign n540 = n539 ^ n532 ;
  assign n583 = n554 ^ n540 ;
  assign n584 = n555 & ~n583 ;
  assign n585 = n584 ^ n553 ;
  assign n579 = n544 ^ n542 ;
  assign n580 = n543 & ~n579 ;
  assign n581 = n580 ^ n541 ;
  assign n575 = n549 ^ n547 ;
  assign n576 = n548 & ~n575 ;
  assign n577 = n576 ^ n546 ;
  assign n572 = n550 ^ n545 ;
  assign n573 = ~n552 & n572 ;
  assign n574 = n573 ^ n545 ;
  assign n578 = n577 ^ n574 ;
  assign n582 = n581 ^ n578 ;
  assign n586 = n585 ^ n582 ;
  assign n568 = n531 ^ n529 ;
  assign n569 = n530 & ~n568 ;
  assign n570 = n569 ^ n528 ;
  assign n564 = n537 ^ n532 ;
  assign n565 = ~n539 & n564 ;
  assign n566 = n565 ^ n532 ;
  assign n561 = n536 ^ n534 ;
  assign n562 = n535 & ~n561 ;
  assign n563 = n562 ^ n533 ;
  assign n567 = n566 ^ n563 ;
  assign n571 = n570 ^ n567 ;
  assign n598 = n585 ^ n571 ;
  assign n599 = n586 & ~n598 ;
  assign n600 = n599 ^ n582 ;
  assign n595 = n581 ^ n577 ;
  assign n596 = n578 & ~n595 ;
  assign n597 = n596 ^ n574 ;
  assign n601 = n600 ^ n597 ;
  assign n592 = n570 ^ n566 ;
  assign n593 = n567 & ~n592 ;
  assign n594 = n593 ^ n563 ;
  assign n607 = n597 ^ n594 ;
  assign n608 = ~n601 & n607 ;
  assign n609 = n608 ^ n594 ;
  assign n526 = x257 ^ x65 ;
  assign n492 = x277 ^ x85 ;
  assign n490 = x275 ^ x83 ;
  assign n489 = x276 ^ x84 ;
  assign n491 = n490 ^ n489 ;
  assign n493 = n492 ^ n491 ;
  assign n487 = x274 ^ x82 ;
  assign n485 = x280 ^ x88 ;
  assign n483 = x278 ^ x86 ;
  assign n482 = x279 ^ x87 ;
  assign n484 = n483 ^ n482 ;
  assign n486 = n485 ^ n484 ;
  assign n488 = n487 ^ n486 ;
  assign n494 = n493 ^ n488 ;
  assign n465 = x282 ^ x90 ;
  assign n464 = x283 ^ x91 ;
  assign n466 = n465 ^ n464 ;
  assign n463 = x284 ^ x92 ;
  assign n467 = n466 ^ n463 ;
  assign n461 = x281 ^ x89 ;
  assign n458 = x285 ^ x93 ;
  assign n457 = x286 ^ x94 ;
  assign n459 = n458 ^ n457 ;
  assign n456 = x287 ^ x95 ;
  assign n460 = n459 ^ n456 ;
  assign n462 = n461 ^ n460 ;
  assign n480 = n467 ^ n462 ;
  assign n479 = x273 ^ x81 ;
  assign n481 = n480 ^ n479 ;
  assign n525 = n494 ^ n481 ;
  assign n527 = n526 ^ n525 ;
  assign n556 = n555 ^ n540 ;
  assign n557 = n556 ^ n526 ;
  assign n558 = n527 & ~n557 ;
  assign n559 = n558 ^ n525 ;
  assign n506 = n492 ^ n490 ;
  assign n507 = n491 & ~n506 ;
  assign n508 = n507 ^ n489 ;
  assign n502 = n485 ^ n483 ;
  assign n503 = n484 & ~n502 ;
  assign n504 = n503 ^ n482 ;
  assign n499 = n493 ^ n487 ;
  assign n500 = n488 & ~n499 ;
  assign n501 = n500 ^ n486 ;
  assign n505 = n504 ^ n501 ;
  assign n509 = n508 ^ n505 ;
  assign n495 = n494 ^ n480 ;
  assign n496 = n481 & ~n495 ;
  assign n497 = n496 ^ n479 ;
  assign n475 = n464 ^ n463 ;
  assign n476 = ~n466 & n475 ;
  assign n477 = n476 ^ n463 ;
  assign n471 = n457 ^ n456 ;
  assign n472 = ~n459 & n471 ;
  assign n473 = n472 ^ n456 ;
  assign n468 = n467 ^ n461 ;
  assign n469 = n462 & ~n468 ;
  assign n470 = n469 ^ n460 ;
  assign n474 = n473 ^ n470 ;
  assign n478 = n477 ^ n474 ;
  assign n498 = n497 ^ n478 ;
  assign n524 = n509 ^ n498 ;
  assign n560 = n559 ^ n524 ;
  assign n587 = n586 ^ n571 ;
  assign n588 = n587 ^ n524 ;
  assign n589 = n560 & ~n588 ;
  assign n590 = n589 ^ n559 ;
  assign n517 = n508 ^ n504 ;
  assign n518 = n505 & ~n517 ;
  assign n519 = n518 ^ n501 ;
  assign n513 = n477 ^ n473 ;
  assign n514 = n474 & ~n513 ;
  assign n515 = n514 ^ n470 ;
  assign n510 = n509 ^ n497 ;
  assign n511 = n498 & ~n510 ;
  assign n512 = n511 ^ n478 ;
  assign n516 = n515 ^ n512 ;
  assign n523 = n519 ^ n516 ;
  assign n591 = n590 ^ n523 ;
  assign n602 = n601 ^ n594 ;
  assign n603 = n602 ^ n590 ;
  assign n604 = n591 & ~n603 ;
  assign n605 = n604 ^ n523 ;
  assign n520 = n519 ^ n515 ;
  assign n521 = n516 & ~n520 ;
  assign n522 = n521 ^ n512 ;
  assign n606 = n605 ^ n522 ;
  assign n610 = n609 ^ n606 ;
  assign n611 = n556 ^ n527 ;
  assign n612 = x256 ^ x64 ;
  assign n613 = n611 & n612 ;
  assign n614 = n587 ^ n560 ;
  assign n615 = n613 & n614 ;
  assign n616 = n602 ^ n591 ;
  assign n617 = n615 & n616 ;
  assign n618 = n610 & n617 ;
  assign n619 = n609 ^ n605 ;
  assign n620 = n606 & ~n619 ;
  assign n621 = n620 ^ n522 ;
  assign n622 = n618 & n621 ;
  assign n721 = x258 ^ x98 ;
  assign n718 = x266 ^ x106 ;
  assign n716 = x272 ^ x112 ;
  assign n714 = x270 ^ x110 ;
  assign n713 = x271 ^ x111 ;
  assign n715 = n714 ^ n713 ;
  assign n717 = n716 ^ n715 ;
  assign n719 = n718 ^ n717 ;
  assign n711 = x269 ^ x109 ;
  assign n709 = x267 ^ x107 ;
  assign n708 = x268 ^ x108 ;
  assign n710 = n709 ^ n708 ;
  assign n712 = n711 ^ n710 ;
  assign n720 = n719 ^ n712 ;
  assign n722 = n721 ^ n720 ;
  assign n705 = x259 ^ x99 ;
  assign n703 = x265 ^ x105 ;
  assign n701 = x263 ^ x103 ;
  assign n700 = x264 ^ x104 ;
  assign n702 = n701 ^ n700 ;
  assign n704 = n703 ^ n702 ;
  assign n706 = n705 ^ n704 ;
  assign n698 = x262 ^ x102 ;
  assign n696 = x260 ^ x100 ;
  assign n695 = x261 ^ x101 ;
  assign n697 = n696 ^ n695 ;
  assign n699 = n698 ^ n697 ;
  assign n707 = n706 ^ n699 ;
  assign n750 = n721 ^ n707 ;
  assign n751 = n722 & ~n750 ;
  assign n752 = n751 ^ n720 ;
  assign n746 = n711 ^ n709 ;
  assign n747 = n710 & ~n746 ;
  assign n748 = n747 ^ n708 ;
  assign n742 = n716 ^ n714 ;
  assign n743 = n715 & ~n742 ;
  assign n744 = n743 ^ n713 ;
  assign n739 = n717 ^ n712 ;
  assign n740 = ~n719 & n739 ;
  assign n741 = n740 ^ n712 ;
  assign n745 = n744 ^ n741 ;
  assign n749 = n748 ^ n745 ;
  assign n753 = n752 ^ n749 ;
  assign n735 = n698 ^ n696 ;
  assign n736 = n697 & ~n735 ;
  assign n737 = n736 ^ n695 ;
  assign n731 = n704 ^ n699 ;
  assign n732 = ~n706 & n731 ;
  assign n733 = n732 ^ n699 ;
  assign n728 = n703 ^ n701 ;
  assign n729 = n702 & ~n728 ;
  assign n730 = n729 ^ n700 ;
  assign n734 = n733 ^ n730 ;
  assign n738 = n737 ^ n734 ;
  assign n765 = n752 ^ n738 ;
  assign n766 = n753 & ~n765 ;
  assign n767 = n766 ^ n749 ;
  assign n762 = n748 ^ n744 ;
  assign n763 = n745 & ~n762 ;
  assign n764 = n763 ^ n741 ;
  assign n768 = n767 ^ n764 ;
  assign n759 = n737 ^ n733 ;
  assign n760 = n734 & ~n759 ;
  assign n761 = n760 ^ n730 ;
  assign n774 = n764 ^ n761 ;
  assign n775 = ~n768 & n774 ;
  assign n776 = n775 ^ n761 ;
  assign n693 = x257 ^ x97 ;
  assign n659 = x277 ^ x117 ;
  assign n657 = x275 ^ x115 ;
  assign n656 = x276 ^ x116 ;
  assign n658 = n657 ^ n656 ;
  assign n660 = n659 ^ n658 ;
  assign n654 = x274 ^ x114 ;
  assign n652 = x280 ^ x120 ;
  assign n650 = x278 ^ x118 ;
  assign n649 = x279 ^ x119 ;
  assign n651 = n650 ^ n649 ;
  assign n653 = n652 ^ n651 ;
  assign n655 = n654 ^ n653 ;
  assign n661 = n660 ^ n655 ;
  assign n632 = x282 ^ x122 ;
  assign n631 = x283 ^ x123 ;
  assign n633 = n632 ^ n631 ;
  assign n630 = x284 ^ x124 ;
  assign n634 = n633 ^ n630 ;
  assign n628 = x281 ^ x121 ;
  assign n625 = x285 ^ x125 ;
  assign n624 = x286 ^ x126 ;
  assign n626 = n625 ^ n624 ;
  assign n623 = x287 ^ x127 ;
  assign n627 = n626 ^ n623 ;
  assign n629 = n628 ^ n627 ;
  assign n647 = n634 ^ n629 ;
  assign n646 = x273 ^ x113 ;
  assign n648 = n647 ^ n646 ;
  assign n692 = n661 ^ n648 ;
  assign n694 = n693 ^ n692 ;
  assign n723 = n722 ^ n707 ;
  assign n724 = n723 ^ n693 ;
  assign n725 = n694 & ~n724 ;
  assign n726 = n725 ^ n692 ;
  assign n673 = n659 ^ n657 ;
  assign n674 = n658 & ~n673 ;
  assign n675 = n674 ^ n656 ;
  assign n669 = n652 ^ n650 ;
  assign n670 = n651 & ~n669 ;
  assign n671 = n670 ^ n649 ;
  assign n666 = n660 ^ n654 ;
  assign n667 = n655 & ~n666 ;
  assign n668 = n667 ^ n653 ;
  assign n672 = n671 ^ n668 ;
  assign n676 = n675 ^ n672 ;
  assign n662 = n661 ^ n647 ;
  assign n663 = n648 & ~n662 ;
  assign n664 = n663 ^ n646 ;
  assign n642 = n631 ^ n630 ;
  assign n643 = ~n633 & n642 ;
  assign n644 = n643 ^ n630 ;
  assign n638 = n624 ^ n623 ;
  assign n639 = ~n626 & n638 ;
  assign n640 = n639 ^ n623 ;
  assign n635 = n634 ^ n628 ;
  assign n636 = n629 & ~n635 ;
  assign n637 = n636 ^ n627 ;
  assign n641 = n640 ^ n637 ;
  assign n645 = n644 ^ n641 ;
  assign n665 = n664 ^ n645 ;
  assign n691 = n676 ^ n665 ;
  assign n727 = n726 ^ n691 ;
  assign n754 = n753 ^ n738 ;
  assign n755 = n754 ^ n691 ;
  assign n756 = n727 & ~n755 ;
  assign n757 = n756 ^ n726 ;
  assign n684 = n675 ^ n671 ;
  assign n685 = n672 & ~n684 ;
  assign n686 = n685 ^ n668 ;
  assign n680 = n644 ^ n640 ;
  assign n681 = n641 & ~n680 ;
  assign n682 = n681 ^ n637 ;
  assign n677 = n676 ^ n664 ;
  assign n678 = n665 & ~n677 ;
  assign n679 = n678 ^ n645 ;
  assign n683 = n682 ^ n679 ;
  assign n690 = n686 ^ n683 ;
  assign n758 = n757 ^ n690 ;
  assign n769 = n768 ^ n761 ;
  assign n770 = n769 ^ n757 ;
  assign n771 = n758 & ~n770 ;
  assign n772 = n771 ^ n690 ;
  assign n687 = n686 ^ n682 ;
  assign n688 = n683 & ~n687 ;
  assign n689 = n688 ^ n679 ;
  assign n773 = n772 ^ n689 ;
  assign n777 = n776 ^ n773 ;
  assign n778 = n754 ^ n727 ;
  assign n779 = n723 ^ n694 ;
  assign n780 = x256 ^ x96 ;
  assign n781 = n779 & n780 ;
  assign n782 = n778 & n781 ;
  assign n783 = n769 ^ n758 ;
  assign n784 = n782 & n783 ;
  assign n785 = n777 & n784 ;
  assign n786 = n776 ^ n772 ;
  assign n787 = n773 & ~n786 ;
  assign n788 = n787 ^ n689 ;
  assign n789 = n785 & n788 ;
  assign n888 = x258 ^ x162 ;
  assign n885 = x266 ^ x170 ;
  assign n883 = x272 ^ x176 ;
  assign n881 = x270 ^ x174 ;
  assign n880 = x271 ^ x175 ;
  assign n882 = n881 ^ n880 ;
  assign n884 = n883 ^ n882 ;
  assign n886 = n885 ^ n884 ;
  assign n878 = x269 ^ x173 ;
  assign n876 = x267 ^ x171 ;
  assign n875 = x268 ^ x172 ;
  assign n877 = n876 ^ n875 ;
  assign n879 = n878 ^ n877 ;
  assign n887 = n886 ^ n879 ;
  assign n889 = n888 ^ n887 ;
  assign n872 = x259 ^ x163 ;
  assign n870 = x265 ^ x169 ;
  assign n868 = x263 ^ x167 ;
  assign n867 = x264 ^ x168 ;
  assign n869 = n868 ^ n867 ;
  assign n871 = n870 ^ n869 ;
  assign n873 = n872 ^ n871 ;
  assign n865 = x262 ^ x166 ;
  assign n863 = x260 ^ x164 ;
  assign n862 = x261 ^ x165 ;
  assign n864 = n863 ^ n862 ;
  assign n866 = n865 ^ n864 ;
  assign n874 = n873 ^ n866 ;
  assign n917 = n888 ^ n874 ;
  assign n918 = n889 & ~n917 ;
  assign n919 = n918 ^ n887 ;
  assign n913 = n878 ^ n876 ;
  assign n914 = n877 & ~n913 ;
  assign n915 = n914 ^ n875 ;
  assign n909 = n883 ^ n881 ;
  assign n910 = n882 & ~n909 ;
  assign n911 = n910 ^ n880 ;
  assign n906 = n884 ^ n879 ;
  assign n907 = ~n886 & n906 ;
  assign n908 = n907 ^ n879 ;
  assign n912 = n911 ^ n908 ;
  assign n916 = n915 ^ n912 ;
  assign n920 = n919 ^ n916 ;
  assign n902 = n865 ^ n863 ;
  assign n903 = n864 & ~n902 ;
  assign n904 = n903 ^ n862 ;
  assign n898 = n871 ^ n866 ;
  assign n899 = ~n873 & n898 ;
  assign n900 = n899 ^ n866 ;
  assign n895 = n870 ^ n868 ;
  assign n896 = n869 & ~n895 ;
  assign n897 = n896 ^ n867 ;
  assign n901 = n900 ^ n897 ;
  assign n905 = n904 ^ n901 ;
  assign n932 = n919 ^ n905 ;
  assign n933 = n920 & ~n932 ;
  assign n934 = n933 ^ n916 ;
  assign n929 = n915 ^ n911 ;
  assign n930 = n912 & ~n929 ;
  assign n931 = n930 ^ n908 ;
  assign n935 = n934 ^ n931 ;
  assign n926 = n904 ^ n900 ;
  assign n927 = n901 & ~n926 ;
  assign n928 = n927 ^ n897 ;
  assign n941 = n931 ^ n928 ;
  assign n942 = ~n935 & n941 ;
  assign n943 = n942 ^ n928 ;
  assign n860 = x257 ^ x161 ;
  assign n826 = x277 ^ x181 ;
  assign n824 = x275 ^ x179 ;
  assign n823 = x276 ^ x180 ;
  assign n825 = n824 ^ n823 ;
  assign n827 = n826 ^ n825 ;
  assign n821 = x274 ^ x178 ;
  assign n819 = x280 ^ x184 ;
  assign n817 = x278 ^ x182 ;
  assign n816 = x279 ^ x183 ;
  assign n818 = n817 ^ n816 ;
  assign n820 = n819 ^ n818 ;
  assign n822 = n821 ^ n820 ;
  assign n828 = n827 ^ n822 ;
  assign n799 = x282 ^ x186 ;
  assign n798 = x283 ^ x187 ;
  assign n800 = n799 ^ n798 ;
  assign n797 = x284 ^ x188 ;
  assign n801 = n800 ^ n797 ;
  assign n795 = x281 ^ x185 ;
  assign n792 = x285 ^ x189 ;
  assign n791 = x286 ^ x190 ;
  assign n793 = n792 ^ n791 ;
  assign n790 = x287 ^ x191 ;
  assign n794 = n793 ^ n790 ;
  assign n796 = n795 ^ n794 ;
  assign n814 = n801 ^ n796 ;
  assign n813 = x273 ^ x177 ;
  assign n815 = n814 ^ n813 ;
  assign n859 = n828 ^ n815 ;
  assign n861 = n860 ^ n859 ;
  assign n890 = n889 ^ n874 ;
  assign n891 = n890 ^ n860 ;
  assign n892 = n861 & ~n891 ;
  assign n893 = n892 ^ n859 ;
  assign n840 = n826 ^ n824 ;
  assign n841 = n825 & ~n840 ;
  assign n842 = n841 ^ n823 ;
  assign n836 = n819 ^ n817 ;
  assign n837 = n818 & ~n836 ;
  assign n838 = n837 ^ n816 ;
  assign n833 = n827 ^ n821 ;
  assign n834 = n822 & ~n833 ;
  assign n835 = n834 ^ n820 ;
  assign n839 = n838 ^ n835 ;
  assign n843 = n842 ^ n839 ;
  assign n829 = n828 ^ n814 ;
  assign n830 = n815 & ~n829 ;
  assign n831 = n830 ^ n813 ;
  assign n809 = n798 ^ n797 ;
  assign n810 = ~n800 & n809 ;
  assign n811 = n810 ^ n797 ;
  assign n805 = n791 ^ n790 ;
  assign n806 = ~n793 & n805 ;
  assign n807 = n806 ^ n790 ;
  assign n802 = n801 ^ n795 ;
  assign n803 = n796 & ~n802 ;
  assign n804 = n803 ^ n794 ;
  assign n808 = n807 ^ n804 ;
  assign n812 = n811 ^ n808 ;
  assign n832 = n831 ^ n812 ;
  assign n858 = n843 ^ n832 ;
  assign n894 = n893 ^ n858 ;
  assign n921 = n920 ^ n905 ;
  assign n922 = n921 ^ n858 ;
  assign n923 = n894 & ~n922 ;
  assign n924 = n923 ^ n893 ;
  assign n851 = n842 ^ n838 ;
  assign n852 = n839 & ~n851 ;
  assign n853 = n852 ^ n835 ;
  assign n847 = n811 ^ n807 ;
  assign n848 = n808 & ~n847 ;
  assign n849 = n848 ^ n804 ;
  assign n844 = n843 ^ n831 ;
  assign n845 = n832 & ~n844 ;
  assign n846 = n845 ^ n812 ;
  assign n850 = n849 ^ n846 ;
  assign n857 = n853 ^ n850 ;
  assign n925 = n924 ^ n857 ;
  assign n936 = n935 ^ n928 ;
  assign n937 = n936 ^ n924 ;
  assign n938 = n925 & ~n937 ;
  assign n939 = n938 ^ n857 ;
  assign n854 = n853 ^ n849 ;
  assign n855 = n850 & ~n854 ;
  assign n856 = n855 ^ n846 ;
  assign n940 = n939 ^ n856 ;
  assign n944 = n943 ^ n940 ;
  assign n945 = n921 ^ n894 ;
  assign n946 = n890 ^ n861 ;
  assign n947 = x256 ^ x160 ;
  assign n948 = n946 & n947 ;
  assign n949 = n945 & n948 ;
  assign n950 = n936 ^ n925 ;
  assign n951 = n949 & n950 ;
  assign n952 = n944 & n951 ;
  assign n953 = n943 ^ n939 ;
  assign n954 = n940 & ~n953 ;
  assign n955 = n954 ^ n856 ;
  assign n956 = n952 & n955 ;
  assign n1032 = x280 ^ x216 ;
  assign n1030 = x279 ^ x215 ;
  assign n1029 = x278 ^ x214 ;
  assign n1031 = n1030 ^ n1029 ;
  assign n1037 = n1032 ^ n1031 ;
  assign n1036 = x274 ^ x210 ;
  assign n1038 = n1037 ^ n1036 ;
  assign n1025 = x277 ^ x213 ;
  assign n1023 = x275 ^ x211 ;
  assign n1022 = x276 ^ x212 ;
  assign n1024 = n1023 ^ n1022 ;
  assign n1039 = n1025 ^ n1024 ;
  assign n1040 = n1039 ^ n1037 ;
  assign n1041 = n1038 & ~n1040 ;
  assign n1042 = n1041 ^ n1036 ;
  assign n1033 = n1032 ^ n1030 ;
  assign n1034 = n1031 & ~n1033 ;
  assign n1035 = n1034 ^ n1029 ;
  assign n1043 = n1042 ^ n1035 ;
  assign n1026 = n1025 ^ n1023 ;
  assign n1027 = n1024 & ~n1026 ;
  assign n1028 = n1027 ^ n1022 ;
  assign n1096 = n1042 ^ n1028 ;
  assign n1097 = n1043 & n1096 ;
  assign n1098 = n1097 ^ n1042 ;
  assign n1057 = x283 ^ x219 ;
  assign n1056 = x282 ^ x218 ;
  assign n1058 = n1057 ^ n1056 ;
  assign n1055 = x284 ^ x220 ;
  assign n1059 = n1058 ^ n1055 ;
  assign n1048 = x287 ^ x223 ;
  assign n1046 = x286 ^ x222 ;
  assign n1045 = x285 ^ x221 ;
  assign n1047 = n1046 ^ n1045 ;
  assign n1053 = n1048 ^ n1047 ;
  assign n1052 = x281 ^ x217 ;
  assign n1054 = n1053 ^ n1052 ;
  assign n1069 = n1059 ^ n1054 ;
  assign n1068 = x273 ^ x209 ;
  assign n1070 = n1069 ^ n1068 ;
  assign n1071 = n1039 ^ n1038 ;
  assign n1072 = n1071 ^ n1068 ;
  assign n1073 = ~n1070 & n1072 ;
  assign n1074 = n1073 ^ n1071 ;
  assign n1064 = n1057 ^ n1055 ;
  assign n1065 = n1058 & ~n1064 ;
  assign n1066 = n1065 ^ n1056 ;
  assign n1060 = n1059 ^ n1052 ;
  assign n1061 = ~n1054 & n1060 ;
  assign n1062 = n1061 ^ n1059 ;
  assign n1049 = n1048 ^ n1046 ;
  assign n1050 = n1047 & ~n1049 ;
  assign n1051 = n1050 ^ n1045 ;
  assign n1063 = n1062 ^ n1051 ;
  assign n1067 = n1066 ^ n1063 ;
  assign n1075 = n1074 ^ n1067 ;
  assign n1044 = n1043 ^ n1028 ;
  assign n1092 = n1067 ^ n1044 ;
  assign n1093 = ~n1075 & n1092 ;
  assign n1094 = n1093 ^ n1044 ;
  assign n1089 = n1066 ^ n1051 ;
  assign n1090 = ~n1063 & n1089 ;
  assign n1091 = n1090 ^ n1066 ;
  assign n1095 = n1094 ^ n1091 ;
  assign n1099 = n1098 ^ n1095 ;
  assign n1078 = n1071 ^ n1070 ;
  assign n1077 = x257 ^ x193 ;
  assign n1079 = n1078 ^ n1077 ;
  assign n993 = x262 ^ x198 ;
  assign n991 = x260 ^ x196 ;
  assign n990 = x261 ^ x197 ;
  assign n992 = n991 ^ n990 ;
  assign n994 = n993 ^ n992 ;
  assign n988 = x259 ^ x195 ;
  assign n983 = x265 ^ x201 ;
  assign n981 = x263 ^ x199 ;
  assign n980 = x264 ^ x200 ;
  assign n982 = n981 ^ n980 ;
  assign n987 = n983 ^ n982 ;
  assign n989 = n988 ^ n987 ;
  assign n1007 = n994 ^ n989 ;
  assign n967 = x269 ^ x205 ;
  assign n965 = x267 ^ x203 ;
  assign n964 = x268 ^ x204 ;
  assign n966 = n965 ^ n964 ;
  assign n968 = n967 ^ n966 ;
  assign n962 = x266 ^ x202 ;
  assign n960 = x272 ^ x208 ;
  assign n958 = x270 ^ x206 ;
  assign n957 = x271 ^ x207 ;
  assign n959 = n958 ^ n957 ;
  assign n961 = n960 ^ n959 ;
  assign n963 = n962 ^ n961 ;
  assign n1005 = n968 ^ n963 ;
  assign n1004 = x258 ^ x194 ;
  assign n1006 = n1005 ^ n1004 ;
  assign n1080 = n1007 ^ n1006 ;
  assign n1081 = n1080 ^ n1078 ;
  assign n1082 = n1079 & ~n1081 ;
  assign n1083 = n1082 ^ n1077 ;
  assign n1076 = n1075 ^ n1044 ;
  assign n1084 = n1083 ^ n1076 ;
  assign n1008 = n1007 ^ n1005 ;
  assign n1009 = n1006 & ~n1008 ;
  assign n1010 = n1009 ^ n1004 ;
  assign n999 = n993 ^ n991 ;
  assign n1000 = n992 & ~n999 ;
  assign n1001 = n1000 ^ n990 ;
  assign n995 = n994 ^ n987 ;
  assign n996 = ~n989 & n995 ;
  assign n997 = n996 ^ n994 ;
  assign n984 = n983 ^ n981 ;
  assign n985 = n982 & ~n984 ;
  assign n986 = n985 ^ n980 ;
  assign n998 = n997 ^ n986 ;
  assign n1002 = n1001 ^ n998 ;
  assign n976 = n967 ^ n965 ;
  assign n977 = n966 & ~n976 ;
  assign n978 = n977 ^ n964 ;
  assign n972 = n960 ^ n958 ;
  assign n973 = n959 & ~n972 ;
  assign n974 = n973 ^ n957 ;
  assign n969 = n968 ^ n961 ;
  assign n970 = ~n963 & n969 ;
  assign n971 = n970 ^ n968 ;
  assign n975 = n974 ^ n971 ;
  assign n979 = n978 ^ n975 ;
  assign n1003 = n1002 ^ n979 ;
  assign n1085 = n1010 ^ n1003 ;
  assign n1086 = n1085 ^ n1076 ;
  assign n1087 = n1084 & ~n1086 ;
  assign n1088 = n1087 ^ n1083 ;
  assign n1100 = n1099 ^ n1088 ;
  assign n1018 = n1001 ^ n997 ;
  assign n1019 = n998 & n1018 ;
  assign n1020 = n1019 ^ n997 ;
  assign n1014 = n978 ^ n974 ;
  assign n1015 = n975 & ~n1014 ;
  assign n1016 = n1015 ^ n971 ;
  assign n1011 = n1010 ^ n979 ;
  assign n1012 = ~n1003 & n1011 ;
  assign n1013 = n1012 ^ n1010 ;
  assign n1017 = n1016 ^ n1013 ;
  assign n1021 = n1020 ^ n1017 ;
  assign n1101 = n1100 ^ n1021 ;
  assign n1102 = n1085 ^ n1084 ;
  assign n1103 = x256 ^ x192 ;
  assign n1104 = n1080 ^ n1079 ;
  assign n1105 = n1103 & n1104 ;
  assign n1106 = n1102 & n1105 ;
  assign n1107 = n1101 & n1106 ;
  assign n1114 = n1088 ^ n1021 ;
  assign n1115 = ~n1100 & n1114 ;
  assign n1116 = n1115 ^ n1021 ;
  assign n1111 = n1098 ^ n1094 ;
  assign n1112 = n1095 & ~n1111 ;
  assign n1113 = n1112 ^ n1091 ;
  assign n1117 = n1116 ^ n1113 ;
  assign n1108 = n1020 ^ n1016 ;
  assign n1109 = n1017 & ~n1108 ;
  assign n1110 = n1109 ^ n1013 ;
  assign n1118 = n1117 ^ n1110 ;
  assign n1119 = n1107 & n1118 ;
  assign n1120 = n1116 ^ n1110 ;
  assign n1121 = n1117 & ~n1120 ;
  assign n1122 = n1121 ^ n1113 ;
  assign n1124 = ~n1119 & ~n1122 ;
  assign n1123 = n1122 ^ n1119 ;
  assign n1125 = n1124 ^ n1123 ;
  assign n1201 = x278 ^ x246 ;
  assign n1200 = x279 ^ x247 ;
  assign n1202 = n1201 ^ n1200 ;
  assign n1199 = x280 ^ x248 ;
  assign n1209 = n1201 ^ n1199 ;
  assign n1210 = n1202 & ~n1209 ;
  assign n1211 = n1210 ^ n1200 ;
  assign n1203 = n1202 ^ n1199 ;
  assign n1198 = x274 ^ x242 ;
  assign n1204 = n1203 ^ n1198 ;
  assign n1194 = x277 ^ x245 ;
  assign n1192 = x275 ^ x243 ;
  assign n1191 = x276 ^ x244 ;
  assign n1193 = n1192 ^ n1191 ;
  assign n1205 = n1194 ^ n1193 ;
  assign n1206 = n1205 ^ n1203 ;
  assign n1207 = n1204 & ~n1206 ;
  assign n1208 = n1207 ^ n1198 ;
  assign n1212 = n1211 ^ n1208 ;
  assign n1195 = n1194 ^ n1192 ;
  assign n1196 = n1193 & ~n1195 ;
  assign n1197 = n1196 ^ n1191 ;
  assign n1265 = n1211 ^ n1197 ;
  assign n1266 = n1212 & ~n1265 ;
  assign n1267 = n1266 ^ n1208 ;
  assign n1238 = x273 ^ x241 ;
  assign n1224 = x284 ^ x252 ;
  assign n1222 = x282 ^ x250 ;
  assign n1221 = x283 ^ x251 ;
  assign n1223 = n1222 ^ n1221 ;
  assign n1225 = n1224 ^ n1223 ;
  assign n1218 = x287 ^ x255 ;
  assign n1216 = x285 ^ x253 ;
  assign n1215 = x286 ^ x254 ;
  assign n1217 = n1216 ^ n1215 ;
  assign n1219 = n1218 ^ n1217 ;
  assign n1214 = x281 ^ x249 ;
  assign n1220 = n1219 ^ n1214 ;
  assign n1237 = n1225 ^ n1220 ;
  assign n1239 = n1238 ^ n1237 ;
  assign n1240 = n1205 ^ n1204 ;
  assign n1241 = n1240 ^ n1238 ;
  assign n1242 = n1239 & ~n1241 ;
  assign n1243 = n1242 ^ n1237 ;
  assign n1233 = n1224 ^ n1222 ;
  assign n1234 = n1223 & ~n1233 ;
  assign n1235 = n1234 ^ n1221 ;
  assign n1229 = n1218 ^ n1216 ;
  assign n1230 = n1217 & ~n1229 ;
  assign n1231 = n1230 ^ n1215 ;
  assign n1226 = n1225 ^ n1219 ;
  assign n1227 = n1220 & ~n1226 ;
  assign n1228 = n1227 ^ n1214 ;
  assign n1232 = n1231 ^ n1228 ;
  assign n1236 = n1235 ^ n1232 ;
  assign n1244 = n1243 ^ n1236 ;
  assign n1213 = n1212 ^ n1197 ;
  assign n1261 = n1243 ^ n1213 ;
  assign n1262 = ~n1244 & n1261 ;
  assign n1263 = n1262 ^ n1213 ;
  assign n1258 = n1235 ^ n1231 ;
  assign n1259 = n1232 & ~n1258 ;
  assign n1260 = n1259 ^ n1228 ;
  assign n1264 = n1263 ^ n1260 ;
  assign n1268 = n1267 ^ n1264 ;
  assign n1247 = x257 ^ x225 ;
  assign n1246 = n1240 ^ n1239 ;
  assign n1248 = n1247 ^ n1246 ;
  assign n1162 = x259 ^ x227 ;
  assign n1160 = x265 ^ x233 ;
  assign n1158 = x263 ^ x231 ;
  assign n1157 = x264 ^ x232 ;
  assign n1159 = n1158 ^ n1157 ;
  assign n1161 = n1160 ^ n1159 ;
  assign n1163 = n1162 ^ n1161 ;
  assign n1155 = x262 ^ x230 ;
  assign n1153 = x260 ^ x228 ;
  assign n1152 = x261 ^ x229 ;
  assign n1154 = n1153 ^ n1152 ;
  assign n1156 = n1155 ^ n1154 ;
  assign n1164 = n1163 ^ n1156 ;
  assign n1136 = x269 ^ x237 ;
  assign n1134 = x267 ^ x235 ;
  assign n1133 = x268 ^ x236 ;
  assign n1135 = n1134 ^ n1133 ;
  assign n1137 = n1136 ^ n1135 ;
  assign n1131 = x266 ^ x234 ;
  assign n1129 = x272 ^ x240 ;
  assign n1127 = x270 ^ x238 ;
  assign n1126 = x271 ^ x239 ;
  assign n1128 = n1127 ^ n1126 ;
  assign n1130 = n1129 ^ n1128 ;
  assign n1132 = n1131 ^ n1130 ;
  assign n1150 = n1137 ^ n1132 ;
  assign n1149 = x258 ^ x226 ;
  assign n1151 = n1150 ^ n1149 ;
  assign n1249 = n1164 ^ n1151 ;
  assign n1250 = n1249 ^ n1247 ;
  assign n1251 = n1248 & ~n1250 ;
  assign n1252 = n1251 ^ n1246 ;
  assign n1245 = n1244 ^ n1213 ;
  assign n1253 = n1252 ^ n1245 ;
  assign n1176 = n1155 ^ n1153 ;
  assign n1177 = n1154 & ~n1176 ;
  assign n1178 = n1177 ^ n1152 ;
  assign n1172 = n1161 ^ n1156 ;
  assign n1173 = ~n1163 & n1172 ;
  assign n1174 = n1173 ^ n1156 ;
  assign n1169 = n1160 ^ n1158 ;
  assign n1170 = n1159 & ~n1169 ;
  assign n1171 = n1170 ^ n1157 ;
  assign n1175 = n1174 ^ n1171 ;
  assign n1179 = n1178 ^ n1175 ;
  assign n1165 = n1164 ^ n1150 ;
  assign n1166 = n1151 & ~n1165 ;
  assign n1167 = n1166 ^ n1149 ;
  assign n1145 = n1136 ^ n1134 ;
  assign n1146 = n1135 & ~n1145 ;
  assign n1147 = n1146 ^ n1133 ;
  assign n1141 = n1129 ^ n1127 ;
  assign n1142 = n1128 & ~n1141 ;
  assign n1143 = n1142 ^ n1126 ;
  assign n1138 = n1137 ^ n1130 ;
  assign n1139 = ~n1132 & n1138 ;
  assign n1140 = n1139 ^ n1137 ;
  assign n1144 = n1143 ^ n1140 ;
  assign n1148 = n1147 ^ n1144 ;
  assign n1168 = n1167 ^ n1148 ;
  assign n1254 = n1179 ^ n1168 ;
  assign n1255 = n1254 ^ n1245 ;
  assign n1256 = n1253 & ~n1255 ;
  assign n1257 = n1256 ^ n1252 ;
  assign n1269 = n1268 ^ n1257 ;
  assign n1187 = n1178 ^ n1174 ;
  assign n1188 = n1175 & ~n1187 ;
  assign n1189 = n1188 ^ n1171 ;
  assign n1183 = n1147 ^ n1143 ;
  assign n1184 = n1144 & ~n1183 ;
  assign n1185 = n1184 ^ n1140 ;
  assign n1180 = n1179 ^ n1148 ;
  assign n1181 = n1168 & ~n1180 ;
  assign n1182 = n1181 ^ n1167 ;
  assign n1186 = n1185 ^ n1182 ;
  assign n1190 = n1189 ^ n1186 ;
  assign n1270 = n1269 ^ n1190 ;
  assign n1271 = n1249 ^ n1248 ;
  assign n1272 = x256 ^ x224 ;
  assign n1273 = n1271 & n1272 ;
  assign n1274 = n1254 ^ n1253 ;
  assign n1275 = n1273 & n1274 ;
  assign n1276 = n1270 & n1275 ;
  assign n1283 = n1257 ^ n1190 ;
  assign n1284 = ~n1269 & n1283 ;
  assign n1285 = n1284 ^ n1190 ;
  assign n1280 = n1267 ^ n1260 ;
  assign n1281 = n1264 & n1280 ;
  assign n1282 = n1281 ^ n1260 ;
  assign n1286 = n1285 ^ n1282 ;
  assign n1277 = n1189 ^ n1185 ;
  assign n1278 = n1186 & ~n1277 ;
  assign n1279 = n1278 ^ n1182 ;
  assign n1287 = n1286 ^ n1279 ;
  assign n1288 = n1276 & n1287 ;
  assign n1289 = n1285 ^ n1279 ;
  assign n1290 = n1286 & ~n1289 ;
  assign n1291 = n1290 ^ n1282 ;
  assign n1293 = ~n1288 & ~n1291 ;
  assign n1292 = n1291 ^ n1288 ;
  assign n1294 = n1293 ^ n1292 ;
  assign n1296 = ~n1125 & n1294 ;
  assign n1295 = n1294 ^ n1125 ;
  assign n1297 = n1296 ^ n1295 ;
  assign n1298 = n1297 ^ n1294 ;
  assign n1299 = n956 & ~n1298 ;
  assign n1398 = x258 ^ x130 ;
  assign n1395 = x266 ^ x138 ;
  assign n1393 = x272 ^ x144 ;
  assign n1391 = x270 ^ x142 ;
  assign n1390 = x271 ^ x143 ;
  assign n1392 = n1391 ^ n1390 ;
  assign n1394 = n1393 ^ n1392 ;
  assign n1396 = n1395 ^ n1394 ;
  assign n1388 = x269 ^ x141 ;
  assign n1386 = x267 ^ x139 ;
  assign n1385 = x268 ^ x140 ;
  assign n1387 = n1386 ^ n1385 ;
  assign n1389 = n1388 ^ n1387 ;
  assign n1397 = n1396 ^ n1389 ;
  assign n1399 = n1398 ^ n1397 ;
  assign n1382 = x259 ^ x131 ;
  assign n1380 = x265 ^ x137 ;
  assign n1378 = x263 ^ x135 ;
  assign n1377 = x264 ^ x136 ;
  assign n1379 = n1378 ^ n1377 ;
  assign n1381 = n1380 ^ n1379 ;
  assign n1383 = n1382 ^ n1381 ;
  assign n1375 = x262 ^ x134 ;
  assign n1373 = x260 ^ x132 ;
  assign n1372 = x261 ^ x133 ;
  assign n1374 = n1373 ^ n1372 ;
  assign n1376 = n1375 ^ n1374 ;
  assign n1384 = n1383 ^ n1376 ;
  assign n1427 = n1398 ^ n1384 ;
  assign n1428 = n1399 & ~n1427 ;
  assign n1429 = n1428 ^ n1397 ;
  assign n1423 = n1388 ^ n1386 ;
  assign n1424 = n1387 & ~n1423 ;
  assign n1425 = n1424 ^ n1385 ;
  assign n1419 = n1393 ^ n1391 ;
  assign n1420 = n1392 & ~n1419 ;
  assign n1421 = n1420 ^ n1390 ;
  assign n1416 = n1394 ^ n1389 ;
  assign n1417 = ~n1396 & n1416 ;
  assign n1418 = n1417 ^ n1389 ;
  assign n1422 = n1421 ^ n1418 ;
  assign n1426 = n1425 ^ n1422 ;
  assign n1430 = n1429 ^ n1426 ;
  assign n1412 = n1375 ^ n1373 ;
  assign n1413 = n1374 & ~n1412 ;
  assign n1414 = n1413 ^ n1372 ;
  assign n1408 = n1381 ^ n1376 ;
  assign n1409 = ~n1383 & n1408 ;
  assign n1410 = n1409 ^ n1376 ;
  assign n1405 = n1380 ^ n1378 ;
  assign n1406 = n1379 & ~n1405 ;
  assign n1407 = n1406 ^ n1377 ;
  assign n1411 = n1410 ^ n1407 ;
  assign n1415 = n1414 ^ n1411 ;
  assign n1442 = n1429 ^ n1415 ;
  assign n1443 = n1430 & ~n1442 ;
  assign n1444 = n1443 ^ n1426 ;
  assign n1439 = n1425 ^ n1421 ;
  assign n1440 = n1422 & ~n1439 ;
  assign n1441 = n1440 ^ n1418 ;
  assign n1445 = n1444 ^ n1441 ;
  assign n1436 = n1414 ^ n1410 ;
  assign n1437 = n1411 & ~n1436 ;
  assign n1438 = n1437 ^ n1407 ;
  assign n1451 = n1441 ^ n1438 ;
  assign n1452 = ~n1445 & n1451 ;
  assign n1453 = n1452 ^ n1438 ;
  assign n1370 = x257 ^ x129 ;
  assign n1336 = x277 ^ x149 ;
  assign n1334 = x275 ^ x147 ;
  assign n1333 = x276 ^ x148 ;
  assign n1335 = n1334 ^ n1333 ;
  assign n1337 = n1336 ^ n1335 ;
  assign n1331 = x274 ^ x146 ;
  assign n1329 = x280 ^ x152 ;
  assign n1327 = x278 ^ x150 ;
  assign n1326 = x279 ^ x151 ;
  assign n1328 = n1327 ^ n1326 ;
  assign n1330 = n1329 ^ n1328 ;
  assign n1332 = n1331 ^ n1330 ;
  assign n1338 = n1337 ^ n1332 ;
  assign n1309 = x282 ^ x154 ;
  assign n1308 = x283 ^ x155 ;
  assign n1310 = n1309 ^ n1308 ;
  assign n1307 = x284 ^ x156 ;
  assign n1311 = n1310 ^ n1307 ;
  assign n1305 = x281 ^ x153 ;
  assign n1302 = x285 ^ x157 ;
  assign n1301 = x286 ^ x158 ;
  assign n1303 = n1302 ^ n1301 ;
  assign n1300 = x287 ^ x159 ;
  assign n1304 = n1303 ^ n1300 ;
  assign n1306 = n1305 ^ n1304 ;
  assign n1324 = n1311 ^ n1306 ;
  assign n1323 = x273 ^ x145 ;
  assign n1325 = n1324 ^ n1323 ;
  assign n1369 = n1338 ^ n1325 ;
  assign n1371 = n1370 ^ n1369 ;
  assign n1400 = n1399 ^ n1384 ;
  assign n1401 = n1400 ^ n1370 ;
  assign n1402 = n1371 & ~n1401 ;
  assign n1403 = n1402 ^ n1369 ;
  assign n1350 = n1336 ^ n1334 ;
  assign n1351 = n1335 & ~n1350 ;
  assign n1352 = n1351 ^ n1333 ;
  assign n1346 = n1329 ^ n1327 ;
  assign n1347 = n1328 & ~n1346 ;
  assign n1348 = n1347 ^ n1326 ;
  assign n1343 = n1337 ^ n1331 ;
  assign n1344 = n1332 & ~n1343 ;
  assign n1345 = n1344 ^ n1330 ;
  assign n1349 = n1348 ^ n1345 ;
  assign n1353 = n1352 ^ n1349 ;
  assign n1339 = n1338 ^ n1324 ;
  assign n1340 = n1325 & ~n1339 ;
  assign n1341 = n1340 ^ n1323 ;
  assign n1319 = n1308 ^ n1307 ;
  assign n1320 = ~n1310 & n1319 ;
  assign n1321 = n1320 ^ n1307 ;
  assign n1315 = n1301 ^ n1300 ;
  assign n1316 = ~n1303 & n1315 ;
  assign n1317 = n1316 ^ n1300 ;
  assign n1312 = n1311 ^ n1305 ;
  assign n1313 = n1306 & ~n1312 ;
  assign n1314 = n1313 ^ n1304 ;
  assign n1318 = n1317 ^ n1314 ;
  assign n1322 = n1321 ^ n1318 ;
  assign n1342 = n1341 ^ n1322 ;
  assign n1368 = n1353 ^ n1342 ;
  assign n1404 = n1403 ^ n1368 ;
  assign n1431 = n1430 ^ n1415 ;
  assign n1432 = n1431 ^ n1368 ;
  assign n1433 = n1404 & ~n1432 ;
  assign n1434 = n1433 ^ n1403 ;
  assign n1361 = n1352 ^ n1348 ;
  assign n1362 = n1349 & ~n1361 ;
  assign n1363 = n1362 ^ n1345 ;
  assign n1357 = n1321 ^ n1317 ;
  assign n1358 = n1318 & ~n1357 ;
  assign n1359 = n1358 ^ n1314 ;
  assign n1354 = n1353 ^ n1341 ;
  assign n1355 = n1342 & ~n1354 ;
  assign n1356 = n1355 ^ n1322 ;
  assign n1360 = n1359 ^ n1356 ;
  assign n1367 = n1363 ^ n1360 ;
  assign n1435 = n1434 ^ n1367 ;
  assign n1446 = n1445 ^ n1438 ;
  assign n1447 = n1446 ^ n1434 ;
  assign n1448 = n1435 & ~n1447 ;
  assign n1449 = n1448 ^ n1367 ;
  assign n1364 = n1363 ^ n1359 ;
  assign n1365 = n1360 & ~n1364 ;
  assign n1366 = n1365 ^ n1356 ;
  assign n1450 = n1449 ^ n1366 ;
  assign n1454 = n1453 ^ n1450 ;
  assign n1455 = n1431 ^ n1404 ;
  assign n1456 = n1400 ^ n1371 ;
  assign n1457 = x256 ^ x128 ;
  assign n1458 = n1456 & n1457 ;
  assign n1459 = n1455 & n1458 ;
  assign n1460 = n1446 ^ n1435 ;
  assign n1461 = n1459 & n1460 ;
  assign n1462 = n1454 & n1461 ;
  assign n1463 = n1453 ^ n1449 ;
  assign n1464 = n1450 & ~n1463 ;
  assign n1465 = n1464 ^ n1366 ;
  assign n1466 = n1462 & n1465 ;
  assign n1467 = n1299 & ~n1466 ;
  assign n1468 = n1467 ^ n1299 ;
  assign n1469 = n789 & n1468 ;
  assign n1471 = ~n622 & n1469 ;
  assign n1470 = n1469 ^ n622 ;
  assign n1472 = n1471 ^ n1470 ;
  assign n1473 = n1472 ^ n622 ;
  assign n1474 = n455 & n1473 ;
  assign n1642 = n1641 ^ n1474 ;
  assign n1859 = n1640 ^ n1637 ;
  assign n1649 = n955 ^ n952 ;
  assign n1647 = ~n1124 & ~n1293 ;
  assign n1648 = n1647 ^ n1298 ;
  assign n1650 = n1649 ^ n1648 ;
  assign n1651 = n1298 ^ n956 ;
  assign n1710 = n1649 ^ n956 ;
  assign n1654 = n1287 ^ n1276 ;
  assign n1653 = n1118 ^ n1107 ;
  assign n1655 = n1654 ^ n1653 ;
  assign n1656 = n1292 ^ n1123 ;
  assign n1666 = n1106 ^ n1101 ;
  assign n1658 = n1274 ^ n1273 ;
  assign n1657 = n1105 ^ n1102 ;
  assign n1659 = n1658 ^ n1657 ;
  assign n1660 = n1272 ^ n1271 ;
  assign n1661 = n1104 ^ n1103 ;
  assign n1662 = ~n1660 & n1661 ;
  assign n1663 = n1662 ^ n1657 ;
  assign n1664 = n1659 & n1663 ;
  assign n1665 = n1664 ^ n1662 ;
  assign n1667 = n1666 ^ n1665 ;
  assign n1668 = n1275 ^ n1270 ;
  assign n1669 = n1668 ^ n1665 ;
  assign n1670 = n1667 & n1669 ;
  assign n1671 = n1670 ^ n1666 ;
  assign n1672 = n1671 ^ n1653 ;
  assign n1673 = n1671 ^ n1654 ;
  assign n1674 = n1672 & n1673 ;
  assign n1675 = n1674 ^ n1653 ;
  assign n1676 = n1675 ^ n1292 ;
  assign n1677 = ~n1656 & ~n1676 ;
  assign n1678 = n1677 ^ n1292 ;
  assign n1679 = n1678 ^ n1294 ;
  assign n1680 = ~n1295 & n1679 ;
  assign n1681 = n1680 ^ n1125 ;
  assign n1682 = n1655 & ~n1681 ;
  assign n1683 = n1682 ^ n1653 ;
  assign n1652 = n951 ^ n944 ;
  assign n1684 = n1683 ^ n1652 ;
  assign n1688 = n950 ^ n949 ;
  assign n1685 = n1668 ^ n1666 ;
  assign n1686 = ~n1681 & n1685 ;
  assign n1687 = n1686 ^ n1666 ;
  assign n1689 = n1688 ^ n1687 ;
  assign n1692 = n948 ^ n945 ;
  assign n1690 = n1659 & ~n1681 ;
  assign n1691 = n1690 ^ n1657 ;
  assign n1693 = n1692 ^ n1691 ;
  assign n1694 = n947 ^ n946 ;
  assign n1695 = n1661 ^ n1660 ;
  assign n1696 = n1681 & n1695 ;
  assign n1697 = n1696 ^ n1660 ;
  assign n1698 = n1694 & ~n1697 ;
  assign n1699 = n1698 ^ n1691 ;
  assign n1700 = ~n1693 & ~n1699 ;
  assign n1701 = n1700 ^ n1691 ;
  assign n1702 = n1701 ^ n1687 ;
  assign n1703 = ~n1689 & n1702 ;
  assign n1704 = n1703 ^ n1687 ;
  assign n1705 = n1704 ^ n1652 ;
  assign n1706 = ~n1684 & ~n1705 ;
  assign n1707 = n1706 ^ n1652 ;
  assign n1708 = n1707 ^ n1648 ;
  assign n1709 = n1650 & ~n1708 ;
  assign n1711 = n1710 ^ n1709 ;
  assign n1712 = n1651 & ~n1711 ;
  assign n1713 = n1712 ^ n1298 ;
  assign n1714 = ~n1650 & n1713 ;
  assign n1715 = n1714 ^ n1649 ;
  assign n1646 = n1465 ^ n1462 ;
  assign n1716 = n1715 ^ n1646 ;
  assign n1717 = ~n1646 & n1715 ;
  assign n1718 = n1717 ^ n1467 ;
  assign n1719 = n1717 ^ n1716 ;
  assign n1721 = n1684 & n1713 ;
  assign n1722 = n1721 ^ n1652 ;
  assign n1720 = n1461 ^ n1454 ;
  assign n1723 = n1722 ^ n1720 ;
  assign n1726 = n1460 ^ n1459 ;
  assign n1724 = n1689 & n1713 ;
  assign n1725 = n1724 ^ n1688 ;
  assign n1727 = n1726 ^ n1725 ;
  assign n1730 = n1458 ^ n1455 ;
  assign n1728 = n1693 & n1713 ;
  assign n1729 = n1728 ^ n1692 ;
  assign n1731 = n1730 ^ n1729 ;
  assign n1732 = n1457 ^ n1456 ;
  assign n1733 = n1697 ^ n1694 ;
  assign n1734 = n1713 & n1733 ;
  assign n1735 = n1734 ^ n1694 ;
  assign n1736 = n1732 & ~n1735 ;
  assign n1737 = n1736 ^ n1729 ;
  assign n1738 = ~n1731 & ~n1737 ;
  assign n1739 = n1738 ^ n1729 ;
  assign n1740 = n1739 ^ n1725 ;
  assign n1741 = ~n1727 & n1740 ;
  assign n1742 = n1741 ^ n1725 ;
  assign n1743 = n1742 ^ n1720 ;
  assign n1744 = ~n1723 & ~n1743 ;
  assign n1745 = n1744 ^ n1720 ;
  assign n1746 = ~n1719 & ~n1745 ;
  assign n1747 = ~n1718 & ~n1746 ;
  assign n1748 = n1468 ^ n1466 ;
  assign n1749 = ~n1747 & ~n1748 ;
  assign n1750 = n1716 & n1749 ;
  assign n1751 = n1750 ^ n1715 ;
  assign n1645 = n788 ^ n785 ;
  assign n1752 = n1751 ^ n1645 ;
  assign n1753 = n1468 ^ n789 ;
  assign n1782 = n1645 ^ n789 ;
  assign n1755 = n1723 & ~n1749 ;
  assign n1756 = n1755 ^ n1720 ;
  assign n1754 = n784 ^ n777 ;
  assign n1757 = n1756 ^ n1754 ;
  assign n1760 = n783 ^ n782 ;
  assign n1758 = n1727 & ~n1749 ;
  assign n1759 = n1758 ^ n1726 ;
  assign n1761 = n1760 ^ n1759 ;
  assign n1764 = n781 ^ n778 ;
  assign n1762 = n1731 & ~n1749 ;
  assign n1763 = n1762 ^ n1730 ;
  assign n1765 = n1764 ^ n1763 ;
  assign n1766 = n780 ^ n779 ;
  assign n1767 = n1735 ^ n1732 ;
  assign n1768 = ~n1749 & n1767 ;
  assign n1769 = n1768 ^ n1732 ;
  assign n1770 = n1766 & ~n1769 ;
  assign n1771 = n1770 ^ n1763 ;
  assign n1772 = ~n1765 & ~n1771 ;
  assign n1773 = n1772 ^ n1763 ;
  assign n1774 = n1773 ^ n1759 ;
  assign n1775 = ~n1761 & n1774 ;
  assign n1776 = n1775 ^ n1759 ;
  assign n1777 = n1776 ^ n1754 ;
  assign n1778 = ~n1757 & ~n1777 ;
  assign n1779 = n1778 ^ n1754 ;
  assign n1780 = n1779 ^ n1751 ;
  assign n1781 = ~n1752 & n1780 ;
  assign n1783 = n1782 ^ n1781 ;
  assign n1784 = ~n1753 & ~n1783 ;
  assign n1785 = n1784 ^ n1468 ;
  assign n1786 = n1752 & n1785 ;
  assign n1787 = n1786 ^ n1751 ;
  assign n1644 = n621 ^ n618 ;
  assign n1788 = n1787 ^ n1644 ;
  assign n1789 = ~n1644 & n1787 ;
  assign n1790 = n1789 ^ n1471 ;
  assign n1791 = n1789 ^ n1788 ;
  assign n1793 = n1757 & ~n1785 ;
  assign n1794 = n1793 ^ n1754 ;
  assign n1792 = n617 ^ n610 ;
  assign n1795 = n1794 ^ n1792 ;
  assign n1798 = n616 ^ n615 ;
  assign n1796 = n1761 & ~n1785 ;
  assign n1797 = n1796 ^ n1760 ;
  assign n1799 = n1798 ^ n1797 ;
  assign n1802 = n614 ^ n613 ;
  assign n1800 = n1765 & ~n1785 ;
  assign n1801 = n1800 ^ n1764 ;
  assign n1803 = n1802 ^ n1801 ;
  assign n1804 = n612 ^ n611 ;
  assign n1805 = n1769 ^ n1766 ;
  assign n1806 = ~n1785 & n1805 ;
  assign n1807 = n1806 ^ n1766 ;
  assign n1808 = n1804 & ~n1807 ;
  assign n1809 = n1808 ^ n1801 ;
  assign n1810 = ~n1803 & ~n1809 ;
  assign n1811 = n1810 ^ n1801 ;
  assign n1812 = n1811 ^ n1797 ;
  assign n1813 = ~n1799 & n1812 ;
  assign n1814 = n1813 ^ n1797 ;
  assign n1815 = n1814 ^ n1792 ;
  assign n1816 = ~n1795 & ~n1815 ;
  assign n1817 = n1816 ^ n1792 ;
  assign n1818 = ~n1791 & ~n1817 ;
  assign n1819 = ~n1790 & ~n1818 ;
  assign n1820 = ~n1472 & ~n1819 ;
  assign n1821 = n1788 & n1820 ;
  assign n1822 = n1821 ^ n1787 ;
  assign n1643 = n454 ^ n451 ;
  assign n1823 = n1822 ^ n1643 ;
  assign n1824 = n1473 ^ n455 ;
  assign n1853 = n1643 ^ n455 ;
  assign n1826 = n1795 & ~n1820 ;
  assign n1827 = n1826 ^ n1792 ;
  assign n1825 = n450 ^ n443 ;
  assign n1828 = n1827 ^ n1825 ;
  assign n1831 = n449 ^ n448 ;
  assign n1829 = n1799 & ~n1820 ;
  assign n1830 = n1829 ^ n1798 ;
  assign n1832 = n1831 ^ n1830 ;
  assign n1834 = n1803 & ~n1820 ;
  assign n1835 = n1834 ^ n1802 ;
  assign n1833 = n447 ^ n446 ;
  assign n1836 = n1835 ^ n1833 ;
  assign n1837 = n445 ^ n444 ;
  assign n1838 = n1807 ^ n1804 ;
  assign n1839 = ~n1820 & n1838 ;
  assign n1840 = n1839 ^ n1804 ;
  assign n1841 = n1837 & ~n1840 ;
  assign n1842 = n1841 ^ n1833 ;
  assign n1843 = ~n1836 & n1842 ;
  assign n1844 = n1843 ^ n1833 ;
  assign n1845 = n1844 ^ n1830 ;
  assign n1846 = ~n1832 & ~n1845 ;
  assign n1847 = n1846 ^ n1830 ;
  assign n1848 = n1847 ^ n1825 ;
  assign n1849 = ~n1828 & ~n1848 ;
  assign n1850 = n1849 ^ n1825 ;
  assign n1851 = n1850 ^ n1822 ;
  assign n1852 = ~n1823 & n1851 ;
  assign n1854 = n1853 ^ n1852 ;
  assign n1855 = ~n1824 & ~n1854 ;
  assign n1856 = n1855 ^ n1473 ;
  assign n1857 = n1823 & ~n1856 ;
  assign n1858 = n1857 ^ n1643 ;
  assign n1860 = n1859 ^ n1858 ;
  assign n1862 = n1828 & ~n1856 ;
  assign n1863 = n1862 ^ n1825 ;
  assign n1861 = n1636 ^ n1629 ;
  assign n1864 = n1863 ^ n1861 ;
  assign n1867 = n1635 ^ n1634 ;
  assign n1865 = n1832 & ~n1856 ;
  assign n1866 = n1865 ^ n1831 ;
  assign n1868 = n1867 ^ n1866 ;
  assign n1871 = n1633 ^ n1630 ;
  assign n1869 = n1836 & n1856 ;
  assign n1870 = n1869 ^ n1835 ;
  assign n1872 = n1871 ^ n1870 ;
  assign n1873 = n1632 ^ n1631 ;
  assign n1874 = n1840 ^ n1837 ;
  assign n1875 = n1856 & n1874 ;
  assign n1876 = n1875 ^ n1840 ;
  assign n1877 = n1873 & ~n1876 ;
  assign n1878 = n1877 ^ n1870 ;
  assign n1879 = ~n1872 & ~n1878 ;
  assign n1880 = n1879 ^ n1870 ;
  assign n1881 = n1880 ^ n1866 ;
  assign n1882 = ~n1868 & n1881 ;
  assign n1883 = n1882 ^ n1866 ;
  assign n1884 = n1883 ^ n1863 ;
  assign n1885 = ~n1864 & n1884 ;
  assign n1886 = n1885 ^ n1863 ;
  assign n1887 = n1886 ^ n1859 ;
  assign n1888 = ~n1860 & n1887 ;
  assign n1889 = n1888 ^ n1858 ;
  assign n1890 = n1889 ^ n1474 ;
  assign n1891 = ~n1642 & ~n1890 ;
  assign n1892 = n1891 ^ n1641 ;
  assign n1893 = x224 ^ x192 ;
  assign n1894 = ~n1681 & n1893 ;
  assign n1895 = n1894 ^ x192 ;
  assign n1896 = n1895 ^ x160 ;
  assign n1897 = n1713 & n1896 ;
  assign n1898 = n1897 ^ x160 ;
  assign n1899 = n1898 ^ x128 ;
  assign n1900 = ~n1749 & n1899 ;
  assign n1901 = n1900 ^ x128 ;
  assign n1902 = n1901 ^ x96 ;
  assign n1903 = ~n1785 & n1902 ;
  assign n1904 = n1903 ^ x96 ;
  assign n1905 = n1904 ^ x64 ;
  assign n1906 = ~n1820 & n1905 ;
  assign n1907 = n1906 ^ x64 ;
  assign n1908 = n1907 ^ x32 ;
  assign n1909 = ~n1856 & n1908 ;
  assign n1910 = n1909 ^ x32 ;
  assign n1911 = n1910 ^ x0 ;
  assign n1912 = n1892 & n1911 ;
  assign n1913 = n1912 ^ x0 ;
  assign n1914 = x225 ^ x193 ;
  assign n1915 = ~n1681 & n1914 ;
  assign n1916 = n1915 ^ x193 ;
  assign n1917 = n1916 ^ x161 ;
  assign n1918 = n1713 & n1917 ;
  assign n1919 = n1918 ^ x161 ;
  assign n1920 = n1919 ^ x129 ;
  assign n1921 = ~n1749 & n1920 ;
  assign n1922 = n1921 ^ x129 ;
  assign n1923 = n1922 ^ x97 ;
  assign n1924 = ~n1785 & n1923 ;
  assign n1925 = n1924 ^ x97 ;
  assign n1926 = n1925 ^ x65 ;
  assign n1927 = ~n1820 & n1926 ;
  assign n1928 = n1927 ^ x65 ;
  assign n1929 = n1928 ^ x33 ;
  assign n1930 = ~n1856 & n1929 ;
  assign n1931 = n1930 ^ x33 ;
  assign n1932 = n1931 ^ x1 ;
  assign n1933 = n1892 & n1932 ;
  assign n1934 = n1933 ^ x1 ;
  assign n1935 = x226 ^ x194 ;
  assign n1936 = ~n1681 & n1935 ;
  assign n1937 = n1936 ^ x194 ;
  assign n1938 = n1937 ^ x162 ;
  assign n1939 = n1713 & n1938 ;
  assign n1940 = n1939 ^ x162 ;
  assign n1941 = n1940 ^ x130 ;
  assign n1942 = ~n1749 & n1941 ;
  assign n1943 = n1942 ^ x130 ;
  assign n1944 = n1943 ^ x98 ;
  assign n1945 = ~n1785 & n1944 ;
  assign n1946 = n1945 ^ x98 ;
  assign n1947 = n1946 ^ x66 ;
  assign n1948 = ~n1820 & n1947 ;
  assign n1949 = n1948 ^ x66 ;
  assign n1950 = n1949 ^ x34 ;
  assign n1951 = ~n1856 & n1950 ;
  assign n1952 = n1951 ^ x34 ;
  assign n1953 = n1952 ^ x2 ;
  assign n1954 = n1892 & n1953 ;
  assign n1955 = n1954 ^ x2 ;
  assign n1956 = x227 ^ x195 ;
  assign n1957 = ~n1681 & n1956 ;
  assign n1958 = n1957 ^ x195 ;
  assign n1959 = n1958 ^ x163 ;
  assign n1960 = n1713 & n1959 ;
  assign n1961 = n1960 ^ x163 ;
  assign n1962 = n1961 ^ x131 ;
  assign n1963 = ~n1749 & n1962 ;
  assign n1964 = n1963 ^ x131 ;
  assign n1965 = n1964 ^ x99 ;
  assign n1966 = ~n1785 & n1965 ;
  assign n1967 = n1966 ^ x99 ;
  assign n1968 = n1967 ^ x67 ;
  assign n1969 = ~n1820 & n1968 ;
  assign n1970 = n1969 ^ x67 ;
  assign n1971 = n1970 ^ x35 ;
  assign n1972 = ~n1856 & n1971 ;
  assign n1973 = n1972 ^ x35 ;
  assign n1974 = n1973 ^ x3 ;
  assign n1975 = n1892 & n1974 ;
  assign n1976 = n1975 ^ x3 ;
  assign n1977 = x228 ^ x196 ;
  assign n1978 = ~n1681 & n1977 ;
  assign n1979 = n1978 ^ x196 ;
  assign n1980 = n1979 ^ x164 ;
  assign n1981 = n1713 & n1980 ;
  assign n1982 = n1981 ^ x164 ;
  assign n1983 = n1982 ^ x132 ;
  assign n1984 = ~n1749 & n1983 ;
  assign n1985 = n1984 ^ x132 ;
  assign n1986 = n1985 ^ x100 ;
  assign n1987 = ~n1785 & n1986 ;
  assign n1988 = n1987 ^ x100 ;
  assign n1989 = n1988 ^ x68 ;
  assign n1990 = ~n1820 & n1989 ;
  assign n1991 = n1990 ^ x68 ;
  assign n1992 = n1991 ^ x36 ;
  assign n1993 = ~n1856 & n1992 ;
  assign n1994 = n1993 ^ x36 ;
  assign n1995 = n1994 ^ x4 ;
  assign n1996 = n1892 & n1995 ;
  assign n1997 = n1996 ^ x4 ;
  assign n1998 = x229 ^ x197 ;
  assign n1999 = ~n1681 & n1998 ;
  assign n2000 = n1999 ^ x197 ;
  assign n2001 = n2000 ^ x165 ;
  assign n2002 = n1713 & n2001 ;
  assign n2003 = n2002 ^ x165 ;
  assign n2004 = n2003 ^ x133 ;
  assign n2005 = ~n1749 & n2004 ;
  assign n2006 = n2005 ^ x133 ;
  assign n2007 = n2006 ^ x101 ;
  assign n2008 = ~n1785 & n2007 ;
  assign n2009 = n2008 ^ x101 ;
  assign n2010 = n2009 ^ x69 ;
  assign n2011 = ~n1820 & n2010 ;
  assign n2012 = n2011 ^ x69 ;
  assign n2013 = n2012 ^ x37 ;
  assign n2014 = ~n1856 & n2013 ;
  assign n2015 = n2014 ^ x37 ;
  assign n2016 = n2015 ^ x5 ;
  assign n2017 = n1892 & n2016 ;
  assign n2018 = n2017 ^ x5 ;
  assign n2019 = x230 ^ x198 ;
  assign n2020 = ~n1681 & n2019 ;
  assign n2021 = n2020 ^ x198 ;
  assign n2022 = n2021 ^ x166 ;
  assign n2023 = n1713 & n2022 ;
  assign n2024 = n2023 ^ x166 ;
  assign n2025 = n2024 ^ x134 ;
  assign n2026 = ~n1749 & n2025 ;
  assign n2027 = n2026 ^ x134 ;
  assign n2028 = n2027 ^ x102 ;
  assign n2029 = ~n1785 & n2028 ;
  assign n2030 = n2029 ^ x102 ;
  assign n2031 = n2030 ^ x70 ;
  assign n2032 = ~n1820 & n2031 ;
  assign n2033 = n2032 ^ x70 ;
  assign n2034 = n2033 ^ x38 ;
  assign n2035 = ~n1856 & n2034 ;
  assign n2036 = n2035 ^ x38 ;
  assign n2037 = n2036 ^ x6 ;
  assign n2038 = n1892 & n2037 ;
  assign n2039 = n2038 ^ x6 ;
  assign n2040 = x231 ^ x199 ;
  assign n2041 = ~n1681 & n2040 ;
  assign n2042 = n2041 ^ x199 ;
  assign n2043 = n2042 ^ x167 ;
  assign n2044 = n1713 & n2043 ;
  assign n2045 = n2044 ^ x167 ;
  assign n2046 = n2045 ^ x135 ;
  assign n2047 = ~n1749 & n2046 ;
  assign n2048 = n2047 ^ x135 ;
  assign n2049 = n2048 ^ x103 ;
  assign n2050 = ~n1785 & n2049 ;
  assign n2051 = n2050 ^ x103 ;
  assign n2052 = n2051 ^ x71 ;
  assign n2053 = ~n1820 & n2052 ;
  assign n2054 = n2053 ^ x71 ;
  assign n2055 = n2054 ^ x39 ;
  assign n2056 = ~n1856 & n2055 ;
  assign n2057 = n2056 ^ x39 ;
  assign n2058 = n2057 ^ x7 ;
  assign n2059 = n1892 & n2058 ;
  assign n2060 = n2059 ^ x7 ;
  assign n2061 = x232 ^ x200 ;
  assign n2062 = ~n1681 & n2061 ;
  assign n2063 = n2062 ^ x200 ;
  assign n2064 = n2063 ^ x168 ;
  assign n2065 = n1713 & n2064 ;
  assign n2066 = n2065 ^ x168 ;
  assign n2067 = n2066 ^ x136 ;
  assign n2068 = ~n1749 & n2067 ;
  assign n2069 = n2068 ^ x136 ;
  assign n2070 = n2069 ^ x104 ;
  assign n2071 = ~n1785 & n2070 ;
  assign n2072 = n2071 ^ x104 ;
  assign n2073 = n2072 ^ x72 ;
  assign n2074 = ~n1820 & n2073 ;
  assign n2075 = n2074 ^ x72 ;
  assign n2076 = n2075 ^ x40 ;
  assign n2077 = ~n1856 & n2076 ;
  assign n2078 = n2077 ^ x40 ;
  assign n2079 = n2078 ^ x8 ;
  assign n2080 = n1892 & n2079 ;
  assign n2081 = n2080 ^ x8 ;
  assign n2082 = x233 ^ x201 ;
  assign n2083 = ~n1681 & n2082 ;
  assign n2084 = n2083 ^ x201 ;
  assign n2085 = n2084 ^ x169 ;
  assign n2086 = n1713 & n2085 ;
  assign n2087 = n2086 ^ x169 ;
  assign n2088 = n2087 ^ x137 ;
  assign n2089 = ~n1749 & n2088 ;
  assign n2090 = n2089 ^ x137 ;
  assign n2091 = n2090 ^ x105 ;
  assign n2092 = ~n1785 & n2091 ;
  assign n2093 = n2092 ^ x105 ;
  assign n2094 = n2093 ^ x73 ;
  assign n2095 = ~n1820 & n2094 ;
  assign n2096 = n2095 ^ x73 ;
  assign n2097 = n2096 ^ x41 ;
  assign n2098 = ~n1856 & n2097 ;
  assign n2099 = n2098 ^ x41 ;
  assign n2100 = n2099 ^ x9 ;
  assign n2101 = n1892 & n2100 ;
  assign n2102 = n2101 ^ x9 ;
  assign n2103 = x234 ^ x202 ;
  assign n2104 = ~n1681 & n2103 ;
  assign n2105 = n2104 ^ x202 ;
  assign n2106 = n2105 ^ x170 ;
  assign n2107 = n1713 & n2106 ;
  assign n2108 = n2107 ^ x170 ;
  assign n2109 = n2108 ^ x138 ;
  assign n2110 = ~n1749 & n2109 ;
  assign n2111 = n2110 ^ x138 ;
  assign n2112 = n2111 ^ x106 ;
  assign n2113 = ~n1785 & n2112 ;
  assign n2114 = n2113 ^ x106 ;
  assign n2115 = n2114 ^ x74 ;
  assign n2116 = ~n1820 & n2115 ;
  assign n2117 = n2116 ^ x74 ;
  assign n2118 = n2117 ^ x42 ;
  assign n2119 = ~n1856 & n2118 ;
  assign n2120 = n2119 ^ x42 ;
  assign n2121 = n2120 ^ x10 ;
  assign n2122 = n1892 & n2121 ;
  assign n2123 = n2122 ^ x10 ;
  assign n2124 = x235 ^ x203 ;
  assign n2125 = ~n1681 & n2124 ;
  assign n2126 = n2125 ^ x203 ;
  assign n2127 = n2126 ^ x171 ;
  assign n2128 = n1713 & n2127 ;
  assign n2129 = n2128 ^ x171 ;
  assign n2130 = n2129 ^ x139 ;
  assign n2131 = ~n1749 & n2130 ;
  assign n2132 = n2131 ^ x139 ;
  assign n2133 = n2132 ^ x107 ;
  assign n2134 = ~n1785 & n2133 ;
  assign n2135 = n2134 ^ x107 ;
  assign n2136 = n2135 ^ x75 ;
  assign n2137 = ~n1820 & n2136 ;
  assign n2138 = n2137 ^ x75 ;
  assign n2139 = n2138 ^ x43 ;
  assign n2140 = ~n1856 & n2139 ;
  assign n2141 = n2140 ^ x43 ;
  assign n2142 = n2141 ^ x11 ;
  assign n2143 = n1892 & n2142 ;
  assign n2144 = n2143 ^ x11 ;
  assign n2145 = x236 ^ x204 ;
  assign n2146 = ~n1681 & n2145 ;
  assign n2147 = n2146 ^ x204 ;
  assign n2148 = n2147 ^ x172 ;
  assign n2149 = n1713 & n2148 ;
  assign n2150 = n2149 ^ x172 ;
  assign n2151 = n2150 ^ x140 ;
  assign n2152 = ~n1749 & n2151 ;
  assign n2153 = n2152 ^ x140 ;
  assign n2154 = n2153 ^ x108 ;
  assign n2155 = ~n1785 & n2154 ;
  assign n2156 = n2155 ^ x108 ;
  assign n2157 = n2156 ^ x76 ;
  assign n2158 = ~n1820 & n2157 ;
  assign n2159 = n2158 ^ x76 ;
  assign n2160 = n2159 ^ x44 ;
  assign n2161 = ~n1856 & n2160 ;
  assign n2162 = n2161 ^ x44 ;
  assign n2163 = n2162 ^ x12 ;
  assign n2164 = n1892 & n2163 ;
  assign n2165 = n2164 ^ x12 ;
  assign n2166 = x237 ^ x205 ;
  assign n2167 = ~n1681 & n2166 ;
  assign n2168 = n2167 ^ x205 ;
  assign n2169 = n2168 ^ x173 ;
  assign n2170 = n1713 & n2169 ;
  assign n2171 = n2170 ^ x173 ;
  assign n2172 = n2171 ^ x141 ;
  assign n2173 = ~n1749 & n2172 ;
  assign n2174 = n2173 ^ x141 ;
  assign n2175 = n2174 ^ x109 ;
  assign n2176 = ~n1785 & n2175 ;
  assign n2177 = n2176 ^ x109 ;
  assign n2178 = n2177 ^ x77 ;
  assign n2179 = ~n1820 & n2178 ;
  assign n2180 = n2179 ^ x77 ;
  assign n2181 = n2180 ^ x45 ;
  assign n2182 = ~n1856 & n2181 ;
  assign n2183 = n2182 ^ x45 ;
  assign n2184 = n2183 ^ x13 ;
  assign n2185 = n1892 & n2184 ;
  assign n2186 = n2185 ^ x13 ;
  assign n2187 = x238 ^ x206 ;
  assign n2188 = ~n1681 & n2187 ;
  assign n2189 = n2188 ^ x206 ;
  assign n2190 = n2189 ^ x174 ;
  assign n2191 = n1713 & n2190 ;
  assign n2192 = n2191 ^ x174 ;
  assign n2193 = n2192 ^ x142 ;
  assign n2194 = ~n1749 & n2193 ;
  assign n2195 = n2194 ^ x142 ;
  assign n2196 = n2195 ^ x110 ;
  assign n2197 = ~n1785 & n2196 ;
  assign n2198 = n2197 ^ x110 ;
  assign n2199 = n2198 ^ x78 ;
  assign n2200 = ~n1820 & n2199 ;
  assign n2201 = n2200 ^ x78 ;
  assign n2202 = n2201 ^ x46 ;
  assign n2203 = ~n1856 & n2202 ;
  assign n2204 = n2203 ^ x46 ;
  assign n2205 = n2204 ^ x14 ;
  assign n2206 = n1892 & n2205 ;
  assign n2207 = n2206 ^ x14 ;
  assign n2208 = x239 ^ x207 ;
  assign n2209 = ~n1681 & n2208 ;
  assign n2210 = n2209 ^ x207 ;
  assign n2211 = n2210 ^ x175 ;
  assign n2212 = n1713 & n2211 ;
  assign n2213 = n2212 ^ x175 ;
  assign n2214 = n2213 ^ x143 ;
  assign n2215 = ~n1749 & n2214 ;
  assign n2216 = n2215 ^ x143 ;
  assign n2217 = n2216 ^ x111 ;
  assign n2218 = ~n1785 & n2217 ;
  assign n2219 = n2218 ^ x111 ;
  assign n2220 = n2219 ^ x79 ;
  assign n2221 = ~n1820 & n2220 ;
  assign n2222 = n2221 ^ x79 ;
  assign n2223 = n2222 ^ x47 ;
  assign n2224 = ~n1856 & n2223 ;
  assign n2225 = n2224 ^ x47 ;
  assign n2226 = n2225 ^ x15 ;
  assign n2227 = n1892 & n2226 ;
  assign n2228 = n2227 ^ x15 ;
  assign n2229 = x240 ^ x208 ;
  assign n2230 = ~n1681 & n2229 ;
  assign n2231 = n2230 ^ x208 ;
  assign n2232 = n2231 ^ x176 ;
  assign n2233 = n1713 & n2232 ;
  assign n2234 = n2233 ^ x176 ;
  assign n2235 = n2234 ^ x144 ;
  assign n2236 = ~n1749 & n2235 ;
  assign n2237 = n2236 ^ x144 ;
  assign n2238 = n2237 ^ x112 ;
  assign n2239 = ~n1785 & n2238 ;
  assign n2240 = n2239 ^ x112 ;
  assign n2241 = n2240 ^ x80 ;
  assign n2242 = ~n1820 & n2241 ;
  assign n2243 = n2242 ^ x80 ;
  assign n2244 = n2243 ^ x48 ;
  assign n2245 = ~n1856 & n2244 ;
  assign n2246 = n2245 ^ x48 ;
  assign n2247 = n2246 ^ x16 ;
  assign n2248 = n1892 & n2247 ;
  assign n2249 = n2248 ^ x16 ;
  assign n2250 = x241 ^ x209 ;
  assign n2251 = ~n1681 & n2250 ;
  assign n2252 = n2251 ^ x209 ;
  assign n2253 = n2252 ^ x177 ;
  assign n2254 = n1713 & n2253 ;
  assign n2255 = n2254 ^ x177 ;
  assign n2256 = n2255 ^ x145 ;
  assign n2257 = ~n1749 & n2256 ;
  assign n2258 = n2257 ^ x145 ;
  assign n2259 = n2258 ^ x113 ;
  assign n2260 = ~n1785 & n2259 ;
  assign n2261 = n2260 ^ x113 ;
  assign n2262 = n2261 ^ x81 ;
  assign n2263 = ~n1820 & n2262 ;
  assign n2264 = n2263 ^ x81 ;
  assign n2265 = n2264 ^ x49 ;
  assign n2266 = ~n1856 & n2265 ;
  assign n2267 = n2266 ^ x49 ;
  assign n2268 = n2267 ^ x17 ;
  assign n2269 = n1892 & n2268 ;
  assign n2270 = n2269 ^ x17 ;
  assign n2271 = x242 ^ x210 ;
  assign n2272 = ~n1681 & n2271 ;
  assign n2273 = n2272 ^ x210 ;
  assign n2274 = n2273 ^ x178 ;
  assign n2275 = n1713 & n2274 ;
  assign n2276 = n2275 ^ x178 ;
  assign n2277 = n2276 ^ x146 ;
  assign n2278 = ~n1749 & n2277 ;
  assign n2279 = n2278 ^ x146 ;
  assign n2280 = n2279 ^ x114 ;
  assign n2281 = ~n1785 & n2280 ;
  assign n2282 = n2281 ^ x114 ;
  assign n2283 = n2282 ^ x82 ;
  assign n2284 = ~n1820 & n2283 ;
  assign n2285 = n2284 ^ x82 ;
  assign n2286 = n2285 ^ x50 ;
  assign n2287 = ~n1856 & n2286 ;
  assign n2288 = n2287 ^ x50 ;
  assign n2289 = n2288 ^ x18 ;
  assign n2290 = n1892 & n2289 ;
  assign n2291 = n2290 ^ x18 ;
  assign n2292 = x243 ^ x211 ;
  assign n2293 = ~n1681 & n2292 ;
  assign n2294 = n2293 ^ x211 ;
  assign n2295 = n2294 ^ x179 ;
  assign n2296 = n1713 & n2295 ;
  assign n2297 = n2296 ^ x179 ;
  assign n2298 = n2297 ^ x147 ;
  assign n2299 = ~n1749 & n2298 ;
  assign n2300 = n2299 ^ x147 ;
  assign n2301 = n2300 ^ x115 ;
  assign n2302 = ~n1785 & n2301 ;
  assign n2303 = n2302 ^ x115 ;
  assign n2304 = n2303 ^ x83 ;
  assign n2305 = ~n1820 & n2304 ;
  assign n2306 = n2305 ^ x83 ;
  assign n2307 = n2306 ^ x51 ;
  assign n2308 = ~n1856 & n2307 ;
  assign n2309 = n2308 ^ x51 ;
  assign n2310 = n2309 ^ x19 ;
  assign n2311 = n1892 & n2310 ;
  assign n2312 = n2311 ^ x19 ;
  assign n2313 = x244 ^ x212 ;
  assign n2314 = ~n1681 & n2313 ;
  assign n2315 = n2314 ^ x212 ;
  assign n2316 = n2315 ^ x180 ;
  assign n2317 = n1713 & n2316 ;
  assign n2318 = n2317 ^ x180 ;
  assign n2319 = n2318 ^ x148 ;
  assign n2320 = ~n1749 & n2319 ;
  assign n2321 = n2320 ^ x148 ;
  assign n2322 = n2321 ^ x116 ;
  assign n2323 = ~n1785 & n2322 ;
  assign n2324 = n2323 ^ x116 ;
  assign n2325 = n2324 ^ x84 ;
  assign n2326 = ~n1820 & n2325 ;
  assign n2327 = n2326 ^ x84 ;
  assign n2328 = n2327 ^ x52 ;
  assign n2329 = ~n1856 & n2328 ;
  assign n2330 = n2329 ^ x52 ;
  assign n2331 = n2330 ^ x20 ;
  assign n2332 = n1892 & n2331 ;
  assign n2333 = n2332 ^ x20 ;
  assign n2334 = x245 ^ x213 ;
  assign n2335 = ~n1681 & n2334 ;
  assign n2336 = n2335 ^ x213 ;
  assign n2337 = n2336 ^ x181 ;
  assign n2338 = n1713 & n2337 ;
  assign n2339 = n2338 ^ x181 ;
  assign n2340 = n2339 ^ x149 ;
  assign n2341 = ~n1749 & n2340 ;
  assign n2342 = n2341 ^ x149 ;
  assign n2343 = n2342 ^ x117 ;
  assign n2344 = ~n1785 & n2343 ;
  assign n2345 = n2344 ^ x117 ;
  assign n2346 = n2345 ^ x85 ;
  assign n2347 = ~n1820 & n2346 ;
  assign n2348 = n2347 ^ x85 ;
  assign n2349 = n2348 ^ x53 ;
  assign n2350 = ~n1856 & n2349 ;
  assign n2351 = n2350 ^ x53 ;
  assign n2352 = n2351 ^ x21 ;
  assign n2353 = n1892 & n2352 ;
  assign n2354 = n2353 ^ x21 ;
  assign n2355 = x246 ^ x214 ;
  assign n2356 = ~n1681 & n2355 ;
  assign n2357 = n2356 ^ x214 ;
  assign n2358 = n2357 ^ x182 ;
  assign n2359 = n1713 & n2358 ;
  assign n2360 = n2359 ^ x182 ;
  assign n2361 = n2360 ^ x150 ;
  assign n2362 = ~n1749 & n2361 ;
  assign n2363 = n2362 ^ x150 ;
  assign n2364 = n2363 ^ x118 ;
  assign n2365 = ~n1785 & n2364 ;
  assign n2366 = n2365 ^ x118 ;
  assign n2367 = n2366 ^ x86 ;
  assign n2368 = ~n1820 & n2367 ;
  assign n2369 = n2368 ^ x86 ;
  assign n2370 = n2369 ^ x54 ;
  assign n2371 = ~n1856 & n2370 ;
  assign n2372 = n2371 ^ x54 ;
  assign n2373 = n2372 ^ x22 ;
  assign n2374 = n1892 & n2373 ;
  assign n2375 = n2374 ^ x22 ;
  assign n2376 = x247 ^ x215 ;
  assign n2377 = ~n1681 & n2376 ;
  assign n2378 = n2377 ^ x215 ;
  assign n2379 = n2378 ^ x183 ;
  assign n2380 = n1713 & n2379 ;
  assign n2381 = n2380 ^ x183 ;
  assign n2382 = n2381 ^ x151 ;
  assign n2383 = ~n1749 & n2382 ;
  assign n2384 = n2383 ^ x151 ;
  assign n2385 = n2384 ^ x119 ;
  assign n2386 = ~n1785 & n2385 ;
  assign n2387 = n2386 ^ x119 ;
  assign n2388 = n2387 ^ x87 ;
  assign n2389 = ~n1820 & n2388 ;
  assign n2390 = n2389 ^ x87 ;
  assign n2391 = n2390 ^ x55 ;
  assign n2392 = ~n1856 & n2391 ;
  assign n2393 = n2392 ^ x55 ;
  assign n2394 = n2393 ^ x23 ;
  assign n2395 = n1892 & n2394 ;
  assign n2396 = n2395 ^ x23 ;
  assign n2397 = x248 ^ x216 ;
  assign n2398 = ~n1681 & n2397 ;
  assign n2399 = n2398 ^ x216 ;
  assign n2400 = n2399 ^ x184 ;
  assign n2401 = n1713 & n2400 ;
  assign n2402 = n2401 ^ x184 ;
  assign n2403 = n2402 ^ x152 ;
  assign n2404 = ~n1749 & n2403 ;
  assign n2405 = n2404 ^ x152 ;
  assign n2406 = n2405 ^ x120 ;
  assign n2407 = ~n1785 & n2406 ;
  assign n2408 = n2407 ^ x120 ;
  assign n2409 = n2408 ^ x88 ;
  assign n2410 = ~n1820 & n2409 ;
  assign n2411 = n2410 ^ x88 ;
  assign n2412 = n2411 ^ x56 ;
  assign n2413 = ~n1856 & n2412 ;
  assign n2414 = n2413 ^ x56 ;
  assign n2415 = n2414 ^ x24 ;
  assign n2416 = n1892 & n2415 ;
  assign n2417 = n2416 ^ x24 ;
  assign n2418 = x249 ^ x217 ;
  assign n2419 = ~n1681 & n2418 ;
  assign n2420 = n2419 ^ x217 ;
  assign n2421 = n2420 ^ x185 ;
  assign n2422 = n1713 & n2421 ;
  assign n2423 = n2422 ^ x185 ;
  assign n2424 = n2423 ^ x153 ;
  assign n2425 = ~n1749 & n2424 ;
  assign n2426 = n2425 ^ x153 ;
  assign n2427 = n2426 ^ x121 ;
  assign n2428 = ~n1785 & n2427 ;
  assign n2429 = n2428 ^ x121 ;
  assign n2430 = n2429 ^ x89 ;
  assign n2431 = ~n1820 & n2430 ;
  assign n2432 = n2431 ^ x89 ;
  assign n2433 = n2432 ^ x57 ;
  assign n2434 = ~n1856 & n2433 ;
  assign n2435 = n2434 ^ x57 ;
  assign n2436 = n2435 ^ x25 ;
  assign n2437 = n1892 & n2436 ;
  assign n2438 = n2437 ^ x25 ;
  assign n2439 = x250 ^ x218 ;
  assign n2440 = ~n1681 & n2439 ;
  assign n2441 = n2440 ^ x218 ;
  assign n2442 = n2441 ^ x186 ;
  assign n2443 = n1713 & n2442 ;
  assign n2444 = n2443 ^ x186 ;
  assign n2445 = n2444 ^ x154 ;
  assign n2446 = ~n1749 & n2445 ;
  assign n2447 = n2446 ^ x154 ;
  assign n2448 = n2447 ^ x122 ;
  assign n2449 = ~n1785 & n2448 ;
  assign n2450 = n2449 ^ x122 ;
  assign n2451 = n2450 ^ x90 ;
  assign n2452 = ~n1820 & n2451 ;
  assign n2453 = n2452 ^ x90 ;
  assign n2454 = n2453 ^ x58 ;
  assign n2455 = ~n1856 & n2454 ;
  assign n2456 = n2455 ^ x58 ;
  assign n2457 = n2456 ^ x26 ;
  assign n2458 = n1892 & n2457 ;
  assign n2459 = n2458 ^ x26 ;
  assign n2460 = x251 ^ x219 ;
  assign n2461 = ~n1681 & n2460 ;
  assign n2462 = n2461 ^ x219 ;
  assign n2463 = n2462 ^ x187 ;
  assign n2464 = n1713 & n2463 ;
  assign n2465 = n2464 ^ x187 ;
  assign n2466 = n2465 ^ x155 ;
  assign n2467 = ~n1749 & n2466 ;
  assign n2468 = n2467 ^ x155 ;
  assign n2469 = n2468 ^ x123 ;
  assign n2470 = ~n1785 & n2469 ;
  assign n2471 = n2470 ^ x123 ;
  assign n2472 = n2471 ^ x91 ;
  assign n2473 = ~n1820 & n2472 ;
  assign n2474 = n2473 ^ x91 ;
  assign n2475 = n2474 ^ x59 ;
  assign n2476 = ~n1856 & n2475 ;
  assign n2477 = n2476 ^ x59 ;
  assign n2478 = n2477 ^ x27 ;
  assign n2479 = n1892 & n2478 ;
  assign n2480 = n2479 ^ x27 ;
  assign n2481 = x252 ^ x220 ;
  assign n2482 = ~n1681 & n2481 ;
  assign n2483 = n2482 ^ x220 ;
  assign n2484 = n2483 ^ x188 ;
  assign n2485 = n1713 & n2484 ;
  assign n2486 = n2485 ^ x188 ;
  assign n2487 = n2486 ^ x156 ;
  assign n2488 = ~n1749 & n2487 ;
  assign n2489 = n2488 ^ x156 ;
  assign n2490 = n2489 ^ x124 ;
  assign n2491 = ~n1785 & n2490 ;
  assign n2492 = n2491 ^ x124 ;
  assign n2493 = n2492 ^ x92 ;
  assign n2494 = ~n1820 & n2493 ;
  assign n2495 = n2494 ^ x92 ;
  assign n2496 = n2495 ^ x60 ;
  assign n2497 = ~n1856 & n2496 ;
  assign n2498 = n2497 ^ x60 ;
  assign n2499 = n2498 ^ x28 ;
  assign n2500 = n1892 & n2499 ;
  assign n2501 = n2500 ^ x28 ;
  assign n2502 = x253 ^ x221 ;
  assign n2503 = ~n1681 & n2502 ;
  assign n2504 = n2503 ^ x221 ;
  assign n2505 = n2504 ^ x189 ;
  assign n2506 = n1713 & n2505 ;
  assign n2507 = n2506 ^ x189 ;
  assign n2508 = n2507 ^ x157 ;
  assign n2509 = ~n1749 & n2508 ;
  assign n2510 = n2509 ^ x157 ;
  assign n2511 = n2510 ^ x125 ;
  assign n2512 = ~n1785 & n2511 ;
  assign n2513 = n2512 ^ x125 ;
  assign n2514 = n2513 ^ x93 ;
  assign n2515 = ~n1820 & n2514 ;
  assign n2516 = n2515 ^ x93 ;
  assign n2517 = n2516 ^ x61 ;
  assign n2518 = ~n1856 & n2517 ;
  assign n2519 = n2518 ^ x61 ;
  assign n2520 = n2519 ^ x29 ;
  assign n2521 = n1892 & n2520 ;
  assign n2522 = n2521 ^ x29 ;
  assign n2523 = x254 ^ x222 ;
  assign n2524 = ~n1681 & n2523 ;
  assign n2525 = n2524 ^ x222 ;
  assign n2526 = n2525 ^ x190 ;
  assign n2527 = n1713 & n2526 ;
  assign n2528 = n2527 ^ x190 ;
  assign n2529 = n2528 ^ x158 ;
  assign n2530 = ~n1749 & n2529 ;
  assign n2531 = n2530 ^ x158 ;
  assign n2532 = n2531 ^ x126 ;
  assign n2533 = ~n1785 & n2532 ;
  assign n2534 = n2533 ^ x126 ;
  assign n2535 = n2534 ^ x94 ;
  assign n2536 = ~n1820 & n2535 ;
  assign n2537 = n2536 ^ x94 ;
  assign n2538 = n2537 ^ x62 ;
  assign n2539 = ~n1856 & n2538 ;
  assign n2540 = n2539 ^ x62 ;
  assign n2541 = n2540 ^ x30 ;
  assign n2542 = n1892 & n2541 ;
  assign n2543 = n2542 ^ x30 ;
  assign n2544 = x255 ^ x223 ;
  assign n2545 = ~n1681 & n2544 ;
  assign n2546 = n2545 ^ x223 ;
  assign n2547 = n2546 ^ x191 ;
  assign n2548 = n1713 & n2547 ;
  assign n2549 = n2548 ^ x191 ;
  assign n2550 = n2549 ^ x159 ;
  assign n2551 = ~n1749 & n2550 ;
  assign n2552 = n2551 ^ x159 ;
  assign n2553 = n2552 ^ x127 ;
  assign n2554 = ~n1785 & n2553 ;
  assign n2555 = n2554 ^ x127 ;
  assign n2556 = n2555 ^ x95 ;
  assign n2557 = ~n1820 & n2556 ;
  assign n2558 = n2557 ^ x95 ;
  assign n2559 = n2558 ^ x63 ;
  assign n2560 = ~n1856 & n2559 ;
  assign n2561 = n2560 ^ x63 ;
  assign n2562 = n2561 ^ x31 ;
  assign n2563 = n1892 & n2562 ;
  assign n2564 = n2563 ^ x31 ;
  assign y0 = n1913 ;
  assign y1 = n1934 ;
  assign y2 = n1955 ;
  assign y3 = n1976 ;
  assign y4 = n1997 ;
  assign y5 = n2018 ;
  assign y6 = n2039 ;
  assign y7 = n2060 ;
  assign y8 = n2081 ;
  assign y9 = n2102 ;
  assign y10 = n2123 ;
  assign y11 = n2144 ;
  assign y12 = n2165 ;
  assign y13 = n2186 ;
  assign y14 = n2207 ;
  assign y15 = n2228 ;
  assign y16 = n2249 ;
  assign y17 = n2270 ;
  assign y18 = n2291 ;
  assign y19 = n2312 ;
  assign y20 = n2333 ;
  assign y21 = n2354 ;
  assign y22 = n2375 ;
  assign y23 = n2396 ;
  assign y24 = n2417 ;
  assign y25 = n2438 ;
  assign y26 = n2459 ;
  assign y27 = n2480 ;
  assign y28 = n2501 ;
  assign y29 = n2522 ;
  assign y30 = n2543 ;
  assign y31 = n2564 ;
endmodule
