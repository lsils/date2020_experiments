module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , y0 , y1 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 ;
  output y0 , y1 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 ;
  assign n40 = x30 & x31 ;
  assign n41 = n40 ^ x31 ;
  assign n36 = x28 & x29 ;
  assign n37 = n36 ^ x29 ;
  assign n221 = n41 ^ n37 ;
  assign n33 = x26 & x27 ;
  assign n34 = n33 ^ x27 ;
  assign n228 = n221 ^ n34 ;
  assign n47 = x18 & x19 ;
  assign n48 = n47 ^ x19 ;
  assign n241 = n228 ^ n48 ;
  assign n58 = x24 & x25 ;
  assign n59 = n58 ^ x25 ;
  assign n51 = x22 & x23 ;
  assign n52 = n51 ^ x23 ;
  assign n225 = n59 ^ n52 ;
  assign n54 = x20 & x21 ;
  assign n55 = n54 ^ x21 ;
  assign n226 = n225 ^ n55 ;
  assign n242 = n241 ^ n226 ;
  assign n74 = x2 & x3 ;
  assign n75 = n74 ^ x3 ;
  assign n243 = n242 ^ n75 ;
  assign n81 = x8 & x9 ;
  assign n82 = n81 ^ x9 ;
  assign n78 = x10 & x11 ;
  assign n79 = n78 ^ x11 ;
  assign n247 = n82 ^ n79 ;
  assign n84 = x6 & x7 ;
  assign n85 = n84 ^ x7 ;
  assign n248 = n247 ^ n85 ;
  assign n95 = x14 & x15 ;
  assign n96 = n95 ^ x15 ;
  assign n92 = x16 & x17 ;
  assign n93 = n92 ^ x17 ;
  assign n244 = n96 ^ n93 ;
  assign n98 = x12 & x13 ;
  assign n99 = n98 ^ x13 ;
  assign n245 = n244 ^ n99 ;
  assign n89 = x4 & x5 ;
  assign n90 = n89 ^ x5 ;
  assign n246 = n245 ^ n90 ;
  assign n249 = n248 ^ n246 ;
  assign n250 = n249 ^ n242 ;
  assign n251 = n243 & ~n250 ;
  assign n252 = n251 ^ n75 ;
  assign n233 = n55 ^ n52 ;
  assign n234 = n59 ^ n55 ;
  assign n235 = n233 & ~n234 ;
  assign n236 = n235 ^ n52 ;
  assign n227 = n226 ^ n48 ;
  assign n229 = n228 ^ n226 ;
  assign n230 = n227 & ~n229 ;
  assign n231 = n230 ^ n48 ;
  assign n222 = n37 ^ n34 ;
  assign n223 = ~n221 & n222 ;
  assign n224 = n223 ^ n34 ;
  assign n232 = n231 ^ n224 ;
  assign n240 = n236 ^ n232 ;
  assign n253 = n252 ^ n240 ;
  assign n261 = n85 ^ n82 ;
  assign n262 = n247 & ~n261 ;
  assign n263 = n262 ^ n79 ;
  assign n257 = n248 ^ n245 ;
  assign n258 = n246 & ~n257 ;
  assign n259 = n258 ^ n90 ;
  assign n254 = n99 ^ n96 ;
  assign n255 = n244 & ~n254 ;
  assign n256 = n255 ^ n93 ;
  assign n260 = n259 ^ n256 ;
  assign n264 = n263 ^ n260 ;
  assign n265 = n264 ^ n240 ;
  assign n266 = ~n253 & n265 ;
  assign n267 = n266 ^ n264 ;
  assign n237 = n236 ^ n231 ;
  assign n238 = n232 & n237 ;
  assign n239 = n238 ^ n231 ;
  assign n268 = n267 ^ n239 ;
  assign n269 = n263 ^ n256 ;
  assign n270 = ~n260 & n269 ;
  assign n271 = n270 ^ n263 ;
  assign n272 = n271 ^ n267 ;
  assign n273 = n268 & ~n272 ;
  assign n274 = n273 ^ n239 ;
  assign n275 = n264 ^ n253 ;
  assign n131 = x0 & x1 ;
  assign n132 = n131 ^ x1 ;
  assign n276 = n249 ^ n243 ;
  assign n277 = n132 & n276 ;
  assign n278 = n275 & n277 ;
  assign n279 = n271 ^ n268 ;
  assign n280 = n278 & n279 ;
  assign n282 = ~n274 & ~n280 ;
  assign n281 = n280 ^ n274 ;
  assign n283 = n282 ^ n281 ;
  assign n287 = n58 ^ n51 ;
  assign n288 = n287 ^ n54 ;
  assign n284 = n40 ^ n36 ;
  assign n285 = n284 ^ n33 ;
  assign n286 = n285 ^ n47 ;
  assign n303 = n288 ^ n286 ;
  assign n304 = n303 ^ n74 ;
  assign n308 = n81 ^ n78 ;
  assign n309 = n308 ^ n84 ;
  assign n305 = n95 ^ n92 ;
  assign n306 = n305 ^ n98 ;
  assign n307 = n306 ^ n89 ;
  assign n310 = n309 ^ n307 ;
  assign n311 = n310 ^ n303 ;
  assign n312 = n304 & ~n311 ;
  assign n313 = n312 ^ n74 ;
  assign n296 = n54 ^ n51 ;
  assign n297 = ~n287 & n296 ;
  assign n298 = n297 ^ n54 ;
  assign n292 = n36 ^ n33 ;
  assign n293 = ~n284 & n292 ;
  assign n294 = n293 ^ n33 ;
  assign n289 = n288 ^ n285 ;
  assign n290 = n286 & ~n289 ;
  assign n291 = n290 ^ n47 ;
  assign n295 = n294 ^ n291 ;
  assign n302 = n298 ^ n295 ;
  assign n314 = n313 ^ n302 ;
  assign n322 = n84 ^ n81 ;
  assign n323 = ~n308 & n322 ;
  assign n324 = n323 ^ n84 ;
  assign n318 = n309 ^ n306 ;
  assign n319 = n307 & ~n318 ;
  assign n320 = n319 ^ n89 ;
  assign n315 = n98 ^ n95 ;
  assign n316 = ~n305 & n315 ;
  assign n317 = n316 ^ n98 ;
  assign n321 = n320 ^ n317 ;
  assign n325 = n324 ^ n321 ;
  assign n326 = n325 ^ n302 ;
  assign n327 = ~n314 & n326 ;
  assign n328 = n327 ^ n325 ;
  assign n299 = n298 ^ n294 ;
  assign n300 = n295 & ~n299 ;
  assign n301 = n300 ^ n291 ;
  assign n329 = n328 ^ n301 ;
  assign n330 = n324 ^ n317 ;
  assign n331 = ~n321 & n330 ;
  assign n332 = n331 ^ n324 ;
  assign n333 = n332 ^ n328 ;
  assign n334 = n329 & ~n333 ;
  assign n335 = n334 ^ n301 ;
  assign n336 = n310 ^ n304 ;
  assign n337 = n131 & n336 ;
  assign n338 = n325 ^ n314 ;
  assign n339 = n337 & n338 ;
  assign n340 = n332 ^ n329 ;
  assign n341 = n339 & n340 ;
  assign n343 = ~n335 & ~n341 ;
  assign n342 = n341 ^ n335 ;
  assign n344 = n343 ^ n342 ;
  assign n346 = ~n283 & n344 ;
  assign n345 = n344 ^ n283 ;
  assign n347 = n346 ^ n345 ;
  assign n348 = n347 ^ n283 ;
  assign n76 = n75 ^ x2 ;
  assign n60 = n59 ^ x24 ;
  assign n56 = n55 ^ x20 ;
  assign n53 = n52 ^ x22 ;
  assign n57 = n56 ^ n53 ;
  assign n61 = n60 ^ n57 ;
  assign n49 = n48 ^ x18 ;
  assign n42 = n41 ^ x30 ;
  assign n38 = n37 ^ x28 ;
  assign n35 = n34 ^ x26 ;
  assign n39 = n38 ^ n35 ;
  assign n46 = n42 ^ n39 ;
  assign n50 = n49 ^ n46 ;
  assign n73 = n61 ^ n50 ;
  assign n77 = n76 ^ n73 ;
  assign n100 = n99 ^ x12 ;
  assign n97 = n96 ^ x14 ;
  assign n101 = n100 ^ n97 ;
  assign n94 = n93 ^ x16 ;
  assign n102 = n101 ^ n94 ;
  assign n91 = n90 ^ x4 ;
  assign n103 = n102 ^ n91 ;
  assign n86 = n85 ^ x6 ;
  assign n83 = n82 ^ x8 ;
  assign n87 = n86 ^ n83 ;
  assign n80 = n79 ^ x10 ;
  assign n88 = n87 ^ n80 ;
  assign n104 = n103 ^ n88 ;
  assign n105 = n104 ^ n76 ;
  assign n106 = n77 & ~n105 ;
  assign n107 = n106 ^ n73 ;
  assign n66 = n60 ^ n56 ;
  assign n67 = n57 & ~n66 ;
  assign n68 = n67 ^ n53 ;
  assign n62 = n61 ^ n46 ;
  assign n63 = ~n50 & n62 ;
  assign n64 = n63 ^ n61 ;
  assign n43 = n42 ^ n38 ;
  assign n44 = n39 & ~n43 ;
  assign n45 = n44 ^ n35 ;
  assign n65 = n64 ^ n45 ;
  assign n72 = n68 ^ n65 ;
  assign n108 = n107 ^ n72 ;
  assign n116 = n83 ^ n80 ;
  assign n117 = ~n87 & n116 ;
  assign n118 = n117 ^ n80 ;
  assign n112 = n97 ^ n94 ;
  assign n113 = ~n101 & n112 ;
  assign n114 = n113 ^ n94 ;
  assign n109 = n91 ^ n88 ;
  assign n110 = ~n103 & n109 ;
  assign n111 = n110 ^ n88 ;
  assign n115 = n114 ^ n111 ;
  assign n119 = n118 ^ n115 ;
  assign n120 = n119 ^ n72 ;
  assign n121 = n108 & ~n120 ;
  assign n122 = n121 ^ n107 ;
  assign n69 = n68 ^ n45 ;
  assign n70 = ~n65 & n69 ;
  assign n71 = n70 ^ n68 ;
  assign n123 = n122 ^ n71 ;
  assign n124 = n118 ^ n114 ;
  assign n125 = n115 & ~n124 ;
  assign n126 = n125 ^ n111 ;
  assign n127 = n126 ^ n71 ;
  assign n128 = ~n123 & n127 ;
  assign n129 = n128 ^ n126 ;
  assign n130 = n104 ^ n77 ;
  assign n133 = n132 ^ x0 ;
  assign n134 = ~n130 & ~n133 ;
  assign n135 = n119 ^ n108 ;
  assign n136 = n134 & ~n135 ;
  assign n137 = n126 ^ n123 ;
  assign n138 = n136 & ~n137 ;
  assign n140 = n129 & ~n138 ;
  assign n139 = n138 ^ n129 ;
  assign n141 = n140 ^ n139 ;
  assign n169 = n74 ^ x2 ;
  assign n151 = n58 ^ x24 ;
  assign n150 = n51 ^ x22 ;
  assign n152 = n151 ^ n150 ;
  assign n149 = n54 ^ x20 ;
  assign n153 = n152 ^ n149 ;
  assign n145 = n40 ^ x30 ;
  assign n144 = n36 ^ x28 ;
  assign n146 = n145 ^ n144 ;
  assign n143 = n33 ^ x26 ;
  assign n147 = n146 ^ n143 ;
  assign n142 = n47 ^ x18 ;
  assign n148 = n147 ^ n142 ;
  assign n168 = n153 ^ n148 ;
  assign n170 = n169 ^ n168 ;
  assign n180 = n78 ^ x10 ;
  assign n179 = n81 ^ x8 ;
  assign n181 = n180 ^ n179 ;
  assign n178 = n84 ^ x6 ;
  assign n182 = n181 ^ n178 ;
  assign n174 = n92 ^ x16 ;
  assign n173 = n95 ^ x14 ;
  assign n175 = n174 ^ n173 ;
  assign n172 = n98 ^ x12 ;
  assign n176 = n175 ^ n172 ;
  assign n171 = n89 ^ x4 ;
  assign n177 = n176 ^ n171 ;
  assign n183 = n182 ^ n177 ;
  assign n184 = n183 ^ n169 ;
  assign n185 = n170 & ~n184 ;
  assign n186 = n185 ^ n168 ;
  assign n161 = n150 ^ n149 ;
  assign n162 = ~n152 & n161 ;
  assign n163 = n162 ^ n149 ;
  assign n157 = n144 ^ n143 ;
  assign n158 = ~n146 & n157 ;
  assign n159 = n158 ^ n143 ;
  assign n154 = n153 ^ n147 ;
  assign n155 = n148 & ~n154 ;
  assign n156 = n155 ^ n142 ;
  assign n160 = n159 ^ n156 ;
  assign n167 = n163 ^ n160 ;
  assign n187 = n186 ^ n167 ;
  assign n195 = n179 ^ n178 ;
  assign n196 = ~n181 & n195 ;
  assign n197 = n196 ^ n178 ;
  assign n191 = n182 ^ n176 ;
  assign n192 = n177 & ~n191 ;
  assign n193 = n192 ^ n171 ;
  assign n188 = n173 ^ n172 ;
  assign n189 = ~n175 & n188 ;
  assign n190 = n189 ^ n172 ;
  assign n194 = n193 ^ n190 ;
  assign n198 = n197 ^ n194 ;
  assign n199 = n198 ^ n167 ;
  assign n200 = ~n187 & n199 ;
  assign n201 = n200 ^ n198 ;
  assign n164 = n163 ^ n159 ;
  assign n165 = n160 & ~n164 ;
  assign n166 = n165 ^ n156 ;
  assign n202 = n201 ^ n166 ;
  assign n203 = n197 ^ n190 ;
  assign n204 = ~n194 & n203 ;
  assign n205 = n204 ^ n197 ;
  assign n206 = n205 ^ n201 ;
  assign n207 = n202 & ~n206 ;
  assign n208 = n207 ^ n166 ;
  assign n209 = n183 ^ n170 ;
  assign n210 = n131 ^ x0 ;
  assign n211 = n209 & n210 ;
  assign n212 = n198 ^ n187 ;
  assign n213 = n211 & n212 ;
  assign n214 = n205 ^ n202 ;
  assign n215 = n213 & n214 ;
  assign n217 = ~n208 & ~n215 ;
  assign n216 = n215 ^ n208 ;
  assign n218 = n217 ^ n216 ;
  assign n219 = n141 & n218 ;
  assign n220 = n219 ^ n218 ;
  assign n349 = n348 ^ n220 ;
  assign n350 = n140 & n217 ;
  assign n351 = n350 ^ n220 ;
  assign n352 = n282 & n343 ;
  assign n353 = n352 ^ n348 ;
  assign n355 = ~n351 & n353 ;
  assign n354 = n353 ^ n351 ;
  assign n356 = n355 ^ n354 ;
  assign n357 = n356 ^ n348 ;
  assign n358 = n357 ^ n348 ;
  assign n386 = n340 ^ n339 ;
  assign n385 = n279 ^ n278 ;
  assign n387 = n386 ^ n385 ;
  assign n388 = n342 ^ n281 ;
  assign n390 = n276 ^ n132 ;
  assign n391 = n336 ^ n131 ;
  assign n392 = n390 & ~n391 ;
  assign n389 = n338 ^ n337 ;
  assign n393 = n392 ^ n389 ;
  assign n394 = n392 ^ n277 ;
  assign n395 = n394 ^ n275 ;
  assign n396 = ~n393 & ~n395 ;
  assign n397 = n396 ^ n389 ;
  assign n398 = n397 ^ n385 ;
  assign n399 = n397 ^ n386 ;
  assign n400 = ~n398 & ~n399 ;
  assign n401 = n400 ^ n385 ;
  assign n402 = n401 ^ n342 ;
  assign n403 = ~n388 & ~n402 ;
  assign n404 = n403 ^ n342 ;
  assign n405 = n404 ^ n283 ;
  assign n406 = ~n345 & ~n405 ;
  assign n407 = n406 ^ n344 ;
  assign n408 = n387 & ~n407 ;
  assign n409 = n408 ^ n385 ;
  assign n359 = n218 ^ n141 ;
  assign n360 = n216 ^ n139 ;
  assign n370 = n137 ^ n136 ;
  assign n362 = n135 ^ n134 ;
  assign n361 = n212 ^ n211 ;
  assign n363 = n362 ^ n361 ;
  assign n364 = n133 ^ n130 ;
  assign n365 = n210 ^ n209 ;
  assign n366 = n364 & ~n365 ;
  assign n367 = n366 ^ n362 ;
  assign n368 = ~n363 & ~n367 ;
  assign n369 = n368 ^ n366 ;
  assign n371 = n370 ^ n369 ;
  assign n372 = n214 ^ n213 ;
  assign n373 = n372 ^ n369 ;
  assign n374 = ~n371 & n373 ;
  assign n375 = n374 ^ n370 ;
  assign n376 = n375 ^ n216 ;
  assign n377 = n360 & n376 ;
  assign n378 = n377 ^ n216 ;
  assign n379 = n378 ^ n141 ;
  assign n380 = n359 & n379 ;
  assign n381 = n380 ^ n218 ;
  assign n382 = n372 ^ n370 ;
  assign n383 = ~n381 & ~n382 ;
  assign n384 = n383 ^ n370 ;
  assign n410 = n409 ^ n384 ;
  assign n413 = n277 ^ n275 ;
  assign n414 = n413 ^ n389 ;
  assign n415 = n407 & n414 ;
  assign n416 = n415 ^ n389 ;
  assign n411 = ~n363 & n381 ;
  assign n412 = n411 ^ n361 ;
  assign n417 = n416 ^ n412 ;
  assign n418 = n391 ^ n390 ;
  assign n419 = ~n407 & n418 ;
  assign n420 = n419 ^ n390 ;
  assign n421 = n365 ^ n364 ;
  assign n422 = ~n381 & n421 ;
  assign n423 = n422 ^ n364 ;
  assign n424 = ~n420 & n423 ;
  assign n425 = n424 ^ n412 ;
  assign n426 = ~n417 & n425 ;
  assign n427 = n426 ^ n412 ;
  assign n428 = n427 ^ n384 ;
  assign n429 = n410 & ~n428 ;
  assign n430 = n429 ^ n384 ;
  assign n431 = ~n355 & ~n430 ;
  assign n432 = n431 ^ n348 ;
  assign n433 = n432 ^ n348 ;
  assign n434 = ~n358 & ~n433 ;
  assign n435 = n434 ^ n348 ;
  assign n436 = ~n349 & n435 ;
  assign n437 = n436 ^ n220 ;
  assign n438 = n407 ^ n381 ;
  assign n439 = n437 & n438 ;
  assign n440 = n439 ^ n381 ;
  assign y0 = ~n440 ;
  assign y1 = n437 ;
endmodule
