module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 ;
  wire n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 ;
  assign n264 = ~x143 & ~x159 ;
  assign n265 = ~x175 & ~x191 ;
  assign n266 = n264 & n265 ;
  assign n267 = ~x207 & ~x223 ;
  assign n268 = ~x239 & ~x255 ;
  assign n269 = n267 & n268 ;
  assign n270 = n266 & n269 ;
  assign n257 = ~x15 & ~x31 ;
  assign n258 = ~x47 & ~x63 ;
  assign n259 = n257 & n258 ;
  assign n260 = ~x79 & ~x95 ;
  assign n261 = ~x111 & ~x127 ;
  assign n262 = n260 & n261 ;
  assign n263 = n259 & n262 ;
  assign n271 = n270 ^ n263 ;
  assign n1246 = x158 ^ x142 ;
  assign n1247 = x159 ^ x143 ;
  assign n1304 = x158 ^ x141 ;
  assign n1248 = x156 ^ x140 ;
  assign n1296 = x156 ^ x139 ;
  assign n1249 = x154 ^ x138 ;
  assign n1288 = x154 ^ x137 ;
  assign n1250 = x152 ^ x136 ;
  assign n1280 = x152 ^ x135 ;
  assign n1251 = x150 ^ x134 ;
  assign n1272 = x150 ^ x133 ;
  assign n1252 = x148 ^ x132 ;
  assign n1264 = x148 ^ x131 ;
  assign n1253 = x146 ^ x130 ;
  assign n1256 = x146 ^ x129 ;
  assign n1254 = x128 & ~x144 ;
  assign n1255 = n1254 ^ x146 ;
  assign n1257 = n1256 ^ n1255 ;
  assign n1258 = x145 ^ x129 ;
  assign n1259 = n1257 & ~n1258 ;
  assign n1260 = n1259 ^ n1256 ;
  assign n1261 = ~n1253 & n1260 ;
  assign n1262 = n1261 ^ x130 ;
  assign n1263 = n1262 ^ x148 ;
  assign n1265 = n1264 ^ n1263 ;
  assign n1266 = x147 ^ x131 ;
  assign n1267 = n1265 & ~n1266 ;
  assign n1268 = n1267 ^ n1264 ;
  assign n1269 = ~n1252 & n1268 ;
  assign n1270 = n1269 ^ x132 ;
  assign n1271 = n1270 ^ x150 ;
  assign n1273 = n1272 ^ n1271 ;
  assign n1274 = x149 ^ x133 ;
  assign n1275 = n1273 & ~n1274 ;
  assign n1276 = n1275 ^ n1272 ;
  assign n1277 = ~n1251 & n1276 ;
  assign n1278 = n1277 ^ x134 ;
  assign n1279 = n1278 ^ x152 ;
  assign n1281 = n1280 ^ n1279 ;
  assign n1282 = x151 ^ x135 ;
  assign n1283 = n1281 & ~n1282 ;
  assign n1284 = n1283 ^ n1280 ;
  assign n1285 = ~n1250 & n1284 ;
  assign n1286 = n1285 ^ x136 ;
  assign n1287 = n1286 ^ x154 ;
  assign n1289 = n1288 ^ n1287 ;
  assign n1290 = x153 ^ x137 ;
  assign n1291 = n1289 & ~n1290 ;
  assign n1292 = n1291 ^ n1288 ;
  assign n1293 = ~n1249 & n1292 ;
  assign n1294 = n1293 ^ x138 ;
  assign n1295 = n1294 ^ x156 ;
  assign n1297 = n1296 ^ n1295 ;
  assign n1298 = x155 ^ x139 ;
  assign n1299 = n1297 & ~n1298 ;
  assign n1300 = n1299 ^ n1296 ;
  assign n1301 = ~n1248 & n1300 ;
  assign n1302 = n1301 ^ x140 ;
  assign n1303 = n1302 ^ x158 ;
  assign n1305 = n1304 ^ n1303 ;
  assign n1306 = x157 ^ x141 ;
  assign n1307 = n1305 & ~n1306 ;
  assign n1308 = n1307 ^ n1304 ;
  assign n1309 = ~n1246 & n1308 ;
  assign n1310 = n1309 ^ x142 ;
  assign n1311 = n1310 ^ x159 ;
  assign n1312 = ~n1247 & n1311 ;
  assign n1313 = n1312 ^ x143 ;
  assign n1314 = n1246 & ~n1313 ;
  assign n1315 = n1314 ^ x142 ;
  assign n1176 = x190 ^ x174 ;
  assign n1177 = x191 ^ x175 ;
  assign n1234 = x190 ^ x173 ;
  assign n1178 = x188 ^ x172 ;
  assign n1226 = x188 ^ x171 ;
  assign n1179 = x186 ^ x170 ;
  assign n1218 = x186 ^ x169 ;
  assign n1180 = x184 ^ x168 ;
  assign n1210 = x184 ^ x167 ;
  assign n1181 = x182 ^ x166 ;
  assign n1202 = x182 ^ x165 ;
  assign n1182 = x180 ^ x164 ;
  assign n1194 = x180 ^ x163 ;
  assign n1183 = x178 ^ x162 ;
  assign n1186 = x178 ^ x161 ;
  assign n1184 = x160 & ~x176 ;
  assign n1185 = n1184 ^ x178 ;
  assign n1187 = n1186 ^ n1185 ;
  assign n1188 = x177 ^ x161 ;
  assign n1189 = n1187 & ~n1188 ;
  assign n1190 = n1189 ^ n1186 ;
  assign n1191 = ~n1183 & n1190 ;
  assign n1192 = n1191 ^ x162 ;
  assign n1193 = n1192 ^ x180 ;
  assign n1195 = n1194 ^ n1193 ;
  assign n1196 = x179 ^ x163 ;
  assign n1197 = n1195 & ~n1196 ;
  assign n1198 = n1197 ^ n1194 ;
  assign n1199 = ~n1182 & n1198 ;
  assign n1200 = n1199 ^ x164 ;
  assign n1201 = n1200 ^ x182 ;
  assign n1203 = n1202 ^ n1201 ;
  assign n1204 = x181 ^ x165 ;
  assign n1205 = n1203 & ~n1204 ;
  assign n1206 = n1205 ^ n1202 ;
  assign n1207 = ~n1181 & n1206 ;
  assign n1208 = n1207 ^ x166 ;
  assign n1209 = n1208 ^ x184 ;
  assign n1211 = n1210 ^ n1209 ;
  assign n1212 = x183 ^ x167 ;
  assign n1213 = n1211 & ~n1212 ;
  assign n1214 = n1213 ^ n1210 ;
  assign n1215 = ~n1180 & n1214 ;
  assign n1216 = n1215 ^ x168 ;
  assign n1217 = n1216 ^ x186 ;
  assign n1219 = n1218 ^ n1217 ;
  assign n1220 = x185 ^ x169 ;
  assign n1221 = n1219 & ~n1220 ;
  assign n1222 = n1221 ^ n1218 ;
  assign n1223 = ~n1179 & n1222 ;
  assign n1224 = n1223 ^ x170 ;
  assign n1225 = n1224 ^ x188 ;
  assign n1227 = n1226 ^ n1225 ;
  assign n1228 = x187 ^ x171 ;
  assign n1229 = n1227 & ~n1228 ;
  assign n1230 = n1229 ^ n1226 ;
  assign n1231 = ~n1178 & n1230 ;
  assign n1232 = n1231 ^ x172 ;
  assign n1233 = n1232 ^ x190 ;
  assign n1235 = n1234 ^ n1233 ;
  assign n1236 = x189 ^ x173 ;
  assign n1237 = n1235 & ~n1236 ;
  assign n1238 = n1237 ^ n1234 ;
  assign n1239 = ~n1176 & n1238 ;
  assign n1240 = n1239 ^ x174 ;
  assign n1241 = n1240 ^ x191 ;
  assign n1242 = ~n1177 & n1241 ;
  assign n1243 = n1242 ^ x175 ;
  assign n1244 = n1176 & ~n1243 ;
  assign n1245 = n1244 ^ x174 ;
  assign n1316 = n1315 ^ n1245 ;
  assign n1317 = n265 ^ n264 ;
  assign n1320 = n1306 & ~n1313 ;
  assign n1321 = n1320 ^ x141 ;
  assign n1318 = n1236 & ~n1243 ;
  assign n1319 = n1318 ^ x173 ;
  assign n1322 = n1321 ^ n1319 ;
  assign n1325 = n1248 & ~n1313 ;
  assign n1326 = n1325 ^ x140 ;
  assign n1323 = n1178 & ~n1243 ;
  assign n1324 = n1323 ^ x172 ;
  assign n1327 = n1326 ^ n1324 ;
  assign n1330 = n1298 & ~n1313 ;
  assign n1331 = n1330 ^ x139 ;
  assign n1328 = n1228 & ~n1243 ;
  assign n1329 = n1328 ^ x171 ;
  assign n1332 = n1331 ^ n1329 ;
  assign n1335 = n1249 & ~n1313 ;
  assign n1336 = n1335 ^ x138 ;
  assign n1333 = n1179 & ~n1243 ;
  assign n1334 = n1333 ^ x170 ;
  assign n1337 = n1336 ^ n1334 ;
  assign n1340 = n1220 & ~n1243 ;
  assign n1341 = n1340 ^ x169 ;
  assign n1338 = n1290 & ~n1313 ;
  assign n1339 = n1338 ^ x137 ;
  assign n1342 = n1341 ^ n1339 ;
  assign n1345 = n1250 & ~n1313 ;
  assign n1346 = n1345 ^ x136 ;
  assign n1343 = n1180 & ~n1243 ;
  assign n1344 = n1343 ^ x168 ;
  assign n1347 = n1346 ^ n1344 ;
  assign n1350 = n1212 & ~n1243 ;
  assign n1351 = n1350 ^ x167 ;
  assign n1348 = n1282 & ~n1313 ;
  assign n1349 = n1348 ^ x135 ;
  assign n1352 = n1351 ^ n1349 ;
  assign n1355 = n1181 & ~n1243 ;
  assign n1356 = n1355 ^ x166 ;
  assign n1353 = n1251 & ~n1313 ;
  assign n1354 = n1353 ^ x134 ;
  assign n1357 = n1356 ^ n1354 ;
  assign n1360 = n1204 & ~n1243 ;
  assign n1361 = n1360 ^ x165 ;
  assign n1358 = n1274 & ~n1313 ;
  assign n1359 = n1358 ^ x133 ;
  assign n1362 = n1361 ^ n1359 ;
  assign n1365 = n1252 & ~n1313 ;
  assign n1366 = n1365 ^ x132 ;
  assign n1363 = n1182 & ~n1243 ;
  assign n1364 = n1363 ^ x164 ;
  assign n1367 = n1366 ^ n1364 ;
  assign n1370 = n1196 & ~n1243 ;
  assign n1371 = n1370 ^ x163 ;
  assign n1368 = n1266 & ~n1313 ;
  assign n1369 = n1368 ^ x131 ;
  assign n1372 = n1371 ^ n1369 ;
  assign n1375 = n1183 & ~n1243 ;
  assign n1376 = n1375 ^ x162 ;
  assign n1373 = n1253 & ~n1313 ;
  assign n1374 = n1373 ^ x130 ;
  assign n1377 = n1376 ^ n1374 ;
  assign n1380 = n1258 & ~n1313 ;
  assign n1381 = n1380 ^ x129 ;
  assign n1378 = n1188 & ~n1243 ;
  assign n1379 = n1378 ^ x161 ;
  assign n1382 = n1381 ^ n1379 ;
  assign n1383 = x176 ^ x160 ;
  assign n1384 = ~n1243 & n1383 ;
  assign n1385 = n1384 ^ x160 ;
  assign n1386 = x144 ^ x128 ;
  assign n1387 = ~n1313 & n1386 ;
  assign n1388 = n1387 ^ x128 ;
  assign n1389 = ~n1385 & n1388 ;
  assign n1390 = n1389 ^ n1379 ;
  assign n1391 = ~n1382 & ~n1390 ;
  assign n1392 = n1391 ^ n1379 ;
  assign n1393 = n1392 ^ n1374 ;
  assign n1394 = ~n1377 & ~n1393 ;
  assign n1395 = n1394 ^ n1374 ;
  assign n1396 = n1395 ^ n1369 ;
  assign n1397 = ~n1372 & n1396 ;
  assign n1398 = n1397 ^ n1369 ;
  assign n1399 = n1398 ^ n1366 ;
  assign n1400 = ~n1367 & n1399 ;
  assign n1401 = n1400 ^ n1366 ;
  assign n1402 = n1401 ^ n1359 ;
  assign n1403 = ~n1362 & n1402 ;
  assign n1404 = n1403 ^ n1359 ;
  assign n1405 = n1404 ^ n1356 ;
  assign n1406 = ~n1357 & ~n1405 ;
  assign n1407 = n1406 ^ n1356 ;
  assign n1408 = n1407 ^ n1349 ;
  assign n1409 = ~n1352 & ~n1408 ;
  assign n1410 = n1409 ^ n1349 ;
  assign n1411 = n1410 ^ n1346 ;
  assign n1412 = ~n1347 & n1411 ;
  assign n1413 = n1412 ^ n1346 ;
  assign n1414 = n1413 ^ n1339 ;
  assign n1415 = ~n1342 & n1414 ;
  assign n1416 = n1415 ^ n1339 ;
  assign n1417 = n1416 ^ n1336 ;
  assign n1418 = ~n1337 & n1417 ;
  assign n1419 = n1418 ^ n1336 ;
  assign n1420 = n1419 ^ n1329 ;
  assign n1421 = ~n1332 & ~n1420 ;
  assign n1422 = n1421 ^ n1329 ;
  assign n1423 = n1422 ^ n1324 ;
  assign n1424 = ~n1327 & n1423 ;
  assign n1425 = n1424 ^ n1324 ;
  assign n1426 = n1425 ^ n1319 ;
  assign n1427 = ~n1322 & ~n1426 ;
  assign n1428 = n1427 ^ n1321 ;
  assign n1429 = n1428 ^ n1245 ;
  assign n1430 = ~n1316 & n1429 ;
  assign n1431 = n1430 ^ n1315 ;
  assign n1432 = n1431 ^ n265 ;
  assign n1433 = ~n1317 & ~n1432 ;
  assign n1434 = n1433 ^ n264 ;
  assign n1435 = n1316 & n1434 ;
  assign n1436 = n1435 ^ n1315 ;
  assign n985 = x254 ^ x238 ;
  assign n986 = x255 ^ x239 ;
  assign n1043 = x254 ^ x237 ;
  assign n987 = x252 ^ x236 ;
  assign n1035 = x252 ^ x235 ;
  assign n988 = x250 ^ x234 ;
  assign n1027 = x250 ^ x233 ;
  assign n989 = x248 ^ x232 ;
  assign n1019 = x248 ^ x231 ;
  assign n990 = x246 ^ x230 ;
  assign n1011 = x246 ^ x229 ;
  assign n991 = x244 ^ x228 ;
  assign n1003 = x244 ^ x227 ;
  assign n992 = x242 ^ x226 ;
  assign n995 = x242 ^ x225 ;
  assign n993 = x224 & ~x240 ;
  assign n994 = n993 ^ x242 ;
  assign n996 = n995 ^ n994 ;
  assign n997 = x241 ^ x225 ;
  assign n998 = n996 & ~n997 ;
  assign n999 = n998 ^ n995 ;
  assign n1000 = ~n992 & n999 ;
  assign n1001 = n1000 ^ x226 ;
  assign n1002 = n1001 ^ x244 ;
  assign n1004 = n1003 ^ n1002 ;
  assign n1005 = x243 ^ x227 ;
  assign n1006 = n1004 & ~n1005 ;
  assign n1007 = n1006 ^ n1003 ;
  assign n1008 = ~n991 & n1007 ;
  assign n1009 = n1008 ^ x228 ;
  assign n1010 = n1009 ^ x246 ;
  assign n1012 = n1011 ^ n1010 ;
  assign n1013 = x245 ^ x229 ;
  assign n1014 = n1012 & ~n1013 ;
  assign n1015 = n1014 ^ n1011 ;
  assign n1016 = ~n990 & n1015 ;
  assign n1017 = n1016 ^ x230 ;
  assign n1018 = n1017 ^ x248 ;
  assign n1020 = n1019 ^ n1018 ;
  assign n1021 = x247 ^ x231 ;
  assign n1022 = n1020 & ~n1021 ;
  assign n1023 = n1022 ^ n1019 ;
  assign n1024 = ~n989 & n1023 ;
  assign n1025 = n1024 ^ x232 ;
  assign n1026 = n1025 ^ x250 ;
  assign n1028 = n1027 ^ n1026 ;
  assign n1029 = x249 ^ x233 ;
  assign n1030 = n1028 & ~n1029 ;
  assign n1031 = n1030 ^ n1027 ;
  assign n1032 = ~n988 & n1031 ;
  assign n1033 = n1032 ^ x234 ;
  assign n1034 = n1033 ^ x252 ;
  assign n1036 = n1035 ^ n1034 ;
  assign n1037 = x251 ^ x235 ;
  assign n1038 = n1036 & ~n1037 ;
  assign n1039 = n1038 ^ n1035 ;
  assign n1040 = ~n987 & n1039 ;
  assign n1041 = n1040 ^ x236 ;
  assign n1042 = n1041 ^ x254 ;
  assign n1044 = n1043 ^ n1042 ;
  assign n1045 = x253 ^ x237 ;
  assign n1046 = n1044 & ~n1045 ;
  assign n1047 = n1046 ^ n1043 ;
  assign n1048 = ~n985 & n1047 ;
  assign n1049 = n1048 ^ x238 ;
  assign n1050 = n1049 ^ x255 ;
  assign n1051 = ~n986 & n1050 ;
  assign n1052 = n1051 ^ x239 ;
  assign n1053 = n985 & ~n1052 ;
  assign n1054 = n1053 ^ x238 ;
  assign n915 = x222 ^ x206 ;
  assign n916 = x223 ^ x207 ;
  assign n973 = x222 ^ x205 ;
  assign n917 = x220 ^ x204 ;
  assign n965 = x220 ^ x203 ;
  assign n918 = x218 ^ x202 ;
  assign n957 = x218 ^ x201 ;
  assign n919 = x216 ^ x200 ;
  assign n949 = x216 ^ x199 ;
  assign n920 = x214 ^ x198 ;
  assign n941 = x214 ^ x197 ;
  assign n921 = x212 ^ x196 ;
  assign n933 = x212 ^ x195 ;
  assign n922 = x210 ^ x194 ;
  assign n925 = x210 ^ x193 ;
  assign n923 = x192 & ~x208 ;
  assign n924 = n923 ^ x210 ;
  assign n926 = n925 ^ n924 ;
  assign n927 = x209 ^ x193 ;
  assign n928 = n926 & ~n927 ;
  assign n929 = n928 ^ n925 ;
  assign n930 = ~n922 & n929 ;
  assign n931 = n930 ^ x194 ;
  assign n932 = n931 ^ x212 ;
  assign n934 = n933 ^ n932 ;
  assign n935 = x211 ^ x195 ;
  assign n936 = n934 & ~n935 ;
  assign n937 = n936 ^ n933 ;
  assign n938 = ~n921 & n937 ;
  assign n939 = n938 ^ x196 ;
  assign n940 = n939 ^ x214 ;
  assign n942 = n941 ^ n940 ;
  assign n943 = x213 ^ x197 ;
  assign n944 = n942 & ~n943 ;
  assign n945 = n944 ^ n941 ;
  assign n946 = ~n920 & n945 ;
  assign n947 = n946 ^ x198 ;
  assign n948 = n947 ^ x216 ;
  assign n950 = n949 ^ n948 ;
  assign n951 = x215 ^ x199 ;
  assign n952 = n950 & ~n951 ;
  assign n953 = n952 ^ n949 ;
  assign n954 = ~n919 & n953 ;
  assign n955 = n954 ^ x200 ;
  assign n956 = n955 ^ x218 ;
  assign n958 = n957 ^ n956 ;
  assign n959 = x217 ^ x201 ;
  assign n960 = n958 & ~n959 ;
  assign n961 = n960 ^ n957 ;
  assign n962 = ~n918 & n961 ;
  assign n963 = n962 ^ x202 ;
  assign n964 = n963 ^ x220 ;
  assign n966 = n965 ^ n964 ;
  assign n967 = x219 ^ x203 ;
  assign n968 = n966 & ~n967 ;
  assign n969 = n968 ^ n965 ;
  assign n970 = ~n917 & n969 ;
  assign n971 = n970 ^ x204 ;
  assign n972 = n971 ^ x222 ;
  assign n974 = n973 ^ n972 ;
  assign n975 = x221 ^ x205 ;
  assign n976 = n974 & ~n975 ;
  assign n977 = n976 ^ n973 ;
  assign n978 = ~n915 & n977 ;
  assign n979 = n978 ^ x206 ;
  assign n980 = n979 ^ x223 ;
  assign n981 = ~n916 & n980 ;
  assign n982 = n981 ^ x207 ;
  assign n983 = n915 & ~n982 ;
  assign n984 = n983 ^ x206 ;
  assign n1055 = n1054 ^ n984 ;
  assign n1056 = n268 ^ n267 ;
  assign n1059 = n975 & ~n982 ;
  assign n1060 = n1059 ^ x205 ;
  assign n1057 = n1045 & ~n1052 ;
  assign n1058 = n1057 ^ x237 ;
  assign n1061 = n1060 ^ n1058 ;
  assign n1064 = n917 & ~n982 ;
  assign n1065 = n1064 ^ x204 ;
  assign n1062 = n987 & ~n1052 ;
  assign n1063 = n1062 ^ x236 ;
  assign n1066 = n1065 ^ n1063 ;
  assign n1069 = n1037 & ~n1052 ;
  assign n1070 = n1069 ^ x235 ;
  assign n1067 = n967 & ~n982 ;
  assign n1068 = n1067 ^ x203 ;
  assign n1071 = n1070 ^ n1068 ;
  assign n1074 = n918 & ~n982 ;
  assign n1075 = n1074 ^ x202 ;
  assign n1072 = n988 & ~n1052 ;
  assign n1073 = n1072 ^ x234 ;
  assign n1076 = n1075 ^ n1073 ;
  assign n1079 = n959 & ~n982 ;
  assign n1080 = n1079 ^ x201 ;
  assign n1077 = n1029 & ~n1052 ;
  assign n1078 = n1077 ^ x233 ;
  assign n1081 = n1080 ^ n1078 ;
  assign n1084 = n919 & ~n982 ;
  assign n1085 = n1084 ^ x200 ;
  assign n1082 = n989 & ~n1052 ;
  assign n1083 = n1082 ^ x232 ;
  assign n1086 = n1085 ^ n1083 ;
  assign n1089 = n1021 & ~n1052 ;
  assign n1090 = n1089 ^ x231 ;
  assign n1087 = n951 & ~n982 ;
  assign n1088 = n1087 ^ x199 ;
  assign n1091 = n1090 ^ n1088 ;
  assign n1094 = n920 & ~n982 ;
  assign n1095 = n1094 ^ x198 ;
  assign n1092 = n990 & ~n1052 ;
  assign n1093 = n1092 ^ x230 ;
  assign n1096 = n1095 ^ n1093 ;
  assign n1099 = n1013 & ~n1052 ;
  assign n1100 = n1099 ^ x229 ;
  assign n1097 = n943 & ~n982 ;
  assign n1098 = n1097 ^ x197 ;
  assign n1101 = n1100 ^ n1098 ;
  assign n1104 = n921 & ~n982 ;
  assign n1105 = n1104 ^ x196 ;
  assign n1102 = n991 & ~n1052 ;
  assign n1103 = n1102 ^ x228 ;
  assign n1106 = n1105 ^ n1103 ;
  assign n1109 = n1005 & ~n1052 ;
  assign n1110 = n1109 ^ x227 ;
  assign n1107 = n935 & ~n982 ;
  assign n1108 = n1107 ^ x195 ;
  assign n1111 = n1110 ^ n1108 ;
  assign n1114 = n992 & ~n1052 ;
  assign n1115 = n1114 ^ x226 ;
  assign n1112 = n922 & ~n982 ;
  assign n1113 = n1112 ^ x194 ;
  assign n1116 = n1115 ^ n1113 ;
  assign n1119 = n927 & ~n982 ;
  assign n1120 = n1119 ^ x193 ;
  assign n1117 = n997 & ~n1052 ;
  assign n1118 = n1117 ^ x225 ;
  assign n1121 = n1120 ^ n1118 ;
  assign n1122 = x240 ^ x224 ;
  assign n1123 = ~n1052 & n1122 ;
  assign n1124 = n1123 ^ x224 ;
  assign n1125 = x208 ^ x192 ;
  assign n1126 = ~n982 & n1125 ;
  assign n1127 = n1126 ^ x192 ;
  assign n1128 = ~n1124 & n1127 ;
  assign n1129 = n1128 ^ n1118 ;
  assign n1130 = ~n1121 & ~n1129 ;
  assign n1131 = n1130 ^ n1118 ;
  assign n1132 = n1131 ^ n1113 ;
  assign n1133 = ~n1116 & ~n1132 ;
  assign n1134 = n1133 ^ n1113 ;
  assign n1135 = n1134 ^ n1108 ;
  assign n1136 = ~n1111 & n1135 ;
  assign n1137 = n1136 ^ n1108 ;
  assign n1138 = n1137 ^ n1105 ;
  assign n1139 = ~n1106 & n1138 ;
  assign n1140 = n1139 ^ n1105 ;
  assign n1141 = n1140 ^ n1098 ;
  assign n1142 = ~n1101 & n1141 ;
  assign n1143 = n1142 ^ n1098 ;
  assign n1144 = n1143 ^ n1095 ;
  assign n1145 = ~n1096 & n1144 ;
  assign n1146 = n1145 ^ n1095 ;
  assign n1147 = n1146 ^ n1088 ;
  assign n1148 = ~n1091 & n1147 ;
  assign n1149 = n1148 ^ n1088 ;
  assign n1150 = n1149 ^ n1085 ;
  assign n1151 = ~n1086 & n1150 ;
  assign n1152 = n1151 ^ n1085 ;
  assign n1153 = n1152 ^ n1078 ;
  assign n1154 = ~n1081 & ~n1153 ;
  assign n1155 = n1154 ^ n1078 ;
  assign n1156 = n1155 ^ n1075 ;
  assign n1157 = ~n1076 & ~n1156 ;
  assign n1158 = n1157 ^ n1075 ;
  assign n1159 = n1158 ^ n1068 ;
  assign n1160 = ~n1071 & n1159 ;
  assign n1161 = n1160 ^ n1068 ;
  assign n1162 = n1161 ^ n1063 ;
  assign n1163 = ~n1066 & ~n1162 ;
  assign n1164 = n1163 ^ n1063 ;
  assign n1165 = n1164 ^ n1058 ;
  assign n1166 = ~n1061 & ~n1165 ;
  assign n1167 = n1166 ^ n1060 ;
  assign n1168 = n1167 ^ n984 ;
  assign n1169 = ~n1055 & ~n1168 ;
  assign n1170 = n1169 ^ n1054 ;
  assign n1171 = n1170 ^ n268 ;
  assign n1172 = ~n1056 & n1171 ;
  assign n1173 = n1172 ^ n267 ;
  assign n1174 = n1055 & ~n1173 ;
  assign n1175 = n1174 ^ n1054 ;
  assign n1437 = n1436 ^ n1175 ;
  assign n1438 = n269 ^ n266 ;
  assign n1441 = n1322 & ~n1434 ;
  assign n1442 = n1441 ^ n1319 ;
  assign n1439 = n1061 & ~n1173 ;
  assign n1440 = n1439 ^ n1058 ;
  assign n1443 = n1442 ^ n1440 ;
  assign n1446 = n1066 & ~n1173 ;
  assign n1447 = n1446 ^ n1063 ;
  assign n1444 = n1327 & ~n1434 ;
  assign n1445 = n1444 ^ n1324 ;
  assign n1448 = n1447 ^ n1445 ;
  assign n1451 = n1332 & ~n1434 ;
  assign n1452 = n1451 ^ n1329 ;
  assign n1449 = n1071 & n1173 ;
  assign n1450 = n1449 ^ n1068 ;
  assign n1453 = n1452 ^ n1450 ;
  assign n1456 = n1076 & n1173 ;
  assign n1457 = n1456 ^ n1075 ;
  assign n1454 = n1337 & n1434 ;
  assign n1455 = n1454 ^ n1336 ;
  assign n1458 = n1457 ^ n1455 ;
  assign n1461 = n1342 & ~n1434 ;
  assign n1462 = n1461 ^ n1341 ;
  assign n1459 = n1081 & n1173 ;
  assign n1460 = n1459 ^ n1080 ;
  assign n1463 = n1462 ^ n1460 ;
  assign n1466 = n1347 & ~n1434 ;
  assign n1467 = n1466 ^ n1344 ;
  assign n1464 = n1086 & ~n1173 ;
  assign n1465 = n1464 ^ n1083 ;
  assign n1468 = n1467 ^ n1465 ;
  assign n1471 = n1091 & n1173 ;
  assign n1472 = n1471 ^ n1088 ;
  assign n1469 = n1352 & n1434 ;
  assign n1470 = n1469 ^ n1349 ;
  assign n1473 = n1472 ^ n1470 ;
  assign n1476 = n1096 & n1173 ;
  assign n1477 = n1476 ^ n1095 ;
  assign n1474 = n1357 & ~n1434 ;
  assign n1475 = n1474 ^ n1356 ;
  assign n1478 = n1477 ^ n1475 ;
  assign n1481 = n1362 & ~n1434 ;
  assign n1482 = n1481 ^ n1361 ;
  assign n1479 = n1101 & ~n1173 ;
  assign n1480 = n1479 ^ n1100 ;
  assign n1483 = n1482 ^ n1480 ;
  assign n1486 = n1367 & ~n1434 ;
  assign n1487 = n1486 ^ n1364 ;
  assign n1484 = n1106 & ~n1173 ;
  assign n1485 = n1484 ^ n1103 ;
  assign n1488 = n1487 ^ n1485 ;
  assign n1491 = n1372 & n1434 ;
  assign n1492 = n1491 ^ n1369 ;
  assign n1489 = n1111 & n1173 ;
  assign n1490 = n1489 ^ n1108 ;
  assign n1493 = n1492 ^ n1490 ;
  assign n1496 = n1116 & ~n1173 ;
  assign n1497 = n1496 ^ n1115 ;
  assign n1494 = n1377 & ~n1434 ;
  assign n1495 = n1494 ^ n1376 ;
  assign n1498 = n1497 ^ n1495 ;
  assign n1501 = n1382 & n1434 ;
  assign n1502 = n1501 ^ n1381 ;
  assign n1499 = n1121 & n1173 ;
  assign n1500 = n1499 ^ n1120 ;
  assign n1503 = n1502 ^ n1500 ;
  assign n1504 = n1127 ^ n1124 ;
  assign n1505 = ~n1173 & n1504 ;
  assign n1506 = n1505 ^ n1124 ;
  assign n1507 = n1388 ^ n1385 ;
  assign n1508 = ~n1434 & n1507 ;
  assign n1509 = n1508 ^ n1385 ;
  assign n1510 = ~n1506 & n1509 ;
  assign n1511 = n1510 ^ n1500 ;
  assign n1512 = ~n1503 & ~n1511 ;
  assign n1513 = n1512 ^ n1500 ;
  assign n1514 = n1513 ^ n1497 ;
  assign n1515 = ~n1498 & n1514 ;
  assign n1516 = n1515 ^ n1497 ;
  assign n1517 = n1516 ^ n1490 ;
  assign n1518 = ~n1493 & n1517 ;
  assign n1519 = n1518 ^ n1490 ;
  assign n1520 = n1519 ^ n1487 ;
  assign n1521 = ~n1488 & ~n1520 ;
  assign n1522 = n1521 ^ n1487 ;
  assign n1523 = n1522 ^ n1480 ;
  assign n1524 = ~n1483 & ~n1523 ;
  assign n1525 = n1524 ^ n1480 ;
  assign n1526 = n1525 ^ n1477 ;
  assign n1527 = ~n1478 & n1526 ;
  assign n1528 = n1527 ^ n1477 ;
  assign n1529 = n1528 ^ n1470 ;
  assign n1530 = ~n1473 & ~n1529 ;
  assign n1531 = n1530 ^ n1470 ;
  assign n1532 = n1531 ^ n1467 ;
  assign n1533 = ~n1468 & n1532 ;
  assign n1534 = n1533 ^ n1467 ;
  assign n1535 = n1534 ^ n1460 ;
  assign n1536 = ~n1463 & ~n1535 ;
  assign n1537 = n1536 ^ n1460 ;
  assign n1538 = n1537 ^ n1457 ;
  assign n1539 = ~n1458 & n1538 ;
  assign n1540 = n1539 ^ n1457 ;
  assign n1541 = n1540 ^ n1450 ;
  assign n1542 = ~n1453 & n1541 ;
  assign n1543 = n1542 ^ n1450 ;
  assign n1544 = n1543 ^ n1447 ;
  assign n1545 = ~n1448 & n1544 ;
  assign n1546 = n1545 ^ n1447 ;
  assign n1547 = n1546 ^ n1442 ;
  assign n1548 = ~n1443 & ~n1547 ;
  assign n1549 = n1548 ^ n1442 ;
  assign n1550 = n1549 ^ n1436 ;
  assign n1551 = ~n1437 & ~n1550 ;
  assign n1552 = n1551 ^ n1175 ;
  assign n1553 = n1552 ^ n269 ;
  assign n1554 = ~n1438 & n1553 ;
  assign n1555 = n1554 ^ n266 ;
  assign n1556 = n1437 & n1555 ;
  assign n1557 = n1556 ^ n1436 ;
  assign n603 = x30 ^ x14 ;
  assign n604 = x31 ^ x15 ;
  assign n661 = x30 ^ x13 ;
  assign n605 = x28 ^ x12 ;
  assign n653 = x28 ^ x11 ;
  assign n606 = x26 ^ x10 ;
  assign n645 = x26 ^ x9 ;
  assign n607 = x24 ^ x8 ;
  assign n637 = x24 ^ x7 ;
  assign n608 = x22 ^ x6 ;
  assign n629 = x22 ^ x5 ;
  assign n609 = x20 ^ x4 ;
  assign n621 = x20 ^ x3 ;
  assign n610 = x18 ^ x2 ;
  assign n613 = x18 ^ x1 ;
  assign n611 = x0 & ~x16 ;
  assign n612 = n611 ^ x18 ;
  assign n614 = n613 ^ n612 ;
  assign n615 = x17 ^ x1 ;
  assign n616 = n614 & ~n615 ;
  assign n617 = n616 ^ n613 ;
  assign n618 = ~n610 & n617 ;
  assign n619 = n618 ^ x2 ;
  assign n620 = n619 ^ x20 ;
  assign n622 = n621 ^ n620 ;
  assign n623 = x19 ^ x3 ;
  assign n624 = n622 & ~n623 ;
  assign n625 = n624 ^ n621 ;
  assign n626 = ~n609 & n625 ;
  assign n627 = n626 ^ x4 ;
  assign n628 = n627 ^ x22 ;
  assign n630 = n629 ^ n628 ;
  assign n631 = x21 ^ x5 ;
  assign n632 = n630 & ~n631 ;
  assign n633 = n632 ^ n629 ;
  assign n634 = ~n608 & n633 ;
  assign n635 = n634 ^ x6 ;
  assign n636 = n635 ^ x24 ;
  assign n638 = n637 ^ n636 ;
  assign n639 = x23 ^ x7 ;
  assign n640 = n638 & ~n639 ;
  assign n641 = n640 ^ n637 ;
  assign n642 = ~n607 & n641 ;
  assign n643 = n642 ^ x8 ;
  assign n644 = n643 ^ x26 ;
  assign n646 = n645 ^ n644 ;
  assign n647 = x25 ^ x9 ;
  assign n648 = n646 & ~n647 ;
  assign n649 = n648 ^ n645 ;
  assign n650 = ~n606 & n649 ;
  assign n651 = n650 ^ x10 ;
  assign n652 = n651 ^ x28 ;
  assign n654 = n653 ^ n652 ;
  assign n655 = x27 ^ x11 ;
  assign n656 = n654 & ~n655 ;
  assign n657 = n656 ^ n653 ;
  assign n658 = ~n605 & n657 ;
  assign n659 = n658 ^ x12 ;
  assign n660 = n659 ^ x30 ;
  assign n662 = n661 ^ n660 ;
  assign n663 = x29 ^ x13 ;
  assign n664 = n662 & ~n663 ;
  assign n665 = n664 ^ n661 ;
  assign n666 = ~n603 & n665 ;
  assign n667 = n666 ^ x14 ;
  assign n668 = n667 ^ x31 ;
  assign n669 = ~n604 & n668 ;
  assign n670 = n669 ^ x15 ;
  assign n671 = n603 & ~n670 ;
  assign n672 = n671 ^ x14 ;
  assign n533 = x62 ^ x46 ;
  assign n534 = x63 ^ x47 ;
  assign n591 = x62 ^ x45 ;
  assign n535 = x60 ^ x44 ;
  assign n583 = x60 ^ x43 ;
  assign n536 = x58 ^ x42 ;
  assign n575 = x58 ^ x41 ;
  assign n537 = x56 ^ x40 ;
  assign n567 = x56 ^ x39 ;
  assign n538 = x54 ^ x38 ;
  assign n559 = x54 ^ x37 ;
  assign n539 = x52 ^ x36 ;
  assign n551 = x52 ^ x35 ;
  assign n540 = x50 ^ x34 ;
  assign n543 = x50 ^ x33 ;
  assign n541 = x32 & ~x48 ;
  assign n542 = n541 ^ x50 ;
  assign n544 = n543 ^ n542 ;
  assign n545 = x49 ^ x33 ;
  assign n546 = n544 & ~n545 ;
  assign n547 = n546 ^ n543 ;
  assign n548 = ~n540 & n547 ;
  assign n549 = n548 ^ x34 ;
  assign n550 = n549 ^ x52 ;
  assign n552 = n551 ^ n550 ;
  assign n553 = x51 ^ x35 ;
  assign n554 = n552 & ~n553 ;
  assign n555 = n554 ^ n551 ;
  assign n556 = ~n539 & n555 ;
  assign n557 = n556 ^ x36 ;
  assign n558 = n557 ^ x54 ;
  assign n560 = n559 ^ n558 ;
  assign n561 = x53 ^ x37 ;
  assign n562 = n560 & ~n561 ;
  assign n563 = n562 ^ n559 ;
  assign n564 = ~n538 & n563 ;
  assign n565 = n564 ^ x38 ;
  assign n566 = n565 ^ x56 ;
  assign n568 = n567 ^ n566 ;
  assign n569 = x55 ^ x39 ;
  assign n570 = n568 & ~n569 ;
  assign n571 = n570 ^ n567 ;
  assign n572 = ~n537 & n571 ;
  assign n573 = n572 ^ x40 ;
  assign n574 = n573 ^ x58 ;
  assign n576 = n575 ^ n574 ;
  assign n577 = x57 ^ x41 ;
  assign n578 = n576 & ~n577 ;
  assign n579 = n578 ^ n575 ;
  assign n580 = ~n536 & n579 ;
  assign n581 = n580 ^ x42 ;
  assign n582 = n581 ^ x60 ;
  assign n584 = n583 ^ n582 ;
  assign n585 = x59 ^ x43 ;
  assign n586 = n584 & ~n585 ;
  assign n587 = n586 ^ n583 ;
  assign n588 = ~n535 & n587 ;
  assign n589 = n588 ^ x44 ;
  assign n590 = n589 ^ x62 ;
  assign n592 = n591 ^ n590 ;
  assign n593 = x61 ^ x45 ;
  assign n594 = n592 & ~n593 ;
  assign n595 = n594 ^ n591 ;
  assign n596 = ~n533 & n595 ;
  assign n597 = n596 ^ x46 ;
  assign n598 = n597 ^ x63 ;
  assign n599 = ~n534 & n598 ;
  assign n600 = n599 ^ x47 ;
  assign n601 = n533 & ~n600 ;
  assign n602 = n601 ^ x46 ;
  assign n673 = n672 ^ n602 ;
  assign n674 = n258 ^ n257 ;
  assign n677 = n663 & ~n670 ;
  assign n678 = n677 ^ x13 ;
  assign n675 = n593 & ~n600 ;
  assign n676 = n675 ^ x45 ;
  assign n679 = n678 ^ n676 ;
  assign n682 = n605 & ~n670 ;
  assign n683 = n682 ^ x12 ;
  assign n680 = n535 & ~n600 ;
  assign n681 = n680 ^ x44 ;
  assign n684 = n683 ^ n681 ;
  assign n687 = n655 & ~n670 ;
  assign n688 = n687 ^ x11 ;
  assign n685 = n585 & ~n600 ;
  assign n686 = n685 ^ x43 ;
  assign n689 = n688 ^ n686 ;
  assign n692 = n536 & ~n600 ;
  assign n693 = n692 ^ x42 ;
  assign n690 = n606 & ~n670 ;
  assign n691 = n690 ^ x10 ;
  assign n694 = n693 ^ n691 ;
  assign n697 = n647 & ~n670 ;
  assign n698 = n697 ^ x9 ;
  assign n695 = n577 & ~n600 ;
  assign n696 = n695 ^ x41 ;
  assign n699 = n698 ^ n696 ;
  assign n702 = n607 & ~n670 ;
  assign n703 = n702 ^ x8 ;
  assign n700 = n537 & ~n600 ;
  assign n701 = n700 ^ x40 ;
  assign n704 = n703 ^ n701 ;
  assign n707 = n569 & ~n600 ;
  assign n708 = n707 ^ x39 ;
  assign n705 = n639 & ~n670 ;
  assign n706 = n705 ^ x7 ;
  assign n709 = n708 ^ n706 ;
  assign n712 = n538 & ~n600 ;
  assign n713 = n712 ^ x38 ;
  assign n710 = n608 & ~n670 ;
  assign n711 = n710 ^ x6 ;
  assign n714 = n713 ^ n711 ;
  assign n717 = n561 & ~n600 ;
  assign n718 = n717 ^ x37 ;
  assign n715 = n631 & ~n670 ;
  assign n716 = n715 ^ x5 ;
  assign n719 = n718 ^ n716 ;
  assign n722 = n539 & ~n600 ;
  assign n723 = n722 ^ x36 ;
  assign n720 = n609 & ~n670 ;
  assign n721 = n720 ^ x4 ;
  assign n724 = n723 ^ n721 ;
  assign n727 = n553 & ~n600 ;
  assign n728 = n727 ^ x35 ;
  assign n725 = n623 & ~n670 ;
  assign n726 = n725 ^ x3 ;
  assign n729 = n728 ^ n726 ;
  assign n732 = n540 & ~n600 ;
  assign n733 = n732 ^ x34 ;
  assign n730 = n610 & ~n670 ;
  assign n731 = n730 ^ x2 ;
  assign n734 = n733 ^ n731 ;
  assign n737 = n615 & ~n670 ;
  assign n738 = n737 ^ x1 ;
  assign n735 = n545 & ~n600 ;
  assign n736 = n735 ^ x33 ;
  assign n739 = n738 ^ n736 ;
  assign n740 = x16 ^ x0 ;
  assign n741 = ~n670 & n740 ;
  assign n742 = n741 ^ x0 ;
  assign n743 = x48 ^ x32 ;
  assign n744 = ~n600 & n743 ;
  assign n745 = n744 ^ x32 ;
  assign n746 = n742 & ~n745 ;
  assign n747 = n746 ^ n736 ;
  assign n748 = ~n739 & ~n747 ;
  assign n749 = n748 ^ n736 ;
  assign n750 = n749 ^ n731 ;
  assign n751 = ~n734 & ~n750 ;
  assign n752 = n751 ^ n731 ;
  assign n753 = n752 ^ n726 ;
  assign n754 = ~n729 & n753 ;
  assign n755 = n754 ^ n726 ;
  assign n756 = n755 ^ n723 ;
  assign n757 = ~n724 & ~n756 ;
  assign n758 = n757 ^ n723 ;
  assign n759 = n758 ^ n716 ;
  assign n760 = ~n719 & ~n759 ;
  assign n761 = n760 ^ n716 ;
  assign n762 = n761 ^ n713 ;
  assign n763 = ~n714 & ~n762 ;
  assign n764 = n763 ^ n713 ;
  assign n765 = n764 ^ n706 ;
  assign n766 = ~n709 & ~n765 ;
  assign n767 = n766 ^ n706 ;
  assign n768 = n767 ^ n703 ;
  assign n769 = ~n704 & n768 ;
  assign n770 = n769 ^ n703 ;
  assign n771 = n770 ^ n696 ;
  assign n772 = ~n699 & ~n771 ;
  assign n773 = n772 ^ n696 ;
  assign n774 = n773 ^ n693 ;
  assign n775 = ~n694 & n774 ;
  assign n776 = n775 ^ n693 ;
  assign n777 = n776 ^ n686 ;
  assign n778 = ~n689 & n777 ;
  assign n779 = n778 ^ n686 ;
  assign n780 = n779 ^ n681 ;
  assign n781 = ~n684 & n780 ;
  assign n782 = n781 ^ n681 ;
  assign n783 = n782 ^ n676 ;
  assign n784 = ~n679 & ~n783 ;
  assign n785 = n784 ^ n678 ;
  assign n786 = n785 ^ n602 ;
  assign n787 = ~n673 & n786 ;
  assign n788 = n787 ^ n672 ;
  assign n789 = n788 ^ n258 ;
  assign n790 = ~n674 & ~n789 ;
  assign n791 = n790 ^ n257 ;
  assign n792 = n673 & n791 ;
  assign n793 = n792 ^ n672 ;
  assign n342 = x126 ^ x110 ;
  assign n343 = x127 ^ x111 ;
  assign n400 = x126 ^ x109 ;
  assign n344 = x124 ^ x108 ;
  assign n392 = x124 ^ x107 ;
  assign n345 = x122 ^ x106 ;
  assign n384 = x122 ^ x105 ;
  assign n346 = x120 ^ x104 ;
  assign n376 = x120 ^ x103 ;
  assign n347 = x118 ^ x102 ;
  assign n368 = x118 ^ x101 ;
  assign n348 = x116 ^ x100 ;
  assign n360 = x116 ^ x99 ;
  assign n349 = x114 ^ x98 ;
  assign n352 = x114 ^ x97 ;
  assign n350 = x96 & ~x112 ;
  assign n351 = n350 ^ x114 ;
  assign n353 = n352 ^ n351 ;
  assign n354 = x113 ^ x97 ;
  assign n355 = n353 & ~n354 ;
  assign n356 = n355 ^ n352 ;
  assign n357 = ~n349 & n356 ;
  assign n358 = n357 ^ x98 ;
  assign n359 = n358 ^ x116 ;
  assign n361 = n360 ^ n359 ;
  assign n362 = x115 ^ x99 ;
  assign n363 = n361 & ~n362 ;
  assign n364 = n363 ^ n360 ;
  assign n365 = ~n348 & n364 ;
  assign n366 = n365 ^ x100 ;
  assign n367 = n366 ^ x118 ;
  assign n369 = n368 ^ n367 ;
  assign n370 = x117 ^ x101 ;
  assign n371 = n369 & ~n370 ;
  assign n372 = n371 ^ n368 ;
  assign n373 = ~n347 & n372 ;
  assign n374 = n373 ^ x102 ;
  assign n375 = n374 ^ x120 ;
  assign n377 = n376 ^ n375 ;
  assign n378 = x119 ^ x103 ;
  assign n379 = n377 & ~n378 ;
  assign n380 = n379 ^ n376 ;
  assign n381 = ~n346 & n380 ;
  assign n382 = n381 ^ x104 ;
  assign n383 = n382 ^ x122 ;
  assign n385 = n384 ^ n383 ;
  assign n386 = x121 ^ x105 ;
  assign n387 = n385 & ~n386 ;
  assign n388 = n387 ^ n384 ;
  assign n389 = ~n345 & n388 ;
  assign n390 = n389 ^ x106 ;
  assign n391 = n390 ^ x124 ;
  assign n393 = n392 ^ n391 ;
  assign n394 = x123 ^ x107 ;
  assign n395 = n393 & ~n394 ;
  assign n396 = n395 ^ n392 ;
  assign n397 = ~n344 & n396 ;
  assign n398 = n397 ^ x108 ;
  assign n399 = n398 ^ x126 ;
  assign n401 = n400 ^ n399 ;
  assign n402 = x125 ^ x109 ;
  assign n403 = n401 & ~n402 ;
  assign n404 = n403 ^ n400 ;
  assign n405 = ~n342 & n404 ;
  assign n406 = n405 ^ x110 ;
  assign n407 = n406 ^ x127 ;
  assign n408 = ~n343 & n407 ;
  assign n409 = n408 ^ x111 ;
  assign n410 = n342 & ~n409 ;
  assign n411 = n410 ^ x110 ;
  assign n272 = x94 ^ x78 ;
  assign n273 = x95 ^ x79 ;
  assign n330 = x94 ^ x77 ;
  assign n274 = x92 ^ x76 ;
  assign n322 = x92 ^ x75 ;
  assign n275 = x90 ^ x74 ;
  assign n314 = x90 ^ x73 ;
  assign n276 = x88 ^ x72 ;
  assign n306 = x88 ^ x71 ;
  assign n277 = x86 ^ x70 ;
  assign n298 = x86 ^ x69 ;
  assign n278 = x84 ^ x68 ;
  assign n290 = x84 ^ x67 ;
  assign n279 = x82 ^ x66 ;
  assign n282 = x82 ^ x65 ;
  assign n280 = x64 & ~x80 ;
  assign n281 = n280 ^ x82 ;
  assign n283 = n282 ^ n281 ;
  assign n284 = x81 ^ x65 ;
  assign n285 = n283 & ~n284 ;
  assign n286 = n285 ^ n282 ;
  assign n287 = ~n279 & n286 ;
  assign n288 = n287 ^ x66 ;
  assign n289 = n288 ^ x84 ;
  assign n291 = n290 ^ n289 ;
  assign n292 = x83 ^ x67 ;
  assign n293 = n291 & ~n292 ;
  assign n294 = n293 ^ n290 ;
  assign n295 = ~n278 & n294 ;
  assign n296 = n295 ^ x68 ;
  assign n297 = n296 ^ x86 ;
  assign n299 = n298 ^ n297 ;
  assign n300 = x85 ^ x69 ;
  assign n301 = n299 & ~n300 ;
  assign n302 = n301 ^ n298 ;
  assign n303 = ~n277 & n302 ;
  assign n304 = n303 ^ x70 ;
  assign n305 = n304 ^ x88 ;
  assign n307 = n306 ^ n305 ;
  assign n308 = x87 ^ x71 ;
  assign n309 = n307 & ~n308 ;
  assign n310 = n309 ^ n306 ;
  assign n311 = ~n276 & n310 ;
  assign n312 = n311 ^ x72 ;
  assign n313 = n312 ^ x90 ;
  assign n315 = n314 ^ n313 ;
  assign n316 = x89 ^ x73 ;
  assign n317 = n315 & ~n316 ;
  assign n318 = n317 ^ n314 ;
  assign n319 = ~n275 & n318 ;
  assign n320 = n319 ^ x74 ;
  assign n321 = n320 ^ x92 ;
  assign n323 = n322 ^ n321 ;
  assign n324 = x91 ^ x75 ;
  assign n325 = n323 & ~n324 ;
  assign n326 = n325 ^ n322 ;
  assign n327 = ~n274 & n326 ;
  assign n328 = n327 ^ x76 ;
  assign n329 = n328 ^ x94 ;
  assign n331 = n330 ^ n329 ;
  assign n332 = x93 ^ x77 ;
  assign n333 = n331 & ~n332 ;
  assign n334 = n333 ^ n330 ;
  assign n335 = ~n272 & n334 ;
  assign n336 = n335 ^ x78 ;
  assign n337 = n336 ^ x95 ;
  assign n338 = ~n273 & n337 ;
  assign n339 = n338 ^ x79 ;
  assign n340 = n272 & ~n339 ;
  assign n341 = n340 ^ x78 ;
  assign n412 = n411 ^ n341 ;
  assign n413 = n261 ^ n260 ;
  assign n416 = n332 & ~n339 ;
  assign n417 = n416 ^ x77 ;
  assign n414 = n402 & ~n409 ;
  assign n415 = n414 ^ x109 ;
  assign n418 = n417 ^ n415 ;
  assign n421 = n274 & ~n339 ;
  assign n422 = n421 ^ x76 ;
  assign n419 = n344 & ~n409 ;
  assign n420 = n419 ^ x108 ;
  assign n423 = n422 ^ n420 ;
  assign n426 = n394 & ~n409 ;
  assign n427 = n426 ^ x107 ;
  assign n424 = n324 & ~n339 ;
  assign n425 = n424 ^ x75 ;
  assign n428 = n427 ^ n425 ;
  assign n431 = n275 & ~n339 ;
  assign n432 = n431 ^ x74 ;
  assign n429 = n345 & ~n409 ;
  assign n430 = n429 ^ x106 ;
  assign n433 = n432 ^ n430 ;
  assign n436 = n386 & ~n409 ;
  assign n437 = n436 ^ x105 ;
  assign n434 = n316 & ~n339 ;
  assign n435 = n434 ^ x73 ;
  assign n438 = n437 ^ n435 ;
  assign n441 = n276 & ~n339 ;
  assign n442 = n441 ^ x72 ;
  assign n439 = n346 & ~n409 ;
  assign n440 = n439 ^ x104 ;
  assign n443 = n442 ^ n440 ;
  assign n446 = n378 & ~n409 ;
  assign n447 = n446 ^ x103 ;
  assign n444 = n308 & ~n339 ;
  assign n445 = n444 ^ x71 ;
  assign n448 = n447 ^ n445 ;
  assign n451 = n277 & ~n339 ;
  assign n452 = n451 ^ x70 ;
  assign n449 = n347 & ~n409 ;
  assign n450 = n449 ^ x102 ;
  assign n453 = n452 ^ n450 ;
  assign n456 = n370 & ~n409 ;
  assign n457 = n456 ^ x101 ;
  assign n454 = n300 & ~n339 ;
  assign n455 = n454 ^ x69 ;
  assign n458 = n457 ^ n455 ;
  assign n461 = n278 & ~n339 ;
  assign n462 = n461 ^ x68 ;
  assign n459 = n348 & ~n409 ;
  assign n460 = n459 ^ x100 ;
  assign n463 = n462 ^ n460 ;
  assign n466 = n292 & ~n339 ;
  assign n467 = n466 ^ x67 ;
  assign n464 = n362 & ~n409 ;
  assign n465 = n464 ^ x99 ;
  assign n468 = n467 ^ n465 ;
  assign n471 = n349 & ~n409 ;
  assign n472 = n471 ^ x98 ;
  assign n469 = n279 & ~n339 ;
  assign n470 = n469 ^ x66 ;
  assign n473 = n472 ^ n470 ;
  assign n476 = n284 & ~n339 ;
  assign n477 = n476 ^ x65 ;
  assign n474 = n354 & ~n409 ;
  assign n475 = n474 ^ x97 ;
  assign n478 = n477 ^ n475 ;
  assign n479 = x112 ^ x96 ;
  assign n480 = ~n409 & n479 ;
  assign n481 = n480 ^ x96 ;
  assign n482 = x80 ^ x64 ;
  assign n483 = ~n339 & n482 ;
  assign n484 = n483 ^ x64 ;
  assign n485 = ~n481 & n484 ;
  assign n486 = n485 ^ n475 ;
  assign n487 = ~n478 & ~n486 ;
  assign n488 = n487 ^ n475 ;
  assign n489 = n488 ^ n470 ;
  assign n490 = ~n473 & ~n489 ;
  assign n491 = n490 ^ n470 ;
  assign n492 = n491 ^ n465 ;
  assign n493 = ~n468 & ~n492 ;
  assign n494 = n493 ^ n465 ;
  assign n495 = n494 ^ n462 ;
  assign n496 = ~n463 & ~n495 ;
  assign n497 = n496 ^ n462 ;
  assign n498 = n497 ^ n455 ;
  assign n499 = ~n458 & n498 ;
  assign n500 = n499 ^ n455 ;
  assign n501 = n500 ^ n452 ;
  assign n502 = ~n453 & n501 ;
  assign n503 = n502 ^ n452 ;
  assign n504 = n503 ^ n445 ;
  assign n505 = ~n448 & n504 ;
  assign n506 = n505 ^ n445 ;
  assign n507 = n506 ^ n442 ;
  assign n508 = ~n443 & n507 ;
  assign n509 = n508 ^ n442 ;
  assign n510 = n509 ^ n435 ;
  assign n511 = ~n438 & n510 ;
  assign n512 = n511 ^ n435 ;
  assign n513 = n512 ^ n432 ;
  assign n514 = ~n433 & n513 ;
  assign n515 = n514 ^ n432 ;
  assign n516 = n515 ^ n425 ;
  assign n517 = ~n428 & n516 ;
  assign n518 = n517 ^ n425 ;
  assign n519 = n518 ^ n420 ;
  assign n520 = ~n423 & ~n519 ;
  assign n521 = n520 ^ n420 ;
  assign n522 = n521 ^ n415 ;
  assign n523 = ~n418 & ~n522 ;
  assign n524 = n523 ^ n417 ;
  assign n525 = n524 ^ n341 ;
  assign n526 = ~n412 & ~n525 ;
  assign n527 = n526 ^ n411 ;
  assign n528 = n527 ^ n261 ;
  assign n529 = ~n413 & n528 ;
  assign n530 = n529 ^ n260 ;
  assign n531 = n412 & ~n530 ;
  assign n532 = n531 ^ n411 ;
  assign n794 = n793 ^ n532 ;
  assign n795 = n262 ^ n259 ;
  assign n798 = n679 & ~n791 ;
  assign n799 = n798 ^ n676 ;
  assign n796 = n418 & ~n530 ;
  assign n797 = n796 ^ n415 ;
  assign n800 = n799 ^ n797 ;
  assign n803 = n423 & ~n530 ;
  assign n804 = n803 ^ n420 ;
  assign n801 = n684 & ~n791 ;
  assign n802 = n801 ^ n681 ;
  assign n805 = n804 ^ n802 ;
  assign n808 = n689 & ~n791 ;
  assign n809 = n808 ^ n686 ;
  assign n806 = n428 & n530 ;
  assign n807 = n806 ^ n425 ;
  assign n810 = n809 ^ n807 ;
  assign n813 = n433 & n530 ;
  assign n814 = n813 ^ n432 ;
  assign n811 = n694 & ~n791 ;
  assign n812 = n811 ^ n693 ;
  assign n815 = n814 ^ n812 ;
  assign n818 = n699 & n791 ;
  assign n819 = n818 ^ n698 ;
  assign n816 = n438 & ~n530 ;
  assign n817 = n816 ^ n437 ;
  assign n820 = n819 ^ n817 ;
  assign n823 = n704 & ~n791 ;
  assign n824 = n823 ^ n701 ;
  assign n821 = n443 & ~n530 ;
  assign n822 = n821 ^ n440 ;
  assign n825 = n824 ^ n822 ;
  assign n828 = n448 & n530 ;
  assign n829 = n828 ^ n445 ;
  assign n826 = n709 & n791 ;
  assign n827 = n826 ^ n706 ;
  assign n830 = n829 ^ n827 ;
  assign n833 = n453 & n530 ;
  assign n834 = n833 ^ n452 ;
  assign n831 = n714 & ~n791 ;
  assign n832 = n831 ^ n713 ;
  assign n835 = n834 ^ n832 ;
  assign n838 = n719 & ~n791 ;
  assign n839 = n838 ^ n718 ;
  assign n836 = n458 & ~n530 ;
  assign n837 = n836 ^ n457 ;
  assign n840 = n839 ^ n837 ;
  assign n843 = n463 & ~n530 ;
  assign n844 = n843 ^ n460 ;
  assign n841 = n724 & n791 ;
  assign n842 = n841 ^ n721 ;
  assign n845 = n844 ^ n842 ;
  assign n848 = n468 & ~n530 ;
  assign n849 = n848 ^ n465 ;
  assign n846 = n729 & n791 ;
  assign n847 = n846 ^ n726 ;
  assign n850 = n849 ^ n847 ;
  assign n853 = n473 & ~n530 ;
  assign n854 = n853 ^ n472 ;
  assign n851 = n734 & ~n791 ;
  assign n852 = n851 ^ n733 ;
  assign n855 = n854 ^ n852 ;
  assign n858 = n739 & n791 ;
  assign n859 = n858 ^ n738 ;
  assign n856 = n478 & n530 ;
  assign n857 = n856 ^ n477 ;
  assign n860 = n859 ^ n857 ;
  assign n861 = n484 ^ n481 ;
  assign n862 = ~n530 & n861 ;
  assign n863 = n862 ^ n481 ;
  assign n864 = n745 ^ n742 ;
  assign n865 = n791 & n864 ;
  assign n866 = n865 ^ n742 ;
  assign n867 = ~n863 & n866 ;
  assign n868 = n867 ^ n857 ;
  assign n869 = ~n860 & ~n868 ;
  assign n870 = n869 ^ n857 ;
  assign n871 = n870 ^ n854 ;
  assign n872 = ~n855 & n871 ;
  assign n873 = n872 ^ n854 ;
  assign n874 = n873 ^ n847 ;
  assign n875 = ~n850 & ~n874 ;
  assign n876 = n875 ^ n847 ;
  assign n877 = n876 ^ n844 ;
  assign n878 = ~n845 & ~n877 ;
  assign n879 = n878 ^ n844 ;
  assign n880 = n879 ^ n837 ;
  assign n881 = ~n840 & n880 ;
  assign n882 = n881 ^ n837 ;
  assign n883 = n882 ^ n834 ;
  assign n884 = ~n835 & n883 ;
  assign n885 = n884 ^ n834 ;
  assign n886 = n885 ^ n827 ;
  assign n887 = ~n830 & ~n886 ;
  assign n888 = n887 ^ n827 ;
  assign n889 = n888 ^ n824 ;
  assign n890 = ~n825 & n889 ;
  assign n891 = n890 ^ n824 ;
  assign n892 = n891 ^ n817 ;
  assign n893 = ~n820 & ~n892 ;
  assign n894 = n893 ^ n817 ;
  assign n895 = n894 ^ n814 ;
  assign n896 = ~n815 & n895 ;
  assign n897 = n896 ^ n814 ;
  assign n898 = n897 ^ n807 ;
  assign n899 = ~n810 & n898 ;
  assign n900 = n899 ^ n807 ;
  assign n901 = n900 ^ n804 ;
  assign n902 = ~n805 & n901 ;
  assign n903 = n902 ^ n804 ;
  assign n904 = n903 ^ n799 ;
  assign n905 = ~n800 & ~n904 ;
  assign n906 = n905 ^ n799 ;
  assign n907 = n906 ^ n793 ;
  assign n908 = ~n794 & ~n907 ;
  assign n909 = n908 ^ n532 ;
  assign n910 = n909 ^ n262 ;
  assign n911 = ~n795 & n910 ;
  assign n912 = n911 ^ n259 ;
  assign n913 = n794 & n912 ;
  assign n914 = n913 ^ n793 ;
  assign n1558 = n1557 ^ n914 ;
  assign n1561 = n800 & n912 ;
  assign n1562 = n1561 ^ n799 ;
  assign n1559 = n1443 & n1555 ;
  assign n1560 = n1559 ^ n1442 ;
  assign n1563 = n1562 ^ n1560 ;
  assign n1566 = n1448 & n1555 ;
  assign n1567 = n1566 ^ n1445 ;
  assign n1564 = n805 & n912 ;
  assign n1565 = n1564 ^ n802 ;
  assign n1568 = n1567 ^ n1565 ;
  assign n1571 = n1453 & ~n1555 ;
  assign n1572 = n1571 ^ n1450 ;
  assign n1569 = n810 & ~n912 ;
  assign n1570 = n1569 ^ n807 ;
  assign n1573 = n1572 ^ n1570 ;
  assign n1576 = n815 & ~n912 ;
  assign n1577 = n1576 ^ n814 ;
  assign n1574 = n1458 & ~n1555 ;
  assign n1575 = n1574 ^ n1457 ;
  assign n1578 = n1577 ^ n1575 ;
  assign n1581 = n820 & n912 ;
  assign n1582 = n1581 ^ n819 ;
  assign n1579 = n1463 & n1555 ;
  assign n1580 = n1579 ^ n1462 ;
  assign n1583 = n1582 ^ n1580 ;
  assign n1586 = n1468 & ~n1555 ;
  assign n1587 = n1586 ^ n1465 ;
  assign n1584 = n825 & ~n912 ;
  assign n1585 = n1584 ^ n822 ;
  assign n1588 = n1587 ^ n1585 ;
  assign n1591 = n830 & n912 ;
  assign n1592 = n1591 ^ n827 ;
  assign n1589 = n1473 & n1555 ;
  assign n1590 = n1589 ^ n1470 ;
  assign n1593 = n1592 ^ n1590 ;
  assign n1596 = n1478 & ~n1555 ;
  assign n1597 = n1596 ^ n1477 ;
  assign n1594 = n835 & ~n912 ;
  assign n1595 = n1594 ^ n834 ;
  assign n1598 = n1597 ^ n1595 ;
  assign n1601 = n840 & n912 ;
  assign n1602 = n1601 ^ n839 ;
  assign n1599 = n1483 & n1555 ;
  assign n1600 = n1599 ^ n1482 ;
  assign n1603 = n1602 ^ n1600 ;
  assign n1606 = n1488 & ~n1555 ;
  assign n1607 = n1606 ^ n1485 ;
  assign n1604 = n845 & n912 ;
  assign n1605 = n1604 ^ n842 ;
  assign n1608 = n1607 ^ n1605 ;
  assign n1612 = n1493 & ~n1555 ;
  assign n1613 = n1612 ^ n1490 ;
  assign n1609 = n850 & n912 ;
  assign n1610 = n1609 ^ n847 ;
  assign n1614 = n1613 ^ n1610 ;
  assign n1617 = n1498 & ~n1555 ;
  assign n1618 = n1617 ^ n1497 ;
  assign n1615 = n855 & ~n912 ;
  assign n1616 = n1615 ^ n854 ;
  assign n1619 = n1618 ^ n1616 ;
  assign n1622 = n860 & n912 ;
  assign n1623 = n1622 ^ n859 ;
  assign n1620 = n1503 & n1555 ;
  assign n1621 = n1620 ^ n1502 ;
  assign n1624 = n1623 ^ n1621 ;
  assign n1625 = n1509 ^ n1506 ;
  assign n1626 = ~n1555 & n1625 ;
  assign n1627 = n1626 ^ n1506 ;
  assign n1628 = n866 ^ n863 ;
  assign n1629 = ~n912 & n1628 ;
  assign n1630 = n1629 ^ n863 ;
  assign n1631 = ~n1627 & n1630 ;
  assign n1632 = n1631 ^ n1621 ;
  assign n1633 = ~n1624 & ~n1632 ;
  assign n1634 = n1633 ^ n1621 ;
  assign n1635 = n1634 ^ n1616 ;
  assign n1636 = ~n1619 & ~n1635 ;
  assign n1637 = n1636 ^ n1616 ;
  assign n1638 = n1637 ^ n1613 ;
  assign n1639 = ~n1614 & n1638 ;
  assign n1611 = n1610 ^ n1605 ;
  assign n1640 = n1639 ^ n1611 ;
  assign n1641 = ~n1608 & ~n1640 ;
  assign n1642 = n1641 ^ n1607 ;
  assign n1643 = n1642 ^ n1600 ;
  assign n1644 = ~n1603 & ~n1643 ;
  assign n1645 = n1644 ^ n1602 ;
  assign n1646 = n1645 ^ n1595 ;
  assign n1647 = ~n1598 & ~n1646 ;
  assign n1648 = n1647 ^ n1597 ;
  assign n1649 = n1648 ^ n1590 ;
  assign n1650 = ~n1593 & ~n1649 ;
  assign n1651 = n1650 ^ n1592 ;
  assign n1652 = n1651 ^ n1585 ;
  assign n1653 = ~n1588 & n1652 ;
  assign n1654 = n1653 ^ n1585 ;
  assign n1655 = n1654 ^ n1582 ;
  assign n1656 = ~n1583 & n1655 ;
  assign n1657 = n1656 ^ n1582 ;
  assign n1658 = n1657 ^ n1575 ;
  assign n1659 = ~n1578 & ~n1658 ;
  assign n1660 = n1659 ^ n1575 ;
  assign n1661 = n1660 ^ n1572 ;
  assign n1662 = ~n1573 & n1661 ;
  assign n1663 = n1662 ^ n1572 ;
  assign n1664 = n1663 ^ n1565 ;
  assign n1665 = ~n1568 & ~n1664 ;
  assign n1666 = n1665 ^ n1565 ;
  assign n1667 = n1666 ^ n1560 ;
  assign n1668 = ~n1563 & ~n1667 ;
  assign n1669 = n1668 ^ n1560 ;
  assign n1670 = n1669 ^ n914 ;
  assign n1671 = ~n1558 & n1670 ;
  assign n1672 = n1671 ^ n1557 ;
  assign n1673 = n1672 ^ n263 ;
  assign n1674 = ~n271 & ~n1673 ;
  assign n1675 = n1674 ^ n270 ;
  assign n1676 = n1555 ^ n912 ;
  assign n1677 = ~n1675 & n1676 ;
  assign n1678 = n1677 ^ n912 ;
  assign n1682 = n1434 & ~n1678 ;
  assign n1683 = n1173 & n1555 ;
  assign n1684 = ~n1682 & ~n1683 ;
  assign n1679 = n791 & ~n1678 ;
  assign n1680 = n530 & n912 ;
  assign n1681 = ~n1679 & ~n1680 ;
  assign n1685 = n1684 ^ n1681 ;
  assign n1686 = n1675 & n1685 ;
  assign n1687 = n1686 ^ n1684 ;
  assign n1700 = n1052 ^ n982 ;
  assign n1701 = n1687 & n1700 ;
  assign n1702 = n1701 ^ n1052 ;
  assign n1697 = n1313 ^ n1243 ;
  assign n1698 = ~n1687 & n1697 ;
  assign n1699 = n1698 ^ n1313 ;
  assign n1703 = n1702 ^ n1699 ;
  assign n1704 = n1678 & n1703 ;
  assign n1705 = n1704 ^ n1699 ;
  assign n1691 = n409 ^ n339 ;
  assign n1692 = n1687 & n1691 ;
  assign n1693 = n1692 ^ n409 ;
  assign n1688 = n670 ^ n600 ;
  assign n1689 = n1687 & n1688 ;
  assign n1690 = n1689 ^ n600 ;
  assign n1694 = n1693 ^ n1690 ;
  assign n1695 = n1678 & n1694 ;
  assign n1696 = n1695 ^ n1690 ;
  assign n1706 = n1705 ^ n1696 ;
  assign n1707 = n1675 & n1706 ;
  assign n1708 = n1707 ^ n1705 ;
  assign n1709 = n1630 ^ n1627 ;
  assign n1710 = n1675 & n1709 ;
  assign n1711 = n1710 ^ n1627 ;
  assign n1712 = n1624 & ~n1675 ;
  assign n1713 = n1712 ^ n1623 ;
  assign n1714 = n1619 & n1675 ;
  assign n1715 = n1714 ^ n1618 ;
  assign n1716 = n1614 & n1675 ;
  assign n1717 = n1716 ^ n1613 ;
  assign n1718 = n1608 & n1675 ;
  assign n1719 = n1718 ^ n1607 ;
  assign n1720 = n1603 & ~n1675 ;
  assign n1721 = n1720 ^ n1602 ;
  assign n1722 = n1598 & n1675 ;
  assign n1723 = n1722 ^ n1597 ;
  assign n1724 = n1593 & ~n1675 ;
  assign n1725 = n1724 ^ n1592 ;
  assign n1726 = n1588 & n1675 ;
  assign n1727 = n1726 ^ n1587 ;
  assign n1728 = n1583 & ~n1675 ;
  assign n1729 = n1728 ^ n1582 ;
  assign n1730 = n1578 & n1675 ;
  assign n1731 = n1730 ^ n1575 ;
  assign n1732 = n1573 & ~n1675 ;
  assign n1733 = n1732 ^ n1570 ;
  assign n1734 = n1568 & n1675 ;
  assign n1735 = n1734 ^ n1567 ;
  assign n1736 = n1563 & ~n1675 ;
  assign n1737 = n1736 ^ n1562 ;
  assign n1738 = n1558 & n1675 ;
  assign n1739 = n1738 ^ n1557 ;
  assign n1740 = n263 & n270 ;
  assign y0 = ~n1708 ;
  assign y1 = ~n1687 ;
  assign y2 = n1678 ;
  assign y3 = ~n1675 ;
  assign y4 = n1711 ;
  assign y5 = n1713 ;
  assign y6 = n1715 ;
  assign y7 = n1717 ;
  assign y8 = n1719 ;
  assign y9 = n1721 ;
  assign y10 = n1723 ;
  assign y11 = n1725 ;
  assign y12 = n1727 ;
  assign y13 = n1729 ;
  assign y14 = n1731 ;
  assign y15 = n1733 ;
  assign y16 = n1735 ;
  assign y17 = n1737 ;
  assign y18 = n1739 ;
  assign y19 = ~n1740 ;
endmodule
