module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10;
  wire n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671;
  assign n31 = x2 & x3;
  assign n32 = n31 ^ x2;
  assign n33 = n32 ^ x3;
  assign n57 = ~x7 & ~x9;
  assign n58 = ~n33 & ~n57;
  assign n13 = x8 & ~x9;
  assign n12 = x9 ^ x8;
  assign n14 = n13 ^ n12;
  assign n59 = n14 ^ x0;
  assign n60 = n58 & n59;
  assign n62 = x8 ^ x7;
  assign n61 = x7 & ~x8;
  assign n63 = n62 ^ n61;
  assign n64 = n63 ^ x7;
  assign n65 = ~n60 & n64;
  assign n11 = ~x0 & x7;
  assign n19 = ~x2 & x8;
  assign n20 = n19 ^ x2;
  assign n15 = n14 ^ x8;
  assign n16 = n15 ^ n12;
  assign n17 = ~x2 & ~n16;
  assign n18 = n17 ^ n15;
  assign n21 = n20 ^ n18;
  assign n22 = n21 ^ x9;
  assign n23 = n22 ^ n20;
  assign n24 = n11 & n23;
  assign n26 = ~x0 & ~x9;
  assign n25 = x9 ^ x0;
  assign n27 = n26 ^ n25;
  assign n28 = n19 & ~n27;
  assign n29 = ~n24 & ~n28;
  assign n30 = ~x3 & ~n29;
  assign n36 = n16 & ~n32;
  assign n37 = n36 ^ n16;
  assign n34 = n33 ^ x2;
  assign n35 = ~n15 & n34;
  assign n38 = n37 ^ n35;
  assign n39 = ~x0 & n38;
  assign n40 = x3 ^ x2;
  assign n41 = n40 ^ x0;
  assign n42 = ~x3 & x9;
  assign n43 = n42 ^ x3;
  assign n44 = n43 ^ n13;
  assign n45 = n44 ^ x3;
  assign n46 = n45 ^ n40;
  assign n47 = ~n41 & ~n46;
  assign n48 = n47 ^ n44;
  assign n49 = n48 ^ x3;
  assign n50 = n49 ^ x0;
  assign n51 = ~n40 & n50;
  assign n52 = n51 ^ n40;
  assign n53 = ~n39 & n52;
  assign n54 = ~x7 & ~n53;
  assign n55 = ~n30 & ~n54;
  assign n56 = ~x1 & ~n55;
  assign n66 = n65 ^ n56;
  assign n67 = x5 & x6;
  assign n68 = n67 ^ x6;
  assign n69 = n68 ^ x5;
  assign n70 = ~n66 & ~n69;
  assign n71 = ~x1 & x8;
  assign n72 = n71 ^ x1;
  assign n73 = ~x3 & n72;
  assign n77 = x0 & ~x8;
  assign n74 = x0 & ~x1;
  assign n75 = n19 ^ x8;
  assign n76 = n74 & n75;
  assign n78 = n77 ^ n76;
  assign n79 = ~n73 & n78;
  assign n80 = x8 ^ x3;
  assign n81 = x3 ^ x1;
  assign n82 = n80 & ~n81;
  assign n83 = n82 ^ n80;
  assign n84 = n40 & n83;
  assign n85 = n84 ^ n82;
  assign n86 = n85 ^ x8;
  assign n87 = n86 ^ n80;
  assign n88 = ~x0 & ~n87;
  assign n90 = x9 ^ x5;
  assign n89 = x5 & x9;
  assign n91 = n90 ^ n89;
  assign n92 = ~n88 & ~n91;
  assign n93 = ~n79 & n92;
  assign n94 = x1 & ~x2;
  assign n95 = n94 ^ x2;
  assign n96 = n95 ^ x8;
  assign n97 = ~x5 & n96;
  assign n98 = n97 ^ x8;
  assign n99 = n33 & n98;
  assign n103 = n72 ^ x8;
  assign n100 = x8 ^ x0;
  assign n101 = n100 ^ n77;
  assign n102 = x1 & ~n101;
  assign n104 = n103 ^ n102;
  assign n105 = ~n99 & ~n104;
  assign n106 = x5 & x8;
  assign n107 = n106 ^ x8;
  assign n108 = ~n105 & ~n107;
  assign n109 = n27 & ~n89;
  assign n110 = ~n36 & n109;
  assign n111 = n34 ^ x8;
  assign n112 = ~x5 & n111;
  assign n113 = n112 ^ x8;
  assign n114 = n74 ^ x1;
  assign n115 = n113 & ~n114;
  assign n116 = ~n110 & ~n115;
  assign n117 = ~n108 & n116;
  assign n118 = ~n33 & ~n114;
  assign n120 = ~x5 & ~n16;
  assign n121 = n120 ^ n107;
  assign n119 = n89 ^ n13;
  assign n122 = n121 ^ n119;
  assign n123 = ~n118 & ~n122;
  assign n124 = x6 & ~x7;
  assign n125 = ~n123 & n124;
  assign n126 = ~n117 & n125;
  assign n127 = ~n93 & n126;
  assign n128 = ~x3 & ~n75;
  assign n129 = x1 & ~x9;
  assign n130 = n129 ^ x1;
  assign n131 = n130 ^ x9;
  assign n132 = n131 ^ x2;
  assign n133 = n74 & n132;
  assign n134 = n128 & ~n133;
  assign n139 = x2 & n15;
  assign n140 = n139 ^ n75;
  assign n136 = x2 ^ x0;
  assign n135 = ~x0 & x2;
  assign n137 = n136 ^ n135;
  assign n138 = ~x9 & n137;
  assign n141 = n140 ^ n138;
  assign n142 = x1 & n141;
  assign n143 = x3 & ~n19;
  assign n144 = ~n142 & n143;
  assign n145 = ~n134 & ~n144;
  assign n149 = ~x1 & n15;
  assign n150 = n149 ^ n72;
  assign n151 = n150 ^ x1;
  assign n152 = n151 ^ n16;
  assign n147 = n130 ^ n102;
  assign n146 = x9 ^ x1;
  assign n148 = n147 ^ n146;
  assign n153 = n152 ^ n148;
  assign n154 = n153 ^ x8;
  assign n156 = n124 ^ x7;
  assign n155 = ~x7 & ~n69;
  assign n157 = n156 ^ n155;
  assign n158 = ~n154 & ~n157;
  assign n159 = ~n145 & n158;
  assign n160 = ~n127 & ~n159;
  assign n161 = ~n70 & n160;
  assign n163 = n118 ^ x4;
  assign n162 = x6 ^ x5;
  assign n164 = n163 ^ n162;
  assign n165 = n162 ^ n15;
  assign n166 = n162 & ~n165;
  assign n167 = n166 ^ n162;
  assign n168 = ~n164 & n167;
  assign n169 = n168 ^ n166;
  assign n170 = n169 ^ n162;
  assign n171 = n170 ^ n15;
  assign n172 = n118 & ~n171;
  assign n173 = n172 ^ n163;
  assign n174 = ~n161 & ~n173;
  assign n178 = n94 & n101;
  assign n179 = n63 ^ n20;
  assign n180 = n74 & ~n179;
  assign n181 = ~n178 & ~n180;
  assign n182 = ~n43 & ~n181;
  assign n183 = n16 ^ x7;
  assign n184 = ~x3 & ~n95;
  assign n185 = n184 ^ x3;
  assign n186 = n183 & ~n185;
  assign n187 = n137 ^ n114;
  assign n188 = n186 & ~n187;
  assign n189 = ~n182 & ~n188;
  assign n175 = ~n20 & ~n114;
  assign n176 = n57 & ~n175;
  assign n177 = ~n76 & n176;
  assign n190 = n189 ^ n177;
  assign n191 = ~n69 & ~n190;
  assign n192 = ~x1 & ~x5;
  assign n193 = ~x0 & x3;
  assign n194 = n193 ^ x9;
  assign n195 = n194 ^ n42;
  assign n196 = n195 ^ x0;
  assign n197 = n12 & n196;
  assign n198 = n197 ^ x3;
  assign n199 = n192 & ~n198;
  assign n200 = n121 ^ n90;
  assign n201 = x1 & n81;
  assign n202 = n201 ^ n130;
  assign n203 = ~n200 & n202;
  assign n204 = x2 & ~n89;
  assign n205 = ~n203 & n204;
  assign n206 = ~n199 & n205;
  assign n207 = n74 ^ x0;
  assign n208 = ~n33 & n207;
  assign n209 = ~x2 & n91;
  assign n210 = ~n208 & ~n209;
  assign n211 = n89 & n102;
  assign n212 = ~n210 & ~n211;
  assign n213 = ~x3 & n114;
  assign n214 = n14 & n207;
  assign n215 = n213 & ~n214;
  assign n216 = n14 & n74;
  assign n217 = x3 & ~n89;
  assign n218 = ~n216 & n217;
  assign n219 = ~n215 & ~n218;
  assign n220 = n212 & ~n219;
  assign n221 = n124 & ~n220;
  assign n222 = ~n206 & n221;
  assign n223 = ~x3 & n76;
  assign n225 = ~x9 & ~n32;
  assign n224 = n32 ^ x9;
  assign n226 = n225 ^ n224;
  assign n227 = n226 ^ n140;
  assign n228 = n227 ^ n37;
  assign n229 = n228 ^ n43;
  assign n230 = x1 & n229;
  assign n231 = ~n223 & ~n230;
  assign n232 = n42 ^ n32;
  assign n233 = n232 ^ n225;
  assign n234 = ~n152 & n233;
  assign n235 = ~x0 & n234;
  assign n236 = x1 & ~n19;
  assign n237 = n225 & ~n236;
  assign n238 = ~n235 & ~n237;
  assign n239 = n231 & n238;
  assign n240 = ~n157 & ~n239;
  assign n241 = ~n222 & ~n240;
  assign n242 = ~n191 & n241;
  assign n246 = n15 & n118;
  assign n243 = ~x0 & ~x6;
  assign n244 = ~x9 & ~n243;
  assign n245 = n184 & ~n244;
  assign n247 = n246 ^ n245;
  assign n248 = ~x4 & ~n247;
  assign n249 = n248 ^ n245;
  assign n250 = ~n242 & n249;
  assign n253 = ~x6 & x8;
  assign n281 = ~x1 & ~n253;
  assign n282 = n138 & n281;
  assign n277 = n26 ^ n13;
  assign n275 = ~x9 & ~n101;
  assign n276 = n275 ^ x0;
  assign n278 = n277 ^ n276;
  assign n279 = n94 & n278;
  assign n274 = n16 & n135;
  assign n280 = n279 ^ n274;
  assign n283 = n282 ^ n280;
  assign n292 = x8 ^ x6;
  assign n293 = n292 ^ n253;
  assign n288 = ~x8 & ~n243;
  assign n289 = n288 ^ x0;
  assign n251 = ~x2 & x6;
  assign n252 = n251 ^ x2;
  assign n290 = n288 ^ n252;
  assign n291 = ~n289 & ~n290;
  assign n294 = n293 ^ n291;
  assign n295 = n129 & n294;
  assign n284 = ~x6 & n16;
  assign n285 = n284 ^ x6;
  assign n286 = ~n21 & n285;
  assign n287 = ~n114 & n286;
  assign n296 = n295 ^ n287;
  assign n297 = ~n283 & ~n296;
  assign n298 = ~x5 & ~x7;
  assign n299 = x0 & n129;
  assign n300 = ~n14 & ~n69;
  assign n301 = ~n299 & n300;
  assign n302 = ~n298 & ~n301;
  assign n303 = ~x3 & ~n11;
  assign n304 = n43 & ~n303;
  assign n264 = x6 ^ x1;
  assign n263 = ~x1 & ~x6;
  assign n265 = n264 ^ n263;
  assign n266 = n265 ^ x1;
  assign n305 = ~x0 & n57;
  assign n306 = ~n266 & n305;
  assign n307 = ~n304 & ~n306;
  assign n308 = ~n302 & n307;
  assign n309 = ~n297 & n308;
  assign n254 = n253 ^ n252;
  assign n255 = n254 ^ n20;
  assign n256 = n255 ^ x2;
  assign n257 = n130 & ~n256;
  assign n258 = ~x0 & ~n257;
  assign n260 = n135 ^ n19;
  assign n259 = ~x2 & ~n101;
  assign n261 = n260 ^ n259;
  assign n262 = n42 & n261;
  assign n267 = ~n13 & ~n266;
  assign n268 = n252 ^ x6;
  assign n269 = ~x3 & ~n268;
  assign n270 = ~n267 & n269;
  assign n271 = ~n262 & ~n270;
  assign n272 = ~n258 & ~n271;
  assign n273 = ~x7 & ~n272;
  assign n310 = n309 ^ n273;
  assign n343 = ~x2 & ~n114;
  assign n344 = ~x8 & n68;
  assign n345 = n343 & ~n344;
  assign n346 = n345 ^ x4;
  assign n311 = ~x6 & x9;
  assign n312 = n311 ^ n68;
  assign n313 = n71 & n312;
  assign n314 = n22 & n107;
  assign n315 = ~n101 & ~n314;
  assign n316 = ~n313 & n315;
  assign n317 = x2 & ~x5;
  assign n318 = n317 ^ n252;
  assign n319 = ~x1 & n318;
  assign n320 = n129 & n317;
  assign n321 = ~x0 & ~n67;
  assign n322 = ~n209 & n321;
  assign n323 = ~n320 & n322;
  assign n324 = ~n319 & n323;
  assign n325 = ~n316 & ~n324;
  assign n326 = n265 ^ x0;
  assign n327 = n317 ^ x9;
  assign n328 = ~n265 & n327;
  assign n329 = n328 ^ x9;
  assign n330 = ~n326 & n329;
  assign n331 = n318 ^ x8;
  assign n332 = x5 & n129;
  assign n333 = n332 ^ x9;
  assign n334 = ~x0 & n333;
  assign n335 = n334 ^ n332;
  assign n336 = n331 & ~n335;
  assign n337 = n336 ^ n334;
  assign n338 = n337 ^ n332;
  assign n339 = n338 ^ x0;
  assign n340 = ~x8 & n339;
  assign n341 = ~n330 & n340;
  assign n342 = ~n325 & ~n341;
  assign n347 = n346 ^ n342;
  assign n348 = n347 ^ n346;
  assign n349 = ~x4 & ~n348;
  assign n350 = n349 ^ n346;
  assign n351 = x3 & ~n350;
  assign n352 = n351 ^ n346;
  assign n353 = n310 & ~n352;
  assign n354 = ~n67 & ~n132;
  assign n355 = x3 & ~n354;
  assign n366 = x0 & n121;
  assign n364 = n67 ^ x5;
  assign n365 = n74 & ~n364;
  assign n367 = n366 ^ n365;
  assign n368 = ~n311 & n367;
  assign n356 = x0 & x5;
  assign n360 = n284 & ~n356;
  assign n361 = x1 & n360;
  assign n362 = n361 ^ n284;
  assign n357 = n356 ^ x5;
  assign n358 = x1 & n357;
  assign n359 = ~n253 & n358;
  assign n363 = n362 ^ n359;
  assign n369 = n368 ^ n363;
  assign n370 = n355 & n369;
  assign n371 = x1 & ~n18;
  assign n372 = ~n15 & ~n95;
  assign n373 = n372 ^ x1;
  assign n374 = ~x6 & n373;
  assign n375 = n374 ^ x1;
  assign n376 = ~n371 & ~n375;
  assign n377 = n356 & ~n376;
  assign n381 = x1 & ~n276;
  assign n382 = n381 ^ x0;
  assign n383 = n382 ^ n147;
  assign n378 = n101 ^ x9;
  assign n379 = n378 ^ n275;
  assign n380 = n379 ^ n114;
  assign n384 = n383 ^ n380;
  assign n385 = ~x6 & n384;
  assign n386 = ~n268 & ~n385;
  assign n387 = n101 ^ x1;
  assign n388 = n146 ^ n68;
  assign n389 = ~n387 & ~n388;
  assign n390 = n389 ^ n101;
  assign n391 = n68 & n390;
  assign n392 = n391 ^ x5;
  assign n393 = n386 & ~n392;
  assign n394 = n75 & n130;
  assign n395 = ~x6 & ~n394;
  assign n400 = n251 ^ n68;
  assign n397 = x5 ^ x2;
  assign n398 = n397 ^ x6;
  assign n399 = n67 & ~n398;
  assign n401 = n400 ^ n399;
  assign n396 = n265 & n357;
  assign n402 = n401 ^ n396;
  assign n403 = ~n395 & n402;
  assign n404 = ~n101 & n320;
  assign n405 = ~x3 & ~n404;
  assign n406 = ~n403 & n405;
  assign n407 = ~n393 & n406;
  assign n408 = ~n377 & n407;
  assign n409 = ~n162 & n184;
  assign n410 = n409 ^ x4;
  assign n411 = ~x7 & ~n410;
  assign n412 = ~n408 & n411;
  assign n413 = ~n370 & n412;
  assign n414 = n114 ^ x2;
  assign n415 = ~n163 & ~n414;
  assign n416 = n298 ^ x7;
  assign n417 = n416 ^ n157;
  assign n418 = n415 & n417;
  assign n419 = x4 ^ x3;
  assign n420 = n343 ^ x4;
  assign n421 = n419 & ~n420;
  assign n422 = n417 & n421;
  assign n423 = ~x3 & ~x4;
  assign n468 = n106 ^ x5;
  assign n477 = ~n207 & n468;
  assign n478 = ~n94 & n477;
  assign n479 = ~n138 & n478;
  assign n480 = n131 & n135;
  assign n481 = n106 & ~n129;
  assign n482 = ~n480 & n481;
  assign n483 = ~x4 & ~n482;
  assign n484 = ~n479 & n483;
  assign n485 = n484 ^ x5;
  assign n486 = ~n75 & ~n311;
  assign n487 = x0 & ~n486;
  assign n488 = n101 ^ n26;
  assign n489 = n251 & n488;
  assign n490 = n489 ^ n26;
  assign n491 = ~n150 & ~n490;
  assign n492 = ~n487 & n491;
  assign n493 = ~n256 & ~n379;
  assign n494 = n244 & n259;
  assign n495 = x1 & ~n494;
  assign n496 = ~n493 & n495;
  assign n497 = ~n492 & ~n496;
  assign n498 = n497 ^ x6;
  assign n499 = n484 & n498;
  assign n500 = n499 ^ x6;
  assign n501 = n485 & ~n500;
  assign n502 = n501 ^ x5;
  assign n503 = x4 & ~n118;
  assign n504 = n503 ^ x4;
  assign n505 = ~n502 & ~n504;
  assign n452 = ~n91 & n265;
  assign n453 = n63 & ~n452;
  assign n454 = x2 & ~n453;
  assign n456 = n266 ^ x5;
  assign n455 = x1 & ~n69;
  assign n457 = n456 ^ n455;
  assign n458 = ~n130 & n457;
  assign n459 = ~x7 & ~n458;
  assign n460 = ~n63 & n263;
  assign n461 = n120 & n460;
  assign n462 = ~n459 & ~n461;
  assign n463 = n454 & n462;
  assign n464 = ~n64 & ~n265;
  assign n465 = ~x2 & ~n417;
  assign n466 = ~n464 & n465;
  assign n467 = n455 ^ x9;
  assign n469 = n468 ^ n61;
  assign n470 = n469 ^ n344;
  assign n471 = ~n467 & n470;
  assign n472 = n471 ^ n455;
  assign n473 = ~x9 & n472;
  assign n474 = n466 & ~n473;
  assign n475 = ~n463 & ~n474;
  assign n424 = ~x2 & n298;
  assign n425 = n15 & n424;
  assign n426 = x6 & ~n425;
  assign n427 = x0 & ~n426;
  assign n428 = x7 ^ x5;
  assign n429 = n311 ^ x2;
  assign n430 = n311 & ~n429;
  assign n431 = n430 ^ n394;
  assign n432 = n431 ^ n311;
  assign n433 = n428 & ~n432;
  assign n434 = n433 ^ n430;
  assign n435 = n434 ^ n311;
  assign n436 = ~x7 & n435;
  assign n437 = n436 ^ x5;
  assign n438 = n427 & ~n437;
  assign n439 = ~x7 & n15;
  assign n440 = x2 & ~n439;
  assign n441 = n57 & n107;
  assign n442 = x1 & ~n61;
  assign n443 = ~n441 & n442;
  assign n444 = ~n440 & n443;
  assign n445 = ~x2 & ~n57;
  assign n446 = n122 & ~n445;
  assign n447 = x7 & n16;
  assign n448 = ~x1 & ~n447;
  assign n449 = n446 & n448;
  assign n450 = ~n444 & ~n449;
  assign n451 = n438 & ~n450;
  assign n476 = n475 ^ n451;
  assign n506 = n505 ^ n476;
  assign n507 = n506 ^ n476;
  assign n508 = ~x7 & ~n507;
  assign n509 = n508 ^ n476;
  assign n510 = ~n423 & n509;
  assign n511 = n510 ^ n476;
  assign n512 = n201 ^ n71;
  assign n513 = n152 & ~n512;
  assign n514 = ~x3 & ~n153;
  assign n515 = n383 & ~n514;
  assign n516 = ~n513 & n515;
  assign n517 = ~x2 & ~n516;
  assign n521 = ~n42 & n77;
  assign n522 = n521 ^ n22;
  assign n519 = n34 & n77;
  assign n518 = n128 ^ x3;
  assign n520 = n519 ^ n518;
  assign n523 = n522 ^ n520;
  assign n524 = x1 & n523;
  assign n525 = n12 & n263;
  assign n526 = ~x0 & ~n33;
  assign n527 = n526 ^ x3;
  assign n528 = n525 & ~n527;
  assign n529 = n364 & ~n528;
  assign n530 = ~n524 & n529;
  assign n531 = ~n517 & n530;
  assign n549 = n193 ^ n137;
  assign n550 = n549 ^ n34;
  assign n546 = x9 ^ x3;
  assign n551 = n550 ^ n546;
  assign n547 = n546 ^ x1;
  assign n548 = n547 ^ n136;
  assign n552 = n551 ^ n548;
  assign n553 = n552 ^ n136;
  assign n554 = n553 ^ x3;
  assign n555 = n146 & n552;
  assign n556 = n555 ^ n546;
  assign n557 = n556 ^ n548;
  assign n558 = n557 ^ n136;
  assign n559 = n558 ^ x3;
  assign n560 = n554 & n559;
  assign n561 = n560 ^ n201;
  assign n562 = n561 ^ n550;
  assign n563 = n562 ^ n546;
  assign n564 = n563 ^ n548;
  assign n565 = n564 ^ n136;
  assign n566 = n565 ^ x3;
  assign n567 = x8 & n566;
  assign n568 = n80 ^ n40;
  assign n569 = n26 ^ x3;
  assign n570 = n569 ^ n80;
  assign n571 = n80 & ~n570;
  assign n572 = n571 ^ n80;
  assign n573 = n568 & n572;
  assign n574 = n573 ^ n571;
  assign n575 = n574 ^ x3;
  assign n576 = n575 ^ n80;
  assign n577 = n576 ^ n226;
  assign n578 = x1 & n577;
  assign n579 = n578 ^ n576;
  assign n580 = ~n567 & n579;
  assign n532 = ~n131 & n278;
  assign n536 = n13 ^ x1;
  assign n534 = n131 ^ n72;
  assign n535 = n534 ^ x8;
  assign n537 = n536 ^ n535;
  assign n533 = ~n15 & n213;
  assign n538 = n537 ^ n533;
  assign n539 = ~n532 & n538;
  assign n540 = ~x2 & ~n539;
  assign n541 = ~n12 & n193;
  assign n542 = ~n139 & ~n541;
  assign n543 = ~x1 & ~n542;
  assign n544 = ~n37 & ~n543;
  assign n545 = ~n540 & n544;
  assign n581 = n580 ^ n545;
  assign n582 = n581 ^ n545;
  assign n583 = ~x6 & ~n582;
  assign n584 = n583 ^ n545;
  assign n585 = ~x4 & ~n584;
  assign n586 = n585 ^ x6;
  assign n587 = ~x5 & ~n586;
  assign n588 = ~n531 & ~n587;
  assign n589 = x7 & ~n528;
  assign n590 = x0 & n263;
  assign n591 = n19 & n57;
  assign n592 = n591 ^ n61;
  assign n593 = n590 & n592;
  assign n594 = ~n589 & ~n593;
  assign n595 = ~n503 & n594;
  assign n596 = ~n588 & n595;
  assign n597 = n298 & n504;
  assign n599 = n275 ^ n130;
  assign n598 = ~n149 & n383;
  assign n600 = n599 ^ n598;
  assign n601 = n600 ^ x1;
  assign n602 = n332 ^ n27;
  assign n603 = n601 & n602;
  assign n604 = ~x2 & ~n603;
  assign n605 = ~x1 & ~n21;
  assign n606 = ~n120 & n605;
  assign n607 = n405 & ~n606;
  assign n608 = ~n604 & n607;
  assign n609 = ~n16 & ~n69;
  assign n610 = n609 ^ n69;
  assign n611 = n610 ^ n285;
  assign n612 = n608 & n611;
  assign n613 = ~n263 & ~n343;
  assign n614 = ~x9 & ~n288;
  assign n615 = ~n613 & n614;
  assign n616 = x6 ^ x2;
  assign n617 = x9 & n616;
  assign n618 = ~n102 & n617;
  assign n619 = ~n71 & ~n252;
  assign n620 = x3 & ~x5;
  assign n621 = ~n619 & n620;
  assign n622 = ~n618 & n621;
  assign n623 = ~n615 & n622;
  assign n624 = n34 & n364;
  assign n625 = n379 ^ n149;
  assign n626 = n625 ^ n598;
  assign n627 = n626 ^ n537;
  assign n628 = n624 & n627;
  assign n629 = ~n623 & ~n628;
  assign n630 = ~n612 & n629;
  assign n632 = ~x2 & ~n129;
  assign n631 = ~n114 & n139;
  assign n633 = n632 ^ n631;
  assign n634 = n609 & n633;
  assign n635 = x7 & ~n634;
  assign n636 = ~x4 & ~n635;
  assign n637 = ~n630 & n636;
  assign n638 = ~n597 & ~n637;
  assign n639 = n184 ^ x4;
  assign n640 = n399 ^ n398;
  assign n642 = ~n385 & n392;
  assign n641 = ~n69 & n598;
  assign n643 = n642 ^ n641;
  assign n644 = n640 & n643;
  assign n645 = x3 & ~x7;
  assign n646 = ~n644 & n645;
  assign n647 = n268 & ~n537;
  assign n648 = n69 & n95;
  assign n649 = ~n647 & n648;
  assign n650 = x7 ^ x2;
  assign n651 = n382 ^ x7;
  assign n652 = n650 & ~n651;
  assign n653 = n652 ^ n381;
  assign n654 = n653 ^ x0;
  assign n655 = n654 ^ x2;
  assign n656 = ~x7 & ~n655;
  assign n657 = n656 ^ x7;
  assign n658 = n657 ^ x7;
  assign n659 = ~n631 & ~n658;
  assign n660 = ~x3 & ~n131;
  assign n661 = ~n128 & ~n660;
  assign n662 = n661 ^ n409;
  assign n663 = ~n659 & ~n662;
  assign n664 = ~n649 & n663;
  assign n665 = ~n646 & ~n664;
  assign n666 = ~n639 & ~n665;
  assign n667 = n31 & n598;
  assign n668 = n667 ^ n118;
  assign n669 = ~x4 & n668;
  assign n670 = n669 ^ n118;
  assign n671 = n155 & n670;
  assign y0 = n174;
  assign y1 = n250;
  assign y2 = n353;
  assign y3 = n413;
  assign y4 = n418;
  assign y5 = n422;
  assign y6 = ~n511;
  assign y7 = ~n596;
  assign y8 = n638;
  assign y9 = n666;
  assign y10 = n671;
endmodule
