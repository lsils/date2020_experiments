// Benchmark "auction_BMR_3_32" written by ABC on Tue Nov 26 13:54:14 2019

module auction_BMR_3_32 ( 
    \p_input[0] , \p_input[1] , \p_input[2] , \p_input[3] , \p_input[4] ,
    \p_input[5] , \p_input[6] , \p_input[7] , \p_input[8] , \p_input[9] ,
    \p_input[10] , \p_input[11] , \p_input[12] , \p_input[13] ,
    \p_input[14] , \p_input[15] , \p_input[16] , \p_input[17] ,
    \p_input[18] , \p_input[19] , \p_input[20] , \p_input[21] ,
    \p_input[22] , \p_input[23] , \p_input[24] , \p_input[25] ,
    \p_input[26] , \p_input[27] , \p_input[28] , \p_input[29] ,
    \p_input[30] , \p_input[31] , \p_input[32] , \p_input[33] ,
    \p_input[34] , \p_input[35] , \p_input[36] , \p_input[37] ,
    \p_input[38] , \p_input[39] , \p_input[40] , \p_input[41] ,
    \p_input[42] , \p_input[43] , \p_input[44] , \p_input[45] ,
    \p_input[46] , \p_input[47] , \p_input[48] , \p_input[49] ,
    \p_input[50] , \p_input[51] , \p_input[52] , \p_input[53] ,
    \p_input[54] , \p_input[55] , \p_input[56] , \p_input[57] ,
    \p_input[58] , \p_input[59] , \p_input[60] , \p_input[61] ,
    \p_input[62] , \p_input[63] , \p_input[64] , \p_input[65] ,
    \p_input[66] , \p_input[67] , \p_input[68] , \p_input[69] ,
    \p_input[70] , \p_input[71] , \p_input[72] , \p_input[73] ,
    \p_input[74] , \p_input[75] , \p_input[76] , \p_input[77] ,
    \p_input[78] , \p_input[79] , \p_input[80] , \p_input[81] ,
    \p_input[82] , \p_input[83] , \p_input[84] , \p_input[85] ,
    \p_input[86] , \p_input[87] , \p_input[88] , \p_input[89] ,
    \p_input[90] , \p_input[91] , \p_input[92] , \p_input[93] ,
    \p_input[94] , \p_input[95] , \p_input[96] , \p_input[97] ,
    \p_input[98] , \p_input[99] , \p_input[100] , \p_input[101] ,
    \p_input[102] , \p_input[103] , \p_input[104] , \p_input[105] ,
    \p_input[106] , \p_input[107] , \p_input[108] , \p_input[109] ,
    \p_input[110] , \p_input[111] , \p_input[112] , \p_input[113] ,
    \p_input[114] , \p_input[115] , \p_input[116] , \p_input[117] ,
    \p_input[118] , \p_input[119] , \p_input[120] , \p_input[121] ,
    \p_input[122] , \p_input[123] , \p_input[124] , \p_input[125] ,
    \p_input[126] , \p_input[127] , \p_input[128] , \p_input[129] ,
    \p_input[130] , \p_input[131] , \p_input[132] , \p_input[133] ,
    \p_input[134] , \p_input[135] , \p_input[136] , \p_input[137] ,
    \p_input[138] , \p_input[139] , \p_input[140] , \p_input[141] ,
    \p_input[142] , \p_input[143] , \p_input[144] , \p_input[145] ,
    \p_input[146] , \p_input[147] , \p_input[148] , \p_input[149] ,
    \p_input[150] , \p_input[151] , \p_input[152] , \p_input[153] ,
    \p_input[154] , \p_input[155] , \p_input[156] , \p_input[157] ,
    \p_input[158] , \p_input[159] , \p_input[160] , \p_input[161] ,
    \p_input[162] , \p_input[163] , \p_input[164] , \p_input[165] ,
    \p_input[166] , \p_input[167] , \p_input[168] , \p_input[169] ,
    \p_input[170] , \p_input[171] , \p_input[172] , \p_input[173] ,
    \p_input[174] , \p_input[175] , \p_input[176] , \p_input[177] ,
    \p_input[178] , \p_input[179] , \p_input[180] , \p_input[181] ,
    \p_input[182] , \p_input[183] , \p_input[184] , \p_input[185] ,
    \p_input[186] , \p_input[187] , \p_input[188] , \p_input[189] ,
    \p_input[190] , \p_input[191] , \p_input[192] , \p_input[193] ,
    \p_input[194] , \p_input[195] , \p_input[196] , \p_input[197] ,
    \p_input[198] , \p_input[199] , \p_input[200] , \p_input[201] ,
    \p_input[202] , \p_input[203] , \p_input[204] , \p_input[205] ,
    \p_input[206] , \p_input[207] , \p_input[208] , \p_input[209] ,
    \p_input[210] , \p_input[211] , \p_input[212] , \p_input[213] ,
    \p_input[214] , \p_input[215] , \p_input[216] , \p_input[217] ,
    \p_input[218] , \p_input[219] , \p_input[220] , \p_input[221] ,
    \p_input[222] , \p_input[223] , \p_input[224] , \p_input[225] ,
    \p_input[226] , \p_input[227] , \p_input[228] , \p_input[229] ,
    \p_input[230] , \p_input[231] , \p_input[232] , \p_input[233] ,
    \p_input[234] , \p_input[235] , \p_input[236] , \p_input[237] ,
    \p_input[238] , \p_input[239] , \p_input[240] , \p_input[241] ,
    \p_input[242] , \p_input[243] , \p_input[244] , \p_input[245] ,
    \p_input[246] , \p_input[247] , \p_input[248] , \p_input[249] ,
    \p_input[250] , \p_input[251] , \p_input[252] , \p_input[253] ,
    \p_input[254] , \p_input[255] ,
    \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] , \o[8] ,
    \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] , \o[16] ,
    \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] , \o[24] ,
    \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] , \o[32] ,
    \o[33] , \o[34]   );
  input  \p_input[0] , \p_input[1] , \p_input[2] , \p_input[3] ,
    \p_input[4] , \p_input[5] , \p_input[6] , \p_input[7] , \p_input[8] ,
    \p_input[9] , \p_input[10] , \p_input[11] , \p_input[12] ,
    \p_input[13] , \p_input[14] , \p_input[15] , \p_input[16] ,
    \p_input[17] , \p_input[18] , \p_input[19] , \p_input[20] ,
    \p_input[21] , \p_input[22] , \p_input[23] , \p_input[24] ,
    \p_input[25] , \p_input[26] , \p_input[27] , \p_input[28] ,
    \p_input[29] , \p_input[30] , \p_input[31] , \p_input[32] ,
    \p_input[33] , \p_input[34] , \p_input[35] , \p_input[36] ,
    \p_input[37] , \p_input[38] , \p_input[39] , \p_input[40] ,
    \p_input[41] , \p_input[42] , \p_input[43] , \p_input[44] ,
    \p_input[45] , \p_input[46] , \p_input[47] , \p_input[48] ,
    \p_input[49] , \p_input[50] , \p_input[51] , \p_input[52] ,
    \p_input[53] , \p_input[54] , \p_input[55] , \p_input[56] ,
    \p_input[57] , \p_input[58] , \p_input[59] , \p_input[60] ,
    \p_input[61] , \p_input[62] , \p_input[63] , \p_input[64] ,
    \p_input[65] , \p_input[66] , \p_input[67] , \p_input[68] ,
    \p_input[69] , \p_input[70] , \p_input[71] , \p_input[72] ,
    \p_input[73] , \p_input[74] , \p_input[75] , \p_input[76] ,
    \p_input[77] , \p_input[78] , \p_input[79] , \p_input[80] ,
    \p_input[81] , \p_input[82] , \p_input[83] , \p_input[84] ,
    \p_input[85] , \p_input[86] , \p_input[87] , \p_input[88] ,
    \p_input[89] , \p_input[90] , \p_input[91] , \p_input[92] ,
    \p_input[93] , \p_input[94] , \p_input[95] , \p_input[96] ,
    \p_input[97] , \p_input[98] , \p_input[99] , \p_input[100] ,
    \p_input[101] , \p_input[102] , \p_input[103] , \p_input[104] ,
    \p_input[105] , \p_input[106] , \p_input[107] , \p_input[108] ,
    \p_input[109] , \p_input[110] , \p_input[111] , \p_input[112] ,
    \p_input[113] , \p_input[114] , \p_input[115] , \p_input[116] ,
    \p_input[117] , \p_input[118] , \p_input[119] , \p_input[120] ,
    \p_input[121] , \p_input[122] , \p_input[123] , \p_input[124] ,
    \p_input[125] , \p_input[126] , \p_input[127] , \p_input[128] ,
    \p_input[129] , \p_input[130] , \p_input[131] , \p_input[132] ,
    \p_input[133] , \p_input[134] , \p_input[135] , \p_input[136] ,
    \p_input[137] , \p_input[138] , \p_input[139] , \p_input[140] ,
    \p_input[141] , \p_input[142] , \p_input[143] , \p_input[144] ,
    \p_input[145] , \p_input[146] , \p_input[147] , \p_input[148] ,
    \p_input[149] , \p_input[150] , \p_input[151] , \p_input[152] ,
    \p_input[153] , \p_input[154] , \p_input[155] , \p_input[156] ,
    \p_input[157] , \p_input[158] , \p_input[159] , \p_input[160] ,
    \p_input[161] , \p_input[162] , \p_input[163] , \p_input[164] ,
    \p_input[165] , \p_input[166] , \p_input[167] , \p_input[168] ,
    \p_input[169] , \p_input[170] , \p_input[171] , \p_input[172] ,
    \p_input[173] , \p_input[174] , \p_input[175] , \p_input[176] ,
    \p_input[177] , \p_input[178] , \p_input[179] , \p_input[180] ,
    \p_input[181] , \p_input[182] , \p_input[183] , \p_input[184] ,
    \p_input[185] , \p_input[186] , \p_input[187] , \p_input[188] ,
    \p_input[189] , \p_input[190] , \p_input[191] , \p_input[192] ,
    \p_input[193] , \p_input[194] , \p_input[195] , \p_input[196] ,
    \p_input[197] , \p_input[198] , \p_input[199] , \p_input[200] ,
    \p_input[201] , \p_input[202] , \p_input[203] , \p_input[204] ,
    \p_input[205] , \p_input[206] , \p_input[207] , \p_input[208] ,
    \p_input[209] , \p_input[210] , \p_input[211] , \p_input[212] ,
    \p_input[213] , \p_input[214] , \p_input[215] , \p_input[216] ,
    \p_input[217] , \p_input[218] , \p_input[219] , \p_input[220] ,
    \p_input[221] , \p_input[222] , \p_input[223] , \p_input[224] ,
    \p_input[225] , \p_input[226] , \p_input[227] , \p_input[228] ,
    \p_input[229] , \p_input[230] , \p_input[231] , \p_input[232] ,
    \p_input[233] , \p_input[234] , \p_input[235] , \p_input[236] ,
    \p_input[237] , \p_input[238] , \p_input[239] , \p_input[240] ,
    \p_input[241] , \p_input[242] , \p_input[243] , \p_input[244] ,
    \p_input[245] , \p_input[246] , \p_input[247] , \p_input[248] ,
    \p_input[249] , \p_input[250] , \p_input[251] , \p_input[252] ,
    \p_input[253] , \p_input[254] , \p_input[255] ;
  output \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] ,
    \o[8] , \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] ,
    \o[16] , \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] ,
    \o[24] , \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] ,
    \o[32] , \o[33] , \o[34] ;
  wire new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1731_, new_n1732_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1743_, new_n1744_, new_n1746_, new_n1747_,
    new_n1749_, new_n1750_, new_n1752_, new_n1753_, new_n1755_, new_n1756_,
    new_n1758_, new_n1759_, new_n1761_, new_n1762_, new_n1764_, new_n1765_,
    new_n1767_, new_n1768_, new_n1770_, new_n1771_, new_n1773_, new_n1774_,
    new_n1776_, new_n1777_, new_n1779_, new_n1780_, new_n1782_, new_n1783_,
    new_n1785_, new_n1786_, new_n1788_, new_n1789_, new_n1791_, new_n1792_,
    new_n1794_, new_n1795_, new_n1797_, new_n1798_, new_n1800_, new_n1801_,
    new_n1803_, new_n1804_, new_n1806_, new_n1807_, new_n1809_, new_n1810_,
    new_n1812_, new_n1813_, new_n1815_, new_n1816_, new_n1818_, new_n1819_,
    new_n1821_, new_n1822_, new_n1824_, new_n1825_, new_n1827_, new_n1828_,
    new_n1830_, new_n1831_, new_n1833_, new_n1834_;
  assign new_n292_ = ~\p_input[159]  & ~\p_input[191] ;
  assign new_n293_ = ~\p_input[223]  & ~\p_input[255] ;
  assign new_n294_ = new_n292_ & new_n293_;
  assign new_n295_ = ~\p_input[31]  & ~\p_input[63] ;
  assign new_n296_ = ~\p_input[95]  & ~\p_input[127] ;
  assign new_n297_ = new_n295_ & new_n296_;
  assign new_n298_ = new_n294_ & ~new_n297_;
  assign new_n299_ = ~\p_input[31]  & \p_input[63] ;
  assign new_n300_ = \p_input[31]  & ~\p_input[63] ;
  assign new_n301_ = ~\p_input[30]  & \p_input[62] ;
  assign new_n302_ = \p_input[30]  & ~\p_input[62] ;
  assign new_n303_ = ~\p_input[29]  & \p_input[61] ;
  assign new_n304_ = \p_input[29]  & ~\p_input[61] ;
  assign new_n305_ = ~\p_input[28]  & \p_input[60] ;
  assign new_n306_ = \p_input[28]  & ~\p_input[60] ;
  assign new_n307_ = ~\p_input[27]  & \p_input[59] ;
  assign new_n308_ = \p_input[27]  & ~\p_input[59] ;
  assign new_n309_ = ~\p_input[26]  & \p_input[58] ;
  assign new_n310_ = \p_input[26]  & ~\p_input[58] ;
  assign new_n311_ = ~\p_input[25]  & \p_input[57] ;
  assign new_n312_ = \p_input[25]  & ~\p_input[57] ;
  assign new_n313_ = ~\p_input[24]  & \p_input[56] ;
  assign new_n314_ = \p_input[24]  & ~\p_input[56] ;
  assign new_n315_ = ~\p_input[23]  & \p_input[55] ;
  assign new_n316_ = \p_input[23]  & ~\p_input[55] ;
  assign new_n317_ = ~\p_input[22]  & \p_input[54] ;
  assign new_n318_ = \p_input[22]  & ~\p_input[54] ;
  assign new_n319_ = ~\p_input[21]  & \p_input[53] ;
  assign new_n320_ = \p_input[21]  & ~\p_input[53] ;
  assign new_n321_ = ~\p_input[20]  & \p_input[52] ;
  assign new_n322_ = \p_input[20]  & ~\p_input[52] ;
  assign new_n323_ = ~\p_input[19]  & \p_input[51] ;
  assign new_n324_ = \p_input[19]  & ~\p_input[51] ;
  assign new_n325_ = ~\p_input[18]  & \p_input[50] ;
  assign new_n326_ = \p_input[18]  & ~\p_input[50] ;
  assign new_n327_ = ~\p_input[17]  & \p_input[49] ;
  assign new_n328_ = \p_input[17]  & ~\p_input[49] ;
  assign new_n329_ = ~\p_input[16]  & \p_input[48] ;
  assign new_n330_ = \p_input[16]  & ~\p_input[48] ;
  assign new_n331_ = ~\p_input[15]  & \p_input[47] ;
  assign new_n332_ = \p_input[15]  & ~\p_input[47] ;
  assign new_n333_ = ~\p_input[14]  & \p_input[46] ;
  assign new_n334_ = \p_input[14]  & ~\p_input[46] ;
  assign new_n335_ = ~\p_input[13]  & \p_input[45] ;
  assign new_n336_ = \p_input[13]  & ~\p_input[45] ;
  assign new_n337_ = ~\p_input[12]  & \p_input[44] ;
  assign new_n338_ = \p_input[12]  & ~\p_input[44] ;
  assign new_n339_ = ~\p_input[11]  & \p_input[43] ;
  assign new_n340_ = \p_input[11]  & ~\p_input[43] ;
  assign new_n341_ = ~\p_input[10]  & \p_input[42] ;
  assign new_n342_ = \p_input[10]  & ~\p_input[42] ;
  assign new_n343_ = ~\p_input[9]  & \p_input[41] ;
  assign new_n344_ = \p_input[9]  & ~\p_input[41] ;
  assign new_n345_ = ~\p_input[8]  & \p_input[40] ;
  assign new_n346_ = \p_input[8]  & ~\p_input[40] ;
  assign new_n347_ = ~\p_input[7]  & \p_input[39] ;
  assign new_n348_ = \p_input[7]  & ~\p_input[39] ;
  assign new_n349_ = ~\p_input[6]  & \p_input[38] ;
  assign new_n350_ = \p_input[6]  & ~\p_input[38] ;
  assign new_n351_ = ~\p_input[5]  & \p_input[37] ;
  assign new_n352_ = \p_input[5]  & ~\p_input[37] ;
  assign new_n353_ = ~\p_input[4]  & \p_input[36] ;
  assign new_n354_ = \p_input[4]  & ~\p_input[36] ;
  assign new_n355_ = ~\p_input[3]  & \p_input[35] ;
  assign new_n356_ = \p_input[3]  & ~\p_input[35] ;
  assign new_n357_ = ~\p_input[2]  & \p_input[34] ;
  assign new_n358_ = \p_input[2]  & ~\p_input[34] ;
  assign new_n359_ = ~\p_input[1]  & \p_input[33] ;
  assign new_n360_ = \p_input[1]  & ~\p_input[33] ;
  assign new_n361_ = \p_input[0]  & ~\p_input[32] ;
  assign new_n362_ = ~new_n360_ & ~new_n361_;
  assign new_n363_ = ~new_n359_ & ~new_n362_;
  assign new_n364_ = ~new_n358_ & ~new_n363_;
  assign new_n365_ = ~new_n357_ & ~new_n364_;
  assign new_n366_ = ~new_n356_ & ~new_n365_;
  assign new_n367_ = ~new_n355_ & ~new_n366_;
  assign new_n368_ = ~new_n354_ & ~new_n367_;
  assign new_n369_ = ~new_n353_ & ~new_n368_;
  assign new_n370_ = ~new_n352_ & ~new_n369_;
  assign new_n371_ = ~new_n351_ & ~new_n370_;
  assign new_n372_ = ~new_n350_ & ~new_n371_;
  assign new_n373_ = ~new_n349_ & ~new_n372_;
  assign new_n374_ = ~new_n348_ & ~new_n373_;
  assign new_n375_ = ~new_n347_ & ~new_n374_;
  assign new_n376_ = ~new_n346_ & ~new_n375_;
  assign new_n377_ = ~new_n345_ & ~new_n376_;
  assign new_n378_ = ~new_n344_ & ~new_n377_;
  assign new_n379_ = ~new_n343_ & ~new_n378_;
  assign new_n380_ = ~new_n342_ & ~new_n379_;
  assign new_n381_ = ~new_n341_ & ~new_n380_;
  assign new_n382_ = ~new_n340_ & ~new_n381_;
  assign new_n383_ = ~new_n339_ & ~new_n382_;
  assign new_n384_ = ~new_n338_ & ~new_n383_;
  assign new_n385_ = ~new_n337_ & ~new_n384_;
  assign new_n386_ = ~new_n336_ & ~new_n385_;
  assign new_n387_ = ~new_n335_ & ~new_n386_;
  assign new_n388_ = ~new_n334_ & ~new_n387_;
  assign new_n389_ = ~new_n333_ & ~new_n388_;
  assign new_n390_ = ~new_n332_ & ~new_n389_;
  assign new_n391_ = ~new_n331_ & ~new_n390_;
  assign new_n392_ = ~new_n330_ & ~new_n391_;
  assign new_n393_ = ~new_n329_ & ~new_n392_;
  assign new_n394_ = ~new_n328_ & ~new_n393_;
  assign new_n395_ = ~new_n327_ & ~new_n394_;
  assign new_n396_ = ~new_n326_ & ~new_n395_;
  assign new_n397_ = ~new_n325_ & ~new_n396_;
  assign new_n398_ = ~new_n324_ & ~new_n397_;
  assign new_n399_ = ~new_n323_ & ~new_n398_;
  assign new_n400_ = ~new_n322_ & ~new_n399_;
  assign new_n401_ = ~new_n321_ & ~new_n400_;
  assign new_n402_ = ~new_n320_ & ~new_n401_;
  assign new_n403_ = ~new_n319_ & ~new_n402_;
  assign new_n404_ = ~new_n318_ & ~new_n403_;
  assign new_n405_ = ~new_n317_ & ~new_n404_;
  assign new_n406_ = ~new_n316_ & ~new_n405_;
  assign new_n407_ = ~new_n315_ & ~new_n406_;
  assign new_n408_ = ~new_n314_ & ~new_n407_;
  assign new_n409_ = ~new_n313_ & ~new_n408_;
  assign new_n410_ = ~new_n312_ & ~new_n409_;
  assign new_n411_ = ~new_n311_ & ~new_n410_;
  assign new_n412_ = ~new_n310_ & ~new_n411_;
  assign new_n413_ = ~new_n309_ & ~new_n412_;
  assign new_n414_ = ~new_n308_ & ~new_n413_;
  assign new_n415_ = ~new_n307_ & ~new_n414_;
  assign new_n416_ = ~new_n306_ & ~new_n415_;
  assign new_n417_ = ~new_n305_ & ~new_n416_;
  assign new_n418_ = ~new_n304_ & ~new_n417_;
  assign new_n419_ = ~new_n303_ & ~new_n418_;
  assign new_n420_ = ~new_n302_ & ~new_n419_;
  assign new_n421_ = ~new_n301_ & ~new_n420_;
  assign new_n422_ = ~new_n300_ & ~new_n421_;
  assign new_n423_ = ~new_n299_ & ~new_n422_;
  assign new_n424_ = \p_input[33]  & ~new_n423_;
  assign new_n425_ = \p_input[1]  & new_n423_;
  assign new_n426_ = ~new_n424_ & ~new_n425_;
  assign new_n427_ = new_n295_ & ~new_n296_;
  assign new_n428_ = ~new_n295_ & new_n296_;
  assign new_n429_ = ~\p_input[95]  & \p_input[127] ;
  assign new_n430_ = \p_input[95]  & ~\p_input[127] ;
  assign new_n431_ = ~\p_input[94]  & \p_input[126] ;
  assign new_n432_ = \p_input[94]  & ~\p_input[126] ;
  assign new_n433_ = ~\p_input[93]  & \p_input[125] ;
  assign new_n434_ = \p_input[93]  & ~\p_input[125] ;
  assign new_n435_ = ~\p_input[92]  & \p_input[124] ;
  assign new_n436_ = \p_input[92]  & ~\p_input[124] ;
  assign new_n437_ = ~\p_input[91]  & \p_input[123] ;
  assign new_n438_ = \p_input[91]  & ~\p_input[123] ;
  assign new_n439_ = ~\p_input[90]  & \p_input[122] ;
  assign new_n440_ = \p_input[90]  & ~\p_input[122] ;
  assign new_n441_ = ~\p_input[89]  & \p_input[121] ;
  assign new_n442_ = \p_input[89]  & ~\p_input[121] ;
  assign new_n443_ = ~\p_input[88]  & \p_input[120] ;
  assign new_n444_ = \p_input[88]  & ~\p_input[120] ;
  assign new_n445_ = ~\p_input[87]  & \p_input[119] ;
  assign new_n446_ = \p_input[87]  & ~\p_input[119] ;
  assign new_n447_ = ~\p_input[86]  & \p_input[118] ;
  assign new_n448_ = \p_input[86]  & ~\p_input[118] ;
  assign new_n449_ = ~\p_input[85]  & \p_input[117] ;
  assign new_n450_ = \p_input[85]  & ~\p_input[117] ;
  assign new_n451_ = ~\p_input[84]  & \p_input[116] ;
  assign new_n452_ = \p_input[84]  & ~\p_input[116] ;
  assign new_n453_ = ~\p_input[83]  & \p_input[115] ;
  assign new_n454_ = \p_input[83]  & ~\p_input[115] ;
  assign new_n455_ = ~\p_input[82]  & \p_input[114] ;
  assign new_n456_ = \p_input[82]  & ~\p_input[114] ;
  assign new_n457_ = ~\p_input[81]  & \p_input[113] ;
  assign new_n458_ = \p_input[81]  & ~\p_input[113] ;
  assign new_n459_ = ~\p_input[80]  & \p_input[112] ;
  assign new_n460_ = \p_input[80]  & ~\p_input[112] ;
  assign new_n461_ = ~\p_input[79]  & \p_input[111] ;
  assign new_n462_ = \p_input[79]  & ~\p_input[111] ;
  assign new_n463_ = ~\p_input[78]  & \p_input[110] ;
  assign new_n464_ = \p_input[78]  & ~\p_input[110] ;
  assign new_n465_ = ~\p_input[77]  & \p_input[109] ;
  assign new_n466_ = \p_input[77]  & ~\p_input[109] ;
  assign new_n467_ = ~\p_input[76]  & \p_input[108] ;
  assign new_n468_ = \p_input[76]  & ~\p_input[108] ;
  assign new_n469_ = ~\p_input[75]  & \p_input[107] ;
  assign new_n470_ = \p_input[75]  & ~\p_input[107] ;
  assign new_n471_ = ~\p_input[74]  & \p_input[106] ;
  assign new_n472_ = \p_input[74]  & ~\p_input[106] ;
  assign new_n473_ = ~\p_input[73]  & \p_input[105] ;
  assign new_n474_ = \p_input[73]  & ~\p_input[105] ;
  assign new_n475_ = ~\p_input[72]  & \p_input[104] ;
  assign new_n476_ = \p_input[72]  & ~\p_input[104] ;
  assign new_n477_ = ~\p_input[71]  & \p_input[103] ;
  assign new_n478_ = \p_input[71]  & ~\p_input[103] ;
  assign new_n479_ = ~\p_input[70]  & \p_input[102] ;
  assign new_n480_ = \p_input[70]  & ~\p_input[102] ;
  assign new_n481_ = ~\p_input[69]  & \p_input[101] ;
  assign new_n482_ = \p_input[69]  & ~\p_input[101] ;
  assign new_n483_ = ~\p_input[68]  & \p_input[100] ;
  assign new_n484_ = \p_input[68]  & ~\p_input[100] ;
  assign new_n485_ = ~\p_input[67]  & \p_input[99] ;
  assign new_n486_ = \p_input[67]  & ~\p_input[99] ;
  assign new_n487_ = ~\p_input[66]  & \p_input[98] ;
  assign new_n488_ = \p_input[66]  & ~\p_input[98] ;
  assign new_n489_ = ~\p_input[65]  & \p_input[97] ;
  assign new_n490_ = \p_input[65]  & ~\p_input[97] ;
  assign new_n491_ = \p_input[64]  & ~\p_input[96] ;
  assign new_n492_ = ~new_n490_ & ~new_n491_;
  assign new_n493_ = ~new_n489_ & ~new_n492_;
  assign new_n494_ = ~new_n488_ & ~new_n493_;
  assign new_n495_ = ~new_n487_ & ~new_n494_;
  assign new_n496_ = ~new_n486_ & ~new_n495_;
  assign new_n497_ = ~new_n485_ & ~new_n496_;
  assign new_n498_ = ~new_n484_ & ~new_n497_;
  assign new_n499_ = ~new_n483_ & ~new_n498_;
  assign new_n500_ = ~new_n482_ & ~new_n499_;
  assign new_n501_ = ~new_n481_ & ~new_n500_;
  assign new_n502_ = ~new_n480_ & ~new_n501_;
  assign new_n503_ = ~new_n479_ & ~new_n502_;
  assign new_n504_ = ~new_n478_ & ~new_n503_;
  assign new_n505_ = ~new_n477_ & ~new_n504_;
  assign new_n506_ = ~new_n476_ & ~new_n505_;
  assign new_n507_ = ~new_n475_ & ~new_n506_;
  assign new_n508_ = ~new_n474_ & ~new_n507_;
  assign new_n509_ = ~new_n473_ & ~new_n508_;
  assign new_n510_ = ~new_n472_ & ~new_n509_;
  assign new_n511_ = ~new_n471_ & ~new_n510_;
  assign new_n512_ = ~new_n470_ & ~new_n511_;
  assign new_n513_ = ~new_n469_ & ~new_n512_;
  assign new_n514_ = ~new_n468_ & ~new_n513_;
  assign new_n515_ = ~new_n467_ & ~new_n514_;
  assign new_n516_ = ~new_n466_ & ~new_n515_;
  assign new_n517_ = ~new_n465_ & ~new_n516_;
  assign new_n518_ = ~new_n464_ & ~new_n517_;
  assign new_n519_ = ~new_n463_ & ~new_n518_;
  assign new_n520_ = ~new_n462_ & ~new_n519_;
  assign new_n521_ = ~new_n461_ & ~new_n520_;
  assign new_n522_ = ~new_n460_ & ~new_n521_;
  assign new_n523_ = ~new_n459_ & ~new_n522_;
  assign new_n524_ = ~new_n458_ & ~new_n523_;
  assign new_n525_ = ~new_n457_ & ~new_n524_;
  assign new_n526_ = ~new_n456_ & ~new_n525_;
  assign new_n527_ = ~new_n455_ & ~new_n526_;
  assign new_n528_ = ~new_n454_ & ~new_n527_;
  assign new_n529_ = ~new_n453_ & ~new_n528_;
  assign new_n530_ = ~new_n452_ & ~new_n529_;
  assign new_n531_ = ~new_n451_ & ~new_n530_;
  assign new_n532_ = ~new_n450_ & ~new_n531_;
  assign new_n533_ = ~new_n449_ & ~new_n532_;
  assign new_n534_ = ~new_n448_ & ~new_n533_;
  assign new_n535_ = ~new_n447_ & ~new_n534_;
  assign new_n536_ = ~new_n446_ & ~new_n535_;
  assign new_n537_ = ~new_n445_ & ~new_n536_;
  assign new_n538_ = ~new_n444_ & ~new_n537_;
  assign new_n539_ = ~new_n443_ & ~new_n538_;
  assign new_n540_ = ~new_n442_ & ~new_n539_;
  assign new_n541_ = ~new_n441_ & ~new_n540_;
  assign new_n542_ = ~new_n440_ & ~new_n541_;
  assign new_n543_ = ~new_n439_ & ~new_n542_;
  assign new_n544_ = ~new_n438_ & ~new_n543_;
  assign new_n545_ = ~new_n437_ & ~new_n544_;
  assign new_n546_ = ~new_n436_ & ~new_n545_;
  assign new_n547_ = ~new_n435_ & ~new_n546_;
  assign new_n548_ = ~new_n434_ & ~new_n547_;
  assign new_n549_ = ~new_n433_ & ~new_n548_;
  assign new_n550_ = ~new_n432_ & ~new_n549_;
  assign new_n551_ = ~new_n431_ & ~new_n550_;
  assign new_n552_ = ~new_n430_ & ~new_n551_;
  assign new_n553_ = ~new_n429_ & ~new_n552_;
  assign new_n554_ = \p_input[126]  & ~new_n553_;
  assign new_n555_ = \p_input[94]  & new_n553_;
  assign new_n556_ = ~new_n554_ & ~new_n555_;
  assign new_n557_ = \p_input[62]  & ~new_n423_;
  assign new_n558_ = \p_input[30]  & new_n423_;
  assign new_n559_ = ~new_n557_ & ~new_n558_;
  assign new_n560_ = ~new_n556_ & new_n559_;
  assign new_n561_ = \p_input[97]  & ~new_n553_;
  assign new_n562_ = \p_input[65]  & new_n553_;
  assign new_n563_ = ~new_n561_ & ~new_n562_;
  assign new_n564_ = new_n426_ & ~new_n563_;
  assign new_n565_ = \p_input[96]  & ~new_n553_;
  assign new_n566_ = \p_input[64]  & new_n553_;
  assign new_n567_ = ~new_n565_ & ~new_n566_;
  assign new_n568_ = \p_input[32]  & ~new_n423_;
  assign new_n569_ = \p_input[0]  & new_n423_;
  assign new_n570_ = ~new_n568_ & ~new_n569_;
  assign new_n571_ = new_n567_ & ~new_n570_;
  assign new_n572_ = ~new_n564_ & new_n571_;
  assign new_n573_ = \p_input[98]  & ~new_n553_;
  assign new_n574_ = \p_input[66]  & new_n553_;
  assign new_n575_ = ~new_n573_ & ~new_n574_;
  assign new_n576_ = \p_input[34]  & ~new_n423_;
  assign new_n577_ = \p_input[2]  & new_n423_;
  assign new_n578_ = ~new_n576_ & ~new_n577_;
  assign new_n579_ = new_n575_ & ~new_n578_;
  assign new_n580_ = ~new_n426_ & new_n563_;
  assign new_n581_ = ~new_n579_ & ~new_n580_;
  assign new_n582_ = ~new_n572_ & new_n581_;
  assign new_n583_ = \p_input[35]  & ~new_n423_;
  assign new_n584_ = \p_input[3]  & new_n423_;
  assign new_n585_ = ~new_n583_ & ~new_n584_;
  assign new_n586_ = \p_input[99]  & ~new_n553_;
  assign new_n587_ = \p_input[67]  & new_n553_;
  assign new_n588_ = ~new_n586_ & ~new_n587_;
  assign new_n589_ = new_n585_ & ~new_n588_;
  assign new_n590_ = ~new_n575_ & new_n578_;
  assign new_n591_ = ~new_n589_ & ~new_n590_;
  assign new_n592_ = ~new_n582_ & new_n591_;
  assign new_n593_ = \p_input[100]  & ~new_n553_;
  assign new_n594_ = \p_input[68]  & new_n553_;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign new_n596_ = \p_input[36]  & ~new_n423_;
  assign new_n597_ = \p_input[4]  & new_n423_;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = new_n595_ & ~new_n598_;
  assign new_n600_ = ~new_n585_ & new_n588_;
  assign new_n601_ = ~new_n599_ & ~new_n600_;
  assign new_n602_ = ~new_n592_ & new_n601_;
  assign new_n603_ = \p_input[101]  & ~new_n553_;
  assign new_n604_ = \p_input[69]  & new_n553_;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = \p_input[37]  & ~new_n423_;
  assign new_n607_ = \p_input[5]  & new_n423_;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = ~new_n605_ & new_n608_;
  assign new_n610_ = ~new_n595_ & new_n598_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = ~new_n602_ & new_n611_;
  assign new_n613_ = \p_input[38]  & ~new_n423_;
  assign new_n614_ = \p_input[6]  & new_n423_;
  assign new_n615_ = ~new_n613_ & ~new_n614_;
  assign new_n616_ = \p_input[102]  & ~new_n553_;
  assign new_n617_ = \p_input[70]  & new_n553_;
  assign new_n618_ = ~new_n616_ & ~new_n617_;
  assign new_n619_ = ~new_n615_ & new_n618_;
  assign new_n620_ = new_n605_ & ~new_n608_;
  assign new_n621_ = ~new_n619_ & ~new_n620_;
  assign new_n622_ = ~new_n612_ & new_n621_;
  assign new_n623_ = \p_input[39]  & ~new_n423_;
  assign new_n624_ = \p_input[7]  & new_n423_;
  assign new_n625_ = ~new_n623_ & ~new_n624_;
  assign new_n626_ = \p_input[103]  & ~new_n553_;
  assign new_n627_ = \p_input[71]  & new_n553_;
  assign new_n628_ = ~new_n626_ & ~new_n627_;
  assign new_n629_ = new_n625_ & ~new_n628_;
  assign new_n630_ = new_n615_ & ~new_n618_;
  assign new_n631_ = ~new_n629_ & ~new_n630_;
  assign new_n632_ = ~new_n622_ & new_n631_;
  assign new_n633_ = ~new_n625_ & new_n628_;
  assign new_n634_ = \p_input[104]  & ~new_n553_;
  assign new_n635_ = \p_input[72]  & new_n553_;
  assign new_n636_ = ~new_n634_ & ~new_n635_;
  assign new_n637_ = \p_input[40]  & ~new_n423_;
  assign new_n638_ = \p_input[8]  & new_n423_;
  assign new_n639_ = ~new_n637_ & ~new_n638_;
  assign new_n640_ = new_n636_ & ~new_n639_;
  assign new_n641_ = ~new_n633_ & ~new_n640_;
  assign new_n642_ = ~new_n632_ & new_n641_;
  assign new_n643_ = ~new_n636_ & new_n639_;
  assign new_n644_ = \p_input[105]  & ~new_n553_;
  assign new_n645_ = \p_input[73]  & new_n553_;
  assign new_n646_ = ~new_n644_ & ~new_n645_;
  assign new_n647_ = \p_input[41]  & ~new_n423_;
  assign new_n648_ = \p_input[9]  & new_n423_;
  assign new_n649_ = ~new_n647_ & ~new_n648_;
  assign new_n650_ = ~new_n646_ & new_n649_;
  assign new_n651_ = ~new_n643_ & ~new_n650_;
  assign new_n652_ = ~new_n642_ & new_n651_;
  assign new_n653_ = new_n646_ & ~new_n649_;
  assign new_n654_ = \p_input[42]  & ~new_n423_;
  assign new_n655_ = \p_input[10]  & new_n423_;
  assign new_n656_ = ~new_n654_ & ~new_n655_;
  assign new_n657_ = \p_input[106]  & ~new_n553_;
  assign new_n658_ = \p_input[74]  & new_n553_;
  assign new_n659_ = ~new_n657_ & ~new_n658_;
  assign new_n660_ = ~new_n656_ & new_n659_;
  assign new_n661_ = ~new_n653_ & ~new_n660_;
  assign new_n662_ = ~new_n652_ & new_n661_;
  assign new_n663_ = \p_input[43]  & ~new_n423_;
  assign new_n664_ = \p_input[11]  & new_n423_;
  assign new_n665_ = ~new_n663_ & ~new_n664_;
  assign new_n666_ = \p_input[107]  & ~new_n553_;
  assign new_n667_ = \p_input[75]  & new_n553_;
  assign new_n668_ = ~new_n666_ & ~new_n667_;
  assign new_n669_ = new_n665_ & ~new_n668_;
  assign new_n670_ = new_n656_ & ~new_n659_;
  assign new_n671_ = ~new_n669_ & ~new_n670_;
  assign new_n672_ = ~new_n662_ & new_n671_;
  assign new_n673_ = \p_input[108]  & ~new_n553_;
  assign new_n674_ = \p_input[76]  & new_n553_;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = \p_input[44]  & ~new_n423_;
  assign new_n677_ = \p_input[12]  & new_n423_;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign new_n679_ = new_n675_ & ~new_n678_;
  assign new_n680_ = ~new_n665_ & new_n668_;
  assign new_n681_ = ~new_n679_ & ~new_n680_;
  assign new_n682_ = ~new_n672_ & new_n681_;
  assign new_n683_ = ~new_n675_ & new_n678_;
  assign new_n684_ = \p_input[109]  & ~new_n553_;
  assign new_n685_ = \p_input[77]  & new_n553_;
  assign new_n686_ = ~new_n684_ & ~new_n685_;
  assign new_n687_ = \p_input[45]  & ~new_n423_;
  assign new_n688_ = \p_input[13]  & new_n423_;
  assign new_n689_ = ~new_n687_ & ~new_n688_;
  assign new_n690_ = ~new_n686_ & new_n689_;
  assign new_n691_ = ~new_n683_ & ~new_n690_;
  assign new_n692_ = ~new_n682_ & new_n691_;
  assign new_n693_ = new_n686_ & ~new_n689_;
  assign new_n694_ = \p_input[46]  & ~new_n423_;
  assign new_n695_ = \p_input[14]  & new_n423_;
  assign new_n696_ = ~new_n694_ & ~new_n695_;
  assign new_n697_ = \p_input[110]  & ~new_n553_;
  assign new_n698_ = \p_input[78]  & new_n553_;
  assign new_n699_ = ~new_n697_ & ~new_n698_;
  assign new_n700_ = ~new_n696_ & new_n699_;
  assign new_n701_ = ~new_n693_ & ~new_n700_;
  assign new_n702_ = ~new_n692_ & new_n701_;
  assign new_n703_ = \p_input[47]  & ~new_n423_;
  assign new_n704_ = \p_input[15]  & new_n423_;
  assign new_n705_ = ~new_n703_ & ~new_n704_;
  assign new_n706_ = \p_input[111]  & ~new_n553_;
  assign new_n707_ = \p_input[79]  & new_n553_;
  assign new_n708_ = ~new_n706_ & ~new_n707_;
  assign new_n709_ = new_n705_ & ~new_n708_;
  assign new_n710_ = new_n696_ & ~new_n699_;
  assign new_n711_ = ~new_n709_ & ~new_n710_;
  assign new_n712_ = ~new_n702_ & new_n711_;
  assign new_n713_ = \p_input[112]  & ~new_n553_;
  assign new_n714_ = \p_input[80]  & new_n553_;
  assign new_n715_ = ~new_n713_ & ~new_n714_;
  assign new_n716_ = \p_input[48]  & ~new_n423_;
  assign new_n717_ = \p_input[16]  & new_n423_;
  assign new_n718_ = ~new_n716_ & ~new_n717_;
  assign new_n719_ = new_n715_ & ~new_n718_;
  assign new_n720_ = ~new_n705_ & new_n708_;
  assign new_n721_ = ~new_n719_ & ~new_n720_;
  assign new_n722_ = ~new_n712_ & new_n721_;
  assign new_n723_ = ~new_n715_ & new_n718_;
  assign new_n724_ = \p_input[113]  & ~new_n553_;
  assign new_n725_ = \p_input[81]  & new_n553_;
  assign new_n726_ = ~new_n724_ & ~new_n725_;
  assign new_n727_ = \p_input[49]  & ~new_n423_;
  assign new_n728_ = \p_input[17]  & new_n423_;
  assign new_n729_ = ~new_n727_ & ~new_n728_;
  assign new_n730_ = ~new_n726_ & new_n729_;
  assign new_n731_ = ~new_n723_ & ~new_n730_;
  assign new_n732_ = ~new_n722_ & new_n731_;
  assign new_n733_ = new_n726_ & ~new_n729_;
  assign new_n734_ = \p_input[50]  & ~new_n423_;
  assign new_n735_ = \p_input[18]  & new_n423_;
  assign new_n736_ = ~new_n734_ & ~new_n735_;
  assign new_n737_ = \p_input[114]  & ~new_n553_;
  assign new_n738_ = \p_input[82]  & new_n553_;
  assign new_n739_ = ~new_n737_ & ~new_n738_;
  assign new_n740_ = ~new_n736_ & new_n739_;
  assign new_n741_ = ~new_n733_ & ~new_n740_;
  assign new_n742_ = ~new_n732_ & new_n741_;
  assign new_n743_ = \p_input[51]  & ~new_n423_;
  assign new_n744_ = \p_input[19]  & new_n423_;
  assign new_n745_ = ~new_n743_ & ~new_n744_;
  assign new_n746_ = \p_input[115]  & ~new_n553_;
  assign new_n747_ = \p_input[83]  & new_n553_;
  assign new_n748_ = ~new_n746_ & ~new_n747_;
  assign new_n749_ = new_n745_ & ~new_n748_;
  assign new_n750_ = new_n736_ & ~new_n739_;
  assign new_n751_ = ~new_n749_ & ~new_n750_;
  assign new_n752_ = ~new_n742_ & new_n751_;
  assign new_n753_ = \p_input[116]  & ~new_n553_;
  assign new_n754_ = \p_input[84]  & new_n553_;
  assign new_n755_ = ~new_n753_ & ~new_n754_;
  assign new_n756_ = \p_input[52]  & ~new_n423_;
  assign new_n757_ = \p_input[20]  & new_n423_;
  assign new_n758_ = ~new_n756_ & ~new_n757_;
  assign new_n759_ = new_n755_ & ~new_n758_;
  assign new_n760_ = ~new_n745_ & new_n748_;
  assign new_n761_ = ~new_n759_ & ~new_n760_;
  assign new_n762_ = ~new_n752_ & new_n761_;
  assign new_n763_ = ~new_n755_ & new_n758_;
  assign new_n764_ = \p_input[117]  & ~new_n553_;
  assign new_n765_ = \p_input[85]  & new_n553_;
  assign new_n766_ = ~new_n764_ & ~new_n765_;
  assign new_n767_ = \p_input[53]  & ~new_n423_;
  assign new_n768_ = \p_input[21]  & new_n423_;
  assign new_n769_ = ~new_n767_ & ~new_n768_;
  assign new_n770_ = ~new_n766_ & new_n769_;
  assign new_n771_ = ~new_n763_ & ~new_n770_;
  assign new_n772_ = ~new_n762_ & new_n771_;
  assign new_n773_ = new_n766_ & ~new_n769_;
  assign new_n774_ = \p_input[54]  & ~new_n423_;
  assign new_n775_ = \p_input[22]  & new_n423_;
  assign new_n776_ = ~new_n774_ & ~new_n775_;
  assign new_n777_ = \p_input[118]  & ~new_n553_;
  assign new_n778_ = \p_input[86]  & new_n553_;
  assign new_n779_ = ~new_n777_ & ~new_n778_;
  assign new_n780_ = ~new_n776_ & new_n779_;
  assign new_n781_ = ~new_n773_ & ~new_n780_;
  assign new_n782_ = ~new_n772_ & new_n781_;
  assign new_n783_ = \p_input[55]  & ~new_n423_;
  assign new_n784_ = \p_input[23]  & new_n423_;
  assign new_n785_ = ~new_n783_ & ~new_n784_;
  assign new_n786_ = \p_input[119]  & ~new_n553_;
  assign new_n787_ = \p_input[87]  & new_n553_;
  assign new_n788_ = ~new_n786_ & ~new_n787_;
  assign new_n789_ = new_n785_ & ~new_n788_;
  assign new_n790_ = new_n776_ & ~new_n779_;
  assign new_n791_ = ~new_n789_ & ~new_n790_;
  assign new_n792_ = ~new_n782_ & new_n791_;
  assign new_n793_ = \p_input[56]  & ~new_n423_;
  assign new_n794_ = \p_input[24]  & new_n423_;
  assign new_n795_ = ~new_n793_ & ~new_n794_;
  assign new_n796_ = \p_input[120]  & ~new_n553_;
  assign new_n797_ = \p_input[88]  & new_n553_;
  assign new_n798_ = ~new_n796_ & ~new_n797_;
  assign new_n799_ = ~new_n795_ & new_n798_;
  assign new_n800_ = ~new_n785_ & new_n788_;
  assign new_n801_ = ~new_n799_ & ~new_n800_;
  assign new_n802_ = ~new_n792_ & new_n801_;
  assign new_n803_ = new_n795_ & ~new_n798_;
  assign new_n804_ = \p_input[121]  & ~new_n553_;
  assign new_n805_ = \p_input[89]  & new_n553_;
  assign new_n806_ = ~new_n804_ & ~new_n805_;
  assign new_n807_ = \p_input[57]  & ~new_n423_;
  assign new_n808_ = \p_input[25]  & new_n423_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = ~new_n806_ & new_n809_;
  assign new_n811_ = ~new_n803_ & ~new_n810_;
  assign new_n812_ = ~new_n802_ & new_n811_;
  assign new_n813_ = new_n806_ & ~new_n809_;
  assign new_n814_ = \p_input[58]  & ~new_n423_;
  assign new_n815_ = \p_input[26]  & new_n423_;
  assign new_n816_ = ~new_n814_ & ~new_n815_;
  assign new_n817_ = \p_input[122]  & ~new_n553_;
  assign new_n818_ = \p_input[90]  & new_n553_;
  assign new_n819_ = ~new_n817_ & ~new_n818_;
  assign new_n820_ = ~new_n816_ & new_n819_;
  assign new_n821_ = ~new_n813_ & ~new_n820_;
  assign new_n822_ = ~new_n812_ & new_n821_;
  assign new_n823_ = \p_input[59]  & ~new_n423_;
  assign new_n824_ = \p_input[27]  & new_n423_;
  assign new_n825_ = ~new_n823_ & ~new_n824_;
  assign new_n826_ = \p_input[123]  & ~new_n553_;
  assign new_n827_ = \p_input[91]  & new_n553_;
  assign new_n828_ = ~new_n826_ & ~new_n827_;
  assign new_n829_ = new_n825_ & ~new_n828_;
  assign new_n830_ = new_n816_ & ~new_n819_;
  assign new_n831_ = ~new_n829_ & ~new_n830_;
  assign new_n832_ = ~new_n822_ & new_n831_;
  assign new_n833_ = \p_input[124]  & ~new_n553_;
  assign new_n834_ = \p_input[92]  & new_n553_;
  assign new_n835_ = ~new_n833_ & ~new_n834_;
  assign new_n836_ = \p_input[60]  & ~new_n423_;
  assign new_n837_ = \p_input[28]  & new_n423_;
  assign new_n838_ = ~new_n836_ & ~new_n837_;
  assign new_n839_ = new_n835_ & ~new_n838_;
  assign new_n840_ = ~new_n825_ & new_n828_;
  assign new_n841_ = ~new_n839_ & ~new_n840_;
  assign new_n842_ = ~new_n832_ & new_n841_;
  assign new_n843_ = ~new_n835_ & new_n838_;
  assign new_n844_ = \p_input[61]  & ~new_n423_;
  assign new_n845_ = \p_input[29]  & new_n423_;
  assign new_n846_ = ~new_n844_ & ~new_n845_;
  assign new_n847_ = \p_input[125]  & ~new_n553_;
  assign new_n848_ = \p_input[93]  & new_n553_;
  assign new_n849_ = ~new_n847_ & ~new_n848_;
  assign new_n850_ = new_n846_ & ~new_n849_;
  assign new_n851_ = ~new_n843_ & ~new_n850_;
  assign new_n852_ = ~new_n842_ & new_n851_;
  assign new_n853_ = new_n556_ & ~new_n559_;
  assign new_n854_ = ~new_n846_ & new_n849_;
  assign new_n855_ = ~new_n853_ & ~new_n854_;
  assign new_n856_ = ~new_n852_ & new_n855_;
  assign new_n857_ = ~new_n560_ & ~new_n856_;
  assign new_n858_ = ~new_n428_ & ~new_n857_;
  assign new_n859_ = ~new_n427_ & ~new_n858_;
  assign new_n860_ = ~new_n426_ & new_n859_;
  assign new_n861_ = ~new_n563_ & ~new_n859_;
  assign new_n862_ = ~new_n860_ & ~new_n861_;
  assign new_n863_ = ~\p_input[159]  & \p_input[191] ;
  assign new_n864_ = \p_input[159]  & ~\p_input[191] ;
  assign new_n865_ = ~\p_input[158]  & \p_input[190] ;
  assign new_n866_ = \p_input[158]  & ~\p_input[190] ;
  assign new_n867_ = ~\p_input[157]  & \p_input[189] ;
  assign new_n868_ = \p_input[157]  & ~\p_input[189] ;
  assign new_n869_ = ~\p_input[156]  & \p_input[188] ;
  assign new_n870_ = \p_input[156]  & ~\p_input[188] ;
  assign new_n871_ = ~\p_input[155]  & \p_input[187] ;
  assign new_n872_ = \p_input[155]  & ~\p_input[187] ;
  assign new_n873_ = ~\p_input[154]  & \p_input[186] ;
  assign new_n874_ = \p_input[154]  & ~\p_input[186] ;
  assign new_n875_ = ~\p_input[153]  & \p_input[185] ;
  assign new_n876_ = \p_input[153]  & ~\p_input[185] ;
  assign new_n877_ = ~\p_input[152]  & \p_input[184] ;
  assign new_n878_ = \p_input[152]  & ~\p_input[184] ;
  assign new_n879_ = ~\p_input[151]  & \p_input[183] ;
  assign new_n880_ = \p_input[151]  & ~\p_input[183] ;
  assign new_n881_ = ~\p_input[150]  & \p_input[182] ;
  assign new_n882_ = \p_input[150]  & ~\p_input[182] ;
  assign new_n883_ = ~\p_input[149]  & \p_input[181] ;
  assign new_n884_ = \p_input[149]  & ~\p_input[181] ;
  assign new_n885_ = ~\p_input[148]  & \p_input[180] ;
  assign new_n886_ = \p_input[148]  & ~\p_input[180] ;
  assign new_n887_ = ~\p_input[147]  & \p_input[179] ;
  assign new_n888_ = \p_input[147]  & ~\p_input[179] ;
  assign new_n889_ = ~\p_input[146]  & \p_input[178] ;
  assign new_n890_ = \p_input[146]  & ~\p_input[178] ;
  assign new_n891_ = ~\p_input[145]  & \p_input[177] ;
  assign new_n892_ = \p_input[145]  & ~\p_input[177] ;
  assign new_n893_ = ~\p_input[144]  & \p_input[176] ;
  assign new_n894_ = \p_input[144]  & ~\p_input[176] ;
  assign new_n895_ = ~\p_input[143]  & \p_input[175] ;
  assign new_n896_ = \p_input[143]  & ~\p_input[175] ;
  assign new_n897_ = ~\p_input[142]  & \p_input[174] ;
  assign new_n898_ = \p_input[142]  & ~\p_input[174] ;
  assign new_n899_ = ~\p_input[141]  & \p_input[173] ;
  assign new_n900_ = \p_input[141]  & ~\p_input[173] ;
  assign new_n901_ = ~\p_input[140]  & \p_input[172] ;
  assign new_n902_ = \p_input[140]  & ~\p_input[172] ;
  assign new_n903_ = ~\p_input[139]  & \p_input[171] ;
  assign new_n904_ = \p_input[139]  & ~\p_input[171] ;
  assign new_n905_ = ~\p_input[138]  & \p_input[170] ;
  assign new_n906_ = \p_input[138]  & ~\p_input[170] ;
  assign new_n907_ = ~\p_input[137]  & \p_input[169] ;
  assign new_n908_ = \p_input[137]  & ~\p_input[169] ;
  assign new_n909_ = ~\p_input[136]  & \p_input[168] ;
  assign new_n910_ = \p_input[136]  & ~\p_input[168] ;
  assign new_n911_ = ~\p_input[135]  & \p_input[167] ;
  assign new_n912_ = \p_input[135]  & ~\p_input[167] ;
  assign new_n913_ = ~\p_input[134]  & \p_input[166] ;
  assign new_n914_ = \p_input[134]  & ~\p_input[166] ;
  assign new_n915_ = ~\p_input[133]  & \p_input[165] ;
  assign new_n916_ = \p_input[133]  & ~\p_input[165] ;
  assign new_n917_ = ~\p_input[132]  & \p_input[164] ;
  assign new_n918_ = \p_input[132]  & ~\p_input[164] ;
  assign new_n919_ = ~\p_input[131]  & \p_input[163] ;
  assign new_n920_ = \p_input[131]  & ~\p_input[163] ;
  assign new_n921_ = ~\p_input[130]  & \p_input[162] ;
  assign new_n922_ = \p_input[130]  & ~\p_input[162] ;
  assign new_n923_ = ~\p_input[129]  & \p_input[161] ;
  assign new_n924_ = \p_input[129]  & ~\p_input[161] ;
  assign new_n925_ = \p_input[128]  & ~\p_input[160] ;
  assign new_n926_ = ~new_n924_ & ~new_n925_;
  assign new_n927_ = ~new_n923_ & ~new_n926_;
  assign new_n928_ = ~new_n922_ & ~new_n927_;
  assign new_n929_ = ~new_n921_ & ~new_n928_;
  assign new_n930_ = ~new_n920_ & ~new_n929_;
  assign new_n931_ = ~new_n919_ & ~new_n930_;
  assign new_n932_ = ~new_n918_ & ~new_n931_;
  assign new_n933_ = ~new_n917_ & ~new_n932_;
  assign new_n934_ = ~new_n916_ & ~new_n933_;
  assign new_n935_ = ~new_n915_ & ~new_n934_;
  assign new_n936_ = ~new_n914_ & ~new_n935_;
  assign new_n937_ = ~new_n913_ & ~new_n936_;
  assign new_n938_ = ~new_n912_ & ~new_n937_;
  assign new_n939_ = ~new_n911_ & ~new_n938_;
  assign new_n940_ = ~new_n910_ & ~new_n939_;
  assign new_n941_ = ~new_n909_ & ~new_n940_;
  assign new_n942_ = ~new_n908_ & ~new_n941_;
  assign new_n943_ = ~new_n907_ & ~new_n942_;
  assign new_n944_ = ~new_n906_ & ~new_n943_;
  assign new_n945_ = ~new_n905_ & ~new_n944_;
  assign new_n946_ = ~new_n904_ & ~new_n945_;
  assign new_n947_ = ~new_n903_ & ~new_n946_;
  assign new_n948_ = ~new_n902_ & ~new_n947_;
  assign new_n949_ = ~new_n901_ & ~new_n948_;
  assign new_n950_ = ~new_n900_ & ~new_n949_;
  assign new_n951_ = ~new_n899_ & ~new_n950_;
  assign new_n952_ = ~new_n898_ & ~new_n951_;
  assign new_n953_ = ~new_n897_ & ~new_n952_;
  assign new_n954_ = ~new_n896_ & ~new_n953_;
  assign new_n955_ = ~new_n895_ & ~new_n954_;
  assign new_n956_ = ~new_n894_ & ~new_n955_;
  assign new_n957_ = ~new_n893_ & ~new_n956_;
  assign new_n958_ = ~new_n892_ & ~new_n957_;
  assign new_n959_ = ~new_n891_ & ~new_n958_;
  assign new_n960_ = ~new_n890_ & ~new_n959_;
  assign new_n961_ = ~new_n889_ & ~new_n960_;
  assign new_n962_ = ~new_n888_ & ~new_n961_;
  assign new_n963_ = ~new_n887_ & ~new_n962_;
  assign new_n964_ = ~new_n886_ & ~new_n963_;
  assign new_n965_ = ~new_n885_ & ~new_n964_;
  assign new_n966_ = ~new_n884_ & ~new_n965_;
  assign new_n967_ = ~new_n883_ & ~new_n966_;
  assign new_n968_ = ~new_n882_ & ~new_n967_;
  assign new_n969_ = ~new_n881_ & ~new_n968_;
  assign new_n970_ = ~new_n880_ & ~new_n969_;
  assign new_n971_ = ~new_n879_ & ~new_n970_;
  assign new_n972_ = ~new_n878_ & ~new_n971_;
  assign new_n973_ = ~new_n877_ & ~new_n972_;
  assign new_n974_ = ~new_n876_ & ~new_n973_;
  assign new_n975_ = ~new_n875_ & ~new_n974_;
  assign new_n976_ = ~new_n874_ & ~new_n975_;
  assign new_n977_ = ~new_n873_ & ~new_n976_;
  assign new_n978_ = ~new_n872_ & ~new_n977_;
  assign new_n979_ = ~new_n871_ & ~new_n978_;
  assign new_n980_ = ~new_n870_ & ~new_n979_;
  assign new_n981_ = ~new_n869_ & ~new_n980_;
  assign new_n982_ = ~new_n868_ & ~new_n981_;
  assign new_n983_ = ~new_n867_ & ~new_n982_;
  assign new_n984_ = ~new_n866_ & ~new_n983_;
  assign new_n985_ = ~new_n865_ & ~new_n984_;
  assign new_n986_ = ~new_n864_ & ~new_n985_;
  assign new_n987_ = ~new_n863_ & ~new_n986_;
  assign new_n988_ = \p_input[161]  & ~new_n987_;
  assign new_n989_ = \p_input[129]  & new_n987_;
  assign new_n990_ = ~new_n988_ & ~new_n989_;
  assign new_n991_ = new_n292_ & ~new_n293_;
  assign new_n992_ = ~new_n292_ & new_n293_;
  assign new_n993_ = ~\p_input[223]  & \p_input[255] ;
  assign new_n994_ = \p_input[223]  & ~\p_input[255] ;
  assign new_n995_ = ~\p_input[222]  & \p_input[254] ;
  assign new_n996_ = \p_input[222]  & ~\p_input[254] ;
  assign new_n997_ = ~\p_input[221]  & \p_input[253] ;
  assign new_n998_ = \p_input[221]  & ~\p_input[253] ;
  assign new_n999_ = ~\p_input[220]  & \p_input[252] ;
  assign new_n1000_ = \p_input[220]  & ~\p_input[252] ;
  assign new_n1001_ = ~\p_input[219]  & \p_input[251] ;
  assign new_n1002_ = \p_input[219]  & ~\p_input[251] ;
  assign new_n1003_ = ~\p_input[218]  & \p_input[250] ;
  assign new_n1004_ = \p_input[218]  & ~\p_input[250] ;
  assign new_n1005_ = ~\p_input[217]  & \p_input[249] ;
  assign new_n1006_ = \p_input[217]  & ~\p_input[249] ;
  assign new_n1007_ = ~\p_input[216]  & \p_input[248] ;
  assign new_n1008_ = \p_input[216]  & ~\p_input[248] ;
  assign new_n1009_ = ~\p_input[215]  & \p_input[247] ;
  assign new_n1010_ = \p_input[215]  & ~\p_input[247] ;
  assign new_n1011_ = ~\p_input[214]  & \p_input[246] ;
  assign new_n1012_ = \p_input[214]  & ~\p_input[246] ;
  assign new_n1013_ = ~\p_input[213]  & \p_input[245] ;
  assign new_n1014_ = \p_input[213]  & ~\p_input[245] ;
  assign new_n1015_ = ~\p_input[212]  & \p_input[244] ;
  assign new_n1016_ = \p_input[212]  & ~\p_input[244] ;
  assign new_n1017_ = ~\p_input[211]  & \p_input[243] ;
  assign new_n1018_ = \p_input[211]  & ~\p_input[243] ;
  assign new_n1019_ = ~\p_input[210]  & \p_input[242] ;
  assign new_n1020_ = \p_input[210]  & ~\p_input[242] ;
  assign new_n1021_ = ~\p_input[209]  & \p_input[241] ;
  assign new_n1022_ = \p_input[209]  & ~\p_input[241] ;
  assign new_n1023_ = ~\p_input[208]  & \p_input[240] ;
  assign new_n1024_ = \p_input[208]  & ~\p_input[240] ;
  assign new_n1025_ = ~\p_input[207]  & \p_input[239] ;
  assign new_n1026_ = \p_input[207]  & ~\p_input[239] ;
  assign new_n1027_ = ~\p_input[206]  & \p_input[238] ;
  assign new_n1028_ = \p_input[206]  & ~\p_input[238] ;
  assign new_n1029_ = ~\p_input[205]  & \p_input[237] ;
  assign new_n1030_ = \p_input[205]  & ~\p_input[237] ;
  assign new_n1031_ = ~\p_input[204]  & \p_input[236] ;
  assign new_n1032_ = \p_input[204]  & ~\p_input[236] ;
  assign new_n1033_ = ~\p_input[203]  & \p_input[235] ;
  assign new_n1034_ = \p_input[203]  & ~\p_input[235] ;
  assign new_n1035_ = ~\p_input[202]  & \p_input[234] ;
  assign new_n1036_ = \p_input[202]  & ~\p_input[234] ;
  assign new_n1037_ = ~\p_input[201]  & \p_input[233] ;
  assign new_n1038_ = \p_input[201]  & ~\p_input[233] ;
  assign new_n1039_ = ~\p_input[200]  & \p_input[232] ;
  assign new_n1040_ = \p_input[200]  & ~\p_input[232] ;
  assign new_n1041_ = ~\p_input[199]  & \p_input[231] ;
  assign new_n1042_ = \p_input[199]  & ~\p_input[231] ;
  assign new_n1043_ = ~\p_input[198]  & \p_input[230] ;
  assign new_n1044_ = \p_input[198]  & ~\p_input[230] ;
  assign new_n1045_ = ~\p_input[197]  & \p_input[229] ;
  assign new_n1046_ = \p_input[197]  & ~\p_input[229] ;
  assign new_n1047_ = ~\p_input[196]  & \p_input[228] ;
  assign new_n1048_ = \p_input[196]  & ~\p_input[228] ;
  assign new_n1049_ = ~\p_input[195]  & \p_input[227] ;
  assign new_n1050_ = \p_input[195]  & ~\p_input[227] ;
  assign new_n1051_ = ~\p_input[194]  & \p_input[226] ;
  assign new_n1052_ = \p_input[194]  & ~\p_input[226] ;
  assign new_n1053_ = ~\p_input[193]  & \p_input[225] ;
  assign new_n1054_ = \p_input[193]  & ~\p_input[225] ;
  assign new_n1055_ = \p_input[192]  & ~\p_input[224] ;
  assign new_n1056_ = ~new_n1054_ & ~new_n1055_;
  assign new_n1057_ = ~new_n1053_ & ~new_n1056_;
  assign new_n1058_ = ~new_n1052_ & ~new_n1057_;
  assign new_n1059_ = ~new_n1051_ & ~new_n1058_;
  assign new_n1060_ = ~new_n1050_ & ~new_n1059_;
  assign new_n1061_ = ~new_n1049_ & ~new_n1060_;
  assign new_n1062_ = ~new_n1048_ & ~new_n1061_;
  assign new_n1063_ = ~new_n1047_ & ~new_n1062_;
  assign new_n1064_ = ~new_n1046_ & ~new_n1063_;
  assign new_n1065_ = ~new_n1045_ & ~new_n1064_;
  assign new_n1066_ = ~new_n1044_ & ~new_n1065_;
  assign new_n1067_ = ~new_n1043_ & ~new_n1066_;
  assign new_n1068_ = ~new_n1042_ & ~new_n1067_;
  assign new_n1069_ = ~new_n1041_ & ~new_n1068_;
  assign new_n1070_ = ~new_n1040_ & ~new_n1069_;
  assign new_n1071_ = ~new_n1039_ & ~new_n1070_;
  assign new_n1072_ = ~new_n1038_ & ~new_n1071_;
  assign new_n1073_ = ~new_n1037_ & ~new_n1072_;
  assign new_n1074_ = ~new_n1036_ & ~new_n1073_;
  assign new_n1075_ = ~new_n1035_ & ~new_n1074_;
  assign new_n1076_ = ~new_n1034_ & ~new_n1075_;
  assign new_n1077_ = ~new_n1033_ & ~new_n1076_;
  assign new_n1078_ = ~new_n1032_ & ~new_n1077_;
  assign new_n1079_ = ~new_n1031_ & ~new_n1078_;
  assign new_n1080_ = ~new_n1030_ & ~new_n1079_;
  assign new_n1081_ = ~new_n1029_ & ~new_n1080_;
  assign new_n1082_ = ~new_n1028_ & ~new_n1081_;
  assign new_n1083_ = ~new_n1027_ & ~new_n1082_;
  assign new_n1084_ = ~new_n1026_ & ~new_n1083_;
  assign new_n1085_ = ~new_n1025_ & ~new_n1084_;
  assign new_n1086_ = ~new_n1024_ & ~new_n1085_;
  assign new_n1087_ = ~new_n1023_ & ~new_n1086_;
  assign new_n1088_ = ~new_n1022_ & ~new_n1087_;
  assign new_n1089_ = ~new_n1021_ & ~new_n1088_;
  assign new_n1090_ = ~new_n1020_ & ~new_n1089_;
  assign new_n1091_ = ~new_n1019_ & ~new_n1090_;
  assign new_n1092_ = ~new_n1018_ & ~new_n1091_;
  assign new_n1093_ = ~new_n1017_ & ~new_n1092_;
  assign new_n1094_ = ~new_n1016_ & ~new_n1093_;
  assign new_n1095_ = ~new_n1015_ & ~new_n1094_;
  assign new_n1096_ = ~new_n1014_ & ~new_n1095_;
  assign new_n1097_ = ~new_n1013_ & ~new_n1096_;
  assign new_n1098_ = ~new_n1012_ & ~new_n1097_;
  assign new_n1099_ = ~new_n1011_ & ~new_n1098_;
  assign new_n1100_ = ~new_n1010_ & ~new_n1099_;
  assign new_n1101_ = ~new_n1009_ & ~new_n1100_;
  assign new_n1102_ = ~new_n1008_ & ~new_n1101_;
  assign new_n1103_ = ~new_n1007_ & ~new_n1102_;
  assign new_n1104_ = ~new_n1006_ & ~new_n1103_;
  assign new_n1105_ = ~new_n1005_ & ~new_n1104_;
  assign new_n1106_ = ~new_n1004_ & ~new_n1105_;
  assign new_n1107_ = ~new_n1003_ & ~new_n1106_;
  assign new_n1108_ = ~new_n1002_ & ~new_n1107_;
  assign new_n1109_ = ~new_n1001_ & ~new_n1108_;
  assign new_n1110_ = ~new_n1000_ & ~new_n1109_;
  assign new_n1111_ = ~new_n999_ & ~new_n1110_;
  assign new_n1112_ = ~new_n998_ & ~new_n1111_;
  assign new_n1113_ = ~new_n997_ & ~new_n1112_;
  assign new_n1114_ = ~new_n996_ & ~new_n1113_;
  assign new_n1115_ = ~new_n995_ & ~new_n1114_;
  assign new_n1116_ = ~new_n994_ & ~new_n1115_;
  assign new_n1117_ = ~new_n993_ & ~new_n1116_;
  assign new_n1118_ = \p_input[225]  & ~new_n1117_;
  assign new_n1119_ = \p_input[193]  & new_n1117_;
  assign new_n1120_ = ~new_n1118_ & ~new_n1119_;
  assign new_n1121_ = new_n990_ & ~new_n1120_;
  assign new_n1122_ = \p_input[224]  & ~new_n1117_;
  assign new_n1123_ = \p_input[192]  & new_n1117_;
  assign new_n1124_ = ~new_n1122_ & ~new_n1123_;
  assign new_n1125_ = \p_input[160]  & ~new_n987_;
  assign new_n1126_ = \p_input[128]  & new_n987_;
  assign new_n1127_ = ~new_n1125_ & ~new_n1126_;
  assign new_n1128_ = new_n1124_ & ~new_n1127_;
  assign new_n1129_ = ~new_n1121_ & new_n1128_;
  assign new_n1130_ = \p_input[226]  & ~new_n1117_;
  assign new_n1131_ = \p_input[194]  & new_n1117_;
  assign new_n1132_ = ~new_n1130_ & ~new_n1131_;
  assign new_n1133_ = \p_input[162]  & ~new_n987_;
  assign new_n1134_ = \p_input[130]  & new_n987_;
  assign new_n1135_ = ~new_n1133_ & ~new_n1134_;
  assign new_n1136_ = new_n1132_ & ~new_n1135_;
  assign new_n1137_ = ~new_n990_ & new_n1120_;
  assign new_n1138_ = ~new_n1136_ & ~new_n1137_;
  assign new_n1139_ = ~new_n1129_ & new_n1138_;
  assign new_n1140_ = ~new_n1132_ & new_n1135_;
  assign new_n1141_ = \p_input[227]  & ~new_n1117_;
  assign new_n1142_ = \p_input[195]  & new_n1117_;
  assign new_n1143_ = ~new_n1141_ & ~new_n1142_;
  assign new_n1144_ = \p_input[163]  & ~new_n987_;
  assign new_n1145_ = \p_input[131]  & new_n987_;
  assign new_n1146_ = ~new_n1144_ & ~new_n1145_;
  assign new_n1147_ = ~new_n1143_ & new_n1146_;
  assign new_n1148_ = ~new_n1140_ & ~new_n1147_;
  assign new_n1149_ = ~new_n1139_ & new_n1148_;
  assign new_n1150_ = \p_input[164]  & ~new_n987_;
  assign new_n1151_ = \p_input[132]  & new_n987_;
  assign new_n1152_ = ~new_n1150_ & ~new_n1151_;
  assign new_n1153_ = \p_input[228]  & ~new_n1117_;
  assign new_n1154_ = \p_input[196]  & new_n1117_;
  assign new_n1155_ = ~new_n1153_ & ~new_n1154_;
  assign new_n1156_ = ~new_n1152_ & new_n1155_;
  assign new_n1157_ = new_n1143_ & ~new_n1146_;
  assign new_n1158_ = ~new_n1156_ & ~new_n1157_;
  assign new_n1159_ = ~new_n1149_ & new_n1158_;
  assign new_n1160_ = \p_input[229]  & ~new_n1117_;
  assign new_n1161_ = \p_input[197]  & new_n1117_;
  assign new_n1162_ = ~new_n1160_ & ~new_n1161_;
  assign new_n1163_ = \p_input[165]  & ~new_n987_;
  assign new_n1164_ = \p_input[133]  & new_n987_;
  assign new_n1165_ = ~new_n1163_ & ~new_n1164_;
  assign new_n1166_ = ~new_n1162_ & new_n1165_;
  assign new_n1167_ = new_n1152_ & ~new_n1155_;
  assign new_n1168_ = ~new_n1166_ & ~new_n1167_;
  assign new_n1169_ = ~new_n1159_ & new_n1168_;
  assign new_n1170_ = \p_input[230]  & ~new_n1117_;
  assign new_n1171_ = \p_input[198]  & new_n1117_;
  assign new_n1172_ = ~new_n1170_ & ~new_n1171_;
  assign new_n1173_ = \p_input[166]  & ~new_n987_;
  assign new_n1174_ = \p_input[134]  & new_n987_;
  assign new_n1175_ = ~new_n1173_ & ~new_n1174_;
  assign new_n1176_ = new_n1172_ & ~new_n1175_;
  assign new_n1177_ = new_n1162_ & ~new_n1165_;
  assign new_n1178_ = ~new_n1176_ & ~new_n1177_;
  assign new_n1179_ = ~new_n1169_ & new_n1178_;
  assign new_n1180_ = ~new_n1172_ & new_n1175_;
  assign new_n1181_ = \p_input[167]  & ~new_n987_;
  assign new_n1182_ = \p_input[135]  & new_n987_;
  assign new_n1183_ = ~new_n1181_ & ~new_n1182_;
  assign new_n1184_ = \p_input[231]  & ~new_n1117_;
  assign new_n1185_ = \p_input[199]  & new_n1117_;
  assign new_n1186_ = ~new_n1184_ & ~new_n1185_;
  assign new_n1187_ = new_n1183_ & ~new_n1186_;
  assign new_n1188_ = ~new_n1180_ & ~new_n1187_;
  assign new_n1189_ = ~new_n1179_ & new_n1188_;
  assign new_n1190_ = ~new_n1183_ & new_n1186_;
  assign new_n1191_ = \p_input[232]  & ~new_n1117_;
  assign new_n1192_ = \p_input[200]  & new_n1117_;
  assign new_n1193_ = ~new_n1191_ & ~new_n1192_;
  assign new_n1194_ = \p_input[168]  & ~new_n987_;
  assign new_n1195_ = \p_input[136]  & new_n987_;
  assign new_n1196_ = ~new_n1194_ & ~new_n1195_;
  assign new_n1197_ = new_n1193_ & ~new_n1196_;
  assign new_n1198_ = ~new_n1190_ & ~new_n1197_;
  assign new_n1199_ = ~new_n1189_ & new_n1198_;
  assign new_n1200_ = ~new_n1193_ & new_n1196_;
  assign new_n1201_ = \p_input[233]  & ~new_n1117_;
  assign new_n1202_ = \p_input[201]  & new_n1117_;
  assign new_n1203_ = ~new_n1201_ & ~new_n1202_;
  assign new_n1204_ = \p_input[169]  & ~new_n987_;
  assign new_n1205_ = \p_input[137]  & new_n987_;
  assign new_n1206_ = ~new_n1204_ & ~new_n1205_;
  assign new_n1207_ = ~new_n1203_ & new_n1206_;
  assign new_n1208_ = ~new_n1200_ & ~new_n1207_;
  assign new_n1209_ = ~new_n1199_ & new_n1208_;
  assign new_n1210_ = new_n1203_ & ~new_n1206_;
  assign new_n1211_ = \p_input[170]  & ~new_n987_;
  assign new_n1212_ = \p_input[138]  & new_n987_;
  assign new_n1213_ = ~new_n1211_ & ~new_n1212_;
  assign new_n1214_ = \p_input[234]  & ~new_n1117_;
  assign new_n1215_ = \p_input[202]  & new_n1117_;
  assign new_n1216_ = ~new_n1214_ & ~new_n1215_;
  assign new_n1217_ = ~new_n1213_ & new_n1216_;
  assign new_n1218_ = ~new_n1210_ & ~new_n1217_;
  assign new_n1219_ = ~new_n1209_ & new_n1218_;
  assign new_n1220_ = \p_input[171]  & ~new_n987_;
  assign new_n1221_ = \p_input[139]  & new_n987_;
  assign new_n1222_ = ~new_n1220_ & ~new_n1221_;
  assign new_n1223_ = \p_input[235]  & ~new_n1117_;
  assign new_n1224_ = \p_input[203]  & new_n1117_;
  assign new_n1225_ = ~new_n1223_ & ~new_n1224_;
  assign new_n1226_ = new_n1222_ & ~new_n1225_;
  assign new_n1227_ = new_n1213_ & ~new_n1216_;
  assign new_n1228_ = ~new_n1226_ & ~new_n1227_;
  assign new_n1229_ = ~new_n1219_ & new_n1228_;
  assign new_n1230_ = \p_input[236]  & ~new_n1117_;
  assign new_n1231_ = \p_input[204]  & new_n1117_;
  assign new_n1232_ = ~new_n1230_ & ~new_n1231_;
  assign new_n1233_ = \p_input[172]  & ~new_n987_;
  assign new_n1234_ = \p_input[140]  & new_n987_;
  assign new_n1235_ = ~new_n1233_ & ~new_n1234_;
  assign new_n1236_ = new_n1232_ & ~new_n1235_;
  assign new_n1237_ = ~new_n1222_ & new_n1225_;
  assign new_n1238_ = ~new_n1236_ & ~new_n1237_;
  assign new_n1239_ = ~new_n1229_ & new_n1238_;
  assign new_n1240_ = ~new_n1232_ & new_n1235_;
  assign new_n1241_ = \p_input[237]  & ~new_n1117_;
  assign new_n1242_ = \p_input[205]  & new_n1117_;
  assign new_n1243_ = ~new_n1241_ & ~new_n1242_;
  assign new_n1244_ = \p_input[173]  & ~new_n987_;
  assign new_n1245_ = \p_input[141]  & new_n987_;
  assign new_n1246_ = ~new_n1244_ & ~new_n1245_;
  assign new_n1247_ = ~new_n1243_ & new_n1246_;
  assign new_n1248_ = ~new_n1240_ & ~new_n1247_;
  assign new_n1249_ = ~new_n1239_ & new_n1248_;
  assign new_n1250_ = new_n1243_ & ~new_n1246_;
  assign new_n1251_ = \p_input[174]  & ~new_n987_;
  assign new_n1252_ = \p_input[142]  & new_n987_;
  assign new_n1253_ = ~new_n1251_ & ~new_n1252_;
  assign new_n1254_ = \p_input[238]  & ~new_n1117_;
  assign new_n1255_ = \p_input[206]  & new_n1117_;
  assign new_n1256_ = ~new_n1254_ & ~new_n1255_;
  assign new_n1257_ = ~new_n1253_ & new_n1256_;
  assign new_n1258_ = ~new_n1250_ & ~new_n1257_;
  assign new_n1259_ = ~new_n1249_ & new_n1258_;
  assign new_n1260_ = \p_input[175]  & ~new_n987_;
  assign new_n1261_ = \p_input[143]  & new_n987_;
  assign new_n1262_ = ~new_n1260_ & ~new_n1261_;
  assign new_n1263_ = \p_input[239]  & ~new_n1117_;
  assign new_n1264_ = \p_input[207]  & new_n1117_;
  assign new_n1265_ = ~new_n1263_ & ~new_n1264_;
  assign new_n1266_ = new_n1262_ & ~new_n1265_;
  assign new_n1267_ = new_n1253_ & ~new_n1256_;
  assign new_n1268_ = ~new_n1266_ & ~new_n1267_;
  assign new_n1269_ = ~new_n1259_ & new_n1268_;
  assign new_n1270_ = \p_input[240]  & ~new_n1117_;
  assign new_n1271_ = \p_input[208]  & new_n1117_;
  assign new_n1272_ = ~new_n1270_ & ~new_n1271_;
  assign new_n1273_ = \p_input[176]  & ~new_n987_;
  assign new_n1274_ = \p_input[144]  & new_n987_;
  assign new_n1275_ = ~new_n1273_ & ~new_n1274_;
  assign new_n1276_ = new_n1272_ & ~new_n1275_;
  assign new_n1277_ = ~new_n1262_ & new_n1265_;
  assign new_n1278_ = ~new_n1276_ & ~new_n1277_;
  assign new_n1279_ = ~new_n1269_ & new_n1278_;
  assign new_n1280_ = ~new_n1272_ & new_n1275_;
  assign new_n1281_ = \p_input[241]  & ~new_n1117_;
  assign new_n1282_ = \p_input[209]  & new_n1117_;
  assign new_n1283_ = ~new_n1281_ & ~new_n1282_;
  assign new_n1284_ = \p_input[177]  & ~new_n987_;
  assign new_n1285_ = \p_input[145]  & new_n987_;
  assign new_n1286_ = ~new_n1284_ & ~new_n1285_;
  assign new_n1287_ = ~new_n1283_ & new_n1286_;
  assign new_n1288_ = ~new_n1280_ & ~new_n1287_;
  assign new_n1289_ = ~new_n1279_ & new_n1288_;
  assign new_n1290_ = new_n1283_ & ~new_n1286_;
  assign new_n1291_ = \p_input[178]  & ~new_n987_;
  assign new_n1292_ = \p_input[146]  & new_n987_;
  assign new_n1293_ = ~new_n1291_ & ~new_n1292_;
  assign new_n1294_ = \p_input[242]  & ~new_n1117_;
  assign new_n1295_ = \p_input[210]  & new_n1117_;
  assign new_n1296_ = ~new_n1294_ & ~new_n1295_;
  assign new_n1297_ = ~new_n1293_ & new_n1296_;
  assign new_n1298_ = ~new_n1290_ & ~new_n1297_;
  assign new_n1299_ = ~new_n1289_ & new_n1298_;
  assign new_n1300_ = \p_input[179]  & ~new_n987_;
  assign new_n1301_ = \p_input[147]  & new_n987_;
  assign new_n1302_ = ~new_n1300_ & ~new_n1301_;
  assign new_n1303_ = \p_input[243]  & ~new_n1117_;
  assign new_n1304_ = \p_input[211]  & new_n1117_;
  assign new_n1305_ = ~new_n1303_ & ~new_n1304_;
  assign new_n1306_ = new_n1302_ & ~new_n1305_;
  assign new_n1307_ = new_n1293_ & ~new_n1296_;
  assign new_n1308_ = ~new_n1306_ & ~new_n1307_;
  assign new_n1309_ = ~new_n1299_ & new_n1308_;
  assign new_n1310_ = \p_input[244]  & ~new_n1117_;
  assign new_n1311_ = \p_input[212]  & new_n1117_;
  assign new_n1312_ = ~new_n1310_ & ~new_n1311_;
  assign new_n1313_ = \p_input[180]  & ~new_n987_;
  assign new_n1314_ = \p_input[148]  & new_n987_;
  assign new_n1315_ = ~new_n1313_ & ~new_n1314_;
  assign new_n1316_ = new_n1312_ & ~new_n1315_;
  assign new_n1317_ = ~new_n1302_ & new_n1305_;
  assign new_n1318_ = ~new_n1316_ & ~new_n1317_;
  assign new_n1319_ = ~new_n1309_ & new_n1318_;
  assign new_n1320_ = ~new_n1312_ & new_n1315_;
  assign new_n1321_ = \p_input[245]  & ~new_n1117_;
  assign new_n1322_ = \p_input[213]  & new_n1117_;
  assign new_n1323_ = ~new_n1321_ & ~new_n1322_;
  assign new_n1324_ = \p_input[181]  & ~new_n987_;
  assign new_n1325_ = \p_input[149]  & new_n987_;
  assign new_n1326_ = ~new_n1324_ & ~new_n1325_;
  assign new_n1327_ = ~new_n1323_ & new_n1326_;
  assign new_n1328_ = ~new_n1320_ & ~new_n1327_;
  assign new_n1329_ = ~new_n1319_ & new_n1328_;
  assign new_n1330_ = new_n1323_ & ~new_n1326_;
  assign new_n1331_ = \p_input[182]  & ~new_n987_;
  assign new_n1332_ = \p_input[150]  & new_n987_;
  assign new_n1333_ = ~new_n1331_ & ~new_n1332_;
  assign new_n1334_ = \p_input[246]  & ~new_n1117_;
  assign new_n1335_ = \p_input[214]  & new_n1117_;
  assign new_n1336_ = ~new_n1334_ & ~new_n1335_;
  assign new_n1337_ = ~new_n1333_ & new_n1336_;
  assign new_n1338_ = ~new_n1330_ & ~new_n1337_;
  assign new_n1339_ = ~new_n1329_ & new_n1338_;
  assign new_n1340_ = \p_input[183]  & ~new_n987_;
  assign new_n1341_ = \p_input[151]  & new_n987_;
  assign new_n1342_ = ~new_n1340_ & ~new_n1341_;
  assign new_n1343_ = \p_input[247]  & ~new_n1117_;
  assign new_n1344_ = \p_input[215]  & new_n1117_;
  assign new_n1345_ = ~new_n1343_ & ~new_n1344_;
  assign new_n1346_ = new_n1342_ & ~new_n1345_;
  assign new_n1347_ = new_n1333_ & ~new_n1336_;
  assign new_n1348_ = ~new_n1346_ & ~new_n1347_;
  assign new_n1349_ = ~new_n1339_ & new_n1348_;
  assign new_n1350_ = \p_input[248]  & ~new_n1117_;
  assign new_n1351_ = \p_input[216]  & new_n1117_;
  assign new_n1352_ = ~new_n1350_ & ~new_n1351_;
  assign new_n1353_ = \p_input[184]  & ~new_n987_;
  assign new_n1354_ = \p_input[152]  & new_n987_;
  assign new_n1355_ = ~new_n1353_ & ~new_n1354_;
  assign new_n1356_ = new_n1352_ & ~new_n1355_;
  assign new_n1357_ = ~new_n1342_ & new_n1345_;
  assign new_n1358_ = ~new_n1356_ & ~new_n1357_;
  assign new_n1359_ = ~new_n1349_ & new_n1358_;
  assign new_n1360_ = ~new_n1352_ & new_n1355_;
  assign new_n1361_ = \p_input[249]  & ~new_n1117_;
  assign new_n1362_ = \p_input[217]  & new_n1117_;
  assign new_n1363_ = ~new_n1361_ & ~new_n1362_;
  assign new_n1364_ = \p_input[185]  & ~new_n987_;
  assign new_n1365_ = \p_input[153]  & new_n987_;
  assign new_n1366_ = ~new_n1364_ & ~new_n1365_;
  assign new_n1367_ = ~new_n1363_ & new_n1366_;
  assign new_n1368_ = ~new_n1360_ & ~new_n1367_;
  assign new_n1369_ = ~new_n1359_ & new_n1368_;
  assign new_n1370_ = new_n1363_ & ~new_n1366_;
  assign new_n1371_ = \p_input[186]  & ~new_n987_;
  assign new_n1372_ = \p_input[154]  & new_n987_;
  assign new_n1373_ = ~new_n1371_ & ~new_n1372_;
  assign new_n1374_ = \p_input[250]  & ~new_n1117_;
  assign new_n1375_ = \p_input[218]  & new_n1117_;
  assign new_n1376_ = ~new_n1374_ & ~new_n1375_;
  assign new_n1377_ = ~new_n1373_ & new_n1376_;
  assign new_n1378_ = ~new_n1370_ & ~new_n1377_;
  assign new_n1379_ = ~new_n1369_ & new_n1378_;
  assign new_n1380_ = \p_input[251]  & ~new_n1117_;
  assign new_n1381_ = \p_input[219]  & new_n1117_;
  assign new_n1382_ = ~new_n1380_ & ~new_n1381_;
  assign new_n1383_ = \p_input[187]  & ~new_n987_;
  assign new_n1384_ = \p_input[155]  & new_n987_;
  assign new_n1385_ = ~new_n1383_ & ~new_n1384_;
  assign new_n1386_ = ~new_n1382_ & new_n1385_;
  assign new_n1387_ = new_n1373_ & ~new_n1376_;
  assign new_n1388_ = ~new_n1386_ & ~new_n1387_;
  assign new_n1389_ = ~new_n1379_ & new_n1388_;
  assign new_n1390_ = \p_input[188]  & ~new_n987_;
  assign new_n1391_ = \p_input[156]  & new_n987_;
  assign new_n1392_ = ~new_n1390_ & ~new_n1391_;
  assign new_n1393_ = \p_input[252]  & ~new_n1117_;
  assign new_n1394_ = \p_input[220]  & new_n1117_;
  assign new_n1395_ = ~new_n1393_ & ~new_n1394_;
  assign new_n1396_ = ~new_n1392_ & new_n1395_;
  assign new_n1397_ = new_n1382_ & ~new_n1385_;
  assign new_n1398_ = ~new_n1396_ & ~new_n1397_;
  assign new_n1399_ = ~new_n1389_ & new_n1398_;
  assign new_n1400_ = new_n1392_ & ~new_n1395_;
  assign new_n1401_ = \p_input[189]  & ~new_n987_;
  assign new_n1402_ = \p_input[157]  & new_n987_;
  assign new_n1403_ = ~new_n1401_ & ~new_n1402_;
  assign new_n1404_ = \p_input[253]  & ~new_n1117_;
  assign new_n1405_ = \p_input[221]  & new_n1117_;
  assign new_n1406_ = ~new_n1404_ & ~new_n1405_;
  assign new_n1407_ = new_n1403_ & ~new_n1406_;
  assign new_n1408_ = ~new_n1400_ & ~new_n1407_;
  assign new_n1409_ = ~new_n1399_ & new_n1408_;
  assign new_n1410_ = ~new_n1403_ & new_n1406_;
  assign new_n1411_ = \p_input[190]  & ~new_n987_;
  assign new_n1412_ = \p_input[158]  & new_n987_;
  assign new_n1413_ = ~new_n1411_ & ~new_n1412_;
  assign new_n1414_ = \p_input[254]  & ~new_n1117_;
  assign new_n1415_ = \p_input[222]  & new_n1117_;
  assign new_n1416_ = ~new_n1414_ & ~new_n1415_;
  assign new_n1417_ = ~new_n1413_ & new_n1416_;
  assign new_n1418_ = ~new_n1410_ & ~new_n1417_;
  assign new_n1419_ = ~new_n1409_ & new_n1418_;
  assign new_n1420_ = new_n1413_ & ~new_n1416_;
  assign new_n1421_ = ~new_n1419_ & ~new_n1420_;
  assign new_n1422_ = ~new_n992_ & ~new_n1421_;
  assign new_n1423_ = ~new_n991_ & ~new_n1422_;
  assign new_n1424_ = ~new_n990_ & new_n1423_;
  assign new_n1425_ = ~new_n1120_ & ~new_n1423_;
  assign new_n1426_ = ~new_n1424_ & ~new_n1425_;
  assign new_n1427_ = new_n862_ & ~new_n1426_;
  assign new_n1428_ = ~new_n1127_ & new_n1423_;
  assign new_n1429_ = ~new_n1124_ & ~new_n1423_;
  assign new_n1430_ = ~new_n1428_ & ~new_n1429_;
  assign new_n1431_ = ~new_n570_ & new_n859_;
  assign new_n1432_ = ~new_n567_ & ~new_n859_;
  assign new_n1433_ = ~new_n1431_ & ~new_n1432_;
  assign new_n1434_ = new_n1430_ & ~new_n1433_;
  assign new_n1435_ = ~new_n1427_ & new_n1434_;
  assign new_n1436_ = ~new_n1135_ & new_n1423_;
  assign new_n1437_ = ~new_n1132_ & ~new_n1423_;
  assign new_n1438_ = ~new_n1436_ & ~new_n1437_;
  assign new_n1439_ = ~new_n578_ & new_n859_;
  assign new_n1440_ = ~new_n575_ & ~new_n859_;
  assign new_n1441_ = ~new_n1439_ & ~new_n1440_;
  assign new_n1442_ = new_n1438_ & ~new_n1441_;
  assign new_n1443_ = ~new_n862_ & new_n1426_;
  assign new_n1444_ = ~new_n1442_ & ~new_n1443_;
  assign new_n1445_ = ~new_n1435_ & new_n1444_;
  assign new_n1446_ = ~new_n1438_ & new_n1441_;
  assign new_n1447_ = ~new_n585_ & new_n859_;
  assign new_n1448_ = ~new_n588_ & ~new_n859_;
  assign new_n1449_ = ~new_n1447_ & ~new_n1448_;
  assign new_n1450_ = ~new_n1146_ & new_n1423_;
  assign new_n1451_ = ~new_n1143_ & ~new_n1423_;
  assign new_n1452_ = ~new_n1450_ & ~new_n1451_;
  assign new_n1453_ = new_n1449_ & ~new_n1452_;
  assign new_n1454_ = ~new_n1446_ & ~new_n1453_;
  assign new_n1455_ = ~new_n1445_ & new_n1454_;
  assign new_n1456_ = ~new_n1152_ & new_n1423_;
  assign new_n1457_ = ~new_n1155_ & ~new_n1423_;
  assign new_n1458_ = ~new_n1456_ & ~new_n1457_;
  assign new_n1459_ = ~new_n598_ & new_n859_;
  assign new_n1460_ = ~new_n595_ & ~new_n859_;
  assign new_n1461_ = ~new_n1459_ & ~new_n1460_;
  assign new_n1462_ = new_n1458_ & ~new_n1461_;
  assign new_n1463_ = ~new_n1449_ & new_n1452_;
  assign new_n1464_ = ~new_n1462_ & ~new_n1463_;
  assign new_n1465_ = ~new_n1455_ & new_n1464_;
  assign new_n1466_ = ~new_n608_ & new_n859_;
  assign new_n1467_ = ~new_n605_ & ~new_n859_;
  assign new_n1468_ = ~new_n1466_ & ~new_n1467_;
  assign new_n1469_ = ~new_n1165_ & new_n1423_;
  assign new_n1470_ = ~new_n1162_ & ~new_n1423_;
  assign new_n1471_ = ~new_n1469_ & ~new_n1470_;
  assign new_n1472_ = new_n1468_ & ~new_n1471_;
  assign new_n1473_ = ~new_n1458_ & new_n1461_;
  assign new_n1474_ = ~new_n1472_ & ~new_n1473_;
  assign new_n1475_ = ~new_n1465_ & new_n1474_;
  assign new_n1476_ = ~new_n615_ & new_n859_;
  assign new_n1477_ = ~new_n618_ & ~new_n859_;
  assign new_n1478_ = ~new_n1476_ & ~new_n1477_;
  assign new_n1479_ = ~new_n1175_ & new_n1423_;
  assign new_n1480_ = ~new_n1172_ & ~new_n1423_;
  assign new_n1481_ = ~new_n1479_ & ~new_n1480_;
  assign new_n1482_ = ~new_n1478_ & new_n1481_;
  assign new_n1483_ = ~new_n1468_ & new_n1471_;
  assign new_n1484_ = ~new_n1482_ & ~new_n1483_;
  assign new_n1485_ = ~new_n1475_ & new_n1484_;
  assign new_n1486_ = ~new_n625_ & new_n859_;
  assign new_n1487_ = ~new_n628_ & ~new_n859_;
  assign new_n1488_ = ~new_n1486_ & ~new_n1487_;
  assign new_n1489_ = ~new_n1183_ & new_n1423_;
  assign new_n1490_ = ~new_n1186_ & ~new_n1423_;
  assign new_n1491_ = ~new_n1489_ & ~new_n1490_;
  assign new_n1492_ = new_n1488_ & ~new_n1491_;
  assign new_n1493_ = new_n1478_ & ~new_n1481_;
  assign new_n1494_ = ~new_n1492_ & ~new_n1493_;
  assign new_n1495_ = ~new_n1485_ & new_n1494_;
  assign new_n1496_ = ~new_n1196_ & new_n1423_;
  assign new_n1497_ = ~new_n1193_ & ~new_n1423_;
  assign new_n1498_ = ~new_n1496_ & ~new_n1497_;
  assign new_n1499_ = ~new_n639_ & new_n859_;
  assign new_n1500_ = ~new_n636_ & ~new_n859_;
  assign new_n1501_ = ~new_n1499_ & ~new_n1500_;
  assign new_n1502_ = new_n1498_ & ~new_n1501_;
  assign new_n1503_ = ~new_n1488_ & new_n1491_;
  assign new_n1504_ = ~new_n1502_ & ~new_n1503_;
  assign new_n1505_ = ~new_n1495_ & new_n1504_;
  assign new_n1506_ = ~new_n649_ & new_n859_;
  assign new_n1507_ = ~new_n646_ & ~new_n859_;
  assign new_n1508_ = ~new_n1506_ & ~new_n1507_;
  assign new_n1509_ = ~new_n1206_ & new_n1423_;
  assign new_n1510_ = ~new_n1203_ & ~new_n1423_;
  assign new_n1511_ = ~new_n1509_ & ~new_n1510_;
  assign new_n1512_ = new_n1508_ & ~new_n1511_;
  assign new_n1513_ = ~new_n1498_ & new_n1501_;
  assign new_n1514_ = ~new_n1512_ & ~new_n1513_;
  assign new_n1515_ = ~new_n1505_ & new_n1514_;
  assign new_n1516_ = ~new_n1213_ & new_n1423_;
  assign new_n1517_ = ~new_n1216_ & ~new_n1423_;
  assign new_n1518_ = ~new_n1516_ & ~new_n1517_;
  assign new_n1519_ = ~new_n656_ & new_n859_;
  assign new_n1520_ = ~new_n659_ & ~new_n859_;
  assign new_n1521_ = ~new_n1519_ & ~new_n1520_;
  assign new_n1522_ = new_n1518_ & ~new_n1521_;
  assign new_n1523_ = ~new_n1508_ & new_n1511_;
  assign new_n1524_ = ~new_n1522_ & ~new_n1523_;
  assign new_n1525_ = ~new_n1515_ & new_n1524_;
  assign new_n1526_ = ~new_n665_ & new_n859_;
  assign new_n1527_ = ~new_n668_ & ~new_n859_;
  assign new_n1528_ = ~new_n1526_ & ~new_n1527_;
  assign new_n1529_ = ~new_n1222_ & new_n1423_;
  assign new_n1530_ = ~new_n1225_ & ~new_n1423_;
  assign new_n1531_ = ~new_n1529_ & ~new_n1530_;
  assign new_n1532_ = new_n1528_ & ~new_n1531_;
  assign new_n1533_ = ~new_n1518_ & new_n1521_;
  assign new_n1534_ = ~new_n1532_ & ~new_n1533_;
  assign new_n1535_ = ~new_n1525_ & new_n1534_;
  assign new_n1536_ = ~new_n1235_ & new_n1423_;
  assign new_n1537_ = ~new_n1232_ & ~new_n1423_;
  assign new_n1538_ = ~new_n1536_ & ~new_n1537_;
  assign new_n1539_ = ~new_n678_ & new_n859_;
  assign new_n1540_ = ~new_n675_ & ~new_n859_;
  assign new_n1541_ = ~new_n1539_ & ~new_n1540_;
  assign new_n1542_ = new_n1538_ & ~new_n1541_;
  assign new_n1543_ = ~new_n1528_ & new_n1531_;
  assign new_n1544_ = ~new_n1542_ & ~new_n1543_;
  assign new_n1545_ = ~new_n1535_ & new_n1544_;
  assign new_n1546_ = ~new_n689_ & new_n859_;
  assign new_n1547_ = ~new_n686_ & ~new_n859_;
  assign new_n1548_ = ~new_n1546_ & ~new_n1547_;
  assign new_n1549_ = ~new_n1246_ & new_n1423_;
  assign new_n1550_ = ~new_n1243_ & ~new_n1423_;
  assign new_n1551_ = ~new_n1549_ & ~new_n1550_;
  assign new_n1552_ = new_n1548_ & ~new_n1551_;
  assign new_n1553_ = ~new_n1538_ & new_n1541_;
  assign new_n1554_ = ~new_n1552_ & ~new_n1553_;
  assign new_n1555_ = ~new_n1545_ & new_n1554_;
  assign new_n1556_ = ~new_n1253_ & new_n1423_;
  assign new_n1557_ = ~new_n1256_ & ~new_n1423_;
  assign new_n1558_ = ~new_n1556_ & ~new_n1557_;
  assign new_n1559_ = ~new_n696_ & new_n859_;
  assign new_n1560_ = ~new_n699_ & ~new_n859_;
  assign new_n1561_ = ~new_n1559_ & ~new_n1560_;
  assign new_n1562_ = new_n1558_ & ~new_n1561_;
  assign new_n1563_ = ~new_n1548_ & new_n1551_;
  assign new_n1564_ = ~new_n1562_ & ~new_n1563_;
  assign new_n1565_ = ~new_n1555_ & new_n1564_;
  assign new_n1566_ = ~new_n705_ & new_n859_;
  assign new_n1567_ = ~new_n708_ & ~new_n859_;
  assign new_n1568_ = ~new_n1566_ & ~new_n1567_;
  assign new_n1569_ = ~new_n1262_ & new_n1423_;
  assign new_n1570_ = ~new_n1265_ & ~new_n1423_;
  assign new_n1571_ = ~new_n1569_ & ~new_n1570_;
  assign new_n1572_ = new_n1568_ & ~new_n1571_;
  assign new_n1573_ = ~new_n1558_ & new_n1561_;
  assign new_n1574_ = ~new_n1572_ & ~new_n1573_;
  assign new_n1575_ = ~new_n1565_ & new_n1574_;
  assign new_n1576_ = ~new_n1275_ & new_n1423_;
  assign new_n1577_ = ~new_n1272_ & ~new_n1423_;
  assign new_n1578_ = ~new_n1576_ & ~new_n1577_;
  assign new_n1579_ = ~new_n718_ & new_n859_;
  assign new_n1580_ = ~new_n715_ & ~new_n859_;
  assign new_n1581_ = ~new_n1579_ & ~new_n1580_;
  assign new_n1582_ = new_n1578_ & ~new_n1581_;
  assign new_n1583_ = ~new_n1568_ & new_n1571_;
  assign new_n1584_ = ~new_n1582_ & ~new_n1583_;
  assign new_n1585_ = ~new_n1575_ & new_n1584_;
  assign new_n1586_ = ~new_n729_ & new_n859_;
  assign new_n1587_ = ~new_n726_ & ~new_n859_;
  assign new_n1588_ = ~new_n1586_ & ~new_n1587_;
  assign new_n1589_ = ~new_n1286_ & new_n1423_;
  assign new_n1590_ = ~new_n1283_ & ~new_n1423_;
  assign new_n1591_ = ~new_n1589_ & ~new_n1590_;
  assign new_n1592_ = new_n1588_ & ~new_n1591_;
  assign new_n1593_ = ~new_n1578_ & new_n1581_;
  assign new_n1594_ = ~new_n1592_ & ~new_n1593_;
  assign new_n1595_ = ~new_n1585_ & new_n1594_;
  assign new_n1596_ = ~new_n1293_ & new_n1423_;
  assign new_n1597_ = ~new_n1296_ & ~new_n1423_;
  assign new_n1598_ = ~new_n1596_ & ~new_n1597_;
  assign new_n1599_ = ~new_n736_ & new_n859_;
  assign new_n1600_ = ~new_n739_ & ~new_n859_;
  assign new_n1601_ = ~new_n1599_ & ~new_n1600_;
  assign new_n1602_ = new_n1598_ & ~new_n1601_;
  assign new_n1603_ = ~new_n1588_ & new_n1591_;
  assign new_n1604_ = ~new_n1602_ & ~new_n1603_;
  assign new_n1605_ = ~new_n1595_ & new_n1604_;
  assign new_n1606_ = ~new_n745_ & new_n859_;
  assign new_n1607_ = ~new_n748_ & ~new_n859_;
  assign new_n1608_ = ~new_n1606_ & ~new_n1607_;
  assign new_n1609_ = ~new_n1302_ & new_n1423_;
  assign new_n1610_ = ~new_n1305_ & ~new_n1423_;
  assign new_n1611_ = ~new_n1609_ & ~new_n1610_;
  assign new_n1612_ = new_n1608_ & ~new_n1611_;
  assign new_n1613_ = ~new_n1598_ & new_n1601_;
  assign new_n1614_ = ~new_n1612_ & ~new_n1613_;
  assign new_n1615_ = ~new_n1605_ & new_n1614_;
  assign new_n1616_ = ~new_n1315_ & new_n1423_;
  assign new_n1617_ = ~new_n1312_ & ~new_n1423_;
  assign new_n1618_ = ~new_n1616_ & ~new_n1617_;
  assign new_n1619_ = ~new_n758_ & new_n859_;
  assign new_n1620_ = ~new_n755_ & ~new_n859_;
  assign new_n1621_ = ~new_n1619_ & ~new_n1620_;
  assign new_n1622_ = new_n1618_ & ~new_n1621_;
  assign new_n1623_ = ~new_n1608_ & new_n1611_;
  assign new_n1624_ = ~new_n1622_ & ~new_n1623_;
  assign new_n1625_ = ~new_n1615_ & new_n1624_;
  assign new_n1626_ = ~new_n769_ & new_n859_;
  assign new_n1627_ = ~new_n766_ & ~new_n859_;
  assign new_n1628_ = ~new_n1626_ & ~new_n1627_;
  assign new_n1629_ = ~new_n1326_ & new_n1423_;
  assign new_n1630_ = ~new_n1323_ & ~new_n1423_;
  assign new_n1631_ = ~new_n1629_ & ~new_n1630_;
  assign new_n1632_ = new_n1628_ & ~new_n1631_;
  assign new_n1633_ = ~new_n1618_ & new_n1621_;
  assign new_n1634_ = ~new_n1632_ & ~new_n1633_;
  assign new_n1635_ = ~new_n1625_ & new_n1634_;
  assign new_n1636_ = ~new_n1333_ & new_n1423_;
  assign new_n1637_ = ~new_n1336_ & ~new_n1423_;
  assign new_n1638_ = ~new_n1636_ & ~new_n1637_;
  assign new_n1639_ = ~new_n776_ & new_n859_;
  assign new_n1640_ = ~new_n779_ & ~new_n859_;
  assign new_n1641_ = ~new_n1639_ & ~new_n1640_;
  assign new_n1642_ = new_n1638_ & ~new_n1641_;
  assign new_n1643_ = ~new_n1628_ & new_n1631_;
  assign new_n1644_ = ~new_n1642_ & ~new_n1643_;
  assign new_n1645_ = ~new_n1635_ & new_n1644_;
  assign new_n1646_ = ~new_n785_ & new_n859_;
  assign new_n1647_ = ~new_n788_ & ~new_n859_;
  assign new_n1648_ = ~new_n1646_ & ~new_n1647_;
  assign new_n1649_ = ~new_n1342_ & new_n1423_;
  assign new_n1650_ = ~new_n1345_ & ~new_n1423_;
  assign new_n1651_ = ~new_n1649_ & ~new_n1650_;
  assign new_n1652_ = new_n1648_ & ~new_n1651_;
  assign new_n1653_ = ~new_n1638_ & new_n1641_;
  assign new_n1654_ = ~new_n1652_ & ~new_n1653_;
  assign new_n1655_ = ~new_n1645_ & new_n1654_;
  assign new_n1656_ = ~new_n795_ & new_n859_;
  assign new_n1657_ = ~new_n798_ & ~new_n859_;
  assign new_n1658_ = ~new_n1656_ & ~new_n1657_;
  assign new_n1659_ = ~new_n1355_ & new_n1423_;
  assign new_n1660_ = ~new_n1352_ & ~new_n1423_;
  assign new_n1661_ = ~new_n1659_ & ~new_n1660_;
  assign new_n1662_ = ~new_n1658_ & new_n1661_;
  assign new_n1663_ = ~new_n1648_ & new_n1651_;
  assign new_n1664_ = ~new_n1662_ & ~new_n1663_;
  assign new_n1665_ = ~new_n1655_ & new_n1664_;
  assign new_n1666_ = ~new_n809_ & new_n859_;
  assign new_n1667_ = ~new_n806_ & ~new_n859_;
  assign new_n1668_ = ~new_n1666_ & ~new_n1667_;
  assign new_n1669_ = ~new_n1366_ & new_n1423_;
  assign new_n1670_ = ~new_n1363_ & ~new_n1423_;
  assign new_n1671_ = ~new_n1669_ & ~new_n1670_;
  assign new_n1672_ = new_n1668_ & ~new_n1671_;
  assign new_n1673_ = new_n1658_ & ~new_n1661_;
  assign new_n1674_ = ~new_n1672_ & ~new_n1673_;
  assign new_n1675_ = ~new_n1665_ & new_n1674_;
  assign new_n1676_ = ~new_n1373_ & new_n1423_;
  assign new_n1677_ = ~new_n1376_ & ~new_n1423_;
  assign new_n1678_ = ~new_n1676_ & ~new_n1677_;
  assign new_n1679_ = ~new_n816_ & new_n859_;
  assign new_n1680_ = ~new_n819_ & ~new_n859_;
  assign new_n1681_ = ~new_n1679_ & ~new_n1680_;
  assign new_n1682_ = new_n1678_ & ~new_n1681_;
  assign new_n1683_ = ~new_n1668_ & new_n1671_;
  assign new_n1684_ = ~new_n1682_ & ~new_n1683_;
  assign new_n1685_ = ~new_n1675_ & new_n1684_;
  assign new_n1686_ = ~new_n1678_ & new_n1681_;
  assign new_n1687_ = ~new_n825_ & new_n859_;
  assign new_n1688_ = ~new_n828_ & ~new_n859_;
  assign new_n1689_ = ~new_n1687_ & ~new_n1688_;
  assign new_n1690_ = ~new_n1385_ & new_n1423_;
  assign new_n1691_ = ~new_n1382_ & ~new_n1423_;
  assign new_n1692_ = ~new_n1690_ & ~new_n1691_;
  assign new_n1693_ = new_n1689_ & ~new_n1692_;
  assign new_n1694_ = ~new_n1686_ & ~new_n1693_;
  assign new_n1695_ = ~new_n1685_ & new_n1694_;
  assign new_n1696_ = ~new_n1689_ & new_n1692_;
  assign new_n1697_ = ~new_n1392_ & new_n1423_;
  assign new_n1698_ = ~new_n1395_ & ~new_n1423_;
  assign new_n1699_ = ~new_n1697_ & ~new_n1698_;
  assign new_n1700_ = ~new_n838_ & new_n859_;
  assign new_n1701_ = ~new_n835_ & ~new_n859_;
  assign new_n1702_ = ~new_n1700_ & ~new_n1701_;
  assign new_n1703_ = new_n1699_ & ~new_n1702_;
  assign new_n1704_ = ~new_n1696_ & ~new_n1703_;
  assign new_n1705_ = ~new_n1695_ & new_n1704_;
  assign new_n1706_ = ~new_n1699_ & new_n1702_;
  assign new_n1707_ = ~new_n1403_ & new_n1423_;
  assign new_n1708_ = ~new_n1406_ & ~new_n1423_;
  assign new_n1709_ = ~new_n1707_ & ~new_n1708_;
  assign new_n1710_ = ~new_n846_ & new_n859_;
  assign new_n1711_ = ~new_n849_ & ~new_n859_;
  assign new_n1712_ = ~new_n1710_ & ~new_n1711_;
  assign new_n1713_ = ~new_n1709_ & new_n1712_;
  assign new_n1714_ = ~new_n1706_ & ~new_n1713_;
  assign new_n1715_ = ~new_n1705_ & new_n1714_;
  assign new_n1716_ = new_n1709_ & ~new_n1712_;
  assign new_n1717_ = ~new_n1413_ & new_n1423_;
  assign new_n1718_ = ~new_n1416_ & ~new_n1423_;
  assign new_n1719_ = ~new_n1717_ & ~new_n1718_;
  assign new_n1720_ = ~new_n559_ & new_n859_;
  assign new_n1721_ = ~new_n556_ & ~new_n859_;
  assign new_n1722_ = ~new_n1720_ & ~new_n1721_;
  assign new_n1723_ = new_n1719_ & ~new_n1722_;
  assign new_n1724_ = ~new_n1716_ & ~new_n1723_;
  assign new_n1725_ = ~new_n1715_ & new_n1724_;
  assign new_n1726_ = ~new_n294_ & new_n297_;
  assign new_n1727_ = ~new_n1719_ & new_n1722_;
  assign new_n1728_ = ~new_n1726_ & ~new_n1727_;
  assign new_n1729_ = ~new_n1725_ & new_n1728_;
  assign \o[2]  = ~new_n298_ & ~new_n1729_;
  assign new_n1731_ = ~new_n1423_ & \o[2] ;
  assign new_n1732_ = ~new_n859_ & ~\o[2] ;
  assign \o[1]  = new_n1731_ | new_n1732_;
  assign new_n1734_ = new_n987_ & ~\o[1] ;
  assign new_n1735_ = new_n1117_ & ~new_n1423_;
  assign new_n1736_ = ~new_n1734_ & ~new_n1735_;
  assign new_n1737_ = \o[2]  & ~new_n1736_;
  assign new_n1738_ = new_n423_ & ~\o[1] ;
  assign new_n1739_ = new_n553_ & ~new_n859_;
  assign new_n1740_ = ~new_n1738_ & ~new_n1739_;
  assign new_n1741_ = ~\o[2]  & ~new_n1740_;
  assign \o[0]  = ~new_n1737_ & ~new_n1741_;
  assign new_n1743_ = ~new_n1433_ & ~\o[2] ;
  assign new_n1744_ = ~new_n1430_ & \o[2] ;
  assign \o[3]  = new_n1743_ | new_n1744_;
  assign new_n1746_ = ~new_n862_ & ~\o[2] ;
  assign new_n1747_ = ~new_n1426_ & \o[2] ;
  assign \o[4]  = new_n1746_ | new_n1747_;
  assign new_n1749_ = ~new_n1441_ & ~\o[2] ;
  assign new_n1750_ = ~new_n1438_ & \o[2] ;
  assign \o[5]  = new_n1749_ | new_n1750_;
  assign new_n1752_ = ~new_n1452_ & \o[2] ;
  assign new_n1753_ = ~new_n1449_ & ~\o[2] ;
  assign \o[6]  = new_n1752_ | new_n1753_;
  assign new_n1755_ = ~new_n1461_ & ~\o[2] ;
  assign new_n1756_ = ~new_n1458_ & \o[2] ;
  assign \o[7]  = new_n1755_ | new_n1756_;
  assign new_n1758_ = ~new_n1468_ & ~\o[2] ;
  assign new_n1759_ = ~new_n1471_ & \o[2] ;
  assign \o[8]  = new_n1758_ | new_n1759_;
  assign new_n1761_ = ~new_n1481_ & \o[2] ;
  assign new_n1762_ = ~new_n1478_ & ~\o[2] ;
  assign \o[9]  = new_n1761_ | new_n1762_;
  assign new_n1764_ = ~new_n1488_ & ~\o[2] ;
  assign new_n1765_ = ~new_n1491_ & \o[2] ;
  assign \o[10]  = new_n1764_ | new_n1765_;
  assign new_n1767_ = ~new_n1501_ & ~\o[2] ;
  assign new_n1768_ = ~new_n1498_ & \o[2] ;
  assign \o[11]  = new_n1767_ | new_n1768_;
  assign new_n1770_ = ~new_n1508_ & ~\o[2] ;
  assign new_n1771_ = ~new_n1511_ & \o[2] ;
  assign \o[12]  = new_n1770_ | new_n1771_;
  assign new_n1773_ = new_n1521_ & ~\o[2] ;
  assign new_n1774_ = new_n1518_ & \o[2] ;
  assign \o[13]  = ~new_n1773_ & ~new_n1774_;
  assign new_n1776_ = ~new_n1528_ & ~\o[2] ;
  assign new_n1777_ = ~new_n1531_ & \o[2] ;
  assign \o[14]  = new_n1776_ | new_n1777_;
  assign new_n1779_ = ~new_n1541_ & ~\o[2] ;
  assign new_n1780_ = ~new_n1538_ & \o[2] ;
  assign \o[15]  = new_n1779_ | new_n1780_;
  assign new_n1782_ = ~new_n1548_ & ~\o[2] ;
  assign new_n1783_ = ~new_n1551_ & \o[2] ;
  assign \o[16]  = new_n1782_ | new_n1783_;
  assign new_n1785_ = new_n1561_ & ~\o[2] ;
  assign new_n1786_ = new_n1558_ & \o[2] ;
  assign \o[17]  = ~new_n1785_ & ~new_n1786_;
  assign new_n1788_ = ~new_n1568_ & ~\o[2] ;
  assign new_n1789_ = ~new_n1571_ & \o[2] ;
  assign \o[18]  = new_n1788_ | new_n1789_;
  assign new_n1791_ = ~new_n1581_ & ~\o[2] ;
  assign new_n1792_ = ~new_n1578_ & \o[2] ;
  assign \o[19]  = new_n1791_ | new_n1792_;
  assign new_n1794_ = ~new_n1588_ & ~\o[2] ;
  assign new_n1795_ = ~new_n1591_ & \o[2] ;
  assign \o[20]  = new_n1794_ | new_n1795_;
  assign new_n1797_ = new_n1601_ & ~\o[2] ;
  assign new_n1798_ = new_n1598_ & \o[2] ;
  assign \o[21]  = ~new_n1797_ & ~new_n1798_;
  assign new_n1800_ = ~new_n1608_ & ~\o[2] ;
  assign new_n1801_ = ~new_n1611_ & \o[2] ;
  assign \o[22]  = new_n1800_ | new_n1801_;
  assign new_n1803_ = ~new_n1621_ & ~\o[2] ;
  assign new_n1804_ = ~new_n1618_ & \o[2] ;
  assign \o[23]  = new_n1803_ | new_n1804_;
  assign new_n1806_ = ~new_n1628_ & ~\o[2] ;
  assign new_n1807_ = ~new_n1631_ & \o[2] ;
  assign \o[24]  = new_n1806_ | new_n1807_;
  assign new_n1809_ = new_n1641_ & ~\o[2] ;
  assign new_n1810_ = new_n1638_ & \o[2] ;
  assign \o[25]  = ~new_n1809_ & ~new_n1810_;
  assign new_n1812_ = ~new_n1648_ & ~\o[2] ;
  assign new_n1813_ = ~new_n1651_ & \o[2] ;
  assign \o[26]  = new_n1812_ | new_n1813_;
  assign new_n1815_ = ~new_n1661_ & \o[2] ;
  assign new_n1816_ = ~new_n1658_ & ~\o[2] ;
  assign \o[27]  = new_n1815_ | new_n1816_;
  assign new_n1818_ = ~new_n1668_ & ~\o[2] ;
  assign new_n1819_ = ~new_n1671_ & \o[2] ;
  assign \o[28]  = new_n1818_ | new_n1819_;
  assign new_n1821_ = new_n1681_ & ~\o[2] ;
  assign new_n1822_ = new_n1678_ & \o[2] ;
  assign \o[29]  = ~new_n1821_ & ~new_n1822_;
  assign new_n1824_ = ~new_n1692_ & \o[2] ;
  assign new_n1825_ = ~new_n1689_ & ~\o[2] ;
  assign \o[30]  = new_n1824_ | new_n1825_;
  assign new_n1827_ = ~new_n1702_ & ~\o[2] ;
  assign new_n1828_ = ~new_n1699_ & \o[2] ;
  assign \o[31]  = new_n1827_ | new_n1828_;
  assign new_n1830_ = new_n1712_ & ~\o[2] ;
  assign new_n1831_ = new_n1709_ & \o[2] ;
  assign \o[32]  = ~new_n1830_ & ~new_n1831_;
  assign new_n1833_ = ~new_n1722_ & ~\o[2] ;
  assign new_n1834_ = ~new_n1719_ & \o[2] ;
  assign \o[33]  = new_n1833_ | new_n1834_;
  assign \o[34]  = ~new_n294_ | ~new_n297_;
endmodule


