// Benchmark "auction_BMR_3_16" written by ABC on Tue Nov 26 14:00:42 2019

module auction_BMR_3_16 ( 
    \p_input[0] , \p_input[1] , \p_input[2] , \p_input[3] , \p_input[4] ,
    \p_input[5] , \p_input[6] , \p_input[7] , \p_input[8] , \p_input[9] ,
    \p_input[10] , \p_input[11] , \p_input[12] , \p_input[13] ,
    \p_input[14] , \p_input[15] , \p_input[16] , \p_input[17] ,
    \p_input[18] , \p_input[19] , \p_input[20] , \p_input[21] ,
    \p_input[22] , \p_input[23] , \p_input[24] , \p_input[25] ,
    \p_input[26] , \p_input[27] , \p_input[28] , \p_input[29] ,
    \p_input[30] , \p_input[31] , \p_input[32] , \p_input[33] ,
    \p_input[34] , \p_input[35] , \p_input[36] , \p_input[37] ,
    \p_input[38] , \p_input[39] , \p_input[40] , \p_input[41] ,
    \p_input[42] , \p_input[43] , \p_input[44] , \p_input[45] ,
    \p_input[46] , \p_input[47] , \p_input[48] , \p_input[49] ,
    \p_input[50] , \p_input[51] , \p_input[52] , \p_input[53] ,
    \p_input[54] , \p_input[55] , \p_input[56] , \p_input[57] ,
    \p_input[58] , \p_input[59] , \p_input[60] , \p_input[61] ,
    \p_input[62] , \p_input[63] , \p_input[64] , \p_input[65] ,
    \p_input[66] , \p_input[67] , \p_input[68] , \p_input[69] ,
    \p_input[70] , \p_input[71] , \p_input[72] , \p_input[73] ,
    \p_input[74] , \p_input[75] , \p_input[76] , \p_input[77] ,
    \p_input[78] , \p_input[79] , \p_input[80] , \p_input[81] ,
    \p_input[82] , \p_input[83] , \p_input[84] , \p_input[85] ,
    \p_input[86] , \p_input[87] , \p_input[88] , \p_input[89] ,
    \p_input[90] , \p_input[91] , \p_input[92] , \p_input[93] ,
    \p_input[94] , \p_input[95] , \p_input[96] , \p_input[97] ,
    \p_input[98] , \p_input[99] , \p_input[100] , \p_input[101] ,
    \p_input[102] , \p_input[103] , \p_input[104] , \p_input[105] ,
    \p_input[106] , \p_input[107] , \p_input[108] , \p_input[109] ,
    \p_input[110] , \p_input[111] , \p_input[112] , \p_input[113] ,
    \p_input[114] , \p_input[115] , \p_input[116] , \p_input[117] ,
    \p_input[118] , \p_input[119] , \p_input[120] , \p_input[121] ,
    \p_input[122] , \p_input[123] , \p_input[124] , \p_input[125] ,
    \p_input[126] , \p_input[127] ,
    \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] , \o[8] ,
    \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] , \o[16] ,
    \o[17] , \o[18]   );
  input  \p_input[0] , \p_input[1] , \p_input[2] , \p_input[3] ,
    \p_input[4] , \p_input[5] , \p_input[6] , \p_input[7] , \p_input[8] ,
    \p_input[9] , \p_input[10] , \p_input[11] , \p_input[12] ,
    \p_input[13] , \p_input[14] , \p_input[15] , \p_input[16] ,
    \p_input[17] , \p_input[18] , \p_input[19] , \p_input[20] ,
    \p_input[21] , \p_input[22] , \p_input[23] , \p_input[24] ,
    \p_input[25] , \p_input[26] , \p_input[27] , \p_input[28] ,
    \p_input[29] , \p_input[30] , \p_input[31] , \p_input[32] ,
    \p_input[33] , \p_input[34] , \p_input[35] , \p_input[36] ,
    \p_input[37] , \p_input[38] , \p_input[39] , \p_input[40] ,
    \p_input[41] , \p_input[42] , \p_input[43] , \p_input[44] ,
    \p_input[45] , \p_input[46] , \p_input[47] , \p_input[48] ,
    \p_input[49] , \p_input[50] , \p_input[51] , \p_input[52] ,
    \p_input[53] , \p_input[54] , \p_input[55] , \p_input[56] ,
    \p_input[57] , \p_input[58] , \p_input[59] , \p_input[60] ,
    \p_input[61] , \p_input[62] , \p_input[63] , \p_input[64] ,
    \p_input[65] , \p_input[66] , \p_input[67] , \p_input[68] ,
    \p_input[69] , \p_input[70] , \p_input[71] , \p_input[72] ,
    \p_input[73] , \p_input[74] , \p_input[75] , \p_input[76] ,
    \p_input[77] , \p_input[78] , \p_input[79] , \p_input[80] ,
    \p_input[81] , \p_input[82] , \p_input[83] , \p_input[84] ,
    \p_input[85] , \p_input[86] , \p_input[87] , \p_input[88] ,
    \p_input[89] , \p_input[90] , \p_input[91] , \p_input[92] ,
    \p_input[93] , \p_input[94] , \p_input[95] , \p_input[96] ,
    \p_input[97] , \p_input[98] , \p_input[99] , \p_input[100] ,
    \p_input[101] , \p_input[102] , \p_input[103] , \p_input[104] ,
    \p_input[105] , \p_input[106] , \p_input[107] , \p_input[108] ,
    \p_input[109] , \p_input[110] , \p_input[111] , \p_input[112] ,
    \p_input[113] , \p_input[114] , \p_input[115] , \p_input[116] ,
    \p_input[117] , \p_input[118] , \p_input[119] , \p_input[120] ,
    \p_input[121] , \p_input[122] , \p_input[123] , \p_input[124] ,
    \p_input[125] , \p_input[126] , \p_input[127] ;
  output \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] ,
    \o[8] , \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] ,
    \o[16] , \o[17] , \o[18] ;
  wire new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_;
  assign new_n148_ = ~\p_input[79]  & ~\p_input[95] ;
  assign new_n149_ = ~\p_input[111]  & ~\p_input[127] ;
  assign new_n150_ = new_n148_ & new_n149_;
  assign new_n151_ = ~\p_input[15]  & ~\p_input[31] ;
  assign new_n152_ = ~\p_input[47]  & ~\p_input[63] ;
  assign new_n153_ = new_n151_ & new_n152_;
  assign new_n154_ = new_n150_ & ~new_n153_;
  assign new_n155_ = ~\p_input[15]  & \p_input[31] ;
  assign new_n156_ = \p_input[15]  & ~\p_input[31] ;
  assign new_n157_ = ~\p_input[14]  & \p_input[30] ;
  assign new_n158_ = \p_input[14]  & ~\p_input[30] ;
  assign new_n159_ = ~\p_input[13]  & \p_input[29] ;
  assign new_n160_ = \p_input[13]  & ~\p_input[29] ;
  assign new_n161_ = ~\p_input[12]  & \p_input[28] ;
  assign new_n162_ = \p_input[12]  & ~\p_input[28] ;
  assign new_n163_ = ~\p_input[11]  & \p_input[27] ;
  assign new_n164_ = \p_input[11]  & ~\p_input[27] ;
  assign new_n165_ = ~\p_input[10]  & \p_input[26] ;
  assign new_n166_ = \p_input[10]  & ~\p_input[26] ;
  assign new_n167_ = ~\p_input[9]  & \p_input[25] ;
  assign new_n168_ = \p_input[9]  & ~\p_input[25] ;
  assign new_n169_ = ~\p_input[8]  & \p_input[24] ;
  assign new_n170_ = \p_input[8]  & ~\p_input[24] ;
  assign new_n171_ = ~\p_input[7]  & \p_input[23] ;
  assign new_n172_ = \p_input[7]  & ~\p_input[23] ;
  assign new_n173_ = ~\p_input[6]  & \p_input[22] ;
  assign new_n174_ = \p_input[6]  & ~\p_input[22] ;
  assign new_n175_ = ~\p_input[5]  & \p_input[21] ;
  assign new_n176_ = \p_input[5]  & ~\p_input[21] ;
  assign new_n177_ = ~\p_input[4]  & \p_input[20] ;
  assign new_n178_ = \p_input[4]  & ~\p_input[20] ;
  assign new_n179_ = ~\p_input[3]  & \p_input[19] ;
  assign new_n180_ = \p_input[3]  & ~\p_input[19] ;
  assign new_n181_ = ~\p_input[2]  & \p_input[18] ;
  assign new_n182_ = \p_input[2]  & ~\p_input[18] ;
  assign new_n183_ = ~\p_input[1]  & \p_input[17] ;
  assign new_n184_ = \p_input[1]  & ~\p_input[17] ;
  assign new_n185_ = \p_input[0]  & ~\p_input[16] ;
  assign new_n186_ = ~new_n184_ & ~new_n185_;
  assign new_n187_ = ~new_n183_ & ~new_n186_;
  assign new_n188_ = ~new_n182_ & ~new_n187_;
  assign new_n189_ = ~new_n181_ & ~new_n188_;
  assign new_n190_ = ~new_n180_ & ~new_n189_;
  assign new_n191_ = ~new_n179_ & ~new_n190_;
  assign new_n192_ = ~new_n178_ & ~new_n191_;
  assign new_n193_ = ~new_n177_ & ~new_n192_;
  assign new_n194_ = ~new_n176_ & ~new_n193_;
  assign new_n195_ = ~new_n175_ & ~new_n194_;
  assign new_n196_ = ~new_n174_ & ~new_n195_;
  assign new_n197_ = ~new_n173_ & ~new_n196_;
  assign new_n198_ = ~new_n172_ & ~new_n197_;
  assign new_n199_ = ~new_n171_ & ~new_n198_;
  assign new_n200_ = ~new_n170_ & ~new_n199_;
  assign new_n201_ = ~new_n169_ & ~new_n200_;
  assign new_n202_ = ~new_n168_ & ~new_n201_;
  assign new_n203_ = ~new_n167_ & ~new_n202_;
  assign new_n204_ = ~new_n166_ & ~new_n203_;
  assign new_n205_ = ~new_n165_ & ~new_n204_;
  assign new_n206_ = ~new_n164_ & ~new_n205_;
  assign new_n207_ = ~new_n163_ & ~new_n206_;
  assign new_n208_ = ~new_n162_ & ~new_n207_;
  assign new_n209_ = ~new_n161_ & ~new_n208_;
  assign new_n210_ = ~new_n160_ & ~new_n209_;
  assign new_n211_ = ~new_n159_ & ~new_n210_;
  assign new_n212_ = ~new_n158_ & ~new_n211_;
  assign new_n213_ = ~new_n157_ & ~new_n212_;
  assign new_n214_ = ~new_n156_ & ~new_n213_;
  assign new_n215_ = ~new_n155_ & ~new_n214_;
  assign new_n216_ = \p_input[17]  & ~new_n215_;
  assign new_n217_ = \p_input[1]  & new_n215_;
  assign new_n218_ = ~new_n216_ & ~new_n217_;
  assign new_n219_ = new_n151_ & ~new_n152_;
  assign new_n220_ = ~new_n151_ & new_n152_;
  assign new_n221_ = ~\p_input[47]  & \p_input[63] ;
  assign new_n222_ = \p_input[47]  & ~\p_input[63] ;
  assign new_n223_ = ~\p_input[46]  & \p_input[62] ;
  assign new_n224_ = \p_input[46]  & ~\p_input[62] ;
  assign new_n225_ = ~\p_input[45]  & \p_input[61] ;
  assign new_n226_ = \p_input[45]  & ~\p_input[61] ;
  assign new_n227_ = ~\p_input[44]  & \p_input[60] ;
  assign new_n228_ = \p_input[44]  & ~\p_input[60] ;
  assign new_n229_ = ~\p_input[43]  & \p_input[59] ;
  assign new_n230_ = \p_input[43]  & ~\p_input[59] ;
  assign new_n231_ = ~\p_input[42]  & \p_input[58] ;
  assign new_n232_ = \p_input[42]  & ~\p_input[58] ;
  assign new_n233_ = ~\p_input[41]  & \p_input[57] ;
  assign new_n234_ = \p_input[41]  & ~\p_input[57] ;
  assign new_n235_ = ~\p_input[40]  & \p_input[56] ;
  assign new_n236_ = \p_input[40]  & ~\p_input[56] ;
  assign new_n237_ = ~\p_input[39]  & \p_input[55] ;
  assign new_n238_ = \p_input[39]  & ~\p_input[55] ;
  assign new_n239_ = ~\p_input[38]  & \p_input[54] ;
  assign new_n240_ = \p_input[38]  & ~\p_input[54] ;
  assign new_n241_ = ~\p_input[37]  & \p_input[53] ;
  assign new_n242_ = \p_input[37]  & ~\p_input[53] ;
  assign new_n243_ = ~\p_input[36]  & \p_input[52] ;
  assign new_n244_ = \p_input[36]  & ~\p_input[52] ;
  assign new_n245_ = ~\p_input[35]  & \p_input[51] ;
  assign new_n246_ = \p_input[35]  & ~\p_input[51] ;
  assign new_n247_ = ~\p_input[34]  & \p_input[50] ;
  assign new_n248_ = \p_input[34]  & ~\p_input[50] ;
  assign new_n249_ = ~\p_input[33]  & \p_input[49] ;
  assign new_n250_ = \p_input[33]  & ~\p_input[49] ;
  assign new_n251_ = \p_input[32]  & ~\p_input[48] ;
  assign new_n252_ = ~new_n250_ & ~new_n251_;
  assign new_n253_ = ~new_n249_ & ~new_n252_;
  assign new_n254_ = ~new_n248_ & ~new_n253_;
  assign new_n255_ = ~new_n247_ & ~new_n254_;
  assign new_n256_ = ~new_n246_ & ~new_n255_;
  assign new_n257_ = ~new_n245_ & ~new_n256_;
  assign new_n258_ = ~new_n244_ & ~new_n257_;
  assign new_n259_ = ~new_n243_ & ~new_n258_;
  assign new_n260_ = ~new_n242_ & ~new_n259_;
  assign new_n261_ = ~new_n241_ & ~new_n260_;
  assign new_n262_ = ~new_n240_ & ~new_n261_;
  assign new_n263_ = ~new_n239_ & ~new_n262_;
  assign new_n264_ = ~new_n238_ & ~new_n263_;
  assign new_n265_ = ~new_n237_ & ~new_n264_;
  assign new_n266_ = ~new_n236_ & ~new_n265_;
  assign new_n267_ = ~new_n235_ & ~new_n266_;
  assign new_n268_ = ~new_n234_ & ~new_n267_;
  assign new_n269_ = ~new_n233_ & ~new_n268_;
  assign new_n270_ = ~new_n232_ & ~new_n269_;
  assign new_n271_ = ~new_n231_ & ~new_n270_;
  assign new_n272_ = ~new_n230_ & ~new_n271_;
  assign new_n273_ = ~new_n229_ & ~new_n272_;
  assign new_n274_ = ~new_n228_ & ~new_n273_;
  assign new_n275_ = ~new_n227_ & ~new_n274_;
  assign new_n276_ = ~new_n226_ & ~new_n275_;
  assign new_n277_ = ~new_n225_ & ~new_n276_;
  assign new_n278_ = ~new_n224_ & ~new_n277_;
  assign new_n279_ = ~new_n223_ & ~new_n278_;
  assign new_n280_ = ~new_n222_ & ~new_n279_;
  assign new_n281_ = ~new_n221_ & ~new_n280_;
  assign new_n282_ = \p_input[62]  & ~new_n281_;
  assign new_n283_ = \p_input[46]  & new_n281_;
  assign new_n284_ = ~new_n282_ & ~new_n283_;
  assign new_n285_ = \p_input[30]  & ~new_n215_;
  assign new_n286_ = \p_input[14]  & new_n215_;
  assign new_n287_ = ~new_n285_ & ~new_n286_;
  assign new_n288_ = ~new_n284_ & new_n287_;
  assign new_n289_ = \p_input[49]  & ~new_n281_;
  assign new_n290_ = \p_input[33]  & new_n281_;
  assign new_n291_ = ~new_n289_ & ~new_n290_;
  assign new_n292_ = new_n218_ & ~new_n291_;
  assign new_n293_ = \p_input[48]  & ~new_n281_;
  assign new_n294_ = \p_input[32]  & new_n281_;
  assign new_n295_ = ~new_n293_ & ~new_n294_;
  assign new_n296_ = \p_input[16]  & ~new_n215_;
  assign new_n297_ = \p_input[0]  & new_n215_;
  assign new_n298_ = ~new_n296_ & ~new_n297_;
  assign new_n299_ = new_n295_ & ~new_n298_;
  assign new_n300_ = ~new_n292_ & new_n299_;
  assign new_n301_ = \p_input[50]  & ~new_n281_;
  assign new_n302_ = \p_input[34]  & new_n281_;
  assign new_n303_ = ~new_n301_ & ~new_n302_;
  assign new_n304_ = \p_input[18]  & ~new_n215_;
  assign new_n305_ = \p_input[2]  & new_n215_;
  assign new_n306_ = ~new_n304_ & ~new_n305_;
  assign new_n307_ = new_n303_ & ~new_n306_;
  assign new_n308_ = ~new_n218_ & new_n291_;
  assign new_n309_ = ~new_n307_ & ~new_n308_;
  assign new_n310_ = ~new_n300_ & new_n309_;
  assign new_n311_ = \p_input[19]  & ~new_n215_;
  assign new_n312_ = \p_input[3]  & new_n215_;
  assign new_n313_ = ~new_n311_ & ~new_n312_;
  assign new_n314_ = \p_input[51]  & ~new_n281_;
  assign new_n315_ = \p_input[35]  & new_n281_;
  assign new_n316_ = ~new_n314_ & ~new_n315_;
  assign new_n317_ = new_n313_ & ~new_n316_;
  assign new_n318_ = ~new_n303_ & new_n306_;
  assign new_n319_ = ~new_n317_ & ~new_n318_;
  assign new_n320_ = ~new_n310_ & new_n319_;
  assign new_n321_ = \p_input[52]  & ~new_n281_;
  assign new_n322_ = \p_input[36]  & new_n281_;
  assign new_n323_ = ~new_n321_ & ~new_n322_;
  assign new_n324_ = \p_input[20]  & ~new_n215_;
  assign new_n325_ = \p_input[4]  & new_n215_;
  assign new_n326_ = ~new_n324_ & ~new_n325_;
  assign new_n327_ = new_n323_ & ~new_n326_;
  assign new_n328_ = ~new_n313_ & new_n316_;
  assign new_n329_ = ~new_n327_ & ~new_n328_;
  assign new_n330_ = ~new_n320_ & new_n329_;
  assign new_n331_ = \p_input[53]  & ~new_n281_;
  assign new_n332_ = \p_input[37]  & new_n281_;
  assign new_n333_ = ~new_n331_ & ~new_n332_;
  assign new_n334_ = \p_input[21]  & ~new_n215_;
  assign new_n335_ = \p_input[5]  & new_n215_;
  assign new_n336_ = ~new_n334_ & ~new_n335_;
  assign new_n337_ = ~new_n333_ & new_n336_;
  assign new_n338_ = ~new_n323_ & new_n326_;
  assign new_n339_ = ~new_n337_ & ~new_n338_;
  assign new_n340_ = ~new_n330_ & new_n339_;
  assign new_n341_ = \p_input[22]  & ~new_n215_;
  assign new_n342_ = \p_input[6]  & new_n215_;
  assign new_n343_ = ~new_n341_ & ~new_n342_;
  assign new_n344_ = \p_input[54]  & ~new_n281_;
  assign new_n345_ = \p_input[38]  & new_n281_;
  assign new_n346_ = ~new_n344_ & ~new_n345_;
  assign new_n347_ = ~new_n343_ & new_n346_;
  assign new_n348_ = new_n333_ & ~new_n336_;
  assign new_n349_ = ~new_n347_ & ~new_n348_;
  assign new_n350_ = ~new_n340_ & new_n349_;
  assign new_n351_ = \p_input[23]  & ~new_n215_;
  assign new_n352_ = \p_input[7]  & new_n215_;
  assign new_n353_ = ~new_n351_ & ~new_n352_;
  assign new_n354_ = \p_input[55]  & ~new_n281_;
  assign new_n355_ = \p_input[39]  & new_n281_;
  assign new_n356_ = ~new_n354_ & ~new_n355_;
  assign new_n357_ = new_n353_ & ~new_n356_;
  assign new_n358_ = new_n343_ & ~new_n346_;
  assign new_n359_ = ~new_n357_ & ~new_n358_;
  assign new_n360_ = ~new_n350_ & new_n359_;
  assign new_n361_ = ~new_n353_ & new_n356_;
  assign new_n362_ = \p_input[24]  & ~new_n215_;
  assign new_n363_ = \p_input[8]  & new_n215_;
  assign new_n364_ = ~new_n362_ & ~new_n363_;
  assign new_n365_ = \p_input[56]  & ~new_n281_;
  assign new_n366_ = \p_input[40]  & new_n281_;
  assign new_n367_ = ~new_n365_ & ~new_n366_;
  assign new_n368_ = ~new_n364_ & new_n367_;
  assign new_n369_ = ~new_n361_ & ~new_n368_;
  assign new_n370_ = ~new_n360_ & new_n369_;
  assign new_n371_ = new_n364_ & ~new_n367_;
  assign new_n372_ = \p_input[57]  & ~new_n281_;
  assign new_n373_ = \p_input[41]  & new_n281_;
  assign new_n374_ = ~new_n372_ & ~new_n373_;
  assign new_n375_ = \p_input[25]  & ~new_n215_;
  assign new_n376_ = \p_input[9]  & new_n215_;
  assign new_n377_ = ~new_n375_ & ~new_n376_;
  assign new_n378_ = ~new_n374_ & new_n377_;
  assign new_n379_ = ~new_n371_ & ~new_n378_;
  assign new_n380_ = ~new_n370_ & new_n379_;
  assign new_n381_ = new_n374_ & ~new_n377_;
  assign new_n382_ = \p_input[26]  & ~new_n215_;
  assign new_n383_ = \p_input[10]  & new_n215_;
  assign new_n384_ = ~new_n382_ & ~new_n383_;
  assign new_n385_ = \p_input[58]  & ~new_n281_;
  assign new_n386_ = \p_input[42]  & new_n281_;
  assign new_n387_ = ~new_n385_ & ~new_n386_;
  assign new_n388_ = ~new_n384_ & new_n387_;
  assign new_n389_ = ~new_n381_ & ~new_n388_;
  assign new_n390_ = ~new_n380_ & new_n389_;
  assign new_n391_ = \p_input[27]  & ~new_n215_;
  assign new_n392_ = \p_input[11]  & new_n215_;
  assign new_n393_ = ~new_n391_ & ~new_n392_;
  assign new_n394_ = \p_input[59]  & ~new_n281_;
  assign new_n395_ = \p_input[43]  & new_n281_;
  assign new_n396_ = ~new_n394_ & ~new_n395_;
  assign new_n397_ = new_n393_ & ~new_n396_;
  assign new_n398_ = new_n384_ & ~new_n387_;
  assign new_n399_ = ~new_n397_ & ~new_n398_;
  assign new_n400_ = ~new_n390_ & new_n399_;
  assign new_n401_ = \p_input[60]  & ~new_n281_;
  assign new_n402_ = \p_input[44]  & new_n281_;
  assign new_n403_ = ~new_n401_ & ~new_n402_;
  assign new_n404_ = \p_input[28]  & ~new_n215_;
  assign new_n405_ = \p_input[12]  & new_n215_;
  assign new_n406_ = ~new_n404_ & ~new_n405_;
  assign new_n407_ = new_n403_ & ~new_n406_;
  assign new_n408_ = ~new_n393_ & new_n396_;
  assign new_n409_ = ~new_n407_ & ~new_n408_;
  assign new_n410_ = ~new_n400_ & new_n409_;
  assign new_n411_ = ~new_n403_ & new_n406_;
  assign new_n412_ = \p_input[29]  & ~new_n215_;
  assign new_n413_ = \p_input[13]  & new_n215_;
  assign new_n414_ = ~new_n412_ & ~new_n413_;
  assign new_n415_ = \p_input[61]  & ~new_n281_;
  assign new_n416_ = \p_input[45]  & new_n281_;
  assign new_n417_ = ~new_n415_ & ~new_n416_;
  assign new_n418_ = new_n414_ & ~new_n417_;
  assign new_n419_ = ~new_n411_ & ~new_n418_;
  assign new_n420_ = ~new_n410_ & new_n419_;
  assign new_n421_ = new_n284_ & ~new_n287_;
  assign new_n422_ = ~new_n414_ & new_n417_;
  assign new_n423_ = ~new_n421_ & ~new_n422_;
  assign new_n424_ = ~new_n420_ & new_n423_;
  assign new_n425_ = ~new_n288_ & ~new_n424_;
  assign new_n426_ = ~new_n220_ & ~new_n425_;
  assign new_n427_ = ~new_n219_ & ~new_n426_;
  assign new_n428_ = ~new_n218_ & new_n427_;
  assign new_n429_ = ~new_n291_ & ~new_n427_;
  assign new_n430_ = ~new_n428_ & ~new_n429_;
  assign new_n431_ = ~\p_input[79]  & \p_input[95] ;
  assign new_n432_ = \p_input[79]  & ~\p_input[95] ;
  assign new_n433_ = ~\p_input[78]  & \p_input[94] ;
  assign new_n434_ = \p_input[78]  & ~\p_input[94] ;
  assign new_n435_ = ~\p_input[77]  & \p_input[93] ;
  assign new_n436_ = \p_input[77]  & ~\p_input[93] ;
  assign new_n437_ = ~\p_input[76]  & \p_input[92] ;
  assign new_n438_ = \p_input[76]  & ~\p_input[92] ;
  assign new_n439_ = ~\p_input[75]  & \p_input[91] ;
  assign new_n440_ = \p_input[75]  & ~\p_input[91] ;
  assign new_n441_ = ~\p_input[74]  & \p_input[90] ;
  assign new_n442_ = \p_input[74]  & ~\p_input[90] ;
  assign new_n443_ = ~\p_input[73]  & \p_input[89] ;
  assign new_n444_ = \p_input[73]  & ~\p_input[89] ;
  assign new_n445_ = ~\p_input[72]  & \p_input[88] ;
  assign new_n446_ = \p_input[72]  & ~\p_input[88] ;
  assign new_n447_ = ~\p_input[71]  & \p_input[87] ;
  assign new_n448_ = \p_input[71]  & ~\p_input[87] ;
  assign new_n449_ = ~\p_input[70]  & \p_input[86] ;
  assign new_n450_ = \p_input[70]  & ~\p_input[86] ;
  assign new_n451_ = ~\p_input[69]  & \p_input[85] ;
  assign new_n452_ = \p_input[69]  & ~\p_input[85] ;
  assign new_n453_ = ~\p_input[68]  & \p_input[84] ;
  assign new_n454_ = \p_input[68]  & ~\p_input[84] ;
  assign new_n455_ = ~\p_input[67]  & \p_input[83] ;
  assign new_n456_ = \p_input[67]  & ~\p_input[83] ;
  assign new_n457_ = ~\p_input[66]  & \p_input[82] ;
  assign new_n458_ = \p_input[66]  & ~\p_input[82] ;
  assign new_n459_ = ~\p_input[65]  & \p_input[81] ;
  assign new_n460_ = \p_input[65]  & ~\p_input[81] ;
  assign new_n461_ = \p_input[64]  & ~\p_input[80] ;
  assign new_n462_ = ~new_n460_ & ~new_n461_;
  assign new_n463_ = ~new_n459_ & ~new_n462_;
  assign new_n464_ = ~new_n458_ & ~new_n463_;
  assign new_n465_ = ~new_n457_ & ~new_n464_;
  assign new_n466_ = ~new_n456_ & ~new_n465_;
  assign new_n467_ = ~new_n455_ & ~new_n466_;
  assign new_n468_ = ~new_n454_ & ~new_n467_;
  assign new_n469_ = ~new_n453_ & ~new_n468_;
  assign new_n470_ = ~new_n452_ & ~new_n469_;
  assign new_n471_ = ~new_n451_ & ~new_n470_;
  assign new_n472_ = ~new_n450_ & ~new_n471_;
  assign new_n473_ = ~new_n449_ & ~new_n472_;
  assign new_n474_ = ~new_n448_ & ~new_n473_;
  assign new_n475_ = ~new_n447_ & ~new_n474_;
  assign new_n476_ = ~new_n446_ & ~new_n475_;
  assign new_n477_ = ~new_n445_ & ~new_n476_;
  assign new_n478_ = ~new_n444_ & ~new_n477_;
  assign new_n479_ = ~new_n443_ & ~new_n478_;
  assign new_n480_ = ~new_n442_ & ~new_n479_;
  assign new_n481_ = ~new_n441_ & ~new_n480_;
  assign new_n482_ = ~new_n440_ & ~new_n481_;
  assign new_n483_ = ~new_n439_ & ~new_n482_;
  assign new_n484_ = ~new_n438_ & ~new_n483_;
  assign new_n485_ = ~new_n437_ & ~new_n484_;
  assign new_n486_ = ~new_n436_ & ~new_n485_;
  assign new_n487_ = ~new_n435_ & ~new_n486_;
  assign new_n488_ = ~new_n434_ & ~new_n487_;
  assign new_n489_ = ~new_n433_ & ~new_n488_;
  assign new_n490_ = ~new_n432_ & ~new_n489_;
  assign new_n491_ = ~new_n431_ & ~new_n490_;
  assign new_n492_ = \p_input[81]  & ~new_n491_;
  assign new_n493_ = \p_input[65]  & new_n491_;
  assign new_n494_ = ~new_n492_ & ~new_n493_;
  assign new_n495_ = new_n148_ & ~new_n149_;
  assign new_n496_ = ~new_n148_ & new_n149_;
  assign new_n497_ = ~\p_input[111]  & \p_input[127] ;
  assign new_n498_ = \p_input[111]  & ~\p_input[127] ;
  assign new_n499_ = ~\p_input[110]  & \p_input[126] ;
  assign new_n500_ = \p_input[110]  & ~\p_input[126] ;
  assign new_n501_ = ~\p_input[109]  & \p_input[125] ;
  assign new_n502_ = \p_input[109]  & ~\p_input[125] ;
  assign new_n503_ = ~\p_input[108]  & \p_input[124] ;
  assign new_n504_ = \p_input[108]  & ~\p_input[124] ;
  assign new_n505_ = ~\p_input[107]  & \p_input[123] ;
  assign new_n506_ = \p_input[107]  & ~\p_input[123] ;
  assign new_n507_ = ~\p_input[106]  & \p_input[122] ;
  assign new_n508_ = \p_input[106]  & ~\p_input[122] ;
  assign new_n509_ = ~\p_input[105]  & \p_input[121] ;
  assign new_n510_ = \p_input[105]  & ~\p_input[121] ;
  assign new_n511_ = ~\p_input[104]  & \p_input[120] ;
  assign new_n512_ = \p_input[104]  & ~\p_input[120] ;
  assign new_n513_ = ~\p_input[103]  & \p_input[119] ;
  assign new_n514_ = \p_input[103]  & ~\p_input[119] ;
  assign new_n515_ = ~\p_input[102]  & \p_input[118] ;
  assign new_n516_ = \p_input[102]  & ~\p_input[118] ;
  assign new_n517_ = ~\p_input[101]  & \p_input[117] ;
  assign new_n518_ = \p_input[101]  & ~\p_input[117] ;
  assign new_n519_ = ~\p_input[100]  & \p_input[116] ;
  assign new_n520_ = \p_input[100]  & ~\p_input[116] ;
  assign new_n521_ = ~\p_input[99]  & \p_input[115] ;
  assign new_n522_ = \p_input[99]  & ~\p_input[115] ;
  assign new_n523_ = ~\p_input[98]  & \p_input[114] ;
  assign new_n524_ = \p_input[98]  & ~\p_input[114] ;
  assign new_n525_ = ~\p_input[97]  & \p_input[113] ;
  assign new_n526_ = \p_input[97]  & ~\p_input[113] ;
  assign new_n527_ = \p_input[96]  & ~\p_input[112] ;
  assign new_n528_ = ~new_n526_ & ~new_n527_;
  assign new_n529_ = ~new_n525_ & ~new_n528_;
  assign new_n530_ = ~new_n524_ & ~new_n529_;
  assign new_n531_ = ~new_n523_ & ~new_n530_;
  assign new_n532_ = ~new_n522_ & ~new_n531_;
  assign new_n533_ = ~new_n521_ & ~new_n532_;
  assign new_n534_ = ~new_n520_ & ~new_n533_;
  assign new_n535_ = ~new_n519_ & ~new_n534_;
  assign new_n536_ = ~new_n518_ & ~new_n535_;
  assign new_n537_ = ~new_n517_ & ~new_n536_;
  assign new_n538_ = ~new_n516_ & ~new_n537_;
  assign new_n539_ = ~new_n515_ & ~new_n538_;
  assign new_n540_ = ~new_n514_ & ~new_n539_;
  assign new_n541_ = ~new_n513_ & ~new_n540_;
  assign new_n542_ = ~new_n512_ & ~new_n541_;
  assign new_n543_ = ~new_n511_ & ~new_n542_;
  assign new_n544_ = ~new_n510_ & ~new_n543_;
  assign new_n545_ = ~new_n509_ & ~new_n544_;
  assign new_n546_ = ~new_n508_ & ~new_n545_;
  assign new_n547_ = ~new_n507_ & ~new_n546_;
  assign new_n548_ = ~new_n506_ & ~new_n547_;
  assign new_n549_ = ~new_n505_ & ~new_n548_;
  assign new_n550_ = ~new_n504_ & ~new_n549_;
  assign new_n551_ = ~new_n503_ & ~new_n550_;
  assign new_n552_ = ~new_n502_ & ~new_n551_;
  assign new_n553_ = ~new_n501_ & ~new_n552_;
  assign new_n554_ = ~new_n500_ & ~new_n553_;
  assign new_n555_ = ~new_n499_ & ~new_n554_;
  assign new_n556_ = ~new_n498_ & ~new_n555_;
  assign new_n557_ = ~new_n497_ & ~new_n556_;
  assign new_n558_ = \p_input[113]  & ~new_n557_;
  assign new_n559_ = \p_input[97]  & new_n557_;
  assign new_n560_ = ~new_n558_ & ~new_n559_;
  assign new_n561_ = new_n494_ & ~new_n560_;
  assign new_n562_ = \p_input[112]  & ~new_n557_;
  assign new_n563_ = \p_input[96]  & new_n557_;
  assign new_n564_ = ~new_n562_ & ~new_n563_;
  assign new_n565_ = \p_input[80]  & ~new_n491_;
  assign new_n566_ = \p_input[64]  & new_n491_;
  assign new_n567_ = ~new_n565_ & ~new_n566_;
  assign new_n568_ = new_n564_ & ~new_n567_;
  assign new_n569_ = ~new_n561_ & new_n568_;
  assign new_n570_ = \p_input[114]  & ~new_n557_;
  assign new_n571_ = \p_input[98]  & new_n557_;
  assign new_n572_ = ~new_n570_ & ~new_n571_;
  assign new_n573_ = \p_input[82]  & ~new_n491_;
  assign new_n574_ = \p_input[66]  & new_n491_;
  assign new_n575_ = ~new_n573_ & ~new_n574_;
  assign new_n576_ = new_n572_ & ~new_n575_;
  assign new_n577_ = ~new_n494_ & new_n560_;
  assign new_n578_ = ~new_n576_ & ~new_n577_;
  assign new_n579_ = ~new_n569_ & new_n578_;
  assign new_n580_ = ~new_n572_ & new_n575_;
  assign new_n581_ = \p_input[115]  & ~new_n557_;
  assign new_n582_ = \p_input[99]  & new_n557_;
  assign new_n583_ = ~new_n581_ & ~new_n582_;
  assign new_n584_ = \p_input[83]  & ~new_n491_;
  assign new_n585_ = \p_input[67]  & new_n491_;
  assign new_n586_ = ~new_n584_ & ~new_n585_;
  assign new_n587_ = ~new_n583_ & new_n586_;
  assign new_n588_ = ~new_n580_ & ~new_n587_;
  assign new_n589_ = ~new_n579_ & new_n588_;
  assign new_n590_ = \p_input[84]  & ~new_n491_;
  assign new_n591_ = \p_input[68]  & new_n491_;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign new_n593_ = \p_input[116]  & ~new_n557_;
  assign new_n594_ = \p_input[100]  & new_n557_;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign new_n596_ = ~new_n592_ & new_n595_;
  assign new_n597_ = new_n583_ & ~new_n586_;
  assign new_n598_ = ~new_n596_ & ~new_n597_;
  assign new_n599_ = ~new_n589_ & new_n598_;
  assign new_n600_ = \p_input[117]  & ~new_n557_;
  assign new_n601_ = \p_input[101]  & new_n557_;
  assign new_n602_ = ~new_n600_ & ~new_n601_;
  assign new_n603_ = \p_input[85]  & ~new_n491_;
  assign new_n604_ = \p_input[69]  & new_n491_;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = ~new_n602_ & new_n605_;
  assign new_n607_ = new_n592_ & ~new_n595_;
  assign new_n608_ = ~new_n606_ & ~new_n607_;
  assign new_n609_ = ~new_n599_ & new_n608_;
  assign new_n610_ = \p_input[118]  & ~new_n557_;
  assign new_n611_ = \p_input[102]  & new_n557_;
  assign new_n612_ = ~new_n610_ & ~new_n611_;
  assign new_n613_ = \p_input[86]  & ~new_n491_;
  assign new_n614_ = \p_input[70]  & new_n491_;
  assign new_n615_ = ~new_n613_ & ~new_n614_;
  assign new_n616_ = new_n612_ & ~new_n615_;
  assign new_n617_ = new_n602_ & ~new_n605_;
  assign new_n618_ = ~new_n616_ & ~new_n617_;
  assign new_n619_ = ~new_n609_ & new_n618_;
  assign new_n620_ = ~new_n612_ & new_n615_;
  assign new_n621_ = \p_input[87]  & ~new_n491_;
  assign new_n622_ = \p_input[71]  & new_n491_;
  assign new_n623_ = ~new_n621_ & ~new_n622_;
  assign new_n624_ = \p_input[119]  & ~new_n557_;
  assign new_n625_ = \p_input[103]  & new_n557_;
  assign new_n626_ = ~new_n624_ & ~new_n625_;
  assign new_n627_ = new_n623_ & ~new_n626_;
  assign new_n628_ = ~new_n620_ & ~new_n627_;
  assign new_n629_ = ~new_n619_ & new_n628_;
  assign new_n630_ = ~new_n623_ & new_n626_;
  assign new_n631_ = \p_input[120]  & ~new_n557_;
  assign new_n632_ = \p_input[104]  & new_n557_;
  assign new_n633_ = ~new_n631_ & ~new_n632_;
  assign new_n634_ = \p_input[88]  & ~new_n491_;
  assign new_n635_ = \p_input[72]  & new_n491_;
  assign new_n636_ = ~new_n634_ & ~new_n635_;
  assign new_n637_ = new_n633_ & ~new_n636_;
  assign new_n638_ = ~new_n630_ & ~new_n637_;
  assign new_n639_ = ~new_n629_ & new_n638_;
  assign new_n640_ = ~new_n633_ & new_n636_;
  assign new_n641_ = \p_input[121]  & ~new_n557_;
  assign new_n642_ = \p_input[105]  & new_n557_;
  assign new_n643_ = ~new_n641_ & ~new_n642_;
  assign new_n644_ = \p_input[89]  & ~new_n491_;
  assign new_n645_ = \p_input[73]  & new_n491_;
  assign new_n646_ = ~new_n644_ & ~new_n645_;
  assign new_n647_ = ~new_n643_ & new_n646_;
  assign new_n648_ = ~new_n640_ & ~new_n647_;
  assign new_n649_ = ~new_n639_ & new_n648_;
  assign new_n650_ = new_n643_ & ~new_n646_;
  assign new_n651_ = \p_input[90]  & ~new_n491_;
  assign new_n652_ = \p_input[74]  & new_n491_;
  assign new_n653_ = ~new_n651_ & ~new_n652_;
  assign new_n654_ = \p_input[122]  & ~new_n557_;
  assign new_n655_ = \p_input[106]  & new_n557_;
  assign new_n656_ = ~new_n654_ & ~new_n655_;
  assign new_n657_ = ~new_n653_ & new_n656_;
  assign new_n658_ = ~new_n650_ & ~new_n657_;
  assign new_n659_ = ~new_n649_ & new_n658_;
  assign new_n660_ = \p_input[123]  & ~new_n557_;
  assign new_n661_ = \p_input[107]  & new_n557_;
  assign new_n662_ = ~new_n660_ & ~new_n661_;
  assign new_n663_ = \p_input[91]  & ~new_n491_;
  assign new_n664_ = \p_input[75]  & new_n491_;
  assign new_n665_ = ~new_n663_ & ~new_n664_;
  assign new_n666_ = ~new_n662_ & new_n665_;
  assign new_n667_ = new_n653_ & ~new_n656_;
  assign new_n668_ = ~new_n666_ & ~new_n667_;
  assign new_n669_ = ~new_n659_ & new_n668_;
  assign new_n670_ = \p_input[92]  & ~new_n491_;
  assign new_n671_ = \p_input[76]  & new_n491_;
  assign new_n672_ = ~new_n670_ & ~new_n671_;
  assign new_n673_ = \p_input[124]  & ~new_n557_;
  assign new_n674_ = \p_input[108]  & new_n557_;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = ~new_n672_ & new_n675_;
  assign new_n677_ = new_n662_ & ~new_n665_;
  assign new_n678_ = ~new_n676_ & ~new_n677_;
  assign new_n679_ = ~new_n669_ & new_n678_;
  assign new_n680_ = new_n672_ & ~new_n675_;
  assign new_n681_ = \p_input[93]  & ~new_n491_;
  assign new_n682_ = \p_input[77]  & new_n491_;
  assign new_n683_ = ~new_n681_ & ~new_n682_;
  assign new_n684_ = \p_input[125]  & ~new_n557_;
  assign new_n685_ = \p_input[109]  & new_n557_;
  assign new_n686_ = ~new_n684_ & ~new_n685_;
  assign new_n687_ = new_n683_ & ~new_n686_;
  assign new_n688_ = ~new_n680_ & ~new_n687_;
  assign new_n689_ = ~new_n679_ & new_n688_;
  assign new_n690_ = ~new_n683_ & new_n686_;
  assign new_n691_ = \p_input[94]  & ~new_n491_;
  assign new_n692_ = \p_input[78]  & new_n491_;
  assign new_n693_ = ~new_n691_ & ~new_n692_;
  assign new_n694_ = \p_input[126]  & ~new_n557_;
  assign new_n695_ = \p_input[110]  & new_n557_;
  assign new_n696_ = ~new_n694_ & ~new_n695_;
  assign new_n697_ = ~new_n693_ & new_n696_;
  assign new_n698_ = ~new_n690_ & ~new_n697_;
  assign new_n699_ = ~new_n689_ & new_n698_;
  assign new_n700_ = new_n693_ & ~new_n696_;
  assign new_n701_ = ~new_n699_ & ~new_n700_;
  assign new_n702_ = ~new_n496_ & ~new_n701_;
  assign new_n703_ = ~new_n495_ & ~new_n702_;
  assign new_n704_ = ~new_n494_ & new_n703_;
  assign new_n705_ = ~new_n560_ & ~new_n703_;
  assign new_n706_ = ~new_n704_ & ~new_n705_;
  assign new_n707_ = new_n430_ & ~new_n706_;
  assign new_n708_ = ~new_n567_ & new_n703_;
  assign new_n709_ = ~new_n564_ & ~new_n703_;
  assign new_n710_ = ~new_n708_ & ~new_n709_;
  assign new_n711_ = ~new_n298_ & new_n427_;
  assign new_n712_ = ~new_n295_ & ~new_n427_;
  assign new_n713_ = ~new_n711_ & ~new_n712_;
  assign new_n714_ = new_n710_ & ~new_n713_;
  assign new_n715_ = ~new_n707_ & new_n714_;
  assign new_n716_ = ~new_n575_ & new_n703_;
  assign new_n717_ = ~new_n572_ & ~new_n703_;
  assign new_n718_ = ~new_n716_ & ~new_n717_;
  assign new_n719_ = ~new_n306_ & new_n427_;
  assign new_n720_ = ~new_n303_ & ~new_n427_;
  assign new_n721_ = ~new_n719_ & ~new_n720_;
  assign new_n722_ = new_n718_ & ~new_n721_;
  assign new_n723_ = ~new_n430_ & new_n706_;
  assign new_n724_ = ~new_n722_ & ~new_n723_;
  assign new_n725_ = ~new_n715_ & new_n724_;
  assign new_n726_ = ~new_n718_ & new_n721_;
  assign new_n727_ = ~new_n313_ & new_n427_;
  assign new_n728_ = ~new_n316_ & ~new_n427_;
  assign new_n729_ = ~new_n727_ & ~new_n728_;
  assign new_n730_ = ~new_n586_ & new_n703_;
  assign new_n731_ = ~new_n583_ & ~new_n703_;
  assign new_n732_ = ~new_n730_ & ~new_n731_;
  assign new_n733_ = new_n729_ & ~new_n732_;
  assign new_n734_ = ~new_n726_ & ~new_n733_;
  assign new_n735_ = ~new_n725_ & new_n734_;
  assign new_n736_ = ~new_n592_ & new_n703_;
  assign new_n737_ = ~new_n595_ & ~new_n703_;
  assign new_n738_ = ~new_n736_ & ~new_n737_;
  assign new_n739_ = ~new_n326_ & new_n427_;
  assign new_n740_ = ~new_n323_ & ~new_n427_;
  assign new_n741_ = ~new_n739_ & ~new_n740_;
  assign new_n742_ = new_n738_ & ~new_n741_;
  assign new_n743_ = ~new_n729_ & new_n732_;
  assign new_n744_ = ~new_n742_ & ~new_n743_;
  assign new_n745_ = ~new_n735_ & new_n744_;
  assign new_n746_ = ~new_n336_ & new_n427_;
  assign new_n747_ = ~new_n333_ & ~new_n427_;
  assign new_n748_ = ~new_n746_ & ~new_n747_;
  assign new_n749_ = ~new_n605_ & new_n703_;
  assign new_n750_ = ~new_n602_ & ~new_n703_;
  assign new_n751_ = ~new_n749_ & ~new_n750_;
  assign new_n752_ = new_n748_ & ~new_n751_;
  assign new_n753_ = ~new_n738_ & new_n741_;
  assign new_n754_ = ~new_n752_ & ~new_n753_;
  assign new_n755_ = ~new_n745_ & new_n754_;
  assign new_n756_ = ~new_n343_ & new_n427_;
  assign new_n757_ = ~new_n346_ & ~new_n427_;
  assign new_n758_ = ~new_n756_ & ~new_n757_;
  assign new_n759_ = ~new_n615_ & new_n703_;
  assign new_n760_ = ~new_n612_ & ~new_n703_;
  assign new_n761_ = ~new_n759_ & ~new_n760_;
  assign new_n762_ = ~new_n758_ & new_n761_;
  assign new_n763_ = ~new_n748_ & new_n751_;
  assign new_n764_ = ~new_n762_ & ~new_n763_;
  assign new_n765_ = ~new_n755_ & new_n764_;
  assign new_n766_ = ~new_n353_ & new_n427_;
  assign new_n767_ = ~new_n356_ & ~new_n427_;
  assign new_n768_ = ~new_n766_ & ~new_n767_;
  assign new_n769_ = ~new_n623_ & new_n703_;
  assign new_n770_ = ~new_n626_ & ~new_n703_;
  assign new_n771_ = ~new_n769_ & ~new_n770_;
  assign new_n772_ = new_n768_ & ~new_n771_;
  assign new_n773_ = new_n758_ & ~new_n761_;
  assign new_n774_ = ~new_n772_ & ~new_n773_;
  assign new_n775_ = ~new_n765_ & new_n774_;
  assign new_n776_ = ~new_n364_ & new_n427_;
  assign new_n777_ = ~new_n367_ & ~new_n427_;
  assign new_n778_ = ~new_n776_ & ~new_n777_;
  assign new_n779_ = ~new_n636_ & new_n703_;
  assign new_n780_ = ~new_n633_ & ~new_n703_;
  assign new_n781_ = ~new_n779_ & ~new_n780_;
  assign new_n782_ = ~new_n778_ & new_n781_;
  assign new_n783_ = ~new_n768_ & new_n771_;
  assign new_n784_ = ~new_n782_ & ~new_n783_;
  assign new_n785_ = ~new_n775_ & new_n784_;
  assign new_n786_ = ~new_n377_ & new_n427_;
  assign new_n787_ = ~new_n374_ & ~new_n427_;
  assign new_n788_ = ~new_n786_ & ~new_n787_;
  assign new_n789_ = ~new_n646_ & new_n703_;
  assign new_n790_ = ~new_n643_ & ~new_n703_;
  assign new_n791_ = ~new_n789_ & ~new_n790_;
  assign new_n792_ = new_n788_ & ~new_n791_;
  assign new_n793_ = new_n778_ & ~new_n781_;
  assign new_n794_ = ~new_n792_ & ~new_n793_;
  assign new_n795_ = ~new_n785_ & new_n794_;
  assign new_n796_ = ~new_n653_ & new_n703_;
  assign new_n797_ = ~new_n656_ & ~new_n703_;
  assign new_n798_ = ~new_n796_ & ~new_n797_;
  assign new_n799_ = ~new_n384_ & new_n427_;
  assign new_n800_ = ~new_n387_ & ~new_n427_;
  assign new_n801_ = ~new_n799_ & ~new_n800_;
  assign new_n802_ = new_n798_ & ~new_n801_;
  assign new_n803_ = ~new_n788_ & new_n791_;
  assign new_n804_ = ~new_n802_ & ~new_n803_;
  assign new_n805_ = ~new_n795_ & new_n804_;
  assign new_n806_ = ~new_n798_ & new_n801_;
  assign new_n807_ = ~new_n393_ & new_n427_;
  assign new_n808_ = ~new_n396_ & ~new_n427_;
  assign new_n809_ = ~new_n807_ & ~new_n808_;
  assign new_n810_ = ~new_n665_ & new_n703_;
  assign new_n811_ = ~new_n662_ & ~new_n703_;
  assign new_n812_ = ~new_n810_ & ~new_n811_;
  assign new_n813_ = new_n809_ & ~new_n812_;
  assign new_n814_ = ~new_n806_ & ~new_n813_;
  assign new_n815_ = ~new_n805_ & new_n814_;
  assign new_n816_ = ~new_n809_ & new_n812_;
  assign new_n817_ = ~new_n672_ & new_n703_;
  assign new_n818_ = ~new_n675_ & ~new_n703_;
  assign new_n819_ = ~new_n817_ & ~new_n818_;
  assign new_n820_ = ~new_n406_ & new_n427_;
  assign new_n821_ = ~new_n403_ & ~new_n427_;
  assign new_n822_ = ~new_n820_ & ~new_n821_;
  assign new_n823_ = new_n819_ & ~new_n822_;
  assign new_n824_ = ~new_n816_ & ~new_n823_;
  assign new_n825_ = ~new_n815_ & new_n824_;
  assign new_n826_ = ~new_n819_ & new_n822_;
  assign new_n827_ = ~new_n683_ & new_n703_;
  assign new_n828_ = ~new_n686_ & ~new_n703_;
  assign new_n829_ = ~new_n827_ & ~new_n828_;
  assign new_n830_ = ~new_n414_ & new_n427_;
  assign new_n831_ = ~new_n417_ & ~new_n427_;
  assign new_n832_ = ~new_n830_ & ~new_n831_;
  assign new_n833_ = ~new_n829_ & new_n832_;
  assign new_n834_ = ~new_n826_ & ~new_n833_;
  assign new_n835_ = ~new_n825_ & new_n834_;
  assign new_n836_ = new_n829_ & ~new_n832_;
  assign new_n837_ = ~new_n693_ & new_n703_;
  assign new_n838_ = ~new_n696_ & ~new_n703_;
  assign new_n839_ = ~new_n837_ & ~new_n838_;
  assign new_n840_ = ~new_n287_ & new_n427_;
  assign new_n841_ = ~new_n284_ & ~new_n427_;
  assign new_n842_ = ~new_n840_ & ~new_n841_;
  assign new_n843_ = new_n839_ & ~new_n842_;
  assign new_n844_ = ~new_n836_ & ~new_n843_;
  assign new_n845_ = ~new_n835_ & new_n844_;
  assign new_n846_ = ~new_n150_ & new_n153_;
  assign new_n847_ = ~new_n839_ & new_n842_;
  assign new_n848_ = ~new_n846_ & ~new_n847_;
  assign new_n849_ = ~new_n845_ & new_n848_;
  assign \o[2]  = ~new_n154_ & ~new_n849_;
  assign new_n851_ = ~new_n703_ & \o[2] ;
  assign new_n852_ = ~new_n427_ & ~\o[2] ;
  assign \o[1]  = new_n851_ | new_n852_;
  assign new_n854_ = new_n491_ & ~\o[1] ;
  assign new_n855_ = new_n557_ & ~new_n703_;
  assign new_n856_ = ~new_n854_ & ~new_n855_;
  assign new_n857_ = \o[2]  & ~new_n856_;
  assign new_n858_ = new_n215_ & ~\o[1] ;
  assign new_n859_ = new_n281_ & ~new_n427_;
  assign new_n860_ = ~new_n858_ & ~new_n859_;
  assign new_n861_ = ~\o[2]  & ~new_n860_;
  assign \o[0]  = ~new_n857_ & ~new_n861_;
  assign new_n863_ = ~new_n713_ & ~\o[2] ;
  assign new_n864_ = ~new_n710_ & \o[2] ;
  assign \o[3]  = new_n863_ | new_n864_;
  assign new_n866_ = ~new_n430_ & ~\o[2] ;
  assign new_n867_ = ~new_n706_ & \o[2] ;
  assign \o[4]  = new_n866_ | new_n867_;
  assign new_n869_ = ~new_n721_ & ~\o[2] ;
  assign new_n870_ = ~new_n718_ & \o[2] ;
  assign \o[5]  = new_n869_ | new_n870_;
  assign new_n872_ = ~new_n732_ & \o[2] ;
  assign new_n873_ = ~new_n729_ & ~\o[2] ;
  assign \o[6]  = new_n872_ | new_n873_;
  assign new_n875_ = ~new_n741_ & ~\o[2] ;
  assign new_n876_ = ~new_n738_ & \o[2] ;
  assign \o[7]  = new_n875_ | new_n876_;
  assign new_n878_ = ~new_n748_ & ~\o[2] ;
  assign new_n879_ = ~new_n751_ & \o[2] ;
  assign \o[8]  = new_n878_ | new_n879_;
  assign new_n881_ = ~new_n761_ & \o[2] ;
  assign new_n882_ = ~new_n758_ & ~\o[2] ;
  assign \o[9]  = new_n881_ | new_n882_;
  assign new_n884_ = ~new_n768_ & ~\o[2] ;
  assign new_n885_ = ~new_n771_ & \o[2] ;
  assign \o[10]  = new_n884_ | new_n885_;
  assign new_n887_ = ~new_n781_ & \o[2] ;
  assign new_n888_ = ~new_n778_ & ~\o[2] ;
  assign \o[11]  = new_n887_ | new_n888_;
  assign new_n890_ = ~new_n788_ & ~\o[2] ;
  assign new_n891_ = ~new_n791_ & \o[2] ;
  assign \o[12]  = new_n890_ | new_n891_;
  assign new_n893_ = new_n801_ & ~\o[2] ;
  assign new_n894_ = new_n798_ & \o[2] ;
  assign \o[13]  = ~new_n893_ & ~new_n894_;
  assign new_n896_ = ~new_n812_ & \o[2] ;
  assign new_n897_ = ~new_n809_ & ~\o[2] ;
  assign \o[14]  = new_n896_ | new_n897_;
  assign new_n899_ = ~new_n822_ & ~\o[2] ;
  assign new_n900_ = ~new_n819_ & \o[2] ;
  assign \o[15]  = new_n899_ | new_n900_;
  assign new_n902_ = new_n832_ & ~\o[2] ;
  assign new_n903_ = new_n829_ & \o[2] ;
  assign \o[16]  = ~new_n902_ & ~new_n903_;
  assign new_n905_ = ~new_n842_ & ~\o[2] ;
  assign new_n906_ = ~new_n839_ & \o[2] ;
  assign \o[17]  = new_n905_ | new_n906_;
  assign \o[18]  = ~new_n150_ | ~new_n153_;
endmodule


