module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173;
  assign n1209 = x88 ^ x2;
  assign n1210 = x93 ^ x28;
  assign n1214 = x91 ^ x44;
  assign n1215 = x90 ^ x52;
  assign n1216 = ~n1214 & n1215;
  assign n1217 = n1216 ^ n1215;
  assign n1211 = x89 ^ x60;
  assign n1212 = x92 ^ x36;
  assign n1213 = n1211 & ~n1212;
  assign n1220 = n1213 ^ n1212;
  assign n1237 = n1217 & ~n1220;
  assign n1228 = n1220 ^ n1211;
  assign n1218 = n1217 ^ n1214;
  assign n1233 = n1218 ^ n1215;
  assign n1234 = n1228 & ~n1233;
  assign n1238 = n1237 ^ n1234;
  assign n1239 = n1238 ^ n1220;
  assign n1229 = n1216 & n1228;
  assign n1223 = n1213 ^ n1211;
  assign n1224 = n1217 & n1223;
  assign n1230 = n1229 ^ n1224;
  assign n1231 = n1230 ^ n1216;
  assign n1226 = n1216 & n1223;
  assign n1222 = n1213 & n1216;
  assign n1225 = n1224 ^ n1222;
  assign n1227 = n1226 ^ n1225;
  assign n1232 = n1231 ^ n1227;
  assign n1235 = n1234 ^ n1232;
  assign n1221 = n1218 & ~n1220;
  assign n1236 = n1235 ^ n1221;
  assign n1240 = n1239 ^ n1236;
  assign n1871 = n1240 ^ n1229;
  assign n1250 = n1211 & n1214;
  assign n1251 = n1250 ^ n1224;
  assign n1247 = n1223 ^ n1222;
  assign n1242 = n1213 & ~n1233;
  assign n1243 = n1242 ^ n1237;
  assign n1244 = n1243 ^ n1233;
  assign n1241 = n1240 ^ n1238;
  assign n1245 = n1244 ^ n1241;
  assign n1246 = n1245 ^ n1227;
  assign n1248 = n1247 ^ n1246;
  assign n1219 = n1213 & n1218;
  assign n1249 = n1248 ^ n1219;
  assign n1252 = n1251 ^ n1249;
  assign n1266 = n1252 ^ n1226;
  assign n1872 = n1871 ^ n1266;
  assign n1873 = ~n1210 & ~n1872;
  assign n1874 = n1873 ^ n1266;
  assign n1875 = n1209 & n1874;
  assign n2034 = n1209 & n1249;
  assign n1258 = n1209 & ~n1210;
  assign n1267 = n1258 ^ n1210;
  assign n2035 = n1246 & ~n1267;
  assign n1268 = n1267 ^ n1209;
  assign n1269 = n1266 & n1268;
  assign n1259 = n1258 ^ n1209;
  assign n1261 = n1221 ^ n1218;
  assign n1262 = n1261 ^ n1249;
  assign n1263 = n1262 ^ n1228;
  assign n1260 = n1234 ^ n1229;
  assign n1264 = n1263 ^ n1260;
  assign n1265 = n1259 & n1264;
  assign n1270 = n1269 ^ n1265;
  assign n2036 = n1234 & ~n1267;
  assign n1892 = n1210 ^ n1209;
  assign n1283 = n1264 ^ n1245;
  assign n2043 = n1283 ^ n1252;
  assign n2044 = n2043 ^ n1221;
  assign n1285 = n1262 ^ n1232;
  assign n2041 = n1285 ^ n1243;
  assign n2042 = n2041 ^ n1283;
  assign n2045 = n2044 ^ n2042;
  assign n2046 = n1209 & n2045;
  assign n2047 = n2046 ^ n2042;
  assign n1882 = n1262 ^ n1221;
  assign n2037 = n1882 ^ n1242;
  assign n2038 = n2037 ^ n1236;
  assign n2039 = ~n1209 & n2038;
  assign n2040 = n2039 ^ n1236;
  assign n2048 = n2047 ^ n2040;
  assign n2049 = n1892 & n2048;
  assign n2050 = n2049 ^ n2040;
  assign n2051 = ~n2036 & ~n2050;
  assign n2052 = ~n1270 & n2051;
  assign n2053 = ~n2035 & n2052;
  assign n2054 = ~n2034 & n2053;
  assign n2055 = ~n1875 & n2054;
  assign n2056 = n2055 ^ x63;
  assign n2057 = n2056 ^ x147;
  assign n1127 = x82 ^ x34;
  assign n1136 = x83 ^ x26;
  assign n1132 = x85 ^ x10;
  assign n1165 = n1136 ^ n1132;
  assign n1129 = x84 ^ x18;
  assign n1166 = n1165 ^ n1129;
  assign n1167 = n1166 ^ n1136;
  assign n1160 = n1129 & ~n1136;
  assign n1168 = n1160 ^ n1129;
  assign n1130 = x86 ^ x2;
  assign n1169 = n1168 ^ n1130;
  assign n1170 = n1167 & ~n1169;
  assign n1171 = n1170 ^ n1165;
  assign n1144 = n1132 ^ n1130;
  assign n1145 = ~n1130 & n1144;
  assign n1146 = n1145 ^ n1129;
  assign n1149 = ~n1136 & ~n1146;
  assign n1150 = n1149 ^ n1144;
  assign n2061 = n1171 ^ n1150;
  assign n2062 = ~n1127 & n2061;
  assign n2063 = n2062 ^ n1150;
  assign n1126 = x87 ^ x60;
  assign n2066 = n2063 ^ n1126;
  assign n1158 = n1136 ^ n1130;
  assign n1133 = n1129 & ~n1132;
  assign n1137 = n1133 ^ n1132;
  assign n1159 = n1137 ^ n1129;
  assign n1161 = n1160 ^ n1159;
  assign n1162 = ~n1158 & n1161;
  assign n1163 = n1162 ^ n1160;
  assign n1152 = n1136 ^ n1129;
  assign n1153 = n1144 ^ n1136;
  assign n1154 = ~n1152 & ~n1153;
  assign n1138 = ~n1130 & ~n1137;
  assign n1139 = n1138 ^ n1137;
  assign n1134 = n1133 ^ n1129;
  assign n1140 = n1139 ^ n1134;
  assign n1141 = n1140 ^ n1133;
  assign n1155 = n1154 ^ n1141;
  assign n1142 = ~n1136 & ~n1141;
  assign n1143 = n1142 ^ n1133;
  assign n1147 = n1146 ^ n1133;
  assign n1148 = ~n1143 & ~n1147;
  assign n1151 = n1150 ^ n1148;
  assign n1156 = n1155 ^ n1151;
  assign n1157 = n1156 ^ n1138;
  assign n1164 = n1163 ^ n1157;
  assign n2058 = n1164 ^ n1148;
  assign n2059 = n1127 & ~n2058;
  assign n2060 = n2059 ^ n1148;
  assign n2064 = n2063 ^ n2060;
  assign n2065 = n1126 & n2064;
  assign n2067 = n2066 ^ n2065;
  assign n2068 = n2067 ^ x37;
  assign n2069 = n2068 ^ x142;
  assign n2070 = ~n2057 & ~n2069;
  assign n2071 = n2070 ^ n2057;
  assign n2072 = n2071 ^ n2069;
  assign n1517 = x106 ^ x38;
  assign n1518 = x111 ^ x56;
  assign n1519 = n1518 ^ n1517;
  assign n1520 = ~n1517 & ~n1519;
  assign n1521 = n1520 ^ n1517;
  assign n1523 = x109 ^ x14;
  assign n1524 = x108 ^ x22;
  assign n1525 = n1523 & n1524;
  assign n1526 = n1525 ^ n1523;
  assign n1528 = x110 ^ x6;
  assign n1529 = x107 ^ x30;
  assign n1530 = n1528 & ~n1529;
  assign n1547 = n1526 & n1530;
  assign n1531 = n1530 ^ n1529;
  assign n1527 = n1526 ^ n1524;
  assign n1544 = n1527 ^ n1523;
  assign n1545 = ~n1531 & n1544;
  assign n1543 = ~n1527 & n1530;
  assign n1546 = n1545 ^ n1543;
  assign n1548 = n1547 ^ n1546;
  assign n1536 = n1529 ^ n1528;
  assign n1537 = n1536 ^ n1524;
  assign n1538 = n1529 ^ n1523;
  assign n1539 = n1538 ^ n1524;
  assign n1540 = n1523 & n1539;
  assign n1541 = n1540 ^ n1538;
  assign n1542 = n1537 & ~n1541;
  assign n1549 = n1548 ^ n1542;
  assign n1532 = n1531 ^ n1528;
  assign n1550 = n1549 ^ n1532;
  assign n1534 = n1525 & n1532;
  assign n1533 = ~n1527 & n1532;
  assign n1535 = n1534 ^ n1533;
  assign n1551 = n1550 ^ n1535;
  assign n1573 = n1551 ^ n1545;
  assign n2073 = ~n1521 & n1573;
  assign n1561 = n1530 ^ n1528;
  assign n1564 = ~n1527 & n1561;
  assign n1565 = n1564 ^ n1561;
  assign n1562 = n1526 & n1561;
  assign n1555 = n1528 ^ n1524;
  assign n1556 = ~n1536 & ~n1555;
  assign n1557 = ~n1523 & n1556;
  assign n1554 = ~n1527 & ~n1531;
  assign n1558 = n1557 ^ n1554;
  assign n1563 = n1562 ^ n1558;
  assign n1566 = n1565 ^ n1563;
  assign n1567 = n1566 ^ n1549;
  assign n1583 = ~n1521 & n1567;
  assign n1607 = n1562 ^ n1534;
  assign n2074 = ~n1519 & n1607;
  assign n2075 = n1557 ^ n1555;
  assign n2076 = ~n1518 & ~n2075;
  assign n1571 = n1525 & ~n1531;
  assign n2077 = n2076 ^ n1571;
  assign n2078 = n2077 ^ n1564;
  assign n2079 = n2077 ^ n1517;
  assign n2080 = ~n2077 & ~n2079;
  assign n2081 = n2080 ^ n2077;
  assign n2082 = n2078 & ~n2081;
  assign n2083 = n2082 ^ n2080;
  assign n2084 = n2083 ^ n2077;
  assign n2085 = n2084 ^ n1517;
  assign n2086 = ~n2074 & ~n2085;
  assign n2087 = n2086 ^ n2074;
  assign n1587 = n1548 ^ n1529;
  assign n1572 = n1558 ^ n1544;
  assign n1574 = n1573 ^ n1572;
  assign n1577 = n1574 ^ n1530;
  assign n1576 = n1548 ^ n1545;
  assign n1578 = n1577 ^ n1576;
  assign n1579 = n1578 ^ n1554;
  assign n1575 = n1574 ^ n1571;
  assign n1580 = n1579 ^ n1575;
  assign n1588 = n1587 ^ n1580;
  assign n2093 = n1588 ^ n1545;
  assign n2094 = ~n1519 & ~n2093;
  assign n2091 = n1520 & n1576;
  assign n1559 = n1558 ^ n1533;
  assign n2090 = ~n1517 & n1559;
  assign n2092 = n2091 ^ n2090;
  assign n2095 = n2094 ^ n2092;
  assign n1599 = n1578 ^ n1547;
  assign n2088 = ~n1521 & n1599;
  assign n1522 = n1521 ^ n1518;
  assign n1904 = n1574 ^ n1554;
  assign n1905 = ~n1522 & n1904;
  assign n2089 = n2088 ^ n1905;
  assign n2096 = n2095 ^ n2089;
  assign n2097 = ~n2087 & ~n2096;
  assign n2098 = ~n1583 & n2097;
  assign n2099 = ~n2073 & n2098;
  assign n2100 = n2099 ^ x29;
  assign n2101 = n2100 ^ x143;
  assign n1033 = x65 ^ x56;
  assign n1034 = x68 ^ x32;
  assign n1035 = ~n1033 & ~n1034;
  assign n1036 = n1035 ^ n1033;
  assign n1037 = x67 ^ x40;
  assign n1038 = x66 ^ x48;
  assign n1039 = ~n1037 & ~n1038;
  assign n1041 = n1039 ^ n1038;
  assign n1044 = ~n1036 & ~n1041;
  assign n1067 = x69 ^ x24;
  assign n1068 = x64 ^ x6;
  assign n1086 = ~n1067 & n1068;
  assign n1096 = n1086 ^ n1067;
  assign n1101 = n1044 & ~n1096;
  assign n1083 = n1034 & ~n1037;
  assign n1084 = n1083 ^ n1039;
  assign n1062 = n1036 ^ n1034;
  assign n1076 = ~n1041 & ~n1062;
  assign n1069 = n1062 ^ n1033;
  assign n1080 = n1076 ^ n1069;
  assign n1063 = n1041 ^ n1037;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = n1064 ^ n1063;
  assign n1056 = n1035 & n1039;
  assign n1045 = n1039 ^ n1037;
  assign n1046 = ~n1036 & ~n1045;
  assign n1057 = n1056 ^ n1046;
  assign n1042 = n1035 & ~n1041;
  assign n1047 = n1046 ^ n1042;
  assign n1058 = n1057 ^ n1047;
  assign n1059 = n1058 ^ n1035;
  assign n1051 = n1037 ^ n1033;
  assign n1052 = n1051 ^ n1038;
  assign n1053 = ~n1033 & ~n1052;
  assign n1054 = n1053 ^ n1033;
  assign n1048 = n1047 ^ n1044;
  assign n1055 = n1054 ^ n1048;
  assign n1060 = n1059 ^ n1055;
  assign n1049 = n1048 ^ n1036;
  assign n1040 = ~n1036 & n1039;
  assign n1043 = n1042 ^ n1040;
  assign n1050 = n1049 ^ n1043;
  assign n1061 = n1060 ^ n1050;
  assign n1066 = n1065 ^ n1061;
  assign n1077 = n1076 ^ n1066;
  assign n1075 = ~n1045 & ~n1069;
  assign n1078 = n1077 ^ n1075;
  assign n1070 = ~n1041 & ~n1069;
  assign n1079 = n1078 ^ n1070;
  assign n1081 = n1080 ^ n1079;
  assign n1082 = n1081 ^ n1057;
  assign n1085 = n1084 ^ n1082;
  assign n1087 = n1068 ^ n1067;
  assign n1088 = n1087 ^ n1086;
  assign n1089 = n1088 ^ n1067;
  assign n1090 = n1085 & n1089;
  assign n1991 = n1085 ^ n1075;
  assign n2102 = ~n1096 & n1991;
  assign n1091 = n1081 & n1089;
  assign n2103 = n2102 ^ n1091;
  assign n1971 = n1047 & n1089;
  assign n1106 = n1055 ^ n1040;
  assign n2104 = n1068 & ~n1106;
  assign n1093 = n1056 ^ n1044;
  assign n2105 = n1086 & n1093;
  assign n2114 = n1077 ^ n1049;
  assign n2113 = n1064 ^ n1060;
  assign n2115 = n2114 ^ n2113;
  assign n2116 = ~n1068 & ~n2115;
  assign n2117 = n2116 ^ n2113;
  assign n1097 = n1070 ^ n1064;
  assign n1992 = n1991 ^ n1097;
  assign n2108 = n1992 ^ n1056;
  assign n1110 = n1061 ^ n1044;
  assign n2109 = n2108 ^ n1110;
  assign n2106 = n1097 ^ n1066;
  assign n1977 = n1078 ^ n1064;
  assign n1994 = n1977 ^ n1062;
  assign n1985 = n1085 ^ n1066;
  assign n1986 = n1985 ^ n1075;
  assign n1995 = n1994 ^ n1986;
  assign n2107 = n2106 ^ n1995;
  assign n2110 = n2109 ^ n2107;
  assign n2111 = ~n1068 & n2110;
  assign n2112 = n2111 ^ n2107;
  assign n2118 = n2117 ^ n2112;
  assign n2119 = n1087 & ~n2118;
  assign n2120 = n2119 ^ n2117;
  assign n2121 = ~n2105 & n2120;
  assign n2122 = ~n2104 & n2121;
  assign n2123 = ~n1971 & n2122;
  assign n2124 = ~n2103 & n2123;
  assign n2125 = ~n1090 & n2124;
  assign n2126 = ~n1101 & n2125;
  assign n2127 = n2126 ^ x13;
  assign n2128 = n2127 ^ x145;
  assign n2129 = ~n2101 & ~n2128;
  assign n2130 = n2129 ^ n2128;
  assign n833 = x105 ^ x30;
  assign n834 = x100 ^ x4;
  assign n838 = x103 ^ x46;
  assign n839 = x101 ^ x62;
  assign n840 = ~n838 & ~n839;
  assign n835 = x102 ^ x54;
  assign n836 = x104 ^ x38;
  assign n837 = ~n835 & ~n836;
  assign n844 = n837 ^ n835;
  assign n845 = n844 ^ n836;
  assign n849 = n845 ^ n835;
  assign n850 = n840 & ~n849;
  assign n846 = n840 & ~n845;
  assign n843 = n837 & n840;
  assign n847 = n846 ^ n843;
  assign n848 = n847 ^ n840;
  assign n851 = n850 ^ n848;
  assign n841 = n840 ^ n839;
  assign n842 = n837 & ~n841;
  assign n852 = n851 ^ n842;
  assign n853 = ~n834 & n852;
  assign n854 = n853 ^ n851;
  assign n855 = n833 & n854;
  assign n856 = ~n833 & ~n834;
  assign n857 = n856 ^ n834;
  assign n881 = ~n841 & ~n844;
  assign n1710 = ~n857 & n881;
  assign n906 = n846 ^ n842;
  assign n1716 = n906 ^ n848;
  assign n1717 = n834 & n1716;
  assign n1718 = n1717 ^ n848;
  assign n1719 = ~n833 & n1718;
  assign n861 = n841 ^ n838;
  assign n921 = ~n857 & ~n861;
  assign n2132 = ~n845 & n921;
  assign n862 = n861 ^ n839;
  assign n863 = n837 & ~n862;
  assign n864 = n863 ^ n848;
  assign n858 = n839 ^ n835;
  assign n859 = n858 ^ n836;
  assign n860 = ~n838 & n859;
  assign n865 = n864 ^ n860;
  assign n896 = n856 ^ n833;
  assign n897 = n896 ^ n834;
  assign n898 = n865 & ~n897;
  assign n2133 = n2132 ^ n898;
  assign n873 = ~n841 & ~n845;
  assign n874 = n873 ^ n861;
  assign n867 = n839 ^ n838;
  assign n868 = n838 ^ n836;
  assign n869 = ~n835 & ~n868;
  assign n870 = n869 ^ n836;
  assign n871 = n867 & n870;
  assign n872 = n871 ^ n839;
  assign n875 = n874 ^ n872;
  assign n866 = n865 ^ n863;
  assign n876 = n875 ^ n866;
  assign n877 = n876 ^ n862;
  assign n878 = n877 ^ n875;
  assign n879 = ~n857 & ~n878;
  assign n2134 = n873 ^ n843;
  assign n2135 = ~n897 & n2134;
  assign n891 = n834 ^ n833;
  assign n902 = n836 ^ n835;
  assign n903 = ~n861 & n902;
  assign n904 = n903 ^ n861;
  assign n2142 = n904 ^ n877;
  assign n2136 = n866 ^ n833;
  assign n2137 = n891 & n2136;
  assign n2138 = n2137 ^ n833;
  assign n2139 = ~n876 & ~n2138;
  assign n2140 = n2139 ^ n875;
  assign n2141 = ~n903 & n2140;
  assign n2143 = n2142 ^ n2141;
  assign n2144 = n2143 ^ n2141;
  assign n2145 = ~n833 & ~n2144;
  assign n2146 = n2145 ^ n2141;
  assign n2147 = n891 & ~n2146;
  assign n2148 = n2147 ^ n2141;
  assign n2149 = ~n2135 & n2148;
  assign n2150 = n873 ^ n863;
  assign n882 = n881 ^ n842;
  assign n2151 = n2150 ^ n882;
  assign n2152 = n2151 ^ n882;
  assign n2153 = n897 & n2152;
  assign n2154 = n2153 ^ n882;
  assign n2155 = ~n856 & n2154;
  assign n2156 = n2155 ^ n882;
  assign n2157 = n2149 & ~n2156;
  assign n2158 = n833 & n865;
  assign n883 = n882 ^ n838;
  assign n884 = n883 ^ n874;
  assign n2159 = n2158 ^ n884;
  assign n2160 = ~n834 & ~n2159;
  assign n2161 = n2160 ^ n884;
  assign n2162 = n2157 & n2161;
  assign n2163 = ~n879 & n2162;
  assign n2164 = ~n2133 & n2163;
  assign n2165 = ~n1719 & n2164;
  assign n2166 = ~n1710 & n2165;
  assign n2167 = ~n855 & n2166;
  assign n2168 = n2167 ^ x21;
  assign n2169 = n2168 ^ x144;
  assign n1618 = x81 ^ x26;
  assign n1617 = x76 ^ x0;
  assign n1627 = x79 ^ x42;
  assign n1628 = x77 ^ x58;
  assign n1629 = ~n1627 & n1628;
  assign n1630 = n1629 ^ n1627;
  assign n1623 = x78 ^ x50;
  assign n1624 = x80 ^ x34;
  assign n1625 = n1623 & ~n1624;
  assign n1626 = n1625 ^ n1623;
  assign n1635 = n1626 ^ n1624;
  assign n1655 = n1635 ^ n1623;
  assign n1666 = ~n1630 & ~n1655;
  assign n1632 = n1630 ^ n1628;
  assign n1636 = n1632 & n1635;
  assign n1689 = n1666 ^ n1636;
  assign n1667 = n1666 ^ n1655;
  assign n1656 = n1629 & ~n1655;
  assign n1638 = n1626 & n1632;
  assign n1639 = n1638 ^ n1632;
  assign n1633 = n1625 & n1632;
  assign n1637 = n1636 ^ n1633;
  assign n1640 = n1639 ^ n1637;
  assign n1665 = n1656 ^ n1640;
  assign n1668 = n1667 ^ n1665;
  assign n1648 = n1638 ^ n1626;
  assign n1646 = n1626 & n1629;
  assign n1631 = n1626 & ~n1630;
  assign n1647 = n1646 ^ n1631;
  assign n1649 = n1648 ^ n1647;
  assign n1669 = n1668 ^ n1649;
  assign n2170 = n1689 ^ n1669;
  assign n2171 = n1617 & ~n2170;
  assign n2172 = n2171 ^ n1669;
  assign n2173 = n1618 & ~n2172;
  assign n1679 = n1618 ^ n1617;
  assign n2174 = n1656 & ~n1679;
  assign n1619 = ~n1617 & ~n1618;
  assign n1620 = n1619 ^ n1618;
  assign n1621 = n1620 ^ n1617;
  assign n1622 = n1621 ^ n1618;
  assign n1684 = n1620 & n1646;
  assign n1831 = n1684 ^ n1631;
  assign n1832 = n1622 & n1831;
  assign n1833 = n1832 ^ n1631;
  assign n2175 = n2174 ^ n1833;
  assign n1673 = n1656 ^ n1628;
  assign n1670 = n1669 ^ n1646;
  assign n1660 = n1632 ^ n1627;
  assign n1661 = n1625 & n1660;
  assign n1671 = n1670 ^ n1661;
  assign n1657 = n1656 ^ n1646;
  assign n1658 = n1657 ^ n1629;
  assign n1672 = n1671 ^ n1658;
  assign n1674 = n1673 ^ n1672;
  assign n1675 = n1620 & ~n1674;
  assign n1651 = n1624 & ~n1627;
  assign n1652 = n1651 ^ n1626;
  assign n1653 = n1652 ^ n1638;
  assign n1642 = n1627 ^ n1624;
  assign n1643 = ~n1628 & ~n1642;
  assign n1644 = n1643 ^ n1628;
  assign n1634 = n1633 ^ n1631;
  assign n1641 = n1640 ^ n1634;
  assign n1645 = n1644 ^ n1641;
  assign n1650 = n1649 ^ n1645;
  assign n1654 = n1653 ^ n1650;
  assign n1659 = n1658 ^ n1654;
  assign n1662 = n1661 ^ n1659;
  assign n1663 = n1662 ^ n1625;
  assign n1664 = n1663 ^ n1633;
  assign n1676 = n1675 ^ n1664;
  assign n1677 = n1622 & ~n1676;
  assign n1678 = n1677 ^ n1664;
  assign n2176 = n1633 ^ n1622;
  assign n2177 = n1645 ^ n1640;
  assign n2178 = n2177 ^ n1620;
  assign n2179 = ~n1633 & ~n2178;
  assign n2180 = n2179 ^ n1620;
  assign n2181 = ~n2176 & ~n2180;
  assign n2182 = n2181 ^ n1622;
  assign n2184 = n1622 & n1661;
  assign n2183 = n1669 ^ n1658;
  assign n2185 = n2184 ^ n2183;
  assign n2186 = n1620 & ~n2185;
  assign n2187 = n2186 ^ n2183;
  assign n2188 = n2182 & n2187;
  assign n2189 = n1678 & n2188;
  assign n2190 = ~n2175 & n2189;
  assign n2191 = n1656 ^ n1638;
  assign n2192 = n1622 & n2191;
  assign n2193 = n2192 ^ n1656;
  assign n2194 = n2190 & ~n2193;
  assign n2195 = ~n1664 & ~n1679;
  assign n2196 = n1640 ^ n1631;
  assign n2197 = n1617 & n2196;
  assign n2198 = n2197 ^ n1631;
  assign n2199 = n2198 ^ n1645;
  assign n2200 = n2198 ^ n1618;
  assign n2201 = ~n2198 & n2200;
  assign n2202 = n2201 ^ n2198;
  assign n2203 = ~n2199 & ~n2202;
  assign n2204 = n2203 ^ n2201;
  assign n2205 = n2204 ^ n2198;
  assign n2206 = n2205 ^ n1618;
  assign n2207 = ~n2195 & n2206;
  assign n2208 = n2207 ^ n2195;
  assign n2209 = n2194 & ~n2208;
  assign n2210 = ~n2173 & n2209;
  assign n2211 = n2210 ^ x5;
  assign n2212 = n2211 ^ x146;
  assign n2213 = n2169 & n2212;
  assign n2216 = n2213 ^ n2169;
  assign n2219 = ~n2130 & n2216;
  assign n2131 = n2130 ^ n2101;
  assign n2249 = n2219 ^ n2131;
  assign n2240 = n2212 ^ n2169;
  assign n2241 = n2129 & n2240;
  assign n2228 = n2129 ^ n2101;
  assign n2229 = n2216 & ~n2228;
  assign n2242 = n2241 ^ n2229;
  assign n2233 = ~n2131 & n2213;
  assign n2234 = n2233 ^ n2213;
  assign n2231 = n2129 & n2213;
  assign n2221 = ~n2130 & n2213;
  assign n2232 = n2231 ^ n2221;
  assign n2235 = n2234 ^ n2232;
  assign n2214 = n2213 ^ n2212;
  assign n2225 = n2129 & n2214;
  assign n2226 = n2225 ^ n2214;
  assign n2222 = n2221 ^ n2130;
  assign n2217 = n2216 ^ n2212;
  assign n2218 = ~n2130 & ~n2217;
  assign n2220 = n2219 ^ n2218;
  assign n2223 = n2222 ^ n2220;
  assign n2215 = ~n2131 & n2214;
  assign n2224 = n2223 ^ n2215;
  assign n2227 = n2226 ^ n2224;
  assign n2230 = n2229 ^ n2227;
  assign n2236 = n2235 ^ n2230;
  assign n2237 = n2236 ^ n2228;
  assign n2238 = n2237 ^ n2225;
  assign n2239 = n2238 ^ n2219;
  assign n2243 = n2242 ^ n2239;
  assign n2244 = n2243 ^ n2216;
  assign n2245 = n2244 ^ n2237;
  assign n2246 = n2245 ^ n2215;
  assign n2247 = n2246 ^ n2219;
  assign n2248 = n2247 ^ n2233;
  assign n2250 = n2249 ^ n2248;
  assign n2251 = n2250 ^ n2223;
  assign n2252 = ~n2072 & n2251;
  assign n2253 = ~n2072 & n2237;
  assign n2254 = n2072 ^ n2070;
  assign n2257 = n2241 ^ n2129;
  assign n2258 = n2257 ^ n2231;
  assign n2255 = n2241 ^ n2225;
  assign n2256 = ~n2057 & n2255;
  assign n2259 = n2258 ^ n2256;
  assign n2260 = ~n2254 & n2259;
  assign n2261 = n2260 ^ n2258;
  assign n2262 = ~n2253 & ~n2261;
  assign n2289 = n2258 ^ n2227;
  assign n3721 = n2070 & n2289;
  assign n3722 = n2250 & n3721;
  assign n3723 = n3722 ^ n2070;
  assign n2810 = n2221 & ~n2254;
  assign n3724 = n2255 ^ n2235;
  assign n3725 = n3724 ^ n2219;
  assign n3726 = n2069 & n3725;
  assign n3727 = n3726 ^ n2219;
  assign n3728 = n2057 & n3727;
  assign n2263 = n2070 ^ n2069;
  assign n2264 = n2263 ^ n2231;
  assign n2265 = n2245 ^ n2071;
  assign n2266 = ~n2231 & n2265;
  assign n2267 = n2266 ^ n2071;
  assign n2268 = ~n2264 & ~n2267;
  assign n2269 = n2268 ^ n2263;
  assign n3729 = n2218 ^ n2072;
  assign n3730 = n2215 ^ n2070;
  assign n3731 = ~n2218 & ~n3730;
  assign n3732 = n3731 ^ n2070;
  assign n3733 = ~n3729 & n3732;
  assign n3734 = n3733 ^ n2072;
  assign n3735 = n2263 ^ n2230;
  assign n3736 = n2251 ^ n2071;
  assign n3737 = n2230 & n3736;
  assign n3738 = n3737 ^ n2071;
  assign n3739 = n3735 & ~n3738;
  assign n3740 = n3739 ^ n2263;
  assign n3741 = n2069 & n2248;
  assign n3742 = n3741 ^ n2233;
  assign n3743 = n3742 ^ n2225;
  assign n3744 = n3742 ^ n2057;
  assign n3745 = ~n3742 & n3744;
  assign n3746 = n3745 ^ n3742;
  assign n3747 = n3743 & ~n3746;
  assign n3748 = n3747 ^ n3745;
  assign n3749 = n3748 ^ n3742;
  assign n3750 = n3749 ^ n2057;
  assign n3751 = n3740 & n3750;
  assign n3752 = n3751 ^ n3740;
  assign n3753 = n3734 & n3752;
  assign n3754 = n2269 & n3753;
  assign n3755 = ~n3728 & n3754;
  assign n3756 = ~n2810 & n3755;
  assign n3757 = ~n3723 & n3756;
  assign n3758 = n2262 & n3757;
  assign n3759 = ~n2252 & n3758;
  assign n3760 = n3759 ^ x30;
  assign n3761 = n3760 ^ x201;
  assign n1253 = n1252 ^ n1248;
  assign n1254 = n1253 ^ n1240;
  assign n1255 = ~n1210 & ~n1254;
  assign n1256 = n1255 ^ n1240;
  assign n1257 = ~n1209 & ~n1256;
  assign n1271 = ~n1209 & ~n1241;
  assign n1272 = n1271 ^ n1240;
  assign n1273 = n1210 & ~n1272;
  assign n1274 = n1260 ^ n1259;
  assign n1275 = n1267 ^ n1221;
  assign n1276 = ~n1260 & n1275;
  assign n1277 = n1276 ^ n1267;
  assign n1278 = n1274 & ~n1277;
  assign n1279 = n1278 ^ n1259;
  assign n1292 = n1243 ^ n1225;
  assign n1293 = n1292 ^ n1261;
  assign n1294 = ~n1210 & n1293;
  assign n1295 = n1294 ^ n1261;
  assign n1280 = n1248 ^ n1222;
  assign n1281 = ~n1258 & ~n1280;
  assign n1282 = ~n1245 & n1281;
  assign n1288 = n1259 & n1280;
  assign n1286 = n1285 ^ n1219;
  assign n1287 = n1286 ^ n1230;
  assign n1289 = n1288 ^ n1287;
  assign n1284 = n1283 ^ n1242;
  assign n1290 = n1289 ^ n1284;
  assign n1291 = ~n1282 & n1290;
  assign n1296 = n1295 ^ n1291;
  assign n1297 = ~n1209 & n1296;
  assign n1298 = n1297 ^ n1291;
  assign n1299 = ~n1279 & ~n1298;
  assign n1300 = ~n1273 & n1299;
  assign n1301 = ~n1270 & n1300;
  assign n1302 = ~n1257 & n1301;
  assign n1303 = n1302 ^ x1;
  assign n1304 = n1303 ^ x124;
  assign n1305 = x73 ^ x8;
  assign n1306 = x71 ^ x24;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = n1307 ^ n1306;
  assign n1309 = x74 ^ x0;
  assign n1310 = x72 ^ x16;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = n1311 ^ n1309;
  assign n1313 = n1312 ^ n1310;
  assign n1314 = ~n1308 & ~n1313;
  assign n1315 = x75 ^ x58;
  assign n1316 = x70 ^ x32;
  assign n1317 = ~n1315 & n1316;
  assign n1318 = n1317 ^ n1316;
  assign n1319 = n1314 & n1318;
  assign n1320 = n1309 ^ n1305;
  assign n1321 = n1306 & n1320;
  assign n1326 = n1308 ^ n1305;
  assign n1343 = n1311 & ~n1326;
  assign n1344 = n1343 ^ n1326;
  assign n1327 = n1326 ^ n1306;
  assign n1328 = ~n1312 & ~n1327;
  assign n1332 = n1328 ^ n1314;
  assign n1331 = n1311 & ~n1327;
  assign n1333 = n1332 ^ n1331;
  assign n1322 = n1313 ^ n1309;
  assign n1330 = ~n1322 & ~n1326;
  assign n1334 = n1333 ^ n1330;
  assign n1335 = n1334 ^ n1320;
  assign n1324 = n1310 ^ n1306;
  assign n1325 = ~n1320 & ~n1324;
  assign n1329 = n1328 ^ n1325;
  assign n1336 = n1335 ^ n1329;
  assign n1340 = n1336 ^ n1312;
  assign n1338 = ~n1308 & ~n1312;
  assign n1339 = n1338 ^ n1328;
  assign n1341 = n1340 ^ n1339;
  assign n1342 = n1341 ^ n1330;
  assign n1345 = n1344 ^ n1342;
  assign n1323 = ~n1308 & ~n1322;
  assign n1337 = n1336 ^ n1323;
  assign n1346 = n1345 ^ n1337;
  assign n1347 = n1346 ^ n1335;
  assign n1348 = n1347 ^ n1322;
  assign n1349 = ~n1321 & n1348;
  assign n1350 = n1349 ^ n1348;
  assign n1351 = n1350 ^ n1343;
  assign n1352 = n1318 ^ n1315;
  assign n1353 = n1351 & n1352;
  assign n1358 = ~n1308 & n1311;
  assign n1357 = n1307 & ~n1313;
  assign n1359 = n1358 ^ n1357;
  assign n1360 = ~n1316 & n1359;
  assign n1354 = n1342 ^ n1314;
  assign n1355 = n1316 & n1354;
  assign n1356 = n1355 ^ n1314;
  assign n1361 = n1360 ^ n1356;
  assign n1362 = n1315 & n1361;
  assign n1363 = n1362 ^ n1356;
  assign n1364 = n1347 ^ n1314;
  assign n1365 = n1364 ^ n1338;
  assign n1366 = n1316 & ~n1365;
  assign n1367 = n1366 ^ n1338;
  assign n1368 = ~n1315 & n1367;
  assign n1369 = n1316 ^ n1315;
  assign n1371 = n1357 ^ n1347;
  assign n1370 = n1336 ^ n1307;
  assign n1372 = n1371 ^ n1370;
  assign n1373 = n1372 ^ n1337;
  assign n1374 = n1315 & ~n1373;
  assign n1375 = n1374 ^ n1372;
  assign n1376 = ~n1369 & n1375;
  assign n1387 = n1317 ^ n1315;
  assign n1388 = n1336 ^ n1321;
  assign n1389 = ~n1387 & ~n1388;
  assign n1379 = n1351 ^ n1338;
  assign n1380 = n1379 ^ n1371;
  assign n1381 = n1380 ^ n1333;
  assign n1382 = n1381 ^ n1358;
  assign n1377 = n1372 ^ n1342;
  assign n1378 = n1377 ^ n1346;
  assign n1383 = n1382 ^ n1378;
  assign n1384 = n1383 ^ n1359;
  assign n1385 = n1384 ^ n1331;
  assign n1386 = n1317 & n1385;
  assign n1390 = n1389 ^ n1386;
  assign n1391 = n1383 ^ n1328;
  assign n1392 = n1391 ^ n1379;
  assign n1393 = n1392 ^ n1325;
  assign n1394 = ~n1316 & n1393;
  assign n1395 = n1394 ^ n1392;
  assign n1396 = n1315 & n1395;
  assign n1397 = ~n1390 & ~n1396;
  assign n1398 = ~n1376 & n1397;
  assign n1399 = ~n1368 & n1398;
  assign n1400 = ~n1363 & n1399;
  assign n1401 = ~n1353 & n1400;
  assign n1402 = ~n1319 & n1401;
  assign n1403 = n1402 ^ x27;
  assign n1404 = n1403 ^ x129;
  assign n885 = n884 ^ n851;
  assign n880 = ~n836 & ~n861;
  assign n886 = n885 ^ n880;
  assign n887 = ~n834 & ~n886;
  assign n888 = n887 ^ n880;
  assign n889 = n833 & n888;
  assign n890 = ~n879 & ~n889;
  assign n892 = n833 & n846;
  assign n893 = n892 ^ n863;
  assign n894 = n891 & n893;
  assign n895 = n894 ^ n863;
  assign n912 = n863 ^ n846;
  assign n913 = n912 ^ n845;
  assign n911 = n877 ^ n865;
  assign n914 = n913 ^ n911;
  assign n915 = n914 ^ n859;
  assign n916 = ~n833 & n915;
  assign n901 = n885 ^ n865;
  assign n905 = n904 ^ n901;
  assign n907 = n906 ^ n905;
  assign n899 = n884 ^ n850;
  assign n900 = n899 ^ n881;
  assign n908 = n907 ^ n900;
  assign n909 = ~n833 & ~n908;
  assign n910 = n909 ^ n900;
  assign n917 = n916 ^ n910;
  assign n918 = n891 & ~n917;
  assign n919 = n918 ^ n910;
  assign n922 = ~n849 & n921;
  assign n920 = ~n857 & n873;
  assign n923 = n922 ^ n920;
  assign n924 = n919 & ~n923;
  assign n925 = ~n898 & n924;
  assign n926 = ~n895 & n925;
  assign n927 = n890 & n926;
  assign n928 = ~n855 & n927;
  assign n929 = n928 ^ x35;
  assign n930 = n929 ^ x128;
  assign n931 = x94 ^ x36;
  assign n932 = x99 ^ x62;
  assign n933 = n931 & ~n932;
  assign n934 = n933 ^ n932;
  assign n935 = n934 ^ n931;
  assign n940 = x98 ^ x4;
  assign n941 = x97 ^ x12;
  assign n942 = n940 & n941;
  assign n943 = n942 ^ n940;
  assign n936 = x95 ^ x28;
  assign n937 = x96 ^ x20;
  assign n938 = ~n936 & n937;
  assign n939 = n938 ^ n937;
  assign n952 = n939 ^ n936;
  assign n953 = n952 ^ n937;
  assign n954 = n943 & ~n953;
  assign n944 = n943 ^ n941;
  assign n951 = n938 & ~n944;
  assign n955 = n954 ^ n951;
  assign n947 = n936 & n943;
  assign n948 = ~n937 & n947;
  assign n949 = n948 ^ n947;
  assign n945 = n944 ^ n940;
  assign n946 = n939 & n945;
  assign n950 = n949 ^ n946;
  assign n956 = n955 ^ n950;
  assign n957 = n935 & n956;
  assign n959 = n947 ^ n943;
  assign n960 = n959 ^ n954;
  assign n958 = ~n944 & ~n953;
  assign n961 = n960 ^ n958;
  assign n962 = n932 & n961;
  assign n963 = n962 ^ n960;
  assign n964 = ~n931 & n963;
  assign n966 = n940 ^ n937;
  assign n967 = n966 ^ n936;
  assign n968 = n967 ^ n941;
  assign n969 = ~n936 & n968;
  assign n970 = ~n940 & n969;
  assign n971 = n970 ^ n951;
  assign n965 = n935 ^ n932;
  assign n972 = n971 ^ n965;
  assign n975 = n951 ^ n938;
  assign n973 = n938 & n945;
  assign n974 = n973 ^ n960;
  assign n976 = n975 ^ n974;
  assign n977 = n976 ^ n934;
  assign n978 = n965 & n977;
  assign n979 = n978 ^ n934;
  assign n980 = n972 & n979;
  assign n981 = n980 ^ n971;
  assign n985 = n954 ^ n953;
  assign n984 = n971 ^ n958;
  assign n986 = n985 ^ n984;
  assign n987 = ~n931 & ~n986;
  assign n982 = n965 ^ n934;
  assign n983 = n973 & ~n982;
  assign n988 = n987 ^ n983;
  assign n1013 = n970 ^ n967;
  assign n1014 = n1013 ^ n953;
  assign n989 = n939 & n942;
  assign n993 = n989 ^ n939;
  assign n994 = n993 ^ n950;
  assign n995 = n994 ^ n948;
  assign n1010 = n995 ^ n946;
  assign n1001 = n976 ^ n971;
  assign n1008 = n1001 ^ n986;
  assign n1009 = n1008 ^ n951;
  assign n1011 = n1010 ^ n1009;
  assign n1012 = n1011 ^ n959;
  assign n1015 = n1014 ^ n1012;
  assign n1007 = ~n944 & n952;
  assign n1016 = n1015 ^ n1007;
  assign n1006 = n952 ^ n948;
  assign n1017 = n1016 ^ n1006;
  assign n1018 = n1017 ^ n949;
  assign n1019 = n1018 ^ n994;
  assign n1020 = n934 & n1016;
  assign n1021 = n1019 & ~n1020;
  assign n990 = ~n933 & ~n989;
  assign n1005 = ~n946 & ~n990;
  assign n1022 = n1021 ^ n1005;
  assign n1002 = n1001 ^ n935;
  assign n1003 = ~n990 & n1002;
  assign n1004 = n1003 ^ n932;
  assign n1023 = n1022 ^ n1004;
  assign n998 = n955 & ~n990;
  assign n991 = n990 ^ n931;
  assign n992 = n990 ^ n954;
  assign n996 = n995 ^ n992;
  assign n997 = ~n991 & ~n996;
  assign n999 = n998 ^ n997;
  assign n1000 = n999 ^ n989;
  assign n1024 = n1023 ^ n1000;
  assign n1025 = ~n988 & n1024;
  assign n1026 = ~n981 & n1025;
  assign n1027 = ~n964 & n1026;
  assign n1028 = ~n957 & n1027;
  assign n1029 = n1028 ^ x43;
  assign n1030 = n1029 ^ x127;
  assign n1031 = ~n930 & n1030;
  assign n1071 = n1070 ^ n1050;
  assign n1072 = n1068 & ~n1071;
  assign n1073 = n1072 ^ n1050;
  assign n1074 = n1067 & ~n1073;
  assign n1092 = n1083 ^ n1043;
  assign n1094 = n1093 ^ n1092;
  assign n1095 = n1088 & n1094;
  assign n1098 = n1097 ^ n1075;
  assign n1099 = ~n1096 & n1098;
  assign n1100 = n1081 & ~n1096;
  assign n1111 = n1110 ^ n1055;
  assign n1112 = n1068 & ~n1111;
  assign n1104 = n1075 ^ n1055;
  assign n1102 = n1071 ^ n1065;
  assign n1103 = n1102 ^ n1051;
  assign n1105 = n1104 ^ n1103;
  assign n1107 = n1106 ^ n1105;
  assign n1108 = n1068 & ~n1107;
  assign n1109 = n1108 ^ n1106;
  assign n1113 = n1112 ^ n1109;
  assign n1114 = n1067 & ~n1113;
  assign n1115 = n1114 ^ n1109;
  assign n1116 = ~n1101 & n1115;
  assign n1117 = ~n1100 & n1116;
  assign n1118 = ~n1099 & n1117;
  assign n1119 = ~n1095 & n1118;
  assign n1120 = ~n1091 & n1119;
  assign n1121 = ~n1090 & n1120;
  assign n1122 = ~n1074 & n1121;
  assign n1123 = n1066 & n1122;
  assign n1124 = n1123 ^ x59;
  assign n1125 = n1124 ^ x125;
  assign n1128 = n1127 ^ n1126;
  assign n1131 = n1129 & ~n1130;
  assign n1135 = n1134 ^ n1131;
  assign n1174 = n1160 ^ n1131;
  assign n1175 = n1174 ^ n1142;
  assign n1172 = n1171 ^ n1164;
  assign n1173 = n1172 ^ n1165;
  assign n1176 = n1175 ^ n1173;
  assign n1177 = ~n1135 & n1176;
  assign n1178 = n1177 ^ n1173;
  assign n1179 = n1178 ^ n1144;
  assign n1180 = n1179 ^ n1177;
  assign n1181 = ~n1126 & n1180;
  assign n1182 = n1181 ^ n1179;
  assign n1183 = n1128 & n1182;
  assign n1185 = n1174 ^ n1130;
  assign n1191 = n1132 & n1185;
  assign n1190 = n1152 ^ n1130;
  assign n1192 = n1191 ^ n1190;
  assign n1193 = ~n1127 & ~n1192;
  assign n1184 = n1163 ^ n1152;
  assign n1186 = n1185 ^ n1184;
  assign n1187 = n1186 ^ n1130;
  assign n1188 = n1127 & ~n1187;
  assign n1189 = n1188 ^ n1156;
  assign n1194 = n1193 ^ n1189;
  assign n1195 = ~n1126 & n1194;
  assign n1196 = n1195 ^ n1189;
  assign n1197 = ~n1183 & ~n1196;
  assign n1198 = n1197 ^ x51;
  assign n1199 = n1198 ^ x126;
  assign n1200 = ~n1125 & n1199;
  assign n1432 = n1031 & n1200;
  assign n3007 = n1404 & n1432;
  assign n1201 = n1200 ^ n1199;
  assign n1202 = n1201 ^ n1125;
  assign n1032 = n1031 ^ n1030;
  assign n1410 = n1032 ^ n930;
  assign n1419 = n1410 ^ n1030;
  assign n1445 = n1202 & ~n1419;
  assign n1446 = n1445 ^ n1419;
  assign n1205 = n1199 ^ n1032;
  assign n1206 = ~n1125 & n1205;
  assign n1442 = n1432 ^ n1206;
  assign n1416 = n1202 ^ n1199;
  assign n1414 = n1200 & n1410;
  assign n1422 = n1416 ^ n1414;
  assign n1420 = ~n1416 & ~n1419;
  assign n1417 = n1410 & ~n1416;
  assign n1412 = n1031 & ~n1199;
  assign n1413 = ~n1125 & n1412;
  assign n1415 = n1414 ^ n1413;
  assign n1418 = n1417 ^ n1415;
  assign n1421 = n1420 ^ n1418;
  assign n1423 = n1422 ^ n1421;
  assign n1441 = n1423 ^ n1414;
  assign n1443 = n1442 ^ n1441;
  assign n1444 = n1443 ^ n1420;
  assign n1447 = n1446 ^ n1444;
  assign n1411 = n1202 & n1410;
  assign n3003 = n1447 ^ n1411;
  assign n3004 = n3003 ^ n1417;
  assign n3005 = n1404 & n3004;
  assign n3006 = n3005 ^ n1417;
  assign n3008 = n3007 ^ n3006;
  assign n3009 = ~n1304 & n3008;
  assign n3010 = n3009 ^ n3006;
  assign n1409 = n1404 ^ n1304;
  assign n1203 = n1032 & n1202;
  assign n1428 = n1203 & ~n1304;
  assign n1207 = n1206 ^ n1200;
  assign n1424 = n1423 ^ n1207;
  assign n1425 = n1424 ^ n1411;
  assign n1426 = ~n1304 & ~n1425;
  assign n1427 = n1426 ^ n1424;
  assign n1429 = n1428 ^ n1427;
  assign n1430 = n1409 & ~n1429;
  assign n1431 = n1430 ^ n1427;
  assign n1449 = n1413 ^ n1412;
  assign n1204 = n1203 ^ n1032;
  assign n1208 = n1207 ^ n1204;
  assign n3014 = n1449 ^ n1208;
  assign n1435 = n1201 & n1410;
  assign n3015 = n3014 ^ n1435;
  assign n3016 = ~n1404 & n3015;
  assign n3017 = n3016 ^ n1435;
  assign n3018 = ~n1304 & n3017;
  assign n1436 = n1435 ^ n1203;
  assign n1437 = n1436 ^ n1424;
  assign n1438 = n1304 & ~n1437;
  assign n1439 = n1438 ^ n1424;
  assign n1440 = ~n1404 & ~n1439;
  assign n1405 = ~n1304 & n1404;
  assign n1406 = n1405 ^ n1304;
  assign n1455 = n1405 ^ n1404;
  assign n3611 = n1445 & ~n1455;
  assign n3610 = n1447 ^ n1417;
  assign n3612 = n3611 ^ n3610;
  assign n3613 = n1406 & n3612;
  assign n3614 = n3613 ^ n3610;
  assign n1456 = n1412 ^ n1032;
  assign n3616 = ~n1405 & ~n1456;
  assign n1407 = n1406 ^ n1404;
  assign n3617 = n1207 & n1407;
  assign n3618 = n3617 ^ n1418;
  assign n3619 = ~n3616 & n3618;
  assign n3615 = n1423 ^ n1413;
  assign n3620 = n3619 ^ n3615;
  assign n3621 = n3620 ^ n3615;
  assign n3622 = n1406 & n3621;
  assign n3623 = n3622 ^ n3615;
  assign n3624 = ~n1455 & ~n3623;
  assign n3625 = n3624 ^ n3615;
  assign n3626 = ~n3614 & n3625;
  assign n1457 = n1456 ^ n1030;
  assign n1458 = n1457 ^ n1432;
  assign n3628 = n1406 & n1458;
  assign n3627 = ~n1409 & ~n1444;
  assign n3629 = n3628 ^ n3627;
  assign n3630 = n3626 & ~n3629;
  assign n3631 = ~n1440 & n3630;
  assign n3632 = ~n3018 & n3631;
  assign n3633 = n1431 & n3632;
  assign n3634 = ~n3010 & n3633;
  assign n3635 = n3634 ^ x4;
  assign n3762 = n3635 ^ x196;
  assign n2388 = n1192 ^ n1187;
  assign n2389 = n1126 & ~n2388;
  assign n2390 = n2389 ^ n1187;
  assign n2385 = n1177 ^ n1126;
  assign n2386 = n2385 ^ n1182;
  assign n2387 = n2386 ^ n1179;
  assign n2391 = n2390 ^ n2387;
  assign n2392 = ~n1128 & ~n2391;
  assign n2393 = n2392 ^ n2390;
  assign n2394 = ~n1156 & n2393;
  assign n2395 = n2394 ^ x57;
  assign n2598 = n2395 ^ x159;
  assign n2599 = n1343 & ~n1387;
  assign n2325 = ~n1316 & n1339;
  assign n2326 = n2325 ^ n1328;
  assign n2327 = n1315 & n2326;
  assign n2600 = n2599 ^ n2327;
  assign n2609 = ~n1316 & n1385;
  assign n2604 = n1350 ^ n1337;
  assign n2603 = n1391 ^ n1341;
  assign n2605 = n2604 ^ n2603;
  assign n2601 = n1383 ^ n1371;
  assign n2602 = n2601 ^ n1342;
  assign n2606 = n2605 ^ n2602;
  assign n2607 = n1316 & n2606;
  assign n2608 = n2607 ^ n2602;
  assign n2610 = n2609 ^ n2608;
  assign n2611 = ~n1369 & ~n2610;
  assign n2612 = n2611 ^ n2608;
  assign n2614 = ~n1345 & ~n1369;
  assign n2331 = n1372 ^ n1358;
  assign n2332 = n2331 ^ n1331;
  assign n2613 = n1318 & n2332;
  assign n2615 = n2614 ^ n2613;
  assign n2616 = n2612 & ~n2615;
  assign n2617 = ~n1376 & n2616;
  assign n2618 = ~n1368 & n2617;
  assign n2619 = ~n2600 & n2618;
  assign n2620 = ~n1353 & n2619;
  assign n2621 = ~n1319 & n2620;
  assign n2622 = n2621 ^ x39;
  assign n2623 = n2622 ^ x154;
  assign n2624 = ~n2598 & ~n2623;
  assign n2490 = ~n931 & n973;
  assign n2491 = n2490 ^ n955;
  assign n2492 = n982 & n2491;
  assign n2493 = n2492 ^ n955;
  assign n1490 = n995 ^ n986;
  assign n1491 = n1490 ^ n989;
  assign n2494 = n1491 ^ n950;
  assign n2495 = n935 & ~n2494;
  assign n2501 = n965 & ~n1007;
  assign n1493 = n1017 ^ n950;
  assign n1495 = n965 & ~n1493;
  assign n2502 = n2501 ^ n1495;
  assign n2503 = n2502 ^ n931;
  assign n1487 = n1017 ^ n976;
  assign n1488 = n1487 ^ n1007;
  assign n2497 = n1488 ^ n932;
  assign n2498 = n1488 ^ n990;
  assign n2499 = ~n2497 & n2498;
  assign n2496 = ~n990 & n1013;
  assign n2500 = n2499 ^ n2496;
  assign n2504 = n2503 ^ n2500;
  assign n2505 = ~n2495 & ~n2504;
  assign n2506 = ~n2493 & n2505;
  assign n2507 = ~n981 & n2506;
  assign n2508 = ~n964 & n2507;
  assign n2509 = n2508 ^ x31;
  assign n2510 = n2509 ^ x155;
  assign n1714 = n877 ^ n873;
  assign n1715 = ~n897 & n1714;
  assign n1712 = n850 & ~n897;
  assign n1711 = n837 & n921;
  assign n1713 = n1712 ^ n1711;
  assign n2305 = n905 ^ n875;
  assign n2306 = ~n896 & ~n2305;
  assign n2307 = n915 ^ n850;
  assign n2308 = ~n833 & n2307;
  assign n2309 = n2308 ^ n850;
  assign n2310 = n2309 ^ n847;
  assign n2311 = ~n834 & n2310;
  assign n2312 = n2311 ^ n847;
  assign n2313 = ~n2306 & ~n2312;
  assign n2314 = ~n1713 & n2313;
  assign n2315 = ~n1715 & n2314;
  assign n2316 = ~n2133 & n2315;
  assign n2317 = n890 & n2316;
  assign n2318 = ~n1710 & n2317;
  assign n2319 = n2318 ^ x7;
  assign n2511 = n2319 ^ x158;
  assign n2512 = n2510 & ~n2511;
  assign n1690 = n1679 & n1689;
  assign n2513 = n1664 ^ n1658;
  assign n2514 = ~n1617 & ~n2513;
  assign n2515 = n2514 ^ n1664;
  assign n2516 = n1679 & ~n2515;
  assign n2520 = n1674 ^ n1658;
  assign n2521 = n2520 ^ n1638;
  assign n2519 = n1649 ^ n1641;
  assign n2522 = n2521 ^ n2519;
  assign n2523 = ~n1618 & ~n2522;
  assign n2524 = n2523 ^ n2519;
  assign n2517 = n1668 ^ n1652;
  assign n2518 = ~n1618 & ~n2517;
  assign n2525 = n2524 ^ n2518;
  assign n2526 = ~n1617 & n2525;
  assign n2527 = n2526 ^ n2524;
  assign n2528 = ~n2516 & ~n2527;
  assign n2529 = ~n1690 & n2528;
  assign n2530 = ~n2173 & n2529;
  assign n2531 = ~n2175 & n2530;
  assign n2532 = ~n1640 & n2531;
  assign n2533 = n2532 ^ x23;
  assign n2534 = n2533 ^ x156;
  assign n2535 = n1991 ^ n1077;
  assign n2536 = n2535 ^ n1050;
  assign n2537 = n2536 ^ n1050;
  assign n2538 = n1067 & ~n2537;
  assign n2539 = n2538 ^ n1050;
  assign n2540 = ~n1068 & ~n2539;
  assign n2541 = n2540 ^ n1050;
  assign n2542 = n1058 & n1068;
  assign n2543 = n2542 ^ n1047;
  assign n2544 = ~n1087 & n2543;
  assign n2545 = n2541 & ~n2544;
  assign n2546 = ~n1060 & ~n1087;
  assign n2561 = n1106 ^ n1079;
  assign n2562 = n1086 & ~n2561;
  assign n2559 = n1043 & n1088;
  assign n2560 = n2559 ^ n1086;
  assign n2563 = n2562 ^ n2560;
  assign n2557 = ~n1060 & ~n1086;
  assign n2558 = n2557 ^ n2546;
  assign n2564 = n2563 ^ n2558;
  assign n2555 = n2103 ^ n1074;
  assign n2551 = n1068 & n1081;
  assign n2552 = n2551 ^ n1091;
  assign n2553 = n2552 ^ n1100;
  assign n2548 = n1068 ^ n1064;
  assign n2549 = ~n1087 & n2548;
  assign n2547 = n1089 & n1995;
  assign n2550 = n2549 ^ n2547;
  assign n2554 = n2553 ^ n2550;
  assign n2556 = n2555 ^ n2554;
  assign n2565 = n2564 ^ n2556;
  assign n2566 = ~n2546 & ~n2565;
  assign n2567 = n2545 & n2566;
  assign n2568 = ~n1101 & n2567;
  assign n2569 = n2568 ^ x15;
  assign n2570 = n2569 ^ x157;
  assign n2571 = n2534 & ~n2570;
  assign n2629 = n2512 & n2571;
  assign n2575 = n2571 ^ n2534;
  assign n2628 = n2512 & n2575;
  assign n2630 = n2629 ^ n2628;
  assign n2631 = n2630 ^ n2512;
  assign n2572 = n2571 ^ n2570;
  assign n2573 = n2572 ^ n2534;
  assign n2574 = n2512 & n2573;
  assign n2632 = n2631 ^ n2574;
  assign n2849 = n2624 & n2632;
  assign n2576 = n2512 ^ n2511;
  assign n2580 = n2576 ^ n2510;
  assign n2581 = n2575 & n2580;
  assign n2589 = n2581 ^ n2580;
  assign n2585 = ~n2510 & ~n2572;
  assign n2586 = ~n2511 & n2585;
  assign n2587 = n2586 ^ n2585;
  assign n2583 = n2571 & n2580;
  assign n2588 = n2587 ^ n2583;
  assign n2590 = n2589 ^ n2588;
  assign n2577 = n2575 & ~n2576;
  assign n2591 = n2590 ^ n2577;
  assign n2592 = n2591 ^ n2585;
  assign n2593 = n2592 ^ n2510;
  assign n2579 = n2571 & ~n2576;
  assign n2582 = n2581 ^ n2579;
  assign n2584 = n2583 ^ n2582;
  assign n2594 = n2593 ^ n2584;
  assign n2850 = ~n2594 & ~n2623;
  assign n2633 = n2580 ^ n2511;
  assign n2634 = ~n2570 & n2633;
  assign n2635 = n2634 ^ n2633;
  assign n2595 = n2594 ^ n2591;
  assign n2596 = n2595 ^ n2573;
  assign n2578 = n2577 ^ n2574;
  assign n2597 = n2596 ^ n2578;
  assign n2636 = n2635 ^ n2597;
  assign n2851 = n2850 ^ n2636;
  assign n2852 = n2598 & ~n2851;
  assign n2853 = n2852 ^ n2636;
  assign n2854 = ~n2849 & n2853;
  assign n2650 = n2578 & n2598;
  assign n2651 = n2650 ^ n2574;
  assign n2652 = ~n2623 & n2651;
  assign n2627 = n2594 ^ n2581;
  assign n2625 = n2624 ^ n2598;
  assign n2662 = n2625 ^ n2623;
  assign n3765 = ~n2627 & ~n2662;
  assign n2653 = n2623 ^ n2598;
  assign n2642 = n2585 ^ n2572;
  assign n2643 = n2642 ^ n2632;
  assign n2654 = n2643 ^ n2634;
  assign n2656 = n2654 ^ n2628;
  assign n2655 = n2654 ^ n2632;
  assign n2657 = n2656 ^ n2655;
  assign n2658 = ~n2623 & n2657;
  assign n2659 = n2658 ^ n2655;
  assign n2660 = n2653 & ~n2659;
  assign n3766 = n2655 ^ n2628;
  assign n3767 = ~n2662 & ~n3766;
  assign n3769 = n2591 ^ n2588;
  assign n3768 = n2590 ^ n2579;
  assign n3770 = n3769 ^ n3768;
  assign n3771 = n3770 ^ n3768;
  assign n3772 = n2623 & n3771;
  assign n3773 = n3772 ^ n3768;
  assign n3774 = n2653 & n3773;
  assign n3775 = n3774 ^ n3768;
  assign n3776 = ~n3767 & ~n3775;
  assign n3783 = n2597 ^ n2583;
  assign n3784 = n3783 ^ n2586;
  assign n3777 = n2570 ^ n2534;
  assign n3778 = n3777 ^ n2511;
  assign n3779 = n2570 ^ n2511;
  assign n3780 = ~n2510 & ~n3779;
  assign n3781 = n3780 ^ n2570;
  assign n3782 = n3778 & ~n3781;
  assign n3785 = n3784 ^ n3782;
  assign n3786 = ~n2598 & ~n3785;
  assign n3787 = n3786 ^ n3782;
  assign n2644 = n2643 ^ n2574;
  assign n2645 = ~n2598 & ~n2644;
  assign n2646 = n2645 ^ n2643;
  assign n3788 = n3787 ^ n2646;
  assign n3789 = ~n2623 & ~n3788;
  assign n3790 = n3789 ^ n2646;
  assign n3791 = n3776 & n3790;
  assign n3792 = ~n2660 & n3791;
  assign n3793 = ~n3765 & n3792;
  assign n3794 = ~n2652 & n3793;
  assign n3795 = n2854 & n3794;
  assign n3796 = n3795 ^ x46;
  assign n3797 = n3796 ^ x199;
  assign n3046 = n2100 ^ x141;
  assign n1680 = ~n1617 & ~n1650;
  assign n1681 = n1680 ^ n1649;
  assign n1682 = n1679 & n1681;
  assign n1834 = ~n1621 & ~n1669;
  assign n1835 = ~n1618 & ~n1674;
  assign n1836 = n1662 ^ n1622;
  assign n1837 = n1627 ^ n1623;
  assign n1838 = n1837 ^ n1628;
  assign n1839 = n1643 ^ n1627;
  assign n1840 = ~n1838 & n1839;
  assign n1841 = n1840 ^ n1620;
  assign n1842 = n1662 & n1841;
  assign n1843 = n1842 ^ n1620;
  assign n1844 = n1836 & ~n1843;
  assign n1845 = n1844 ^ n1622;
  assign n1848 = n1665 ^ n1637;
  assign n1849 = n1637 ^ n1617;
  assign n1850 = n1679 & n1849;
  assign n1851 = n1850 ^ n1617;
  assign n1852 = n1848 & ~n1851;
  assign n1853 = n1852 ^ n1665;
  assign n1854 = n1664 & ~n1853;
  assign n1855 = ~n1638 & n1854;
  assign n1693 = n1666 ^ n1640;
  assign n1694 = n1693 ^ n1631;
  assign n1846 = n1694 ^ n1645;
  assign n1847 = n1617 & ~n1846;
  assign n1856 = n1855 ^ n1847;
  assign n1857 = n1679 & ~n1856;
  assign n1858 = n1857 ^ n1855;
  assign n1859 = n1845 & n1858;
  assign n1860 = ~n1835 & n1859;
  assign n1861 = ~n1834 & n1860;
  assign n1863 = n1619 & ~n1668;
  assign n1862 = ~n1654 & ~n1679;
  assign n1864 = n1863 ^ n1862;
  assign n1865 = n1861 & ~n1864;
  assign n1866 = ~n1833 & n1865;
  assign n1867 = ~n1682 & n1866;
  assign n1868 = n1867 ^ x3;
  assign n3129 = n1868 ^ x136;
  assign n3141 = ~n3046 & ~n3129;
  assign n3142 = n3141 ^ n3129;
  assign n1970 = n1082 & n1088;
  assign n1976 = n1110 ^ n1040;
  assign n1978 = n1977 ^ n1976;
  assign n1979 = n1068 & ~n1978;
  assign n1980 = n1979 ^ n1977;
  assign n1972 = n1060 ^ n1048;
  assign n1973 = n1096 & n1972;
  assign n1974 = ~n1111 & ~n1973;
  assign n1975 = ~n1971 & ~n1974;
  assign n1981 = n1980 ^ n1975;
  assign n1982 = n1087 & n1981;
  assign n1983 = n1982 ^ n1975;
  assign n1984 = ~n1970 & n1983;
  assign n1987 = ~n1068 & ~n1986;
  assign n1988 = n1987 ^ n1075;
  assign n1989 = ~n1087 & n1988;
  assign n1990 = n1984 & ~n1989;
  assign n1993 = n1068 & n1992;
  assign n1996 = n1995 ^ n1993;
  assign n1997 = n1087 & ~n1996;
  assign n1998 = n1997 ^ n1995;
  assign n1999 = n1990 & n1998;
  assign n2000 = ~n1090 & n1999;
  assign n2001 = ~n1100 & n2000;
  assign n2002 = ~n1074 & n2001;
  assign n2003 = n2002 ^ x61;
  assign n3047 = n2003 ^ x137;
  assign n3070 = n2068 ^ x140;
  assign n3048 = ~n934 & ~n986;
  assign n3049 = n965 & n974;
  assign n3051 = n958 ^ n950;
  assign n3050 = n1008 ^ n994;
  assign n3052 = n3051 ^ n3050;
  assign n3053 = n982 & n3052;
  assign n3054 = ~n1007 & n3053;
  assign n1494 = n1493 ^ n965;
  assign n1496 = n1495 ^ n1494;
  assign n3055 = n1017 & n1020;
  assign n3056 = ~n1496 & ~n3055;
  assign n3057 = n990 & ~n3056;
  assign n3058 = ~n3054 & ~n3057;
  assign n3059 = ~n3049 & ~n3058;
  assign n3060 = ~n3048 & n3059;
  assign n3062 = ~n931 & n947;
  assign n3061 = n935 & ~n1487;
  assign n3063 = n3062 ^ n3061;
  assign n3064 = n3060 & ~n3063;
  assign n3065 = ~n957 & n3064;
  assign n3066 = ~n2493 & n3065;
  assign n3067 = n3066 ^ x45;
  assign n3068 = n3067 ^ x139;
  assign n3119 = n3070 ^ n3068;
  assign n2321 = n1391 ^ n1338;
  assign n2322 = ~n1315 & n2321;
  assign n2323 = n2322 ^ n1338;
  assign n2324 = ~n1369 & n2323;
  assign n3073 = n1351 ^ n1307;
  assign n3074 = n3073 ^ n1334;
  assign n3075 = n1315 & n3074;
  assign n3076 = n3075 ^ n3073;
  assign n3071 = ~n1316 & n1378;
  assign n3072 = n3071 ^ n1377;
  assign n3077 = n3076 ^ n3072;
  assign n3078 = ~n1369 & n3077;
  assign n3079 = n3078 ^ n3076;
  assign n3081 = n1358 & ~n1369;
  assign n3080 = n1315 & n1350;
  assign n3082 = n3081 ^ n3080;
  assign n3083 = ~n3079 & ~n3082;
  assign n3084 = ~n2324 & n3083;
  assign n3085 = ~n2600 & n3084;
  assign n3086 = ~n1363 & n3085;
  assign n3087 = ~n1319 & n3086;
  assign n3088 = n3087 ^ x53;
  assign n3089 = n3088 ^ x138;
  assign n3120 = n3119 ^ n3089;
  assign n3121 = ~n3047 & n3120;
  assign n3122 = n3121 ^ n3047;
  assign n3069 = ~n3047 & ~n3068;
  assign n3093 = n3069 ^ n3047;
  assign n3090 = ~n3070 & ~n3089;
  assign n3091 = n3090 ^ n3070;
  assign n3102 = n3091 ^ n3089;
  assign n3108 = n3102 ^ n3070;
  assign n3116 = ~n3093 & ~n3108;
  assign n3094 = ~n3091 & ~n3093;
  assign n3117 = n3116 ^ n3094;
  assign n3103 = n3069 & ~n3102;
  assign n3118 = n3117 ^ n3103;
  assign n3123 = n3122 ^ n3118;
  assign n3124 = n3123 ^ n3090;
  assign n3114 = n3090 & ~n3093;
  assign n3096 = n3093 ^ n3068;
  assign n3111 = ~n3096 & ~n3102;
  assign n3112 = n3111 ^ n3096;
  assign n3109 = ~n3096 & ~n3108;
  assign n3097 = ~n3091 & ~n3096;
  assign n3110 = n3109 ^ n3097;
  assign n3113 = n3112 ^ n3110;
  assign n3115 = n3114 ^ n3113;
  assign n3125 = n3124 ^ n3115;
  assign n3105 = ~n3068 & n3089;
  assign n3098 = n3097 ^ n3091;
  assign n3106 = n3105 ^ n3098;
  assign n3104 = n3103 ^ n3094;
  assign n3107 = n3106 ^ n3104;
  assign n3126 = n3125 ^ n3107;
  assign n3147 = n3126 ^ n3108;
  assign n3146 = n3123 ^ n3110;
  assign n3148 = n3147 ^ n3146;
  assign n3100 = n3069 ^ n3068;
  assign n3092 = n3069 & ~n3091;
  assign n3095 = n3094 ^ n3092;
  assign n3099 = n3098 ^ n3095;
  assign n3101 = n3100 ^ n3099;
  assign n3143 = n3101 ^ n3097;
  assign n3144 = n3143 ^ n3123;
  assign n3145 = n3144 ^ n3116;
  assign n3149 = n3148 ^ n3145;
  assign n3150 = n3149 ^ n3114;
  assign n3151 = ~n3142 & n3150;
  assign n3137 = n3103 & n3129;
  assign n3133 = n3111 ^ n3099;
  assign n3134 = n3133 ^ n3113;
  assign n3135 = n3129 & n3134;
  assign n3136 = n3135 ^ n3113;
  assign n3138 = n3137 ^ n3136;
  assign n3139 = n3046 & ~n3138;
  assign n3140 = n3139 ^ n3136;
  assign n3152 = n3151 ^ n3140;
  assign n3153 = n3141 ^ n3092;
  assign n3154 = n3142 ^ n3094;
  assign n3155 = ~n3092 & n3154;
  assign n3156 = n3155 ^ n3142;
  assign n3157 = n3153 & ~n3156;
  assign n3158 = n3157 ^ n3141;
  assign n3165 = n3114 ^ n3093;
  assign n3166 = n3165 ^ n3117;
  assign n3167 = n3166 ^ n3123;
  assign n3326 = n3167 ^ n3113;
  assign n3516 = n3046 & ~n3326;
  assign n3517 = n3516 ^ n3113;
  assign n3518 = n3129 & ~n3517;
  assign n3322 = n3141 ^ n3046;
  assign n3519 = n3150 ^ n3146;
  assign n3520 = ~n3322 & ~n3519;
  assign n3521 = n3126 & n3141;
  assign n3522 = n3521 ^ n3096;
  assign n3523 = ~n3147 & ~n3522;
  assign n3524 = n3523 ^ n3096;
  assign n3525 = n3521 & ~n3524;
  assign n3526 = n3525 ^ n3141;
  assign n3527 = ~n3520 & ~n3526;
  assign n3529 = n3110 ^ n3107;
  assign n3530 = n3529 ^ n3113;
  assign n3531 = n3530 ^ n3092;
  assign n3528 = n3166 ^ n3143;
  assign n3532 = n3531 ^ n3528;
  assign n3533 = n3129 & ~n3532;
  assign n3534 = n3533 ^ n3528;
  assign n3535 = n3046 & ~n3534;
  assign n3536 = n3527 & ~n3535;
  assign n3537 = ~n3518 & n3536;
  assign n3538 = ~n3158 & n3537;
  assign n3539 = n3152 & n3538;
  assign n3540 = n3539 ^ x62;
  assign n3799 = n3540 ^ x197;
  assign n3834 = n3797 & n3799;
  assign n3838 = n3834 ^ n3799;
  assign n3839 = n3838 ^ n3797;
  assign n3840 = n3839 ^ n3799;
  assign n2004 = n2003 ^ x135;
  assign n1582 = ~n1522 & n1547;
  assign n1584 = n1583 ^ n1582;
  assign n1906 = n1575 ^ n1546;
  assign n1907 = n1520 & n1906;
  assign n1553 = n1520 ^ n1518;
  assign n1908 = n1571 ^ n1543;
  assign n1909 = n1908 ^ n1579;
  assign n1910 = ~n1553 & n1909;
  assign n1552 = ~n1522 & n1551;
  assign n1911 = ~n1521 & n1906;
  assign n1915 = n1520 & n1533;
  assign n1597 = n1564 ^ n1551;
  assign n1912 = n1597 ^ n1558;
  assign n1913 = ~n1553 & n1912;
  assign n1914 = n1913 ^ n1549;
  assign n1916 = n1915 ^ n1914;
  assign n1917 = ~n1518 & n1916;
  assign n1918 = n1562 ^ n1535;
  assign n1919 = n1517 & n1918;
  assign n1920 = n1919 ^ n1562;
  assign n1921 = ~n1566 & ~n1920;
  assign n1922 = ~n1519 & n1921;
  assign n1923 = n1922 ^ n1519;
  assign n1924 = ~n1917 & n1923;
  assign n1925 = ~n1911 & n1924;
  assign n1926 = ~n1552 & n1925;
  assign n1927 = ~n1910 & n1926;
  assign n1928 = ~n1907 & n1927;
  assign n1929 = n1588 ^ n1563;
  assign n1930 = ~n1517 & ~n1929;
  assign n1931 = n1930 ^ n1588;
  assign n1932 = n1518 & ~n1931;
  assign n1933 = n1928 & ~n1932;
  assign n1934 = ~n1584 & n1933;
  assign n1935 = ~n1905 & n1934;
  assign n1936 = n1935 ^ x11;
  assign n1937 = n1936 ^ x133;
  assign n1884 = n1237 ^ n1225;
  assign n1885 = n1884 ^ n1249;
  assign n1883 = n1882 ^ n1229;
  assign n1886 = n1885 ^ n1883;
  assign n1887 = n1210 & n1886;
  assign n1888 = n1887 ^ n1885;
  assign n1878 = n1287 ^ n1243;
  assign n1876 = n1264 ^ n1236;
  assign n1877 = n1876 ^ n1222;
  assign n1879 = n1878 ^ n1877;
  assign n1880 = n1210 & n1879;
  assign n1881 = n1880 ^ n1877;
  assign n1889 = n1888 ^ n1881;
  assign n1890 = n1209 & n1889;
  assign n1891 = n1890 ^ n1881;
  assign n1894 = n1209 & n1242;
  assign n1893 = n1245 & ~n1892;
  assign n1895 = n1894 ^ n1893;
  assign n1896 = ~n1891 & ~n1895;
  assign n1897 = ~n1875 & n1896;
  assign n1898 = ~n1257 & n1897;
  assign n1899 = ~n1265 & n1898;
  assign n1900 = n1899 ^ x19;
  assign n1901 = n1900 ^ x132;
  assign n2010 = n1937 ^ n1901;
  assign n1869 = n1868 ^ x134;
  assign n2014 = n1937 ^ n1869;
  assign n2019 = ~n2010 & ~n2014;
  assign n2020 = n2019 ^ n1901;
  assign n2021 = n2020 ^ n1869;
  assign n1870 = n929 ^ x130;
  assign n2022 = n2021 ^ n1870;
  assign n2023 = ~n2020 & ~n2022;
  assign n1948 = n1869 & ~n1937;
  assign n1949 = n1948 ^ n1869;
  assign n1961 = n1901 & n1949;
  assign n1956 = n1948 ^ n1901;
  assign n1957 = n1956 ^ n1937;
  assign n2006 = n1961 ^ n1957;
  assign n1902 = n1403 ^ x131;
  assign n2017 = n1870 & ~n1902;
  assign n2018 = ~n2006 & n2017;
  assign n2024 = n2023 ^ n2018;
  assign n1903 = ~n1901 & n1902;
  assign n1946 = n1903 ^ n1902;
  assign n1947 = n1946 ^ n1901;
  assign n2015 = n1947 & n2014;
  assign n1950 = n1949 ^ n1937;
  assign n1951 = ~n1870 & n1950;
  assign n1952 = n1947 & n1951;
  assign n2012 = n1952 ^ n1947;
  assign n2011 = n1947 & n2010;
  assign n2013 = n2012 ^ n2011;
  assign n2016 = n2015 ^ n2013;
  assign n2025 = n2024 ^ n2016;
  assign n2007 = n2006 ^ n1903;
  assign n1963 = n1903 & n1948;
  assign n1960 = ~n1902 & ~n1956;
  assign n1962 = n1961 ^ n1960;
  assign n1964 = n1963 ^ n1962;
  assign n2008 = n2007 ^ n1964;
  assign n1939 = n1937 ^ n1902;
  assign n1940 = ~n1902 & ~n1939;
  assign n2009 = n2008 ^ n1940;
  assign n2026 = n2025 ^ n2009;
  assign n1943 = n1903 & n1937;
  assign n1938 = n1937 ^ n1903;
  assign n1941 = n1940 ^ n1938;
  assign n1942 = n1870 & ~n1941;
  assign n1944 = n1943 ^ n1942;
  assign n1945 = ~n1869 & n1944;
  assign n1953 = n1947 ^ n1903;
  assign n1954 = ~n1869 & n1953;
  assign n1955 = n1954 ^ n1902;
  assign n1958 = n1955 & n1957;
  assign n1959 = n1958 ^ n1937;
  assign n1965 = n1964 ^ n1959;
  assign n1966 = n1870 & ~n1965;
  assign n1967 = n1966 ^ n1959;
  assign n1968 = ~n1952 & n1967;
  assign n1969 = ~n1945 & n1968;
  assign n2027 = n2026 ^ n1969;
  assign n2028 = ~n2004 & ~n2027;
  assign n2029 = n2028 ^ n2026;
  assign n3763 = n2029 ^ x54;
  assign n3764 = n3763 ^ x198;
  assign n1483 = n1124 ^ x123;
  assign n1484 = n965 & n984;
  assign n1485 = n1019 ^ n1015;
  assign n1486 = n932 & ~n1485;
  assign n1497 = n1015 & n1496;
  assign n1489 = n1488 ^ n951;
  assign n1492 = n1491 ^ n1489;
  assign n1498 = n1497 ^ n1492;
  assign n1499 = n1498 ^ n1497;
  assign n1500 = n931 & n1499;
  assign n1501 = n1500 ^ n1497;
  assign n1502 = n982 & ~n1501;
  assign n1503 = n1502 ^ n1497;
  assign n1504 = ~n1486 & ~n1503;
  assign n1505 = ~n1484 & ~n1504;
  assign n1506 = ~n931 & ~n1011;
  assign n1507 = n1506 ^ n959;
  assign n1508 = n982 & n1507;
  assign n1509 = n1508 ^ n959;
  assign n1510 = n1505 & ~n1509;
  assign n1512 = ~n934 & n973;
  assign n1511 = ~n931 & n1007;
  assign n1513 = n1512 ^ n1511;
  assign n1514 = n1510 & ~n1513;
  assign n1515 = n1514 ^ x33;
  assign n1516 = n1515 ^ x118;
  assign n1757 = n1483 & ~n1516;
  assign n1560 = ~n1553 & n1559;
  assign n1568 = n1567 ^ n1551;
  assign n1569 = n1520 & n1568;
  assign n1570 = ~n1560 & ~n1569;
  assign n1581 = ~n1521 & n1580;
  assign n1585 = ~n1519 & n1546;
  assign n1586 = n1554 ^ n1553;
  assign n1589 = n1588 ^ n1564;
  assign n1590 = n1589 ^ n1534;
  assign n1591 = n1590 ^ n1522;
  assign n1592 = ~n1554 & ~n1591;
  assign n1593 = n1592 ^ n1522;
  assign n1594 = ~n1586 & ~n1593;
  assign n1595 = n1594 ^ n1553;
  assign n1596 = ~n1585 & n1595;
  assign n1600 = ~n1518 & n1599;
  assign n1598 = ~n1521 & n1597;
  assign n1601 = n1600 ^ n1598;
  assign n1602 = n1596 & ~n1601;
  assign n1603 = ~n1584 & n1602;
  assign n1604 = ~n1581 & n1603;
  assign n1605 = n1570 & n1604;
  assign n1606 = n1558 ^ n1522;
  assign n1608 = n1607 ^ n1520;
  assign n1609 = ~n1558 & ~n1608;
  assign n1610 = n1609 ^ n1520;
  assign n1611 = ~n1606 & n1610;
  assign n1612 = n1611 ^ n1522;
  assign n1613 = n1605 & n1612;
  assign n1614 = ~n1552 & n1613;
  assign n1615 = n1614 ^ x25;
  assign n1616 = n1615 ^ x119;
  assign n1720 = n881 & ~n896;
  assign n1722 = n903 ^ n842;
  assign n1723 = n833 & n1722;
  assign n1721 = n911 ^ n884;
  assign n1724 = n1723 ^ n1721;
  assign n1725 = ~n891 & ~n1724;
  assign n1726 = n1725 ^ n1721;
  assign n1728 = n875 ^ n849;
  assign n1729 = n1728 ^ n899;
  assign n1727 = ~n834 & n872;
  assign n1730 = n1729 ^ n1727;
  assign n1731 = ~n833 & ~n1730;
  assign n1732 = n1726 & ~n1731;
  assign n1733 = ~n1720 & n1732;
  assign n1734 = n843 & n891;
  assign n1735 = n1733 & ~n1734;
  assign n1736 = ~n1719 & n1735;
  assign n1737 = ~n895 & n1736;
  assign n1738 = ~n1715 & n1737;
  assign n1739 = ~n1713 & n1738;
  assign n1740 = ~n855 & n1739;
  assign n1741 = ~n1710 & n1740;
  assign n1742 = n1741 ^ x9;
  assign n1743 = n1742 ^ x121;
  assign n1778 = ~n1616 & n1743;
  assign n1744 = n1303 ^ x122;
  assign n1745 = n1743 & ~n1744;
  assign n1688 = ~n1618 & n1656;
  assign n1691 = n1690 ^ n1688;
  assign n1685 = ~n1617 & n1646;
  assign n1686 = n1685 ^ n1684;
  assign n1683 = ~n1620 & n1634;
  assign n1687 = n1686 ^ n1683;
  assign n1692 = n1691 ^ n1687;
  assign n1700 = ~n1622 & ~n1672;
  assign n1699 = n1619 & n1641;
  assign n1701 = n1700 ^ n1699;
  assign n1696 = n1638 & ~n1679;
  assign n1695 = ~n1621 & n1694;
  assign n1697 = n1696 ^ n1695;
  assign n1698 = n1697 ^ n1658;
  assign n1702 = n1701 ^ n1698;
  assign n1703 = ~n1692 & ~n1702;
  assign n1704 = ~n1682 & n1703;
  assign n1705 = n1678 & n1704;
  assign n1706 = n1705 ^ x17;
  assign n1707 = n1706 ^ x120;
  assign n1708 = ~n1616 & ~n1707;
  assign n1750 = n1708 ^ n1616;
  assign n1767 = n1745 & ~n1750;
  assign n1779 = n1778 ^ n1767;
  assign n1776 = n1708 & n1745;
  assign n1709 = n1708 ^ n1707;
  assign n1746 = n1745 ^ n1744;
  assign n1747 = n1746 ^ n1743;
  assign n1771 = ~n1709 & n1747;
  assign n1751 = n1750 ^ n1707;
  assign n1752 = n1747 & ~n1751;
  assign n1772 = n1771 ^ n1752;
  assign n1773 = n1772 ^ n1747;
  assign n1770 = n1708 & n1747;
  assign n1774 = n1773 ^ n1770;
  assign n1764 = n1750 ^ n1743;
  assign n1765 = ~n1744 & ~n1764;
  assign n1766 = n1765 ^ n1745;
  assign n1769 = n1766 ^ n1750;
  assign n1775 = n1774 ^ n1769;
  assign n1777 = n1776 ^ n1775;
  assign n1780 = n1779 ^ n1777;
  assign n1784 = n1780 ^ n1746;
  assign n1768 = n1767 ^ n1766;
  assign n1781 = n1780 ^ n1768;
  assign n1763 = n1708 & ~n1746;
  assign n1782 = n1781 ^ n1763;
  assign n1762 = ~n1709 & ~n1746;
  assign n1783 = n1782 ^ n1762;
  assign n1785 = n1784 ^ n1783;
  assign n1794 = n1785 ^ n1762;
  assign n1795 = n1794 ^ n1709;
  assign n1790 = n1785 ^ n1771;
  assign n1748 = n1747 ^ n1744;
  assign n1749 = ~n1709 & n1748;
  assign n1791 = n1790 ^ n1749;
  assign n1796 = n1795 ^ n1791;
  assign n1797 = n1796 ^ n1752;
  assign n3361 = n1757 & ~n1797;
  assign n1758 = n1757 ^ n1516;
  assign n1759 = n1758 ^ n1483;
  assign n1760 = n1759 ^ n1516;
  assign n1802 = n1760 & n1767;
  assign n3362 = n3361 ^ n1802;
  assign n3376 = n1770 ^ n1767;
  assign n3801 = ~n1758 & n3376;
  assign n1803 = n1760 & n1763;
  assign n3802 = n3801 ^ n1803;
  assign n3350 = n1516 & n1749;
  assign n1815 = n1745 & ~n1751;
  assign n3349 = n1759 & n1815;
  assign n3351 = n3350 ^ n3349;
  assign n3803 = n1760 & ~n1781;
  assign n1761 = n1760 ^ n1758;
  assign n1786 = ~n1516 & ~n1785;
  assign n1787 = n1786 ^ n1774;
  assign n1788 = n1761 & n1787;
  assign n1789 = n1788 ^ n1774;
  assign n3804 = n1797 ^ n1776;
  assign n3805 = ~n1758 & ~n3804;
  assign n3807 = n1815 ^ n1777;
  assign n3808 = n3807 ^ n1770;
  assign n3352 = n1748 & ~n1751;
  assign n3806 = n3352 ^ n1762;
  assign n3809 = n3808 ^ n3806;
  assign n3810 = n3809 ^ n3806;
  assign n3811 = ~n1516 & ~n3810;
  assign n3812 = n3811 ^ n3806;
  assign n3813 = n1761 & n3812;
  assign n3814 = n3813 ^ n3806;
  assign n3815 = ~n3805 & ~n3814;
  assign n3816 = n1761 & n1771;
  assign n3817 = n1796 ^ n1782;
  assign n3818 = n3817 ^ n1775;
  assign n3819 = n1759 & ~n3818;
  assign n3820 = ~n3816 & ~n3819;
  assign n3821 = n3815 & n3820;
  assign n3822 = ~n1789 & n3821;
  assign n3823 = ~n3803 & n3822;
  assign n3824 = ~n3351 & n3823;
  assign n3825 = ~n3802 & n3824;
  assign n3826 = ~n3362 & n3825;
  assign n3827 = n3826 ^ x38;
  assign n3828 = n3827 ^ x200;
  assign n3835 = ~n3764 & n3828;
  assign n3836 = n3835 ^ n3764;
  assign n3842 = n3836 ^ n3828;
  assign n3853 = n3842 ^ n3764;
  assign n3854 = n3840 & n3853;
  assign n3844 = n3828 ^ n3764;
  assign n3845 = ~n3839 & ~n3844;
  assign n3846 = n3845 ^ n3839;
  assign n3843 = ~n3839 & n3842;
  assign n3847 = n3846 ^ n3843;
  assign n3870 = n3854 ^ n3847;
  assign n3871 = n3870 ^ n3843;
  assign n3858 = n3840 & n3842;
  assign n3872 = n3871 ^ n3858;
  assign n3873 = n3872 ^ n3797;
  assign n3863 = n3838 & n3842;
  assign n3849 = n3834 & n3835;
  assign n3850 = n3849 ^ n3835;
  assign n3841 = n3835 & n3840;
  assign n3848 = n3847 ^ n3841;
  assign n3851 = n3850 ^ n3848;
  assign n3864 = n3863 ^ n3851;
  assign n3857 = n3848 ^ n3843;
  assign n3859 = n3858 ^ n3857;
  assign n3837 = n3834 & ~n3836;
  assign n3852 = n3851 ^ n3837;
  assign n3855 = n3854 ^ n3852;
  assign n3798 = n3797 ^ n3764;
  assign n3800 = n3799 ^ n3797;
  assign n3829 = n3828 ^ n3800;
  assign n3830 = ~n3764 & n3829;
  assign n3831 = n3830 ^ n3828;
  assign n3832 = ~n3798 & ~n3831;
  assign n3833 = n3832 ^ n3829;
  assign n3856 = n3855 ^ n3833;
  assign n3860 = n3859 ^ n3856;
  assign n3862 = n3860 ^ n3838;
  assign n3865 = n3864 ^ n3862;
  assign n3866 = n3865 ^ n3841;
  assign n3867 = n3866 ^ n3800;
  assign n3861 = n3860 ^ n3854;
  assign n3868 = n3867 ^ n3861;
  assign n3869 = n3868 ^ n3844;
  assign n3874 = n3873 ^ n3869;
  assign n3875 = n3874 ^ n3834;
  assign n3876 = n3875 ^ n3849;
  assign n3877 = n3876 ^ n3860;
  assign n3878 = n3877 ^ n3864;
  assign n3879 = ~n3762 & n3878;
  assign n3880 = n3879 ^ n3877;
  assign n3881 = n3761 & ~n3880;
  assign n3883 = n3762 ^ n3761;
  assign n3882 = n3761 & n3762;
  assign n3884 = n3883 ^ n3882;
  assign n3885 = n3865 & ~n3884;
  assign n3887 = n3843 & n3882;
  assign n3886 = n3874 & ~n3884;
  assign n3888 = n3887 ^ n3886;
  assign n3889 = ~n3761 & ~n3861;
  assign n3890 = n3889 ^ n3854;
  assign n3891 = ~n3762 & n3890;
  assign n3897 = n3858 ^ n3847;
  assign n3899 = n3897 ^ n3837;
  assign n3900 = n3899 ^ n3866;
  assign n3895 = ~n3839 & n3853;
  assign n3893 = n3872 ^ n3799;
  assign n3892 = n3845 ^ n3841;
  assign n3894 = n3893 ^ n3892;
  assign n3896 = n3895 ^ n3894;
  assign n3898 = n3897 ^ n3896;
  assign n3901 = n3900 ^ n3898;
  assign n3902 = n3901 ^ n3898;
  assign n3903 = n3761 & ~n3902;
  assign n3904 = n3903 ^ n3898;
  assign n3905 = n3762 & ~n3904;
  assign n3906 = n3905 ^ n3898;
  assign n3907 = n3876 ^ n3833;
  assign n3908 = n3762 & n3907;
  assign n3909 = n3908 ^ n3876;
  assign n3910 = n3883 & n3909;
  assign n3911 = n3906 & ~n3910;
  assign n3912 = ~n3891 & n3911;
  assign n3913 = ~n3888 & n3912;
  assign n3914 = ~n3885 & n3913;
  assign n3915 = ~n3881 & n3914;
  assign n3916 = n3915 ^ n929;
  assign n6044 = n3916 ^ x226;
  assign n2882 = n2509 ^ x153;
  assign n2883 = n2211 ^ x148;
  assign n2889 = n2056 ^ x149;
  assign n2890 = ~n1519 & n1908;
  assign n2891 = n1599 ^ n1546;
  assign n2892 = ~n1553 & n2891;
  assign n2896 = n1559 ^ n1549;
  assign n2897 = n2896 ^ n1564;
  assign n2894 = ~n1522 & n1562;
  assign n2893 = n1567 ^ n1560;
  assign n2895 = n2894 ^ n2893;
  assign n2898 = n2897 ^ n2895;
  assign n2899 = n2898 ^ n2895;
  assign n2900 = ~n1518 & n2899;
  assign n2901 = n2900 ^ n2895;
  assign n2902 = ~n1517 & n2901;
  assign n2903 = n2902 ^ n2895;
  assign n2904 = ~n2892 & ~n2903;
  assign n2905 = ~n2890 & n2904;
  assign n2907 = n1542 ^ n1538;
  assign n2906 = n1588 ^ n1578;
  assign n2908 = n2907 ^ n2906;
  assign n2909 = n1518 & n2908;
  assign n2910 = n2909 ^ n2906;
  assign n2911 = ~n1517 & ~n2910;
  assign n2912 = n2905 & ~n2911;
  assign n2913 = ~n2073 & n2912;
  assign n2914 = ~n1552 & n2913;
  assign n2915 = ~n1905 & n2914;
  assign n2916 = n2915 ^ x47;
  assign n2917 = n2916 ^ x151;
  assign n2918 = ~n2889 & ~n2917;
  assign n2919 = n2918 ^ n2917;
  assign n2884 = n2622 ^ x152;
  assign n2885 = n2065 ^ n2060;
  assign n2886 = n2885 ^ x55;
  assign n2887 = n2886 ^ x150;
  assign n2888 = n2884 & ~n2887;
  assign n2922 = n2888 ^ n2884;
  assign n2923 = ~n2919 & n2922;
  assign n2968 = n2923 ^ n2919;
  assign n2939 = n2887 ^ n2884;
  assign n2940 = n2939 ^ n2889;
  assign n2941 = n2940 ^ n2917;
  assign n2942 = ~n2919 & ~n2941;
  assign n2969 = n2968 ^ n2942;
  assign n3397 = n2969 ^ n2923;
  assign n2920 = n2919 ^ n2889;
  assign n2970 = ~n2920 & n2922;
  assign n2990 = n2970 ^ n2920;
  assign n2951 = n2884 & ~n2917;
  assign n2952 = n2951 ^ n2887;
  assign n2953 = ~n2889 & n2952;
  assign n2954 = n2953 ^ n2889;
  assign n2924 = n2922 ^ n2887;
  assign n2947 = n2918 & n2924;
  assign n2925 = ~n2919 & n2924;
  assign n2943 = n2942 ^ n2925;
  assign n2926 = n2925 ^ n2923;
  assign n2928 = n2926 ^ n2888;
  assign n2944 = n2943 ^ n2928;
  assign n2929 = n2917 ^ n2887;
  assign n2930 = n2928 & n2929;
  assign n2945 = n2944 ^ n2930;
  assign n2935 = n2918 ^ n2889;
  assign n2936 = n2922 & ~n2935;
  assign n2946 = n2945 ^ n2936;
  assign n2948 = n2947 ^ n2946;
  assign n2932 = n2888 ^ n2887;
  assign n2933 = n2918 & ~n2932;
  assign n2937 = n2936 ^ n2933;
  assign n2938 = n2937 ^ n2918;
  assign n2949 = n2948 ^ n2938;
  assign n2921 = n2888 & ~n2920;
  assign n2927 = n2926 ^ n2921;
  assign n2931 = n2930 ^ n2927;
  assign n2934 = n2933 ^ n2931;
  assign n2950 = n2949 ^ n2934;
  assign n2955 = n2954 ^ n2950;
  assign n2977 = n2955 ^ n2947;
  assign n2978 = n2977 ^ n2924;
  assign n2973 = n2953 ^ n2948;
  assign n2974 = n2973 ^ n2949;
  assign n2975 = n2974 ^ n2925;
  assign n2972 = n2955 ^ n2949;
  assign n2976 = n2975 ^ n2972;
  assign n2979 = n2978 ^ n2976;
  assign n2980 = n2979 ^ n2921;
  assign n2991 = n2990 ^ n2980;
  assign n2992 = n2991 ^ n2943;
  assign n3398 = n3397 ^ n2992;
  assign n3399 = n2883 & n3398;
  assign n3400 = n3399 ^ n3397;
  assign n3401 = n2882 & ~n3400;
  assign n2960 = ~n2882 & ~n2883;
  assign n2966 = n2960 ^ n2882;
  assign n3402 = n2966 ^ n2883;
  assign n3403 = n2979 & ~n3402;
  assign n3404 = ~n3401 & ~n3403;
  assign n2965 = n2960 ^ n2883;
  assign n2967 = n2966 ^ n2965;
  assign n3405 = ~n2882 & n2946;
  assign n3406 = n3405 ^ n2936;
  assign n3407 = n2967 & n3406;
  assign n3408 = ~n2882 & ~n2977;
  assign n3409 = n3408 ^ n2947;
  assign n3410 = n2883 & n3409;
  assign n3411 = n2966 ^ n2949;
  assign n2994 = n2979 ^ n2943;
  assign n3412 = n2994 ^ n2921;
  assign n3413 = n3412 ^ n2969;
  assign n3414 = n3413 ^ n2947;
  assign n3415 = n3414 ^ n2965;
  assign n3416 = ~n2966 & ~n3415;
  assign n3417 = n3416 ^ n2965;
  assign n3418 = ~n3411 & n3417;
  assign n3419 = n3418 ^ n2949;
  assign n3427 = n2940 ^ n2930;
  assign n3428 = ~n2883 & n3427;
  assign n3422 = n2980 ^ n2933;
  assign n3423 = n3422 ^ n2955;
  assign n3420 = n2934 ^ n2923;
  assign n3421 = n3420 ^ n2945;
  assign n3424 = n3423 ^ n3421;
  assign n3425 = ~n2883 & ~n3424;
  assign n3426 = n3425 ^ n3421;
  assign n3429 = n3428 ^ n3426;
  assign n3430 = ~n2882 & n3429;
  assign n3431 = n3430 ^ n3426;
  assign n3432 = ~n3419 & ~n3431;
  assign n3433 = ~n3410 & n3432;
  assign n3434 = ~n3407 & n3433;
  assign n3435 = n3404 & n3434;
  assign n3436 = n3435 ^ x6;
  assign n3437 = n3436 ^ x160;
  assign n2626 = ~n2597 & ~n2625;
  assign n2648 = n2586 & ~n2625;
  assign n2647 = n2623 & ~n2646;
  assign n2649 = n2648 ^ n2647;
  assign n2855 = n2630 & ~n2662;
  assign n2856 = ~n2595 & ~n2623;
  assign n2857 = n2856 ^ n2594;
  assign n2858 = ~n2598 & ~n2857;
  assign n2859 = ~n2598 & n2629;
  assign n2860 = n2859 ^ n2656;
  assign n2861 = n2623 & ~n2860;
  assign n2862 = n2861 ^ n2656;
  assign n2866 = n2597 ^ n2584;
  assign n2867 = n2866 ^ n2632;
  assign n2864 = n2594 ^ n2587;
  assign n2863 = n2636 ^ n2591;
  assign n2865 = n2864 ^ n2863;
  assign n2868 = n2867 ^ n2865;
  assign n2869 = ~n2623 & ~n2868;
  assign n2870 = n2869 ^ n2865;
  assign n2871 = n2870 ^ n2588;
  assign n2872 = n2598 & n2871;
  assign n2873 = n2872 ^ n2588;
  assign n2874 = n2862 & ~n2873;
  assign n2875 = ~n2858 & n2874;
  assign n2876 = ~n2855 & n2875;
  assign n2877 = ~n2649 & n2876;
  assign n2878 = n2854 & n2877;
  assign n2879 = ~n2626 & n2878;
  assign n2880 = n2879 ^ x24;
  assign n3438 = n2880 ^ x165;
  assign n3288 = n1901 ^ n1869;
  assign n3297 = n3288 ^ n1955;
  assign n3298 = ~n1901 & n3297;
  assign n3296 = n1869 & n2017;
  assign n3299 = n3298 ^ n3296;
  assign n3293 = n1953 ^ n1951;
  assign n3294 = n1903 ^ n1901;
  assign n3295 = ~n3293 & n3294;
  assign n3300 = n3299 ^ n3295;
  assign n3289 = n3288 ^ n1937;
  assign n3290 = n3289 ^ n2008;
  assign n3291 = n3290 ^ n2010;
  assign n3292 = n1870 & n3291;
  assign n3301 = n3300 ^ n3292;
  assign n3302 = ~n1963 & ~n3301;
  assign n3277 = n1949 & n2017;
  assign n3278 = n2021 ^ n1950;
  assign n3279 = n3278 ^ n2015;
  assign n3280 = n3279 ^ n1960;
  assign n3281 = n3280 ^ n1954;
  assign n3282 = ~n1870 & ~n3281;
  assign n3283 = n3282 ^ n1954;
  assign n3284 = ~n3277 & ~n3283;
  assign n3285 = ~n1945 & n3284;
  assign n3286 = ~n1963 & n3285;
  assign n3303 = n3302 ^ n3286;
  assign n3304 = n2004 & ~n3303;
  assign n3287 = n3286 ^ n2004;
  assign n3305 = n3304 ^ n3287;
  assign n3306 = n3305 ^ x56;
  assign n3307 = n3306 ^ x161;
  assign n3174 = ~n3115 & ~n3129;
  assign n3175 = n3174 ^ n3114;
  assign n3313 = n3046 & n3175;
  assign n3314 = n3111 ^ n3109;
  assign n3315 = n3314 ^ n3126;
  assign n3316 = n3315 ^ n3119;
  assign n3317 = n3316 ^ n3125;
  assign n3318 = ~n3129 & n3317;
  assign n3319 = n3318 ^ n3125;
  assign n3320 = n3046 & n3319;
  assign n3321 = n3320 ^ n3125;
  assign n3127 = n3126 ^ n3101;
  assign n3330 = n3127 ^ n3095;
  assign n3331 = n3330 ^ n3111;
  assign n3323 = n3149 ^ n3123;
  assign n3324 = n3322 & n3323;
  assign n3325 = ~n3104 & n3324;
  assign n3327 = n3326 ^ n3103;
  assign n3328 = ~n3141 & n3327;
  assign n3329 = ~n3325 & ~n3328;
  assign n3332 = n3331 ^ n3329;
  assign n3333 = n3332 ^ n3329;
  assign n3334 = n3129 & ~n3333;
  assign n3335 = n3334 ^ n3329;
  assign n3336 = n3046 & n3335;
  assign n3337 = n3336 ^ n3329;
  assign n3338 = ~n3321 & ~n3337;
  assign n3339 = n3129 ^ n3046;
  assign n3340 = ~n3127 & n3129;
  assign n3341 = n3340 ^ n3110;
  assign n3342 = n3339 & n3341;
  assign n3343 = n3342 ^ n3110;
  assign n3344 = n3338 & ~n3343;
  assign n3345 = ~n3313 & n3344;
  assign n3346 = n3140 & n3345;
  assign n3347 = n3346 ^ x40;
  assign n3348 = n3347 ^ x163;
  assign n1753 = n1752 ^ n1749;
  assign n1754 = n1516 & n1753;
  assign n1755 = n1754 ^ n1749;
  assign n1756 = ~n1483 & n1755;
  assign n3353 = n1761 & n3352;
  assign n1816 = n1815 ^ n1770;
  assign n1817 = n1516 & n1816;
  assign n1821 = n1817 ^ n1815;
  assign n3354 = n1821 ^ n1763;
  assign n3355 = n1483 & n3354;
  assign n3356 = n3355 ^ n1763;
  assign n3357 = n1777 ^ n1762;
  assign n3358 = n1483 & ~n3357;
  assign n3359 = n3358 ^ n1777;
  assign n3360 = n1761 & ~n3359;
  assign n3365 = n1775 ^ n1768;
  assign n3363 = n3352 ^ n1774;
  assign n3364 = n3363 ^ n1767;
  assign n3366 = n3365 ^ n3364;
  assign n3367 = n1516 & ~n3366;
  assign n3368 = n3367 ^ n3364;
  assign n1814 = n1516 & n1770;
  assign n3369 = n3368 ^ n1814;
  assign n3370 = n1761 & n3369;
  assign n3371 = n3370 ^ n3368;
  assign n3372 = ~n3362 & ~n3371;
  assign n3373 = ~n3360 & n3372;
  assign n3374 = ~n3356 & n3373;
  assign n3375 = ~n3353 & n3374;
  assign n3377 = n3376 ^ n1774;
  assign n3378 = n3377 ^ n1794;
  assign n3379 = ~n1516 & ~n3378;
  assign n3380 = n3379 ^ n1794;
  assign n3381 = n1483 & ~n3380;
  assign n3382 = n3375 & ~n3381;
  assign n3383 = n1796 ^ n1758;
  assign n3384 = n1790 ^ n1760;
  assign n3385 = ~n1758 & n3384;
  assign n3386 = n3385 ^ n1760;
  assign n3387 = n3383 & ~n3386;
  assign n3388 = n3387 ^ n1796;
  assign n3389 = n3382 & n3388;
  assign n3390 = ~n3351 & n3389;
  assign n3391 = ~n1756 & n3390;
  assign n3392 = n3391 ^ x48;
  assign n3393 = n3392 ^ x162;
  assign n3394 = ~n3348 & ~n3393;
  assign n3441 = n3307 & n3394;
  assign n3467 = n3441 ^ n3394;
  assign n2811 = ~n2072 & n2258;
  assign n2270 = n2245 ^ n2223;
  assign n2271 = ~n2071 & ~n2270;
  assign n2812 = n2811 ^ n2271;
  assign n2278 = ~n2071 & ~n2250;
  assign n2813 = n2245 ^ n2218;
  assign n2814 = ~n2069 & n2813;
  assign n2815 = n2235 ^ n2219;
  assign n2816 = n2072 & ~n2815;
  assign n2817 = ~n2254 & ~n2816;
  assign n2818 = n2817 ^ n2070;
  assign n2819 = n2250 ^ n2220;
  assign n2820 = n2819 ^ n2289;
  assign n2821 = n2817 & ~n2820;
  assign n2822 = n2821 ^ n2289;
  assign n2823 = n2818 & n2822;
  assign n2824 = n2823 ^ n2070;
  assign n2825 = ~n2814 & ~n2824;
  assign n2833 = n2057 & ~n2236;
  assign n2826 = n2239 ^ n2057;
  assign n2827 = ~n2254 & n2826;
  assign n2828 = n2827 ^ n2057;
  assign n2829 = n2243 & ~n2828;
  assign n2830 = n2829 ^ n2242;
  assign n2831 = ~n2231 & ~n2830;
  assign n2832 = ~n2233 & n2831;
  assign n2834 = n2833 ^ n2832;
  assign n2835 = ~n2254 & ~n2834;
  assign n2836 = n2835 ^ n2832;
  assign n2837 = n2825 & n2836;
  assign n2838 = ~n2057 & ~n2224;
  assign n2839 = n2838 ^ n2223;
  assign n2840 = ~n2069 & ~n2839;
  assign n2841 = n2837 & ~n2840;
  assign n2842 = ~n2278 & n2841;
  assign n2843 = ~n2812 & n2842;
  assign n2844 = ~n2810 & n2843;
  assign n2845 = n2844 ^ x32;
  assign n3308 = n2845 ^ x164;
  assign n3309 = ~n3307 & ~n3308;
  assign n3453 = n3309 & n3394;
  assign n3468 = n3467 ^ n3453;
  assign n3310 = n3309 ^ n3307;
  assign n3311 = n3310 ^ n3308;
  assign n3312 = n3311 ^ n3307;
  assign n3395 = n3394 ^ n3348;
  assign n3444 = n3395 ^ n3393;
  assign n3445 = ~n3312 & ~n3444;
  assign n4494 = n3468 ^ n3445;
  assign n4495 = n3438 & n4494;
  assign n4496 = n4495 ^ n3468;
  assign n4497 = ~n3437 & n4496;
  assign n3456 = ~n3310 & ~n3395;
  assign n3452 = n3309 & ~n3395;
  assign n3454 = n3453 ^ n3452;
  assign n3450 = n3309 & ~n3444;
  assign n3451 = n3450 ^ n3309;
  assign n3455 = n3454 ^ n3451;
  assign n3457 = n3456 ^ n3455;
  assign n3439 = n3437 & ~n3438;
  assign n3440 = n3439 ^ n3437;
  assign n3458 = n3440 ^ n3438;
  assign n3459 = n3457 & n3458;
  assign n3460 = ~n3310 & ~n3444;
  assign n3447 = n3441 ^ n3312;
  assign n3442 = n3308 & n3441;
  assign n3396 = ~n3312 & ~n3395;
  assign n3443 = n3442 ^ n3396;
  assign n3446 = n3445 ^ n3443;
  assign n3448 = n3447 ^ n3446;
  assign n3461 = n3460 ^ n3448;
  assign n3462 = n3438 & ~n3461;
  assign n3463 = n3462 ^ n3448;
  assign n3464 = ~n3437 & ~n3463;
  assign n3465 = ~n3459 & ~n3464;
  assign n3466 = n3438 ^ n3437;
  assign n3475 = n3456 ^ n3452;
  assign n3476 = n3475 ^ n3395;
  assign n3477 = n3476 ^ n3396;
  assign n4502 = n3438 & ~n3477;
  assign n3479 = n3442 ^ n3311;
  assign n3473 = n3444 ^ n3348;
  assign n3474 = ~n3311 & ~n3473;
  assign n3478 = n3477 ^ n3474;
  assign n3480 = n3479 ^ n3478;
  assign n4498 = n3480 ^ n3456;
  assign n4499 = n4498 ^ n3460;
  assign n4500 = ~n3438 & n4499;
  assign n4501 = n4500 ^ n3460;
  assign n4503 = n4502 ^ n4501;
  assign n4504 = n3466 & n4503;
  assign n4505 = n4504 ^ n4501;
  assign n4506 = n3456 ^ n3443;
  assign n4507 = n3438 & n4506;
  assign n4508 = n4507 ^ n3456;
  assign n4509 = n3466 & n4508;
  assign n4510 = n3452 ^ n3440;
  assign n4511 = n3453 ^ n3438;
  assign n4512 = ~n3452 & n4511;
  assign n4513 = n4512 ^ n3438;
  assign n4514 = n4510 & ~n4513;
  assign n4515 = n4514 ^ n3440;
  assign n3492 = ~n3310 & ~n3473;
  assign n4517 = n3439 & n3492;
  assign n4516 = n3437 & n3468;
  assign n4518 = n4517 ^ n4516;
  assign n4519 = ~n4515 & ~n4518;
  assign n4528 = n3474 ^ n3396;
  assign n4529 = n4528 ^ n3450;
  assign n4530 = ~n3438 & n4529;
  assign n4525 = n3440 & n3474;
  assign n3489 = n3442 ^ n3441;
  assign n4526 = n4525 ^ n3489;
  assign n4523 = ~n3439 & ~n3445;
  assign n3500 = n3477 ^ n3445;
  assign n4520 = n3500 ^ n3480;
  assign n4521 = n4520 ^ n3439;
  assign n4522 = n3500 & ~n4521;
  assign n4524 = n4523 ^ n4522;
  assign n4527 = n4526 ^ n4524;
  assign n4531 = n4530 ^ n4527;
  assign n4532 = ~n3437 & ~n4531;
  assign n4533 = n4532 ^ n4527;
  assign n4534 = ~n3438 & ~n3448;
  assign n4535 = n4534 ^ n3448;
  assign n3449 = n3440 & ~n3448;
  assign n4536 = n4535 ^ n3449;
  assign n4537 = n4533 & n4536;
  assign n4538 = n4519 & n4537;
  assign n4539 = ~n4509 & n4538;
  assign n4540 = ~n4505 & n4539;
  assign n4541 = n3465 & n4540;
  assign n4542 = ~n4497 & n4541;
  assign n4543 = n4542 ^ n2003;
  assign n6045 = n4543 ^ x231;
  assign n6046 = n6044 & n6045;
  assign n6047 = n6046 ^ n6045;
  assign n2328 = n1342 & ~n1387;
  assign n2329 = n1383 ^ n1345;
  assign n2330 = n1315 & ~n2329;
  assign n2333 = n2332 ^ n1387;
  assign n2334 = n1352 ^ n1314;
  assign n2335 = ~n2332 & ~n2334;
  assign n2336 = n2335 ^ n1352;
  assign n2337 = ~n2333 & n2336;
  assign n2338 = n2337 ^ n1387;
  assign n2339 = n1381 ^ n1349;
  assign n2340 = ~n1315 & ~n2339;
  assign n2341 = n2340 ^ n1349;
  assign n2342 = n1316 & n2341;
  assign n2343 = n2338 & ~n2342;
  assign n2344 = ~n1353 & n2343;
  assign n2345 = ~n2330 & n2344;
  assign n2346 = ~n2328 & n2345;
  assign n2347 = ~n2327 & n2346;
  assign n2348 = ~n2324 & n2347;
  assign n2349 = n2348 ^ x49;
  assign n2350 = n2349 ^ x114;
  assign n2354 = n1212 ^ n1211;
  assign n2355 = n1884 ^ n1250;
  assign n2356 = n2355 ^ n1254;
  assign n2357 = n2356 ^ n1214;
  assign n2358 = ~n2354 & n2357;
  assign n2352 = n1215 ^ n1214;
  assign n2353 = n2352 ^ n1211;
  assign n2359 = n2358 ^ n2353;
  assign n2360 = ~n1210 & n2359;
  assign n2351 = n1253 ^ n1224;
  assign n2361 = n2360 ^ n2351;
  assign n2362 = n1209 & n2361;
  assign n2364 = n2354 ^ n1280;
  assign n2365 = n2364 ^ n2358;
  assign n2363 = n1215 ^ n1212;
  assign n2366 = n2365 ^ n2363;
  assign n2367 = n2366 ^ n1245;
  assign n2368 = n1268 & n2367;
  assign n2369 = n2368 ^ n1245;
  assign n2370 = ~n2362 & ~n2369;
  assign n2371 = n1285 ^ n1267;
  assign n2372 = n1885 ^ n1259;
  assign n2373 = ~n1267 & ~n2372;
  assign n2374 = n2373 ^ n1259;
  assign n2375 = ~n2371 & ~n2374;
  assign n2376 = n2375 ^ n1285;
  assign n2377 = n2370 & ~n2376;
  assign n2378 = ~n1273 & n2377;
  assign n2379 = ~n1265 & n2378;
  assign n2380 = n2379 ^ x41;
  assign n2381 = n2380 ^ x115;
  assign n2382 = n2350 & ~n2381;
  assign n2383 = n2382 ^ n2381;
  assign n2396 = n2395 ^ x113;
  assign n2397 = n1515 ^ x116;
  assign n2398 = n2396 & ~n2397;
  assign n2399 = n2398 ^ n2396;
  assign n2421 = ~n2383 & n2399;
  assign n2422 = n2421 ^ n2399;
  assign n2384 = n2383 ^ n2350;
  assign n2419 = n2384 & n2399;
  assign n2403 = n2382 ^ n2350;
  assign n2404 = n2399 & n2403;
  assign n2420 = n2419 ^ n2404;
  assign n2423 = n2422 ^ n2420;
  assign n2434 = n2423 ^ n2382;
  assign n2400 = n2399 ^ n2397;
  assign n2418 = n2400 & n2403;
  assign n2431 = n2418 ^ n2400;
  assign n2424 = n2423 ^ n2418;
  assign n2412 = n2384 & n2398;
  assign n2427 = n2424 ^ n2412;
  assign n2428 = n2427 ^ n2384;
  assign n2401 = n2400 ^ n2396;
  assign n2402 = n2384 & ~n2401;
  assign n2425 = n2424 ^ n2402;
  assign n2426 = n2425 ^ n2419;
  assign n2429 = n2428 ^ n2426;
  assign n2417 = ~n2383 & n2400;
  assign n2430 = n2429 ^ n2417;
  assign n2432 = n2431 ^ n2430;
  assign n2416 = n2382 & ~n2401;
  assign n2433 = n2432 ^ n2416;
  assign n2435 = n2434 ^ n2433;
  assign n2304 = n1615 ^ x117;
  assign n2320 = n2319 ^ x112;
  assign n2405 = n2404 ^ n2402;
  assign n2406 = ~n2320 & n2405;
  assign n2407 = n2406 ^ n2404;
  assign n2408 = n2304 & n2407;
  assign n2409 = ~n2304 & n2320;
  assign n2454 = n2409 ^ n2304;
  assign n2455 = n2412 & ~n2454;
  assign n2776 = n2304 & n2404;
  assign n2413 = ~n2383 & n2398;
  assign n2414 = n2413 ^ n2412;
  assign n2415 = n2414 ^ n2398;
  assign n2436 = n2435 ^ n2415;
  assign n2773 = n2436 ^ n2433;
  assign n2774 = n2304 & n2773;
  assign n2775 = n2774 ^ n2436;
  assign n2777 = n2776 ^ n2775;
  assign n2778 = ~n2320 & n2777;
  assign n2779 = n2778 ^ n2775;
  assign n2437 = n2436 ^ n2421;
  assign n2780 = n2320 & n2437;
  assign n2781 = n2780 ^ n2436;
  assign n2782 = ~n2304 & n2781;
  assign n2785 = n2402 & n2409;
  assign n2410 = n2409 ^ n2320;
  assign n2783 = n2410 & n2412;
  assign n2449 = ~n2304 & n2433;
  assign n2442 = n2417 ^ n2416;
  assign n2443 = ~n2304 & n2442;
  assign n2450 = n2449 ^ n2443;
  assign n2451 = n2450 ^ n2432;
  assign n2452 = ~n2320 & n2451;
  assign n2784 = n2783 ^ n2452;
  assign n2786 = n2785 ^ n2784;
  assign n2446 = n2304 & n2430;
  assign n2447 = n2446 ^ n2429;
  assign n2448 = n2320 & n2447;
  assign n2440 = n2410 & n2413;
  assign n2467 = n2320 ^ n2304;
  assign n2469 = ~n2383 & ~n2401;
  assign n2470 = n2469 ^ n2418;
  assign n2471 = n2470 ^ n2419;
  assign n2793 = n2471 ^ n2417;
  assign n2792 = n2424 ^ n2416;
  assign n2794 = n2793 ^ n2792;
  assign n2795 = ~n2320 & n2794;
  assign n2796 = n2795 ^ n2792;
  assign n2468 = ~n2401 & n2403;
  assign n2787 = n2468 ^ n2429;
  assign n2456 = n2423 ^ n2413;
  assign n2788 = n2787 ^ n2456;
  assign n2789 = n2788 ^ n2468;
  assign n2790 = ~n2320 & n2789;
  assign n2791 = n2790 ^ n2468;
  assign n2797 = n2796 ^ n2791;
  assign n2798 = ~n2467 & n2797;
  assign n2799 = n2798 ^ n2796;
  assign n2800 = ~n2440 & ~n2799;
  assign n2801 = ~n2448 & n2800;
  assign n2802 = ~n2786 & n2801;
  assign n2803 = ~n2782 & n2802;
  assign n2804 = ~n2779 & n2803;
  assign n2805 = ~n2455 & n2804;
  assign n2806 = ~n2408 & n2805;
  assign n2807 = ~n2435 & n2806;
  assign n2808 = n2807 ^ x58;
  assign n2809 = n2808 ^ x171;
  assign n2846 = n2845 ^ x166;
  assign n2847 = n2809 & n2846;
  assign n2848 = n2847 ^ n2809;
  assign n2956 = n2955 ^ n2925;
  assign n2957 = ~n2883 & ~n2956;
  assign n2958 = n2957 ^ n2925;
  assign n2959 = n2882 & n2958;
  assign n2961 = n2950 ^ n2925;
  assign n2962 = n2961 ^ n2923;
  assign n2963 = ~n2960 & n2962;
  assign n2964 = n2963 ^ n2961;
  assign n2982 = n2942 ^ n2941;
  assign n2971 = n2970 ^ n2969;
  assign n2981 = n2980 ^ n2971;
  assign n2983 = n2982 ^ n2981;
  assign n2984 = n2882 & n2983;
  assign n2985 = n2984 ^ n2981;
  assign n2986 = n2985 ^ n2953;
  assign n2987 = ~n2967 & ~n2986;
  assign n2988 = n2987 ^ n2953;
  assign n2989 = ~n2964 & ~n2988;
  assign n2993 = n2992 ^ n2955;
  assign n2995 = n2994 ^ n2993;
  assign n2996 = ~n2882 & n2995;
  assign n2997 = n2996 ^ n2994;
  assign n2998 = n2967 & n2997;
  assign n2999 = n2989 & ~n2998;
  assign n3000 = ~n2959 & n2999;
  assign n3001 = n3000 ^ x8;
  assign n3002 = n3001 ^ x169;
  assign n1408 = n1208 & n1407;
  assign n1459 = n1443 ^ n1417;
  assign n1460 = ~n1407 & n1459;
  assign n1461 = ~n1413 & n1460;
  assign n3011 = n1461 ^ n1458;
  assign n1462 = ~n1458 & n1461;
  assign n3012 = n3011 ^ n1462;
  assign n3013 = ~n3010 & ~n3012;
  assign n1433 = ~n1409 & n1432;
  assign n1434 = n1433 ^ n1431;
  assign n1450 = n1449 ^ n1435;
  assign n3019 = n1407 & n1450;
  assign n3020 = n1415 ^ n1203;
  assign n3021 = n3020 ^ n1445;
  assign n3022 = n1455 & n3021;
  assign n3023 = n1405 & n3014;
  assign n3026 = ~n1405 & n1444;
  assign n3027 = ~n1460 & ~n3026;
  assign n3028 = n1423 & ~n3027;
  assign n3024 = n1458 ^ n1420;
  assign n3025 = n3024 ^ n1441;
  assign n3029 = n3028 ^ n3025;
  assign n3030 = n3029 ^ n3025;
  assign n3031 = ~n1455 & ~n3030;
  assign n3032 = n3031 ^ n3025;
  assign n3033 = n1406 & ~n3032;
  assign n3034 = n3033 ^ n3025;
  assign n3035 = ~n3023 & n3034;
  assign n3036 = ~n3022 & n3035;
  assign n3037 = ~n3019 & n3036;
  assign n3038 = ~n3018 & n3037;
  assign n3039 = n1434 & n3038;
  assign n3040 = n3013 & n3039;
  assign n3041 = ~n1408 & n3040;
  assign n3042 = n3041 ^ x16;
  assign n3043 = n3042 ^ x168;
  assign n3044 = n3002 & ~n3043;
  assign n3045 = n3044 ^ n3002;
  assign n2881 = n2880 ^ x167;
  assign n3130 = ~n3100 & n3129;
  assign n3128 = n3127 ^ n3099;
  assign n3131 = n3130 ^ n3128;
  assign n3132 = ~n3046 & n3131;
  assign n3163 = n3125 ^ n3117;
  assign n3164 = n3163 ^ n3111;
  assign n3168 = n3167 ^ n3164;
  assign n3169 = n3046 & n3168;
  assign n3170 = n3169 ^ n3167;
  assign n3159 = n3114 ^ n3104;
  assign n3160 = n3159 ^ n3145;
  assign n3161 = n3046 & ~n3160;
  assign n3162 = n3161 ^ n3159;
  assign n3171 = n3170 ^ n3162;
  assign n3172 = ~n3129 & n3171;
  assign n3173 = n3172 ^ n3162;
  assign n3176 = n3175 ^ n3109;
  assign n3177 = ~n3046 & n3176;
  assign n3178 = n3177 ^ n3175;
  assign n3179 = ~n3173 & ~n3178;
  assign n3180 = ~n3158 & n3179;
  assign n3181 = n3152 & n3180;
  assign n3182 = ~n3132 & n3181;
  assign n3183 = n3182 ^ x0;
  assign n3184 = n3183 ^ x170;
  assign n3187 = n2881 & n3184;
  assign n3195 = n3045 & n3187;
  assign n3188 = n3187 ^ n3184;
  assign n3192 = n3045 & n3188;
  assign n3193 = n3192 ^ n3045;
  assign n3189 = n3188 ^ n2881;
  assign n3190 = n3189 ^ n3184;
  assign n3185 = n3184 ^ n3045;
  assign n3186 = n2881 & ~n3185;
  assign n3191 = n3190 ^ n3186;
  assign n3194 = n3193 ^ n3191;
  assign n3196 = n3195 ^ n3194;
  assign n3197 = n3196 ^ n3193;
  assign n3198 = n2848 & n3197;
  assign n3199 = n2848 ^ n2846;
  assign n3200 = n3199 ^ n2847;
  assign n3206 = n3184 ^ n3002;
  assign n3207 = n3206 ^ n3186;
  assign n3208 = n3207 ^ n3044;
  assign n3203 = n3045 ^ n3043;
  assign n3204 = ~n3189 & n3203;
  assign n3201 = n3044 & ~n3189;
  assign n3202 = n3201 ^ n3192;
  assign n3205 = n3204 ^ n3202;
  assign n3209 = n3208 ^ n3205;
  assign n3210 = n3209 ^ n3194;
  assign n3211 = n2846 & ~n3210;
  assign n3212 = n3211 ^ n3194;
  assign n3213 = ~n3200 & n3212;
  assign n3214 = ~n3198 & ~n3213;
  assign n3215 = n3203 ^ n3002;
  assign n3216 = n3190 & ~n3215;
  assign n3217 = n3216 ^ n3204;
  assign n3218 = ~n2846 & n3217;
  assign n3219 = n3218 ^ n3204;
  assign n3220 = n2809 & n3219;
  assign n3223 = n3044 & n3187;
  assign n3224 = n2848 & n3223;
  assign n3221 = n3199 ^ n2809;
  assign n3222 = n3202 & n3221;
  assign n3225 = n3224 ^ n3222;
  assign n3227 = n2881 & n3203;
  assign n3226 = n3204 ^ n3203;
  assign n3228 = n3227 ^ n3226;
  assign n3229 = n3228 ^ n3209;
  assign n3230 = n3221 & ~n3229;
  assign n3231 = n3187 & ~n3215;
  assign n3232 = n3221 & n3231;
  assign n3234 = n2847 & n3223;
  assign n3233 = ~n3199 & n3231;
  assign n3235 = n3234 ^ n3233;
  assign n3237 = n3228 ^ n3194;
  assign n3238 = ~n2846 & n3237;
  assign n3236 = ~n2846 & n3196;
  assign n3239 = n3238 ^ n3236;
  assign n3240 = n3239 ^ n3195;
  assign n3254 = n3044 & n3188;
  assign n3251 = n3188 & ~n3215;
  assign n3242 = ~n3184 & n3227;
  assign n3249 = n3242 ^ n3227;
  assign n3243 = n3242 ^ n3197;
  assign n3241 = n3216 ^ n3190;
  assign n3244 = n3243 ^ n3241;
  assign n3250 = n3249 ^ n3244;
  assign n3252 = n3251 ^ n3250;
  assign n3253 = n3252 ^ n3197;
  assign n3255 = n3254 ^ n3253;
  assign n3245 = n3244 ^ n3242;
  assign n3246 = n3245 ^ n3205;
  assign n3247 = ~n2846 & n3246;
  assign n3248 = n3247 ^ n3245;
  assign n3256 = n3255 ^ n3248;
  assign n3257 = n3256 ^ n3255;
  assign n3258 = ~n3240 & ~n3257;
  assign n3259 = n3258 ^ n3255;
  assign n3260 = n3200 & ~n3259;
  assign n3261 = n3260 ^ n3255;
  assign n3262 = ~n3235 & ~n3261;
  assign n3263 = ~n3232 & n3262;
  assign n3264 = ~n3230 & n3263;
  assign n3265 = n3249 ^ n3209;
  assign n3266 = n2809 & ~n3265;
  assign n3267 = n3266 ^ n3209;
  assign n3268 = ~n2846 & ~n3267;
  assign n3269 = n3264 & ~n3268;
  assign n3270 = ~n3225 & n3269;
  assign n3271 = ~n3220 & n3270;
  assign n3272 = n3214 & n3271;
  assign n3273 = n3272 ^ n1403;
  assign n6076 = n3273 ^ x227;
  assign n1448 = n1406 & n1447;
  assign n1451 = n1450 ^ n1423;
  assign n1452 = n1451 ^ n1445;
  assign n1453 = ~n1409 & ~n1452;
  assign n1454 = ~n1448 & ~n1453;
  assign n1463 = ~n1405 & ~n1421;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = n1464 ^ n1443;
  assign n1466 = n1465 ^ n1443;
  assign n1467 = ~n1455 & n1466;
  assign n1468 = n1467 ^ n1443;
  assign n1469 = n1406 & ~n1468;
  assign n1470 = n1469 ^ n1443;
  assign n1471 = n1411 ^ n1208;
  assign n1472 = n1471 ^ n1420;
  assign n1473 = ~n1304 & n1472;
  assign n1474 = n1473 ^ n1420;
  assign n1475 = n1404 & n1474;
  assign n1476 = n1470 & ~n1475;
  assign n1477 = n1454 & n1476;
  assign n1478 = ~n1440 & n1477;
  assign n1479 = n1434 & n1478;
  assign n1480 = ~n1408 & n1479;
  assign n1481 = n1480 ^ x2;
  assign n1482 = n1481 ^ x184;
  assign n2637 = n2636 ^ n2632;
  assign n2638 = n2637 ^ n2627;
  assign n2639 = n2623 & n2638;
  assign n2640 = n2639 ^ n2637;
  assign n2641 = n2598 & ~n2640;
  assign n2661 = n2629 & ~n2653;
  assign n2663 = n2597 ^ n2579;
  assign n2664 = ~n2662 & ~n2663;
  assign n2667 = n2576 & ~n2624;
  assign n2668 = n2592 & ~n2667;
  assign n2665 = n2588 ^ n2574;
  assign n2666 = ~n2623 & n2665;
  assign n2669 = n2668 ^ n2666;
  assign n2670 = n2653 & n2669;
  assign n2671 = n2670 ^ n2668;
  assign n2672 = ~n2664 & ~n2671;
  assign n2673 = ~n2661 & n2672;
  assign n2674 = n2643 ^ n2636;
  assign n2675 = n2674 ^ n2584;
  assign n2676 = ~n2623 & n2675;
  assign n2677 = n2676 ^ n2584;
  assign n2678 = ~n2598 & n2677;
  assign n2679 = n2673 & ~n2678;
  assign n2680 = ~n2660 & n2679;
  assign n2681 = ~n2652 & n2680;
  assign n2682 = ~n2649 & n2681;
  assign n2683 = ~n2641 & n2682;
  assign n2684 = ~n2626 & n2683;
  assign n2685 = n2684 ^ x28;
  assign n2686 = n2685 ^ x189;
  assign n2687 = n1482 & n2686;
  assign n2272 = ~n2072 & n2221;
  assign n2273 = ~n2057 & n2235;
  assign n2274 = n2251 ^ n2220;
  assign n2275 = n2274 ^ n2230;
  assign n2276 = n2070 & ~n2275;
  assign n2277 = n2233 & ~n2263;
  assign n2279 = n2278 ^ n2277;
  assign n2280 = n2279 ^ n2215;
  assign n2281 = n2280 ^ n2263;
  assign n2282 = n2239 ^ n2071;
  assign n2283 = ~n2280 & n2282;
  assign n2284 = n2283 ^ n2071;
  assign n2285 = ~n2281 & ~n2284;
  assign n2286 = n2285 ^ n2263;
  assign n2287 = ~n2276 & n2286;
  assign n2288 = ~n2273 & n2287;
  assign n2290 = n2289 ^ n2231;
  assign n2291 = n2290 ^ n2245;
  assign n2292 = n2291 ^ n2221;
  assign n2293 = n2057 & ~n2292;
  assign n2294 = n2293 ^ n2221;
  assign n2295 = n2069 & n2294;
  assign n2296 = n2288 & ~n2295;
  assign n2297 = ~n2272 & n2296;
  assign n2298 = ~n2271 & n2297;
  assign n2299 = n2269 & n2298;
  assign n2300 = n2262 & n2299;
  assign n2301 = ~n2252 & n2300;
  assign n2302 = n2301 ^ x44;
  assign n2303 = n2302 ^ x187;
  assign n2005 = n2004 ^ n1969;
  assign n2030 = n2029 ^ n2005;
  assign n2031 = n2030 ^ n2026;
  assign n2032 = n2031 ^ x36;
  assign n2033 = n2032 ^ x188;
  assign n2411 = n2410 ^ n2304;
  assign n2438 = n2437 ^ n2435;
  assign n2439 = n2411 & n2438;
  assign n2441 = n2440 ^ n2439;
  assign n2444 = n2443 ^ n2416;
  assign n2445 = n2320 & n2444;
  assign n2453 = n2411 & n2427;
  assign n2459 = n2435 ^ n2420;
  assign n2457 = n2456 ^ n2404;
  assign n2458 = n2457 ^ n2436;
  assign n2460 = n2459 ^ n2458;
  assign n2461 = n2320 & n2460;
  assign n2462 = n2461 ^ n2459;
  assign n2463 = ~n2304 & n2462;
  assign n2464 = ~n2455 & ~n2463;
  assign n2465 = ~n2453 & n2464;
  assign n2466 = ~n2449 & n2465;
  assign n2472 = n2471 ^ n2436;
  assign n2473 = n2472 ^ n2468;
  assign n2474 = n2320 & n2473;
  assign n2475 = n2474 ^ n2468;
  assign n2476 = ~n2467 & n2475;
  assign n2477 = n2466 & ~n2476;
  assign n2478 = ~n2452 & n2477;
  assign n2479 = ~n2448 & n2478;
  assign n2480 = ~n2445 & n2479;
  assign n2481 = ~n2441 & n2480;
  assign n2482 = ~n2408 & n2481;
  assign n2483 = n2482 ^ x60;
  assign n2484 = n2483 ^ x185;
  assign n2698 = n2033 & ~n2484;
  assign n2723 = n2698 ^ n2033;
  assign n1798 = ~n1483 & ~n1797;
  assign n1792 = ~n1483 & ~n1791;
  assign n1793 = n1792 ^ n1749;
  assign n1799 = n1798 ^ n1793;
  assign n1800 = ~n1516 & n1799;
  assign n1801 = n1800 ^ n1793;
  assign n1804 = n1760 & ~n1790;
  assign n1808 = n1743 ^ n1616;
  assign n1809 = n1808 ^ n1765;
  assign n1810 = ~n1516 & ~n1809;
  assign n1805 = n1783 ^ n1778;
  assign n1806 = ~n1516 & ~n1805;
  assign n1807 = n1806 ^ n1778;
  assign n1811 = n1810 ^ n1807;
  assign n1812 = n1483 & n1811;
  assign n1813 = n1812 ^ n1807;
  assign n1818 = n1817 ^ n1814;
  assign n1819 = ~n1813 & ~n1818;
  assign n1820 = ~n1804 & n1819;
  assign n1822 = n1483 & n1821;
  assign n1823 = n1820 & ~n1822;
  assign n1824 = ~n1803 & n1823;
  assign n1825 = ~n1802 & n1824;
  assign n1826 = ~n1801 & n1825;
  assign n1827 = ~n1789 & n1826;
  assign n1828 = ~n1756 & n1827;
  assign n1829 = n1828 ^ x52;
  assign n1830 = n1829 ^ x186;
  assign n2691 = n1830 & n2033;
  assign n2692 = ~n2484 & n2691;
  assign n2718 = n2692 ^ n2691;
  assign n2724 = n2723 ^ n2718;
  assign n2732 = n2303 & n2724;
  assign n5138 = n2687 & n2732;
  assign n2699 = n2698 ^ n2692;
  assign n2696 = n2033 ^ n1830;
  assign n2697 = ~n2484 & n2696;
  assign n2700 = n2699 ^ n2697;
  assign n2485 = n2303 & ~n2484;
  assign n2486 = n2033 & n2485;
  assign n2487 = n2486 ^ n2485;
  assign n2488 = n1830 & n2487;
  assign n2701 = n2700 ^ n2488;
  assign n2709 = n2687 ^ n2686;
  assign n2710 = n2701 & n2709;
  assign n5139 = n5138 ^ n2710;
  assign n2702 = ~n2033 & ~n2303;
  assign n2703 = n2484 & n2702;
  assign n2704 = n2703 ^ n2702;
  assign n2705 = n2704 ^ n2701;
  assign n5144 = n2705 ^ n2488;
  assign n6078 = n2709 & n5144;
  assign n2733 = n2732 ^ n2724;
  assign n2720 = ~n1830 & n2484;
  assign n2721 = n2702 & n2720;
  assign n2730 = n2721 ^ n2703;
  assign n2734 = n2733 ^ n2730;
  assign n2693 = n2692 ^ n2486;
  assign n2690 = ~n1830 & n2486;
  assign n2694 = n2693 ^ n2690;
  assign n6079 = n2734 ^ n2694;
  assign n6080 = n2687 & n6079;
  assign n2759 = n2732 ^ n2488;
  assign n2760 = n2759 ^ n2694;
  assign n6087 = n2760 ^ n2690;
  assign n6088 = n6087 ^ n2734;
  assign n2751 = n2730 ^ n2484;
  assign n2725 = n2724 ^ n2720;
  assign n2726 = n2725 ^ n2721;
  assign n2735 = n2734 ^ n2726;
  assign n2736 = n2735 ^ n2732;
  assign n2719 = n2303 & n2718;
  assign n2728 = n2719 ^ n2718;
  assign n2722 = n2721 ^ n2719;
  assign n2729 = n2728 ^ n2722;
  assign n2731 = n2730 ^ n2729;
  assign n2737 = n2736 ^ n2731;
  assign n2752 = n2751 ^ n2737;
  assign n2753 = n2752 ^ n2728;
  assign n4998 = n2753 ^ n2726;
  assign n4999 = n4998 ^ n2732;
  assign n6089 = n6088 ^ n4999;
  assign n6090 = ~n2686 & n6089;
  assign n6091 = n6090 ^ n4999;
  assign n2695 = n2694 ^ n2692;
  assign n2706 = n2705 ^ n2695;
  assign n6082 = n2706 ^ n2488;
  assign n6083 = n6082 ^ n2690;
  assign n6081 = n2728 ^ n2726;
  assign n6084 = n6083 ^ n6081;
  assign n6085 = n2686 & n6084;
  assign n6086 = n6085 ^ n6081;
  assign n6092 = n6091 ^ n6086;
  assign n6093 = ~n1482 & n6092;
  assign n6094 = n6093 ^ n6086;
  assign n6095 = ~n2686 & n2722;
  assign n6096 = ~n6094 & ~n6095;
  assign n6097 = ~n6080 & n6096;
  assign n6098 = ~n6078 & n6097;
  assign n5008 = n2699 ^ n2690;
  assign n2688 = n2687 ^ n1482;
  assign n6099 = n5008 ^ n2688;
  assign n2712 = n2488 ^ n2487;
  assign n5004 = n2712 ^ n2695;
  assign n6100 = n5004 ^ n2701;
  assign n6101 = n6100 ^ n2709;
  assign n6102 = ~n5008 & ~n6101;
  assign n6103 = n6102 ^ n2709;
  assign n6104 = n6099 & n6103;
  assign n6105 = n6104 ^ n2688;
  assign n6106 = n6098 & ~n6105;
  assign n6107 = ~n5139 & n6106;
  assign n6108 = n6107 ^ n1900;
  assign n6109 = n6108 ^ x228;
  assign n6122 = n6076 & n6109;
  assign n6123 = n6122 ^ n6109;
  assign n6124 = n6123 ^ n6076;
  assign n4312 = n3827 ^ x202;
  assign n4311 = n3306 ^ x207;
  assign n4313 = n4312 ^ n4311;
  assign n3550 = ~n2320 & n2404;
  assign n3546 = n2787 ^ n2435;
  assign n3547 = n3546 ^ n2416;
  assign n3548 = n2320 & n3547;
  assign n3549 = n3548 ^ n2416;
  assign n3551 = n3550 ^ n3549;
  assign n3552 = ~n2467 & n3551;
  assign n3553 = n3552 ^ n3549;
  assign n4345 = n2432 ^ n2414;
  assign n4346 = n2409 & n4345;
  assign n4347 = n2470 ^ n2416;
  assign n4348 = ~n2454 & n4347;
  assign n4352 = ~n2320 & n2423;
  assign n3560 = n2469 ^ n2429;
  assign n4349 = n3560 ^ n2426;
  assign n4350 = n2320 & n4349;
  assign n4351 = n4350 ^ n3560;
  assign n4353 = n4352 ^ n4351;
  assign n4354 = ~n2304 & n4353;
  assign n4355 = n4354 ^ n4351;
  assign n4356 = ~n2455 & ~n4355;
  assign n4357 = ~n4348 & n4356;
  assign n4358 = ~n4346 & n4357;
  assign n4359 = ~n3553 & n4358;
  assign n4360 = ~n2784 & n4359;
  assign n4361 = ~n2782 & n4360;
  assign n4362 = ~n2441 & n4361;
  assign n4363 = ~n2779 & n4362;
  assign n4364 = n4363 ^ x14;
  assign n4365 = n4364 ^ x205;
  assign n4366 = n3760 ^ x203;
  assign n4373 = n4365 & ~n4366;
  assign n4412 = n4373 ^ n4366;
  assign n4437 = n4412 ^ n4365;
  assign n4314 = n1432 ^ n1418;
  assign n4315 = n4314 ^ n1435;
  assign n4316 = n4315 ^ n1424;
  assign n4317 = ~n1304 & ~n4316;
  assign n4318 = n4317 ^ n1424;
  assign n4319 = ~n1404 & ~n4318;
  assign n4320 = n3024 ^ n1447;
  assign n4321 = n3024 ^ n1304;
  assign n4322 = ~n1409 & n4321;
  assign n4323 = n4322 ^ n1304;
  assign n4324 = n4320 & ~n4323;
  assign n4325 = n4324 ^ n1447;
  assign n4326 = ~n1411 & ~n4325;
  assign n4327 = ~n1203 & n4326;
  assign n4328 = n4327 ^ n1206;
  assign n4329 = n4328 ^ n1206;
  assign n4330 = n1406 & ~n4329;
  assign n4331 = n4330 ^ n1206;
  assign n4332 = ~n1455 & n4331;
  assign n4333 = n4332 ^ n1206;
  assign n4334 = ~n4319 & ~n4333;
  assign n4335 = ~n1304 & ~n1441;
  assign n4336 = n4335 ^ n3014;
  assign n4337 = n1409 & n4336;
  assign n4338 = n4337 ^ n3014;
  assign n4339 = n4334 & ~n4338;
  assign n4340 = n3013 & n4339;
  assign n4341 = ~n1408 & n4340;
  assign n4342 = n1443 & n4341;
  assign n4343 = n4342 ^ x22;
  assign n4344 = n4343 ^ x204;
  assign n4370 = n3436 ^ x206;
  assign n4374 = ~n4344 & n4370;
  assign n4375 = n4374 ^ n4370;
  assign n4379 = n4373 ^ n4365;
  assign n4383 = n4375 & n4379;
  assign n4421 = n4383 ^ n4375;
  assign n4401 = ~n4366 & n4375;
  assign n4422 = n4421 ^ n4401;
  assign n4417 = n4366 ^ n4344;
  assign n4389 = n4366 & n4374;
  assign n4385 = n4374 & n4379;
  assign n4390 = n4389 ^ n4385;
  assign n4418 = n4417 ^ n4390;
  assign n4367 = n4366 ^ n4365;
  assign n4368 = n4344 & ~n4367;
  assign n4369 = n4368 ^ n4366;
  assign n4409 = n4373 ^ n4369;
  assign n4392 = n4385 ^ n4374;
  assign n4388 = n4373 & n4374;
  assign n4391 = n4390 ^ n4388;
  assign n4393 = n4392 ^ n4391;
  assign n4386 = n4385 ^ n4379;
  assign n4380 = n4375 ^ n4344;
  assign n4381 = n4380 ^ n4370;
  assign n4382 = n4379 & ~n4381;
  assign n4384 = n4383 ^ n4382;
  assign n4387 = n4386 ^ n4384;
  assign n4394 = n4393 ^ n4387;
  assign n4408 = n4394 ^ n4383;
  assign n4410 = n4409 ^ n4408;
  assign n4376 = n4373 & n4375;
  assign n4402 = n4401 ^ n4376;
  assign n4411 = n4410 ^ n4402;
  assign n4413 = n4412 ^ n4411;
  assign n4414 = n4413 ^ n4393;
  assign n4415 = n4414 ^ n4385;
  assign n4416 = n4415 ^ n4376;
  assign n4419 = n4418 ^ n4416;
  assign n4377 = n4376 ^ n4373;
  assign n4371 = n4370 ^ n4344;
  assign n4372 = ~n4369 & n4371;
  assign n4378 = n4377 ^ n4372;
  assign n4395 = n4394 ^ n4378;
  assign n4396 = n4395 ^ n4388;
  assign n4404 = n4396 ^ n4377;
  assign n4400 = n4393 ^ n4384;
  assign n4403 = n4402 ^ n4400;
  assign n4405 = n4404 ^ n4403;
  assign n4406 = n4405 ^ n4382;
  assign n4407 = n4406 ^ n4400;
  assign n4420 = n4419 ^ n4407;
  assign n4423 = n4422 ^ n4420;
  assign n4429 = n4423 ^ n4390;
  assign n4438 = n4437 ^ n4429;
  assign n5271 = n4438 ^ n4423;
  assign n5272 = n4311 & n5271;
  assign n5273 = n5272 ^ n4423;
  assign n5274 = ~n4313 & n5273;
  assign n5020 = n4422 ^ n4387;
  assign n5021 = n5020 ^ n4404;
  assign n5022 = n4312 & n5021;
  assign n5023 = n5022 ^ n4404;
  assign n5024 = n4311 & n5023;
  assign n4425 = ~n4311 & n4312;
  assign n4426 = n4425 ^ n4311;
  assign n4441 = n4390 & ~n4426;
  assign n6050 = n4367 ^ n4344;
  assign n6051 = n6050 ^ n4389;
  assign n6052 = n4425 & n6051;
  assign n6057 = n4429 ^ n4383;
  assign n6054 = n4401 ^ n4366;
  assign n6055 = n4311 & ~n6054;
  assign n5028 = n4388 ^ n4376;
  assign n5029 = n5028 ^ n4414;
  assign n6053 = n5029 ^ n4404;
  assign n6056 = n6055 ^ n6053;
  assign n6058 = n6057 ^ n6056;
  assign n6059 = n6058 ^ n6056;
  assign n6060 = n4311 & n6059;
  assign n6061 = n6060 ^ n6056;
  assign n6062 = n4313 & n6061;
  assign n6063 = n6062 ^ n6056;
  assign n6064 = ~n6052 & ~n6063;
  assign n6065 = ~n4441 & n6064;
  assign n5030 = n5029 ^ n4311;
  assign n5031 = ~n4311 & ~n5030;
  assign n5032 = n5031 ^ n4311;
  assign n6066 = n5032 ^ n5029;
  assign n6067 = n6066 ^ n4382;
  assign n6068 = n4313 & ~n6067;
  assign n6069 = n6068 ^ n4382;
  assign n6070 = n6065 & ~n6069;
  assign n6071 = ~n5024 & n6070;
  assign n6072 = ~n5274 & n6071;
  assign n6073 = n6072 ^ n1936;
  assign n6074 = n6073 ^ x229;
  assign n3938 = n1759 & n3352;
  assign n3951 = n1757 & ~n1780;
  assign n3948 = n1780 ^ n1774;
  assign n3949 = ~n1516 & ~n3948;
  assign n3950 = n3949 ^ n1774;
  assign n3952 = n3951 ^ n3950;
  assign n3945 = n1777 ^ n1753;
  assign n3946 = n1757 & ~n3945;
  assign n3947 = n3946 ^ n3356;
  assign n3953 = n3952 ^ n3947;
  assign n3943 = n3802 ^ n3360;
  assign n3941 = ~n1768 & n3803;
  assign n3939 = n1774 ^ n1768;
  assign n3940 = n1483 & n3939;
  assign n3942 = n3941 ^ n3940;
  assign n3944 = n3943 ^ n3942;
  assign n3954 = n3953 ^ n3944;
  assign n3955 = ~n3938 & ~n3954;
  assign n3956 = n1516 & ~n1796;
  assign n3957 = n3956 ^ n1815;
  assign n3958 = ~n1483 & n1772;
  assign n3959 = n3958 ^ n1752;
  assign n3960 = ~n3957 & ~n3959;
  assign n3961 = n3960 ^ n3956;
  assign n3962 = ~n1761 & ~n3961;
  assign n3963 = n3962 ^ n3956;
  assign n3964 = n3955 & ~n3963;
  assign n3965 = ~n1801 & n3964;
  assign n3966 = n3965 ^ x26;
  assign n4184 = n3966 ^ x177;
  assign n4185 = n3183 ^ x172;
  assign n4186 = n4184 & n4185;
  assign n4187 = n4186 ^ n4184;
  assign n4188 = n4187 ^ n4185;
  assign n4189 = n4188 ^ n4186;
  assign n4220 = n2808 ^ x173;
  assign n4221 = n3304 ^ n3302;
  assign n4222 = n4221 ^ x50;
  assign n4223 = n4222 ^ x174;
  assign n4224 = ~n4220 & n4223;
  assign n3578 = ~n2882 & ~n2976;
  assign n3579 = n3578 ^ n2972;
  assign n3580 = ~n2967 & ~n3579;
  assign n3927 = n3427 ^ n2937;
  assign n3928 = ~n2882 & n3927;
  assign n3929 = n3928 ^ n2937;
  assign n3922 = n3412 ^ n2945;
  assign n3923 = n3922 ^ n2955;
  assign n3920 = n2991 ^ n2931;
  assign n3919 = n2974 ^ n2945;
  assign n3921 = n3920 ^ n3919;
  assign n3924 = n3923 ^ n3921;
  assign n3925 = ~n2882 & n3924;
  assign n3926 = n3925 ^ n3921;
  assign n3930 = n3929 ^ n3926;
  assign n3931 = ~n2883 & ~n3930;
  assign n3932 = n3931 ^ n3929;
  assign n3933 = ~n2959 & ~n3932;
  assign n3934 = ~n3580 & n3933;
  assign n3935 = n3404 & n3934;
  assign n3936 = n3935 ^ x34;
  assign n4190 = n3936 ^ x176;
  assign n4191 = ~n2069 & n2233;
  assign n4202 = ~n2069 & n2231;
  assign n4200 = ~n2228 & ~n2263;
  assign n4199 = ~n2072 & n2233;
  assign n4201 = n4200 ^ n4199;
  assign n4203 = n4202 ^ n4201;
  assign n4196 = n2816 ^ n2815;
  assign n4197 = n4196 ^ n2817;
  assign n4198 = n4197 ^ n2235;
  assign n4204 = n4203 ^ n4198;
  assign n4194 = ~n2071 & n2238;
  assign n4192 = n2229 ^ n2215;
  assign n4193 = ~n2057 & n4192;
  assign n4195 = n4194 ^ n4193;
  assign n4205 = n4204 ^ n4195;
  assign n4206 = ~n3723 & n4205;
  assign n4207 = ~n2252 & n4206;
  assign n4208 = n2218 & n2254;
  assign n4209 = n4207 & ~n4208;
  assign n4210 = ~n4191 & n4209;
  assign n4211 = n2069 & n2232;
  assign n4212 = n4211 ^ n2221;
  assign n4213 = n2057 & n4212;
  assign n4214 = n4210 & ~n4213;
  assign n4215 = ~n3728 & n4214;
  assign n4216 = ~n2812 & n4215;
  assign n4217 = n4216 ^ x42;
  assign n4218 = n4217 ^ x175;
  assign n4219 = ~n4190 & ~n4218;
  assign n4227 = n4219 ^ n4218;
  assign n4228 = n4224 & ~n4227;
  assign n4225 = n4224 ^ n4220;
  assign n4226 = n4219 & ~n4225;
  assign n4229 = n4228 ^ n4226;
  assign n4230 = ~n4184 & n4229;
  assign n4231 = n4230 ^ n4226;
  assign n4232 = n4189 & n4231;
  assign n4237 = n4184 & n4228;
  assign n4235 = n4219 & n4224;
  assign n4233 = n4226 ^ n4219;
  assign n4234 = n4184 & n4233;
  assign n4236 = n4235 ^ n4234;
  assign n4238 = n4237 ^ n4236;
  assign n4239 = ~n4185 & n4238;
  assign n4240 = n4239 ^ n4236;
  assign n4259 = n4235 ^ n4224;
  assign n4242 = n4219 ^ n4190;
  assign n4257 = n4224 & ~n4242;
  assign n4258 = n4257 ^ n4228;
  assign n4260 = n4259 ^ n4258;
  assign n4251 = n4228 ^ n4227;
  assign n4245 = n4225 ^ n4223;
  assign n4246 = n4245 ^ n4220;
  assign n4247 = n4219 & n4246;
  assign n4252 = n4251 ^ n4247;
  assign n4248 = n4247 ^ n4235;
  assign n4249 = n4248 ^ n4233;
  assign n4244 = ~n4218 & n4220;
  assign n4250 = n4249 ^ n4244;
  assign n4253 = n4252 ^ n4250;
  assign n4243 = ~n4225 & ~n4242;
  assign n4254 = n4253 ^ n4243;
  assign n4241 = n4226 ^ n4225;
  assign n4255 = n4254 ^ n4241;
  assign n4256 = n4255 ^ n4226;
  assign n4261 = n4260 ^ n4256;
  assign n4262 = n4261 ^ n4243;
  assign n4263 = ~n4188 & n4262;
  assign n4265 = n4227 ^ n4190;
  assign n4266 = n4246 & ~n4265;
  assign n4267 = n4266 ^ n4265;
  assign n4264 = n4260 ^ n4255;
  assign n4268 = n4267 ^ n4264;
  assign n4269 = n4268 ^ n4266;
  assign n4270 = n4269 ^ n4249;
  assign n4271 = n4186 ^ n4185;
  assign n4272 = ~n4270 & n4271;
  assign n4291 = n4266 ^ n4255;
  assign n4292 = n4291 ^ n4223;
  assign n4273 = n4223 ^ n4218;
  assign n4274 = n4190 & ~n4273;
  assign n4275 = n4274 ^ n4223;
  assign n4276 = n4220 & n4275;
  assign n4277 = n4276 ^ n4220;
  assign n4278 = n4277 ^ n4270;
  assign n4279 = n4278 ^ n4266;
  assign n4280 = n4279 ^ n4245;
  assign n4281 = n4280 ^ n4270;
  assign n4282 = n4281 ^ n4253;
  assign n4283 = n4282 ^ n4251;
  assign n4284 = n4283 ^ n4249;
  assign n4285 = n4284 ^ n4269;
  assign n4286 = n4285 ^ n4282;
  assign n4293 = n4292 ^ n4286;
  assign n4289 = n4220 ^ n4190;
  assign n4290 = n4289 ^ n4218;
  assign n4294 = n4293 ^ n4290;
  assign n4295 = n4294 ^ n4276;
  assign n4296 = n4184 & n4295;
  assign n4297 = n4296 ^ n4276;
  assign n4287 = n4184 & n4286;
  assign n4288 = n4287 ^ n4282;
  assign n4298 = n4297 ^ n4288;
  assign n4299 = n4189 & ~n4298;
  assign n4300 = n4299 ^ n4297;
  assign n4301 = ~n4272 & ~n4300;
  assign n4302 = ~n4263 & n4301;
  assign n4304 = n4189 & n4257;
  assign n4303 = n4187 & ~n4278;
  assign n4305 = n4304 ^ n4303;
  assign n4306 = n4302 & ~n4305;
  assign n4307 = ~n4240 & n4306;
  assign n4308 = ~n4232 & n4307;
  assign n4309 = n4308 ^ n1868;
  assign n6049 = n4309 ^ x230;
  assign n6119 = n6074 ^ n6049;
  assign n6075 = n6049 & ~n6074;
  assign n6137 = n6119 ^ n6075;
  assign n6155 = ~n6124 & n6137;
  assign n6636 = n6047 & n6155;
  assign n6166 = n6137 ^ n6049;
  assign n6169 = n6046 & ~n6076;
  assign n6170 = ~n6166 & n6169;
  assign n6637 = n6636 ^ n6170;
  assign n6173 = n6045 ^ n6044;
  assign n6121 = ~n6049 & ~n6076;
  assign n6125 = n6124 ^ n6121;
  assign n6110 = n6109 ^ n6049;
  assign n6111 = ~n6109 & ~n6110;
  assign n6112 = n6111 ^ n6109;
  assign n6120 = n6112 ^ n6049;
  assign n6126 = n6125 ^ n6120;
  assign n6127 = ~n6119 & n6126;
  assign n6128 = n6127 ^ n6125;
  assign n6153 = ~n6076 & ~n6128;
  assign n6146 = n6076 & n6137;
  assign n6152 = n6146 ^ n6122;
  assign n6154 = n6153 ^ n6152;
  assign n6147 = n6146 ^ n6075;
  assign n6148 = n6147 ^ n6124;
  assign n6731 = n6154 ^ n6148;
  assign n6732 = n6045 & ~n6731;
  assign n6733 = n6732 ^ n6148;
  assign n6113 = n6109 ^ n6074;
  assign n6114 = ~n6112 & ~n6113;
  assign n6115 = n6114 ^ n6111;
  assign n6116 = n6115 ^ n6109;
  assign n6117 = n6116 ^ n6049;
  assign n6077 = n6075 & n6076;
  assign n6118 = n6117 ^ n6077;
  assign n6129 = n6128 ^ n6118;
  assign n6130 = n6129 ^ n6114;
  assign n6158 = n6153 ^ n6130;
  assign n6159 = n6158 ^ n6049;
  assign n6156 = n6155 ^ n6154;
  assign n6150 = n6146 ^ n6077;
  assign n6151 = n6150 ^ n6125;
  assign n6157 = n6156 ^ n6151;
  assign n6160 = n6159 ^ n6157;
  assign n6145 = n6125 ^ n6049;
  assign n6149 = n6148 ^ n6145;
  assign n6161 = n6160 ^ n6149;
  assign n6142 = n6124 ^ n6114;
  assign n6138 = n6137 ^ n6076;
  assign n6139 = n6138 ^ n6109;
  assign n6140 = n6139 ^ n6119;
  assign n6134 = n6122 ^ n6120;
  assign n6135 = n6134 ^ n6049;
  assign n6136 = n6074 & ~n6135;
  assign n6141 = n6140 ^ n6136;
  assign n6143 = n6142 ^ n6141;
  assign n6133 = n6109 ^ n6076;
  assign n6144 = n6143 ^ n6133;
  assign n6162 = n6161 ^ n6144;
  assign n6174 = n6045 & n6162;
  assign n6175 = n6174 ^ n6144;
  assign n6734 = n6733 ^ n6175;
  assign n6735 = ~n6173 & ~n6734;
  assign n6736 = n6735 ^ n6733;
  assign n6737 = ~n6637 & n6736;
  assign n6738 = n6737 ^ n2032;
  assign n7189 = n6738 ^ x284;
  assign n4979 = n2701 ^ n2694;
  assign n4980 = n4979 ^ n2721;
  assign n4981 = n4980 ^ n2721;
  assign n4982 = n2686 & n4981;
  assign n4983 = n4982 ^ n2721;
  assign n4984 = n1482 & n4983;
  assign n4985 = n4984 ^ n2721;
  assign n4986 = n1482 & n2706;
  assign n4987 = n4986 ^ n2726;
  assign n4988 = n2686 & n4987;
  assign n4989 = n4988 ^ n2726;
  assign n4991 = ~n1482 & n2733;
  assign n4990 = n2709 & n2753;
  assign n4992 = n4991 ^ n4990;
  assign n4993 = ~n4989 & ~n4992;
  assign n2689 = n2688 ^ n2686;
  assign n4994 = ~n2689 & n2728;
  assign n4995 = n2752 ^ n2719;
  assign n4996 = n4995 ^ n2730;
  assign n4997 = n2688 & n4996;
  assign n2750 = n2709 ^ n2688;
  assign n5000 = n4999 ^ n2697;
  assign n5001 = n2686 & n5000;
  assign n5002 = n5001 ^ n2697;
  assign n5003 = ~n2750 & n5002;
  assign n5009 = n5008 ^ n5004;
  assign n5010 = n2750 & n5009;
  assign n5005 = n5004 ^ n2732;
  assign n2713 = n2712 ^ n2705;
  assign n2714 = n2713 ^ n2710;
  assign n5006 = n5005 ^ n2714;
  assign n5007 = n2688 & n5006;
  assign n5011 = n5010 ^ n5007;
  assign n5012 = n5011 ^ n2710;
  assign n5013 = ~n5003 & ~n5012;
  assign n5014 = ~n4997 & n5013;
  assign n5015 = ~n4994 & n5014;
  assign n5016 = n4993 & n5015;
  assign n5017 = ~n4985 & n5016;
  assign n5018 = n5017 ^ n2056;
  assign n5353 = n5018 ^ x243;
  assign n3918 = n2483 ^ x183;
  assign n3937 = n3936 ^ x178;
  assign n3997 = n1481 ^ x182;
  assign n3967 = n3966 ^ x179;
  assign n3968 = n2581 & ~n2623;
  assign n3969 = n2585 & ~n2662;
  assign n3970 = n2579 & ~n2598;
  assign n3972 = n2628 ^ n2590;
  assign n3971 = n2637 ^ n2583;
  assign n3973 = n3972 ^ n3971;
  assign n3974 = ~n2625 & ~n3973;
  assign n3975 = ~n3970 & ~n3974;
  assign n3979 = n2656 ^ n2629;
  assign n3980 = ~n2624 & n3979;
  assign n3981 = n2655 ^ n2643;
  assign n3982 = n3981 ^ n2855;
  assign n3983 = ~n3980 & n3982;
  assign n3984 = ~n2574 & ~n3983;
  assign n3976 = n2591 ^ n2579;
  assign n3977 = n3976 ^ n2634;
  assign n3978 = ~n2623 & n3977;
  assign n3985 = n3984 ^ n3978;
  assign n3986 = n2653 & ~n3985;
  assign n3987 = n3986 ^ n3984;
  assign n3988 = n3975 & n3987;
  assign n3989 = ~n3969 & n3988;
  assign n3990 = ~n3968 & n3989;
  assign n3991 = ~n2641 & n3990;
  assign n3992 = ~n2858 & n3991;
  assign n3993 = ~n2626 & n3992;
  assign n3994 = n3993 ^ x10;
  assign n3995 = n3994 ^ x181;
  assign n3996 = ~n3967 & n3995;
  assign n4022 = n3996 ^ n3967;
  assign n4023 = ~n3997 & ~n4022;
  assign n4059 = n4023 ^ n3996;
  assign n4026 = n3996 ^ n3995;
  assign n4032 = n4026 ^ n3967;
  assign n4048 = n4032 ^ n3997;
  assign n4060 = n4059 ^ n4048;
  assign n4040 = ~n3997 & n4026;
  assign n4061 = n4060 ^ n4040;
  assign n3998 = n3118 ^ n3109;
  assign n3999 = ~n3339 & n3998;
  assign n4000 = ~n3095 & n3324;
  assign n4001 = n3121 & ~n3322;
  assign n4002 = n4001 ^ n3142;
  assign n4003 = ~n4000 & ~n4002;
  assign n4004 = ~n3999 & ~n4003;
  assign n4006 = n3125 & n3141;
  assign n4005 = ~n3046 & n3111;
  assign n4007 = n4006 ^ n4005;
  assign n4008 = n4004 & ~n4007;
  assign n4009 = n3530 ^ n3128;
  assign n4010 = ~n3129 & n4009;
  assign n4011 = n4010 ^ n3128;
  assign n4012 = n3046 & n4011;
  assign n4013 = n4008 & ~n4012;
  assign n4014 = ~n3518 & n4013;
  assign n4015 = ~n3132 & n4014;
  assign n4016 = n4015 ^ x18;
  assign n4017 = n4016 ^ x180;
  assign n4031 = n4017 ^ n3967;
  assign n4033 = ~n3997 & n4032;
  assign n4034 = n4033 ^ n3997;
  assign n4035 = ~n4031 & ~n4034;
  assign n4055 = n4035 ^ n3997;
  assign n4056 = n4055 ^ n4040;
  assign n4018 = ~n3997 & ~n4017;
  assign n4019 = n4018 ^ n4017;
  assign n4052 = n3996 & ~n4019;
  assign n4049 = n4048 ^ n3996;
  assign n4045 = ~n3967 & n4018;
  assign n4020 = n4019 ^ n3997;
  assign n4044 = ~n4020 & ~n4022;
  assign n4046 = n4045 ^ n4044;
  assign n4041 = n4040 ^ n3996;
  assign n4039 = n4033 ^ n3995;
  assign n4042 = n4041 ^ n4039;
  assign n4043 = n4017 & n4042;
  assign n4047 = n4046 ^ n4043;
  assign n4050 = n4049 ^ n4047;
  assign n4051 = n4050 ^ n4043;
  assign n4053 = n4052 ^ n4051;
  assign n4036 = n4035 ^ n4033;
  assign n4024 = n4017 ^ n3997;
  assign n4025 = ~n3995 & ~n4017;
  assign n4027 = n4026 ^ n4025;
  assign n4028 = ~n4024 & n4027;
  assign n4029 = n4028 ^ n4026;
  assign n4030 = ~n4023 & ~n4029;
  assign n4037 = n4036 ^ n4030;
  assign n4038 = n4037 ^ n4031;
  assign n4054 = n4053 ^ n4038;
  assign n4057 = n4056 ^ n4054;
  assign n4021 = n3996 & ~n4020;
  assign n4058 = n4057 ^ n4021;
  assign n4062 = n4061 ^ n4058;
  assign n4063 = n4062 ^ n4057;
  assign n4064 = n3937 & ~n4063;
  assign n4065 = n4064 ^ n4057;
  assign n4066 = n3918 & ~n4065;
  assign n4549 = ~n3937 & n4049;
  assign n4082 = n4045 ^ n3997;
  assign n4083 = n4082 ^ n4056;
  assign n4084 = n4083 ^ n4044;
  assign n4085 = n4084 ^ n4021;
  assign n4086 = ~n3937 & n4085;
  assign n4087 = n4086 ^ n4021;
  assign n4548 = n4087 ^ n4047;
  assign n4550 = n4549 ^ n4548;
  assign n4546 = n3937 & ~n4054;
  assign n4547 = n4546 ^ n4038;
  assign n4551 = n4550 ^ n4547;
  assign n4552 = n3918 & n4551;
  assign n4553 = n4552 ^ n4547;
  assign n4554 = ~n4066 & ~n4553;
  assign n4555 = n4554 ^ n2068;
  assign n5354 = n4555 ^ x238;
  assign n4397 = n4311 & n4396;
  assign n4398 = n4397 ^ n4388;
  assign n4399 = ~n4313 & n4398;
  assign n4424 = n4423 ^ n4387;
  assign n4427 = n4426 ^ n4312;
  assign n4428 = n4424 & n4427;
  assign n4430 = n4311 & n4429;
  assign n4431 = n4430 ^ n4423;
  assign n4432 = n4312 & n4431;
  assign n4433 = ~n4311 & ~n4411;
  assign n4434 = n4433 ^ n4404;
  assign n4435 = n4313 & n4434;
  assign n4436 = n4435 ^ n4404;
  assign n4443 = n4312 & n4416;
  assign n4440 = n4400 & ~n4426;
  assign n4442 = n4441 ^ n4440;
  assign n4444 = n4443 ^ n4442;
  assign n4446 = ~n4312 & n4406;
  assign n4447 = n4446 ^ n4382;
  assign n4448 = ~n4444 & ~n4447;
  assign n4439 = n4438 ^ n4410;
  assign n4445 = n4444 ^ n4439;
  assign n4449 = n4448 ^ n4445;
  assign n4450 = n4313 & n4449;
  assign n4451 = n4450 ^ n4445;
  assign n4452 = ~n4436 & n4451;
  assign n4453 = ~n4432 & n4452;
  assign n4454 = ~n4428 & n4453;
  assign n4455 = ~n4399 & n4454;
  assign n4456 = n4455 ^ n2100;
  assign n5424 = n4456 ^ x239;
  assign n4734 = n4276 ^ n4250;
  assign n4735 = n4734 ^ n4268;
  assign n4927 = ~n4184 & ~n4735;
  assign n4928 = n4927 ^ n4281;
  assign n4929 = ~n4189 & n4928;
  assign n4930 = n4929 ^ n4281;
  assign n4931 = n4186 & n4257;
  assign n4731 = n4184 & ~n4279;
  assign n4732 = n4731 ^ n4278;
  assign n4733 = n4189 & ~n4732;
  assign n4932 = n4931 ^ n4733;
  assign n4933 = ~n4188 & n4284;
  assign n4934 = n4266 & n4271;
  assign n4935 = n4186 & n4261;
  assign n4945 = n4284 ^ n4278;
  assign n4944 = n4256 ^ n4228;
  assign n4946 = n4945 ^ n4944;
  assign n4947 = n4189 & ~n4945;
  assign n4948 = n4947 ^ n4188;
  assign n4949 = ~n4946 & n4948;
  assign n4950 = n4949 ^ n4944;
  assign n4951 = ~n4235 & ~n4950;
  assign n4738 = n4258 ^ n4254;
  assign n4936 = n4738 ^ n4264;
  assign n4937 = ~n4187 & ~n4258;
  assign n4938 = n4937 ^ n4271;
  assign n4939 = ~n4738 & n4938;
  assign n4940 = n4939 ^ n4271;
  assign n4941 = ~n4936 & ~n4940;
  assign n4942 = n4941 ^ n4264;
  assign n4943 = ~n4247 & ~n4942;
  assign n4952 = n4951 ^ n4943;
  assign n4953 = ~n4189 & n4952;
  assign n4954 = n4953 ^ n4943;
  assign n4955 = ~n4935 & n4954;
  assign n4956 = ~n4303 & n4955;
  assign n4957 = ~n4934 & n4956;
  assign n4958 = ~n4933 & n4957;
  assign n4959 = ~n4932 & n4958;
  assign n4960 = ~n4930 & n4959;
  assign n4961 = n4960 ^ n2211;
  assign n5425 = n4961 ^ x242;
  assign n5426 = n5424 & n5425;
  assign n5355 = n3884 ^ n3761;
  assign n5356 = n3896 & n5355;
  assign n5357 = n3858 ^ n3854;
  assign n5358 = n3762 & n5357;
  assign n5359 = n3882 ^ n3761;
  assign n5360 = n3894 ^ n3866;
  assign n5361 = n5359 & n5360;
  assign n5368 = n3800 ^ n3764;
  assign n5369 = n3798 & n3828;
  assign n5370 = n5369 ^ n3797;
  assign n5371 = ~n5368 & ~n5370;
  assign n5372 = n5371 ^ n3869;
  assign n5373 = ~n3762 & ~n5372;
  assign n5374 = n5373 ^ n5371;
  assign n5362 = ~n3853 & ~n5355;
  assign n5365 = n3874 ^ n3865;
  assign n5363 = ~n3860 & n5359;
  assign n5364 = n5363 ^ n3851;
  assign n5366 = n5365 ^ n5364;
  assign n5367 = ~n5362 & ~n5366;
  assign n5375 = n5374 ^ n5367;
  assign n5376 = ~n3883 & n5375;
  assign n5377 = n5376 ^ n5367;
  assign n5378 = ~n5361 & ~n5377;
  assign n5379 = ~n3881 & n5378;
  assign n5380 = ~n5358 & n5379;
  assign n5381 = ~n5356 & n5380;
  assign n5382 = ~n3891 & n5381;
  assign n5383 = ~n3885 & n5382;
  assign n5384 = n5383 ^ n2168;
  assign n5385 = n5384 ^ x240;
  assign n3469 = n3468 ^ n3455;
  assign n3470 = n3438 & n3469;
  assign n3471 = n3470 ^ n3455;
  assign n3472 = n3466 & n3471;
  assign n4763 = n3492 ^ n3450;
  assign n4764 = n3439 & n4763;
  assign n5386 = n3492 ^ n3453;
  assign n5387 = ~n3466 & n5386;
  assign n5388 = n3477 ^ n3437;
  assign n5390 = n4528 ^ n3489;
  assign n5389 = n3480 ^ n3452;
  assign n5391 = n5390 ^ n5389;
  assign n5392 = ~n3438 & n5391;
  assign n5393 = n5392 ^ n5389;
  assign n5394 = n5393 ^ n3477;
  assign n5395 = n5388 & ~n5394;
  assign n5396 = n5395 ^ n5392;
  assign n5397 = n5396 ^ n5389;
  assign n5398 = n5397 ^ n3437;
  assign n5399 = n3477 & ~n5398;
  assign n5400 = n5399 ^ n3477;
  assign n5401 = n5400 ^ n3437;
  assign n5402 = ~n5387 & ~n5401;
  assign n5407 = n3468 ^ n3446;
  assign n5408 = ~n3437 & n5407;
  assign n5409 = n5408 ^ n3468;
  assign n3490 = n3489 ^ n3480;
  assign n5403 = n3490 ^ n3452;
  assign n5404 = n5403 ^ n3450;
  assign n5405 = ~n3437 & n5404;
  assign n5406 = n5405 ^ n3450;
  assign n5410 = n5409 ^ n5406;
  assign n5411 = ~n3438 & n5410;
  assign n5412 = n5411 ^ n5406;
  assign n5413 = n5402 & ~n5412;
  assign n5414 = ~n4764 & n5413;
  assign n5415 = ~n3472 & n5414;
  assign n5416 = ~n3459 & n5415;
  assign n5417 = ~n4505 & n5416;
  assign n5418 = ~n3449 & n5417;
  assign n5419 = ~n4497 & n5418;
  assign n5420 = n5419 ^ n2127;
  assign n5421 = n5420 ^ x241;
  assign n5422 = n5385 & n5421;
  assign n5423 = n5422 ^ n5385;
  assign n5429 = n5423 ^ n5421;
  assign n5430 = n5426 & ~n5429;
  assign n5427 = n5426 ^ n5425;
  assign n5428 = n5423 & n5427;
  assign n5431 = n5430 ^ n5428;
  assign n5432 = ~n5354 & n5431;
  assign n5433 = n5432 ^ n5430;
  assign n5434 = n5353 & n5433;
  assign n5461 = n5353 & n5354;
  assign n5979 = n5461 ^ n5354;
  assign n5986 = n5979 ^ n5353;
  assign n5456 = n5422 & n5427;
  assign n5436 = n5427 ^ n5424;
  assign n5448 = ~n5429 & ~n5436;
  assign n5440 = n5429 ^ n5385;
  assign n5441 = ~n5436 & n5440;
  assign n5454 = n5448 ^ n5441;
  assign n7190 = n5456 ^ n5454;
  assign n7191 = ~n5986 & n7190;
  assign n5462 = n5426 ^ n5424;
  assign n5471 = n5423 & n5462;
  assign n5463 = n5385 & n5462;
  assign n5477 = n5471 ^ n5463;
  assign n5439 = n5427 & ~n5429;
  assign n5449 = n5448 ^ n5439;
  assign n5447 = n5430 ^ n5429;
  assign n5450 = n5449 ^ n5447;
  assign n5464 = n5463 ^ n5450;
  assign n5469 = n5464 ^ n5462;
  assign n5468 = n5423 & n5426;
  assign n5470 = n5469 ^ n5468;
  assign n5478 = n5477 ^ n5470;
  assign n5437 = n5422 & ~n5436;
  assign n7197 = n5478 ^ n5437;
  assign n5453 = n5437 ^ n5436;
  assign n5455 = n5454 ^ n5453;
  assign n5457 = n5456 ^ n5455;
  assign n5985 = n5457 ^ n5439;
  assign n7198 = n7197 ^ n5985;
  assign n5482 = n5422 & n5426;
  assign n7193 = n5482 ^ n5478;
  assign n7192 = n5468 ^ n5464;
  assign n7194 = n7193 ^ n7192;
  assign n7195 = n5354 & n7194;
  assign n7196 = n7195 ^ n7192;
  assign n7199 = n7198 ^ n7196;
  assign n7200 = n7199 ^ n7196;
  assign n7201 = n5354 & n7200;
  assign n7202 = n7201 ^ n7196;
  assign n7203 = n5353 & ~n7202;
  assign n7204 = n7203 ^ n7196;
  assign n7205 = ~n7191 & n7204;
  assign n5467 = n5426 & n5440;
  assign n6604 = n5467 ^ n5450;
  assign n7206 = n6604 ^ n5437;
  assign n5483 = n5482 ^ n5469;
  assign n7207 = n7206 ^ n5483;
  assign n5452 = n5427 & n5440;
  assign n7208 = n7207 ^ n5452;
  assign n7209 = n7208 ^ n5452;
  assign n7210 = ~n5354 & n7209;
  assign n7211 = n7210 ^ n5452;
  assign n7212 = n5353 & n7211;
  assign n7213 = n7212 ^ n5452;
  assign n7214 = n7205 & ~n7213;
  assign n5980 = n5455 ^ n5439;
  assign n7215 = n5980 ^ n5979;
  assign n5987 = n5986 ^ n5354;
  assign n7216 = n5987 ^ n5430;
  assign n7217 = n5980 & ~n7216;
  assign n7218 = n7217 ^ n5987;
  assign n7219 = ~n7215 & n7218;
  assign n7220 = n7219 ^ n5979;
  assign n7221 = n7214 & ~n7220;
  assign n7222 = ~n5434 & n7221;
  assign n7223 = n7222 ^ n2302;
  assign n7224 = n7223 ^ x283;
  assign n7225 = n7189 & ~n7224;
  assign n3541 = n3540 ^ x195;
  assign n3542 = n2032 ^ x190;
  assign n3543 = ~n3541 & n3542;
  assign n3544 = n3543 ^ n3541;
  assign n3545 = n3544 ^ n3542;
  assign n3554 = n2456 ^ n2419;
  assign n3555 = n2409 & n3554;
  assign n3556 = n2432 & ~n2454;
  assign n3557 = n2458 ^ n2417;
  assign n3558 = n2411 & n3557;
  assign n3559 = n2787 ^ n2470;
  assign n3561 = ~n2454 & n3560;
  assign n3562 = n3561 ^ n2410;
  assign n3563 = n3559 & n3562;
  assign n3564 = ~n3558 & ~n3563;
  assign n3565 = ~n3556 & n3564;
  assign n3566 = ~n3555 & n3565;
  assign n3567 = n2438 ^ n2423;
  assign n3568 = n2320 & n3567;
  assign n3569 = n3568 ^ n2438;
  assign n3570 = ~n2467 & n3569;
  assign n3571 = n3566 & ~n3570;
  assign n3572 = ~n3553 & n3571;
  assign n3573 = ~n2786 & n3572;
  assign n3574 = ~n2445 & n3573;
  assign n3575 = ~n2408 & n3574;
  assign n3576 = n3575 ^ x12;
  assign n3577 = n3576 ^ x193;
  assign n3581 = n2970 ^ n2937;
  assign n3582 = n3581 ^ n2992;
  assign n3583 = n3582 ^ n2931;
  assign n3584 = ~n2960 & ~n3583;
  assign n3585 = n3584 ^ n3582;
  assign n3586 = n2980 ^ n2926;
  assign n3587 = n2965 & ~n3586;
  assign n3588 = n3412 ^ n2966;
  assign n3589 = ~n2928 & n2966;
  assign n3590 = n3589 ^ n2926;
  assign n3591 = ~n3588 & n3590;
  assign n3592 = n3591 ^ n3412;
  assign n3593 = ~n3587 & n3592;
  assign n3594 = ~n2973 & ~n3593;
  assign n3595 = n2967 & ~n3594;
  assign n3596 = n3585 & ~n3595;
  assign n3597 = n2971 ^ n2925;
  assign n3598 = n2883 & ~n3597;
  assign n3599 = n3598 ^ n2925;
  assign n3600 = n2882 & n3599;
  assign n3601 = n3596 & ~n3600;
  assign n3602 = ~n3410 & n3601;
  assign n3603 = ~n3407 & n3602;
  assign n3604 = ~n3401 & n3603;
  assign n3605 = ~n3580 & n3604;
  assign n3606 = n3605 ^ x20;
  assign n3607 = n3606 ^ x192;
  assign n3608 = ~n3577 & n3607;
  assign n3640 = n3608 ^ n3577;
  assign n3609 = n2685 ^ x191;
  assign n3636 = n3635 ^ x194;
  assign n3637 = n3609 & ~n3636;
  assign n3642 = n3637 ^ n3609;
  assign n3643 = ~n3640 & n3642;
  assign n3676 = n3643 ^ n3642;
  assign n3645 = n3642 ^ n3636;
  assign n3646 = n3645 ^ n3609;
  assign n3647 = n3640 ^ n3607;
  assign n3670 = n3647 ^ n3577;
  assign n3671 = ~n3646 & n3670;
  assign n3649 = n3636 ^ n3577;
  assign n3650 = n3649 ^ n3607;
  assign n3651 = ~n3607 & ~n3609;
  assign n3652 = n3650 & n3651;
  assign n3669 = n3652 ^ n3650;
  assign n3672 = n3671 ^ n3669;
  assign n3673 = n3672 ^ n3607;
  assign n3667 = n3608 & n3645;
  assign n3641 = n3637 & ~n3640;
  assign n3664 = n3641 ^ n3637;
  assign n3659 = n3637 & n3647;
  assign n3638 = n3608 & n3637;
  assign n3663 = n3659 ^ n3638;
  assign n3665 = n3664 ^ n3663;
  assign n3662 = n3659 ^ n3643;
  assign n3666 = n3665 ^ n3662;
  assign n3668 = n3667 ^ n3666;
  assign n3674 = n3673 ^ n3668;
  assign n3660 = n3659 ^ n3647;
  assign n3656 = n3652 ^ n3651;
  assign n3648 = ~n3646 & n3647;
  assign n3653 = n3652 ^ n3648;
  assign n3654 = n3653 ^ n3640;
  assign n3644 = n3643 ^ n3641;
  assign n3655 = n3654 ^ n3644;
  assign n3657 = n3656 ^ n3655;
  assign n3658 = n3657 ^ n3648;
  assign n3661 = n3660 ^ n3658;
  assign n3675 = n3674 ^ n3661;
  assign n3677 = n3676 ^ n3675;
  assign n3678 = n3545 & ~n3677;
  assign n4814 = ~n3544 & n3656;
  assign n3679 = n3542 ^ n3541;
  assign n3680 = n3671 ^ n3667;
  assign n3681 = n3680 ^ n3653;
  assign n3682 = ~n3542 & n3681;
  assign n3683 = n3682 ^ n3653;
  assign n3684 = n3679 & n3683;
  assign n4815 = n4814 ^ n3684;
  assign n4464 = n3665 ^ n3653;
  assign n4465 = n4464 ^ n3656;
  assign n4466 = ~n3542 & n4465;
  assign n4467 = n4466 ^ n3656;
  assign n4468 = n3541 & n4467;
  assign n3690 = n3674 ^ n3641;
  assign n5206 = ~n3679 & n3690;
  assign n4473 = n3668 ^ n3648;
  assign n5208 = n4473 ^ n3677;
  assign n3700 = n3665 ^ n3661;
  assign n3693 = n3645 & n3670;
  assign n5207 = n3700 ^ n3693;
  assign n5209 = n5208 ^ n5207;
  assign n5210 = n3542 & n5209;
  assign n5211 = n5210 ^ n5207;
  assign n5212 = n5211 ^ n3638;
  assign n5213 = n5211 ^ n3541;
  assign n5214 = n5211 & ~n5213;
  assign n5215 = n5214 ^ n5211;
  assign n5216 = ~n5212 & n5215;
  assign n5217 = n5216 ^ n5214;
  assign n5218 = n5217 ^ n5211;
  assign n5219 = n5218 ^ n3541;
  assign n5220 = ~n5206 & ~n5219;
  assign n5221 = n5220 ^ n5206;
  assign n4459 = n3608 & ~n3646;
  assign n4818 = n4459 ^ n3644;
  assign n4469 = n3671 ^ n3638;
  assign n4470 = n4469 ^ n3693;
  assign n4471 = n4470 ^ n3659;
  assign n5222 = n4818 ^ n4471;
  assign n5223 = n3542 & n5222;
  assign n5224 = n5223 ^ n4818;
  assign n5225 = n3541 & n5224;
  assign n5226 = ~n5221 & ~n5225;
  assign n5227 = ~n4468 & n5226;
  assign n5228 = ~n4815 & n5227;
  assign n5229 = ~n3678 & n5228;
  assign n5230 = n5229 ^ n1515;
  assign n5584 = n5230 ^ x214;
  assign n3481 = n3480 ^ n3475;
  assign n3482 = n3437 & n3481;
  assign n3483 = n3482 ^ n3480;
  assign n3484 = n3438 & n3483;
  assign n3485 = n3460 ^ n3452;
  assign n3486 = n3439 & n3485;
  assign n3487 = n3468 ^ n3450;
  assign n3488 = ~n3466 & n3487;
  assign n3491 = n3437 & n3490;
  assign n3493 = n3492 ^ n3491;
  assign n3494 = n3438 & n3493;
  assign n3495 = n3494 ^ n3492;
  assign n3496 = ~n3488 & ~n3495;
  assign n3497 = ~n3486 & n3496;
  assign n3501 = n3437 ^ n3308;
  assign n3502 = ~n3438 & ~n3501;
  assign n3503 = n3441 & n3502;
  assign n3504 = n3500 & ~n3503;
  assign n3498 = n3474 ^ n3453;
  assign n3499 = ~n3437 & n3498;
  assign n3505 = n3504 ^ n3499;
  assign n3506 = n3438 & ~n3505;
  assign n3507 = n3506 ^ n3504;
  assign n3508 = n3497 & n3507;
  assign n3509 = ~n3484 & n3508;
  assign n3510 = ~n3472 & n3509;
  assign n3511 = n3465 & n3510;
  assign n3512 = ~n3449 & n3511;
  assign n3513 = ~n3396 & n3512;
  assign n3514 = n3513 ^ n1124;
  assign n5585 = n3514 ^ x219;
  assign n5275 = n4402 & ~n4426;
  assign n5276 = n4416 ^ n4402;
  assign n5277 = n5276 ^ n4395;
  assign n5278 = n5277 ^ n4408;
  assign n5279 = n5278 ^ n4408;
  assign n5280 = n4311 & n5279;
  assign n5281 = n5280 ^ n4408;
  assign n5282 = n4313 & n5281;
  assign n5283 = n5282 ^ n4408;
  assign n5284 = ~n5275 & ~n5283;
  assign n5285 = n4370 ^ n4367;
  assign n5286 = n5285 ^ n4419;
  assign n5287 = n5286 ^ n4391;
  assign n5288 = ~n4311 & n5287;
  assign n5289 = n5288 ^ n4391;
  assign n5290 = n4312 & n5289;
  assign n5291 = n5284 & ~n5290;
  assign n5292 = ~n4436 & n5291;
  assign n5293 = ~n5274 & n5292;
  assign n5294 = ~n4428 & n5293;
  assign n5295 = ~n4399 & n5294;
  assign n5296 = n5295 ^ n1615;
  assign n5586 = n5296 ^ x215;
  assign n4729 = n4186 & ~n4254;
  assign n4730 = n4729 ^ n4232;
  assign n4750 = n4278 ^ n4235;
  assign n4749 = n4260 ^ n4254;
  assign n4751 = n4750 ^ n4749;
  assign n5588 = ~n4184 & n4751;
  assign n5587 = n4735 ^ n4260;
  assign n5589 = n5588 ^ n5587;
  assign n5590 = ~n4189 & ~n5589;
  assign n5591 = n5590 ^ n5587;
  assign n5592 = n4186 & n4291;
  assign n5593 = n4243 ^ n4226;
  assign n5594 = ~n4185 & n5593;
  assign n5595 = n5594 ^ n4226;
  assign n5596 = n5595 ^ n4283;
  assign n5597 = n4189 & n5596;
  assign n5598 = n5597 ^ n4283;
  assign n5599 = ~n5592 & ~n5598;
  assign n5600 = n5591 & n5599;
  assign n5601 = ~n4240 & n5600;
  assign n5602 = ~n4930 & n5601;
  assign n5603 = ~n4932 & n5602;
  assign n5604 = ~n4730 & n5603;
  assign n5605 = n5604 ^ n1706;
  assign n5606 = n5605 ^ x216;
  assign n5607 = n5586 & ~n5606;
  assign n5608 = n5607 ^ n5586;
  assign n5609 = n5608 ^ n5606;
  assign n2489 = ~n1482 & n2488;
  assign n2707 = n2706 ^ n2701;
  assign n2708 = ~n2689 & n2707;
  assign n2711 = n2710 ^ n2687;
  assign n2715 = n2714 ^ n2694;
  assign n2716 = n2715 ^ n2690;
  assign n2717 = n2711 & n2716;
  assign n2738 = ~n2688 & ~n2737;
  assign n2739 = n2738 ^ n2731;
  assign n2740 = n2739 ^ n1482;
  assign n2727 = n2726 ^ n2722;
  assign n2741 = n2740 ^ n2727;
  assign n2742 = n2741 ^ n2740;
  assign n2743 = ~n1482 & n2742;
  assign n2744 = n2743 ^ n2740;
  assign n2745 = n2686 & ~n2744;
  assign n2746 = n2745 ^ n2740;
  assign n2747 = ~n2717 & n2746;
  assign n2748 = ~n2708 & n2747;
  assign n2749 = ~n2489 & n2748;
  assign n2761 = n2760 ^ n2699;
  assign n2762 = ~n2686 & n2761;
  assign n2763 = n2762 ^ n2699;
  assign n2754 = n2753 ^ n2733;
  assign n2755 = n2754 ^ n2721;
  assign n2756 = n2755 ^ n2712;
  assign n2757 = n2756 ^ n2712;
  assign n2758 = n2686 & n2757;
  assign n2764 = n2763 ^ n2758;
  assign n2765 = n2764 ^ n2758;
  assign n2766 = ~n2712 & ~n2765;
  assign n2767 = n2766 ^ n2758;
  assign n2768 = n2750 & ~n2767;
  assign n2769 = n2768 ^ n2758;
  assign n2770 = n2749 & ~n2769;
  assign n2771 = n2770 ^ n1303;
  assign n5610 = n2771 ^ x218;
  assign n4792 = n3860 ^ n3858;
  assign n4793 = n3762 & ~n4792;
  assign n4794 = n4793 ^ n3858;
  assign n4795 = n3883 & n4794;
  assign n5611 = ~n3852 & n5359;
  assign n5612 = n3876 ^ n3851;
  assign n5613 = n3762 & ~n5612;
  assign n5614 = n3865 ^ n3849;
  assign n5615 = n3882 & n5614;
  assign n5617 = n3892 ^ n3870;
  assign n5618 = n3870 & ~n3884;
  assign n5619 = n5618 ^ n3882;
  assign n5620 = ~n5617 & n5619;
  assign n5621 = n5620 ^ n3892;
  assign n5622 = ~n3894 & ~n5621;
  assign n5616 = n3863 ^ n3849;
  assign n5623 = n5622 ^ n5616;
  assign n5624 = n3884 & ~n5623;
  assign n5625 = n5624 ^ n5616;
  assign n5626 = ~n5615 & ~n5625;
  assign n5627 = ~n3888 & n5626;
  assign n5628 = ~n5613 & n5627;
  assign n5629 = ~n5611 & n5628;
  assign n5630 = ~n3762 & ~n3872;
  assign n5631 = n5630 ^ n3858;
  assign n5632 = ~n3761 & n5631;
  assign n5633 = n5629 & ~n5632;
  assign n5634 = ~n4795 & n5633;
  assign n5635 = ~n5363 & n5634;
  assign n5636 = ~n3885 & n5635;
  assign n5637 = n5636 ^ n1742;
  assign n5638 = n5637 ^ x217;
  assign n5639 = ~n5610 & n5638;
  assign n5640 = n5639 ^ n5610;
  assign n5643 = n5640 ^ n5638;
  assign n5644 = n5609 & n5643;
  assign n5642 = n5609 & n5639;
  assign n5645 = n5644 ^ n5642;
  assign n5652 = ~n5585 & n5645;
  assign n5653 = n5652 ^ n5642;
  assign n5648 = n5607 & n5643;
  assign n5646 = n5645 ^ n5609;
  assign n5641 = n5609 & ~n5640;
  assign n5647 = n5646 ^ n5641;
  assign n5649 = n5648 ^ n5647;
  assign n5650 = n5585 & n5649;
  assign n5651 = n5650 ^ n5647;
  assign n5654 = n5653 ^ n5651;
  assign n5655 = n5584 & n5654;
  assign n5656 = n5655 ^ n5651;
  assign n5657 = n5607 ^ n5606;
  assign n5658 = ~n5640 & ~n5657;
  assign n5659 = ~n5584 & ~n5585;
  assign n5660 = n5659 ^ n5584;
  assign n5661 = n5660 ^ n5585;
  assign n5662 = n5661 ^ n5584;
  assign n5663 = n5658 & ~n5662;
  assign n6192 = n5641 & ~n5662;
  assign n5696 = n5639 & ~n5657;
  assign n6189 = n5585 ^ n5584;
  assign n6190 = n5696 & ~n6189;
  assign n5670 = n5643 & ~n5657;
  assign n6188 = ~n5661 & n5670;
  assign n6191 = n6190 ^ n6188;
  assign n6193 = n6192 ^ n6191;
  assign n5673 = n5608 & n5639;
  assign n5672 = n5608 & n5643;
  assign n5674 = n5673 ^ n5672;
  assign n5685 = n5674 ^ n5608;
  assign n5664 = n5643 ^ n5610;
  assign n5682 = n5607 & n5664;
  assign n5683 = n5682 ^ n5664;
  assign n5665 = ~n5657 & n5664;
  assign n5666 = n5665 ^ n5647;
  assign n5684 = n5683 ^ n5666;
  assign n5686 = n5685 ^ n5684;
  assign n5692 = n5686 ^ n5647;
  assign n5693 = ~n5584 & n5692;
  assign n5694 = n5693 ^ n5647;
  assign n5695 = n5585 & n5694;
  assign n5687 = n5686 ^ n5644;
  assign n5688 = n5584 & n5687;
  assign n5689 = n5688 ^ n5644;
  assign n5690 = n5585 & n5689;
  assign n6194 = n5673 ^ n5648;
  assign n6195 = n6194 ^ n5682;
  assign n5698 = n5607 & ~n5640;
  assign n5699 = n5698 ^ n5682;
  assign n5705 = n5699 ^ n5607;
  assign n5706 = n5705 ^ n5648;
  assign n6196 = n6195 ^ n5706;
  assign n7173 = n6196 ^ n5670;
  assign n6456 = n5698 ^ n5696;
  assign n6463 = n6456 ^ n5642;
  assign n7171 = n6463 ^ n5647;
  assign n7172 = n7171 ^ n5682;
  assign n7174 = n7173 ^ n7172;
  assign n7175 = n5584 & n7174;
  assign n7176 = n7175 ^ n7172;
  assign n6208 = n5686 ^ n5665;
  assign n7166 = n6208 ^ n5641;
  assign n5707 = n5706 ^ n5684;
  assign n6202 = n5707 ^ n5672;
  assign n7167 = n7166 ^ n6202;
  assign n7168 = n7167 ^ n6195;
  assign n7169 = ~n5584 & n7168;
  assign n7170 = n7169 ^ n6195;
  assign n7177 = n7176 ^ n7170;
  assign n7178 = n6189 & n7177;
  assign n7179 = n7178 ^ n7170;
  assign n7180 = ~n5690 & ~n7179;
  assign n7181 = ~n5695 & n7180;
  assign n7182 = ~n6193 & n7181;
  assign n7183 = ~n5663 & n7182;
  assign n7184 = ~n5656 & n7183;
  assign n7185 = n7184 ^ n1829;
  assign n7186 = n7185 ^ x282;
  assign n5297 = n5296 ^ x213;
  assign n4800 = ~n3762 & ~n3856;
  assign n4801 = n4800 ^ n3855;
  assign n4796 = n3897 ^ n3863;
  assign n4797 = n4796 ^ n3857;
  assign n4798 = ~n3762 & n4797;
  assign n4799 = n4798 ^ n4796;
  assign n4802 = n4801 ^ n4799;
  assign n4803 = ~n3883 & n4802;
  assign n4804 = n4803 ^ n4799;
  assign n4806 = n3762 & n3845;
  assign n4805 = n3874 & n3883;
  assign n4807 = n4806 ^ n4805;
  assign n4808 = n4804 & ~n4807;
  assign n4809 = ~n3887 & n4808;
  assign n4810 = ~n4795 & n4809;
  assign n4811 = ~n3881 & n4810;
  assign n4812 = n4811 ^ n2319;
  assign n5298 = n4812 ^ x208;
  assign n5135 = n2709 & n2728;
  assign n5136 = n2752 ^ n2732;
  assign n5137 = ~n2689 & n5136;
  assign n5140 = n2706 ^ n2694;
  assign n5141 = n5140 ^ n2726;
  assign n5142 = n2688 & n5141;
  assign n5150 = n4995 ^ n2733;
  assign n5145 = n5144 ^ n5008;
  assign n5146 = n5145 ^ n2694;
  assign n5143 = n2706 ^ n2690;
  assign n5147 = n5146 ^ n5143;
  assign n5148 = ~n2686 & n5147;
  assign n5149 = n5148 ^ n5143;
  assign n5151 = n5150 ^ n5149;
  assign n5152 = n5151 ^ n5149;
  assign n5153 = n2686 & n5152;
  assign n5154 = n5153 ^ n5149;
  assign n5155 = n1482 & n5154;
  assign n5156 = n5155 ^ n5149;
  assign n5157 = ~n5142 & ~n5156;
  assign n5158 = ~n5139 & n5157;
  assign n5159 = ~n5137 & n5158;
  assign n5160 = ~n5135 & n5159;
  assign n5161 = n2730 & n2750;
  assign n5162 = n2733 ^ n2722;
  assign n5163 = n5162 ^ n2487;
  assign n5164 = ~n2686 & n5163;
  assign n5165 = n5164 ^ n2487;
  assign n5166 = n5165 ^ n2726;
  assign n5167 = n1482 & n5166;
  assign n5168 = n5167 ^ n2726;
  assign n5169 = ~n5161 & ~n5168;
  assign n5170 = n5160 & n5169;
  assign n5171 = ~n4985 & n5170;
  assign n5172 = n5171 ^ n2380;
  assign n5173 = n5172 ^ x211;
  assign n4712 = ~n3937 & ~n4058;
  assign n4713 = n4712 ^ n4021;
  assign n4715 = n4084 ^ n4050;
  assign n4714 = n4062 ^ n4047;
  assign n4716 = n4715 ^ n4714;
  assign n4717 = ~n3937 & n4716;
  assign n4718 = n4717 ^ n4549;
  assign n4078 = n4062 ^ n4035;
  assign n4079 = n4078 ^ n4055;
  assign n4080 = ~n3937 & ~n4079;
  assign n4719 = n4718 ^ n4080;
  assign n4720 = n4719 ^ n4055;
  assign n4721 = n4720 ^ n4713;
  assign n4722 = ~n4713 & n4721;
  assign n4069 = n4030 ^ n4021;
  assign n4070 = ~n4046 & n4069;
  assign n4067 = n4044 ^ n4030;
  assign n4709 = n4070 ^ n4067;
  assign n4710 = n3937 & ~n4709;
  assign n4711 = n4710 ^ n4070;
  assign n4723 = n4722 ^ n4711;
  assign n4724 = n3918 & ~n4723;
  assign n4725 = n4724 ^ n4722;
  assign n4726 = ~n4062 & n4725;
  assign n4727 = n4726 ^ n2395;
  assign n5232 = n4727 ^ x209;
  assign n5240 = n5173 & n5232;
  assign n5249 = n5240 ^ n5173;
  assign n4568 = n3251 ^ n3197;
  assign n4569 = ~n2846 & n4568;
  assign n4570 = n4569 ^ n3197;
  assign n4571 = n3200 & n4570;
  assign n5174 = n3200 & n3240;
  assign n5175 = ~n3200 & n3245;
  assign n5186 = n3250 ^ n3192;
  assign n5187 = n2847 & ~n5186;
  assign n5188 = n5187 ^ n2846;
  assign n5184 = n3221 & ~n3251;
  assign n5185 = n5184 ^ n3220;
  assign n5189 = n5188 ^ n5185;
  assign n5181 = n3196 & ~n3199;
  assign n4561 = n2847 & n3251;
  assign n4562 = n4561 ^ n3198;
  assign n5182 = n5181 ^ n4562;
  assign n5176 = n3250 ^ n3209;
  assign n5177 = n2809 & ~n5176;
  assign n5178 = n5177 ^ n3209;
  assign n5179 = n5178 ^ n3222;
  assign n4557 = n3238 ^ n3194;
  assign n4558 = ~n3200 & n4557;
  assign n5180 = n5179 ^ n4558;
  assign n5183 = n5182 ^ n5180;
  assign n5190 = n5189 ^ n5183;
  assign n5191 = ~n5175 & n5190;
  assign n5192 = n3236 ^ n3223;
  assign n5193 = n2809 & n5192;
  assign n5194 = n5193 ^ n3223;
  assign n5195 = n5191 & ~n5194;
  assign n5196 = n3249 ^ n3216;
  assign n5197 = ~n2809 & n5196;
  assign n5198 = n5197 ^ n3216;
  assign n5199 = n2846 & n5198;
  assign n5200 = n5195 & ~n5199;
  assign n5201 = ~n3235 & n5200;
  assign n5202 = ~n5174 & n5201;
  assign n5203 = ~n4571 & n5202;
  assign n5204 = n5203 ^ n2349;
  assign n5205 = n5204 ^ x210;
  assign n5231 = n5230 ^ x212;
  assign n5239 = n5205 & n5231;
  assign n5244 = n5239 ^ n5231;
  assign n5245 = n5244 ^ n5205;
  assign n5259 = n5245 ^ n5231;
  assign n5260 = n5249 & n5259;
  assign n5250 = n5249 ^ n5232;
  assign n5254 = n5244 & ~n5250;
  assign n5261 = n5260 ^ n5254;
  assign n5258 = n5244 & n5249;
  assign n5262 = n5261 ^ n5258;
  assign n5233 = n5232 ^ n5231;
  assign n5234 = n5233 ^ n5205;
  assign n5263 = n5262 ^ n5234;
  assign n5255 = n5254 ^ n5250;
  assign n5252 = ~n5245 & ~n5250;
  assign n5251 = n5239 & ~n5250;
  assign n5253 = n5252 ^ n5251;
  assign n5256 = n5255 ^ n5253;
  assign n5246 = n5240 & ~n5245;
  assign n5243 = n5239 & n5240;
  assign n5247 = n5246 ^ n5243;
  assign n5241 = n5240 ^ n5232;
  assign n5242 = n5239 & n5241;
  assign n5248 = n5247 ^ n5242;
  assign n5257 = n5256 ^ n5248;
  assign n5264 = n5263 ^ n5257;
  assign n5265 = n5264 ^ n5253;
  assign n5266 = n5265 ^ n5250;
  assign n5235 = n5234 ^ n5231;
  assign n5236 = n5205 & ~n5235;
  assign n5237 = n5236 ^ n5234;
  assign n5238 = ~n5173 & n5237;
  assign n5267 = n5266 ^ n5238;
  assign n5299 = n5267 ^ n5264;
  assign n5300 = ~n5298 & ~n5299;
  assign n5301 = n5300 ^ n5267;
  assign n5302 = ~n5297 & n5301;
  assign n5308 = ~n5297 & n5298;
  assign n5309 = n5308 ^ n5298;
  assign n5314 = n5260 & n5309;
  assign n5914 = n5258 & n5308;
  assign n5322 = n5264 ^ n5246;
  assign n5321 = n5252 ^ n5245;
  assign n5323 = n5322 ^ n5321;
  assign n5915 = n5323 ^ n5251;
  assign n5268 = n5267 ^ n5242;
  assign n5269 = n5268 ^ n5243;
  assign n5310 = n5269 ^ n5251;
  assign n5311 = n5310 ^ n5239;
  assign n5312 = n5311 ^ n5267;
  assign n5916 = n5915 ^ n5312;
  assign n5917 = n5916 ^ n5312;
  assign n5918 = n5297 & n5917;
  assign n5919 = n5918 ^ n5312;
  assign n5920 = n5298 & n5919;
  assign n5921 = n5920 ^ n5312;
  assign n5922 = ~n5914 & ~n5921;
  assign n5303 = n5298 ^ n5297;
  assign n5304 = n5261 & n5298;
  assign n5305 = n5304 ^ n5258;
  assign n5306 = n5303 & n5305;
  assign n5307 = n5306 ^ n5258;
  assign n5923 = n5312 ^ n5260;
  assign n5924 = n5298 & n5923;
  assign n5925 = n5924 ^ n5260;
  assign n5926 = ~n5297 & n5925;
  assign n5316 = n5309 ^ n5297;
  assign n5325 = n5242 ^ n5241;
  assign n5326 = n5325 ^ n5299;
  assign n5335 = n5326 ^ n5240;
  assign n5333 = n5326 ^ n5247;
  assign n5270 = n5269 ^ n5236;
  assign n5334 = n5333 ^ n5270;
  assign n5336 = n5335 ^ n5334;
  assign n5927 = n5336 ^ n5270;
  assign n5928 = n5927 ^ n5267;
  assign n5929 = n5316 & n5928;
  assign n5930 = ~n5257 & n5298;
  assign n5931 = n5930 ^ n5256;
  assign n5932 = ~n5297 & ~n5931;
  assign n5935 = n5270 ^ n5242;
  assign n5936 = ~n5309 & ~n5935;
  assign n5938 = n5270 & ~n5297;
  assign n5939 = ~n5298 & n5938;
  assign n5937 = n5268 ^ n5246;
  assign n5940 = n5939 ^ n5937;
  assign n5941 = ~n5936 & n5940;
  assign n5942 = n5326 & ~n5941;
  assign n5933 = n5265 ^ n5243;
  assign n5934 = ~n5298 & ~n5933;
  assign n5943 = n5942 ^ n5934;
  assign n5944 = n5303 & ~n5943;
  assign n5945 = n5944 ^ n5942;
  assign n5946 = ~n5932 & n5945;
  assign n5947 = ~n5929 & n5946;
  assign n5948 = ~n5926 & n5947;
  assign n5949 = ~n5307 & n5948;
  assign n5950 = n5922 & n5949;
  assign n5951 = ~n5314 & n5950;
  assign n5952 = ~n5302 & n5951;
  assign n5953 = n5952 ^ n2483;
  assign n7187 = n5953 ^ x281;
  assign n7188 = ~n7186 & ~n7187;
  assign n7228 = n7188 ^ n7186;
  assign n7246 = n7225 & ~n7228;
  assign n7247 = n7246 ^ n7228;
  assign n7226 = n7225 ^ n7189;
  assign n7232 = n7226 ^ n7224;
  assign n7243 = n7232 ^ n7189;
  assign n7244 = ~n7228 & ~n7243;
  assign n7238 = ~n7228 & n7232;
  assign n7245 = n7244 ^ n7238;
  assign n7248 = n7247 ^ n7245;
  assign n7257 = n7248 ^ n7226;
  assign n7229 = n7228 ^ n7187;
  assign n7251 = ~n7229 & ~n7243;
  assign n7252 = n7251 ^ n7246;
  assign n7253 = n7252 ^ n7244;
  assign n7254 = n7253 ^ n7187;
  assign n7236 = n7188 & n7232;
  assign n7231 = n7188 & n7225;
  assign n7237 = n7236 ^ n7231;
  assign n7239 = n7238 ^ n7237;
  assign n7240 = n7239 ^ n7232;
  assign n7233 = n7229 ^ n7186;
  assign n7234 = n7232 & ~n7233;
  assign n7235 = n7234 ^ n7231;
  assign n7241 = n7240 ^ n7235;
  assign n7230 = n7225 & ~n7229;
  assign n7242 = n7241 ^ n7230;
  assign n7249 = n7248 ^ n7242;
  assign n7250 = n7249 ^ n7238;
  assign n7255 = n7254 ^ n7250;
  assign n7227 = n7188 & n7226;
  assign n7256 = n7255 ^ n7227;
  assign n7258 = n7257 ^ n7256;
  assign n7259 = n7258 ^ n7248;
  assign n4559 = n2848 & n3242;
  assign n4560 = n4559 ^ n4558;
  assign n4686 = n3216 ^ n3195;
  assign n4687 = ~n3200 & n4686;
  assign n4563 = n3254 ^ n3204;
  assign n4694 = n4563 ^ n3228;
  assign n4695 = n4694 ^ n3207;
  assign n4696 = ~n2809 & ~n4695;
  assign n4697 = n4696 ^ n4694;
  assign n4690 = n3252 ^ n3201;
  assign n4688 = n3250 ^ n3231;
  assign n4689 = n4688 ^ n3202;
  assign n4691 = n4690 ^ n4689;
  assign n4692 = ~n2809 & n4691;
  assign n4693 = n4692 ^ n4689;
  assign n4698 = n4697 ^ n4693;
  assign n4699 = n2846 & n4698;
  assign n4700 = n4699 ^ n4693;
  assign n4701 = ~n4687 & ~n4700;
  assign n4702 = n3214 & n4701;
  assign n4703 = ~n4560 & n4702;
  assign n4704 = ~n3232 & n4703;
  assign n4705 = ~n3234 & n4704;
  assign n4706 = ~n4571 & n4705;
  assign n4707 = n4706 ^ n2622;
  assign n4708 = n4707 ^ x250;
  assign n4728 = n4727 ^ x255;
  assign n4894 = ~n4708 & n4728;
  assign n4895 = n4894 ^ n4728;
  assign n4736 = n4735 ^ n4226;
  assign n4737 = ~n4189 & ~n4736;
  assign n4739 = n4738 ^ n4281;
  assign n4740 = ~n4188 & ~n4739;
  assign n4741 = ~n4737 & ~n4740;
  assign n4742 = n4284 ^ n4260;
  assign n4743 = n4742 ^ n4256;
  assign n4744 = n4184 & n4743;
  assign n4745 = n4744 ^ n4256;
  assign n4746 = n4185 & n4745;
  assign n4747 = n4741 & ~n4746;
  assign n4748 = n4283 ^ n4187;
  assign n4752 = n4751 ^ n4271;
  assign n4753 = ~n4283 & ~n4752;
  assign n4754 = n4753 ^ n4271;
  assign n4755 = n4748 & n4754;
  assign n4756 = n4755 ^ n4187;
  assign n4757 = n4747 & ~n4756;
  assign n4758 = ~n4733 & n4757;
  assign n4759 = ~n4272 & n4758;
  assign n4760 = ~n4730 & n4759;
  assign n4761 = n4760 ^ n2533;
  assign n4762 = n4761 ^ x252;
  assign n4770 = n3456 ^ n3454;
  assign n4771 = n4770 ^ n3492;
  assign n4772 = n3438 & n4771;
  assign n4766 = n4520 ^ n3454;
  assign n4765 = n3478 ^ n3455;
  assign n4767 = n4766 ^ n4765;
  assign n4768 = ~n3438 & n4767;
  assign n4769 = n4768 ^ n4765;
  assign n4773 = n4772 ^ n4769;
  assign n4774 = n3466 & ~n4773;
  assign n4775 = n4774 ^ n4769;
  assign n4777 = n3437 & n3489;
  assign n4776 = n3460 & ~n3466;
  assign n4778 = n4777 ^ n4776;
  assign n4779 = n4775 & ~n4778;
  assign n4780 = n3439 & n3446;
  assign n4781 = n4780 ^ n4534;
  assign n4782 = n4779 & ~n4781;
  assign n4783 = ~n3484 & n4782;
  assign n4784 = ~n4509 & n4783;
  assign n4785 = ~n4764 & n4784;
  assign n4786 = ~n3449 & n4785;
  assign n4787 = ~n4497 & n4786;
  assign n4788 = n4787 ^ n2569;
  assign n4789 = n4788 ^ x253;
  assign n4790 = ~n4762 & n4789;
  assign n4844 = n4790 ^ n4789;
  assign n4813 = n4812 ^ x254;
  assign n3639 = n3545 & n3638;
  assign n3688 = n3667 ^ n3655;
  assign n4460 = n4459 ^ n3688;
  assign n4461 = n3542 & ~n4460;
  assign n4462 = n4461 ^ n4459;
  assign n4463 = ~n3541 & n4462;
  assign n4816 = n3659 & ~n3679;
  assign n4826 = n3690 ^ n3677;
  assign n4827 = n4826 ^ n3653;
  assign n4824 = n4469 ^ n3657;
  assign n4825 = n4824 ^ n3700;
  assign n4828 = n4827 ^ n4825;
  assign n4829 = ~n3542 & ~n4828;
  assign n4830 = n4829 ^ n4825;
  assign n4479 = n3693 ^ n3675;
  assign n4819 = n4479 ^ n3648;
  assign n4820 = n4819 ^ n4818;
  assign n4817 = n3666 ^ n3656;
  assign n4821 = n4820 ^ n4817;
  assign n4822 = n3542 & ~n4821;
  assign n4823 = n4822 ^ n4817;
  assign n4831 = n4830 ^ n4823;
  assign n4832 = ~n3541 & n4831;
  assign n4833 = n4832 ^ n4823;
  assign n4834 = ~n4816 & ~n4833;
  assign n4835 = ~n4463 & n4834;
  assign n4836 = ~n4815 & n4835;
  assign n4837 = ~n3639 & n4836;
  assign n4838 = n4837 ^ n2509;
  assign n4839 = n4838 ^ x251;
  assign n4840 = n4813 & n4839;
  assign n4859 = n4840 ^ n4813;
  assign n4864 = n4844 & n4859;
  assign n4860 = n4790 & n4859;
  assign n4865 = n4864 ^ n4860;
  assign n4866 = n4865 ^ n4859;
  assign n4791 = n4790 ^ n4762;
  assign n4853 = ~n4791 & n4840;
  assign n4841 = n4840 ^ n4839;
  assign n4845 = n4841 ^ n4813;
  assign n4850 = n4790 & ~n4845;
  assign n4851 = n4850 ^ n4845;
  assign n4847 = n4844 ^ n4762;
  assign n4848 = ~n4845 & n4847;
  assign n4846 = n4844 & ~n4845;
  assign n4849 = n4848 ^ n4846;
  assign n4852 = n4851 ^ n4849;
  assign n4854 = n4853 ^ n4852;
  assign n4842 = ~n4791 & n4841;
  assign n4843 = n4842 ^ n4791;
  assign n4855 = n4854 ^ n4843;
  assign n4867 = n4866 ^ n4855;
  assign n5779 = n4867 ^ n4852;
  assign n5780 = n4895 & ~n5779;
  assign n4872 = n4853 ^ n4840;
  assign n4869 = n4848 ^ n4847;
  assign n4863 = n4841 & n4847;
  assign n4868 = n4867 ^ n4863;
  assign n4870 = n4869 ^ n4868;
  assign n4857 = n4790 & n4840;
  assign n4871 = n4870 ^ n4857;
  assign n4873 = n4872 ^ n4871;
  assign n4861 = n4860 ^ n4850;
  assign n4858 = n4857 ^ n4790;
  assign n4862 = n4861 ^ n4858;
  assign n4874 = n4873 ^ n4862;
  assign n4856 = n4855 ^ n4848;
  assign n4875 = n4874 ^ n4856;
  assign n4876 = ~n4728 & n4875;
  assign n4877 = n4876 ^ n4874;
  assign n4878 = ~n4708 & n4877;
  assign n4896 = n4895 ^ n4708;
  assign n6229 = n4874 & n4896;
  assign n4897 = n4842 & n4896;
  assign n6230 = n6229 ^ n4897;
  assign n4881 = n4870 ^ n4863;
  assign n4882 = n4881 ^ n4862;
  assign n4879 = n4870 ^ n4842;
  assign n4880 = n4879 ^ n4841;
  assign n4883 = n4882 ^ n4880;
  assign n4884 = n4883 ^ n4857;
  assign n4885 = n4884 ^ n4850;
  assign n4886 = n4728 & n4885;
  assign n4887 = n4886 ^ n4850;
  assign n4888 = n4708 & n4887;
  assign n4889 = n4728 ^ n4708;
  assign n5773 = n4853 ^ n4848;
  assign n5774 = n4708 & n5773;
  assign n5775 = n5774 ^ n4848;
  assign n5776 = n4889 & n5775;
  assign n4901 = n4896 ^ n4728;
  assign n6231 = n4879 & ~n4901;
  assign n6806 = n4881 ^ n4842;
  assign n6807 = n6806 ^ n4865;
  assign n6808 = n6807 ^ n4850;
  assign n6809 = n6808 ^ n4850;
  assign n6810 = ~n4708 & n6809;
  assign n6811 = n6810 ^ n4850;
  assign n6812 = n4889 & n6811;
  assign n6813 = n6812 ^ n4850;
  assign n4898 = n4867 ^ n4846;
  assign n4899 = n4898 ^ n4864;
  assign n6819 = n4708 & n4899;
  assign n6815 = n4853 ^ n4849;
  assign n6814 = n4884 ^ n4860;
  assign n6816 = n6815 ^ n6814;
  assign n6817 = n4708 & n6816;
  assign n6818 = n6817 ^ n6814;
  assign n6820 = n6819 ^ n6818;
  assign n6821 = n4889 & n6820;
  assign n6822 = n6821 ^ n6818;
  assign n6823 = ~n6813 & ~n6822;
  assign n6824 = ~n6231 & n6823;
  assign n6825 = ~n5776 & n6824;
  assign n6826 = ~n4888 & n6825;
  assign n6827 = ~n6230 & n6826;
  assign n6828 = ~n4878 & n6827;
  assign n6829 = ~n5780 & n6828;
  assign n6830 = n6829 ^ n2685;
  assign n7260 = n6830 ^ x285;
  assign n3917 = n3916 ^ x224;
  assign n4071 = ~n3918 & ~n4070;
  assign n4068 = ~n3918 & ~n4062;
  assign n4072 = n4071 ^ n4068;
  assign n4073 = n4072 ^ n4071;
  assign n4074 = n4067 & n4073;
  assign n4075 = n4074 ^ n4071;
  assign n4076 = n3937 & n4075;
  assign n4077 = n4076 ^ n4071;
  assign n4081 = n4080 ^ n4055;
  assign n4088 = n4087 ^ n4081;
  assign n4089 = n4081 ^ n3918;
  assign n4090 = n4081 & n4089;
  assign n4091 = n4090 ^ n4081;
  assign n4092 = ~n4088 & n4091;
  assign n4093 = n4092 ^ n4090;
  assign n4094 = n4093 ^ n4081;
  assign n4095 = n4094 ^ n3918;
  assign n4096 = ~n4077 & n4095;
  assign n4097 = n4096 ^ n4077;
  assign n4098 = ~n4066 & ~n4097;
  assign n4099 = n4098 ^ n1198;
  assign n4100 = n4099 ^ x222;
  assign n4101 = ~n3917 & ~n4100;
  assign n3515 = n3514 ^ x221;
  assign n3685 = ~n3541 & ~n3658;
  assign n3686 = n3685 ^ n3648;
  assign n3687 = ~n3542 & n3686;
  assign n3689 = ~n3679 & ~n3688;
  assign n3691 = n3690 ^ n3657;
  assign n3692 = n3545 & ~n3691;
  assign n3694 = n3693 ^ n3648;
  assign n3695 = n3543 & n3694;
  assign n3696 = n3677 ^ n3663;
  assign n3697 = ~n3544 & ~n3696;
  assign n3698 = n3696 ^ n3661;
  assign n3699 = ~n3543 & ~n3698;
  assign n3701 = n3700 ^ n3644;
  assign n3702 = ~n3699 & ~n3701;
  assign n3703 = ~n3697 & ~n3702;
  assign n3704 = ~n3541 & ~n3703;
  assign n3705 = ~n3695 & ~n3704;
  assign n3706 = ~n3692 & n3705;
  assign n3707 = ~n3689 & n3706;
  assign n3708 = n3542 & n3669;
  assign n3709 = n3708 ^ n3671;
  assign n3710 = n3541 & n3709;
  assign n3711 = n3710 ^ n3671;
  assign n3712 = n3707 & ~n3711;
  assign n3713 = ~n3687 & n3712;
  assign n3714 = ~n3684 & n3713;
  assign n3715 = ~n3678 & n3714;
  assign n3716 = ~n3639 & n3715;
  assign n3717 = n3716 ^ n1029;
  assign n3718 = n3717 ^ x223;
  assign n3719 = ~n3515 & n3718;
  assign n3720 = n3719 ^ n3718;
  assign n4105 = n3720 ^ n3515;
  assign n4106 = n4101 & n4105;
  assign n4124 = n4106 ^ n4105;
  assign n4119 = n4101 ^ n4100;
  assign n4122 = n4105 & ~n4119;
  assign n4111 = n4101 ^ n3917;
  assign n4113 = n4105 & ~n4111;
  assign n4123 = n4122 ^ n4113;
  assign n4125 = n4124 ^ n4123;
  assign n2772 = n2771 ^ x220;
  assign n3274 = n3273 ^ x225;
  assign n3275 = n2772 & n3274;
  assign n4110 = n3275 ^ n3274;
  assign n4156 = n4110 ^ n2772;
  assign n5726 = n4125 & ~n4156;
  assign n3276 = n3275 ^ n2772;
  assign n4104 = n3719 & n4101;
  assign n4107 = n4106 ^ n4104;
  assign n4102 = n3720 & n4101;
  assign n4103 = n4102 ^ n4101;
  assign n4108 = n4107 ^ n4103;
  assign n4109 = n3276 & n4108;
  assign n4131 = n4119 ^ n3917;
  assign n4134 = n3720 & ~n4131;
  assign n5727 = n3275 & n4134;
  assign n4152 = n4108 & n4110;
  assign n5728 = n5727 ^ n4152;
  assign n4148 = n4134 ^ n4122;
  assign n4149 = ~n2772 & n4148;
  assign n4150 = n4149 ^ n4134;
  assign n4151 = ~n3274 & n4150;
  assign n4120 = n3719 ^ n3515;
  assign n4121 = ~n4119 & ~n4120;
  assign n4126 = n4125 ^ n4121;
  assign n4127 = ~n2772 & n4126;
  assign n4128 = n4127 ^ n4125;
  assign n4129 = n3274 & n4128;
  assign n5729 = n3275 & n4122;
  assign n4141 = n3274 ^ n2772;
  assign n5733 = n3275 & n4107;
  assign n4115 = n3719 & ~n4111;
  assign n4116 = n4115 ^ n4111;
  assign n4112 = n3720 & ~n4111;
  assign n4114 = n4113 ^ n4112;
  assign n4117 = n4116 ^ n4114;
  assign n5734 = n5733 ^ n4117;
  assign n5735 = n5734 ^ n4102;
  assign n4142 = ~n4120 & ~n4131;
  assign n4143 = n4142 ^ n4104;
  assign n4132 = n3719 & ~n4131;
  assign n4144 = n4143 ^ n4132;
  assign n4171 = n4144 ^ n3719;
  assign n4160 = n4142 ^ n4115;
  assign n4172 = n4171 ^ n4160;
  assign n5730 = n4172 ^ n4115;
  assign n5731 = ~n4156 & n5730;
  assign n5732 = n5731 ^ n4132;
  assign n5736 = n5735 ^ n5732;
  assign n5737 = ~n4141 & ~n5736;
  assign n5738 = ~n5729 & ~n5737;
  assign n4153 = n4112 ^ n3720;
  assign n4135 = n4134 ^ n4102;
  assign n4154 = n4153 ^ n4135;
  assign n5739 = n4154 ^ n4112;
  assign n5740 = n5739 ^ n4102;
  assign n5741 = n5740 ^ n4113;
  assign n5742 = n4110 & n5741;
  assign n5743 = n4143 ^ n4121;
  assign n5744 = n5743 ^ n4114;
  assign n5745 = n4114 ^ n3276;
  assign n5746 = ~n4114 & ~n5745;
  assign n5747 = n5746 ^ n4114;
  assign n5748 = n5744 & ~n5747;
  assign n5749 = n5748 ^ n5746;
  assign n5750 = n5749 ^ n4114;
  assign n5751 = n5750 ^ n3276;
  assign n5752 = ~n5742 & ~n5751;
  assign n5753 = n5752 ^ n5742;
  assign n5754 = n5738 & ~n5753;
  assign n5755 = ~n2772 & n4160;
  assign n5756 = n5755 ^ n4154;
  assign n5757 = n3274 & n5756;
  assign n5758 = n5757 ^ n4154;
  assign n5759 = n5754 & ~n5758;
  assign n5760 = ~n4129 & n5759;
  assign n5761 = ~n4151 & n5760;
  assign n5762 = ~n5728 & n5761;
  assign n5763 = ~n4109 & n5762;
  assign n5764 = ~n5726 & n5763;
  assign n5765 = n5764 ^ n1481;
  assign n7261 = n5765 ^ x280;
  assign n7262 = ~n7260 & n7261;
  assign n7263 = n7262 ^ n7261;
  assign n7264 = n7263 ^ n7260;
  assign n7265 = ~n7259 & n7264;
  assign n7307 = n7245 & n7263;
  assign n7273 = n7253 ^ n7233;
  assign n7269 = n7225 & ~n7233;
  assign n7270 = n7269 ^ n7244;
  assign n7271 = n7270 ^ n7234;
  assign n7268 = n7258 ^ n7252;
  assign n7272 = n7271 ^ n7268;
  assign n7274 = n7273 ^ n7272;
  assign n7275 = n7262 & ~n7274;
  assign n7266 = n7262 ^ n7260;
  assign n7267 = n7258 & ~n7266;
  assign n7276 = n7275 ^ n7267;
  assign n7573 = ~n7255 & n7260;
  assign n7570 = n7274 ^ n7244;
  assign n7571 = ~n7260 & ~n7570;
  assign n7572 = n7571 ^ n7274;
  assign n7574 = n7573 ^ n7572;
  assign n7575 = n7261 & ~n7574;
  assign n7576 = n7575 ^ n7572;
  assign n7277 = n7227 ^ n7188;
  assign n7278 = n7277 ^ n7237;
  assign n7291 = n7260 & n7278;
  assign n7289 = n7237 & ~n7260;
  assign n7290 = n7289 ^ n7231;
  assign n7292 = n7291 ^ n7290;
  assign n7293 = ~n7261 & n7292;
  assign n7294 = n7293 ^ n7290;
  assign n7577 = n7234 ^ n7227;
  assign n7578 = ~n7260 & n7577;
  assign n7579 = n7578 ^ n7234;
  assign n7580 = n7261 & n7579;
  assign n7581 = ~n7250 & ~n7266;
  assign n7279 = n7266 ^ n7263;
  assign n7583 = n7234 ^ n7230;
  assign n7584 = n7583 ^ n7252;
  assign n7582 = n7269 ^ n7236;
  assign n7585 = n7584 ^ n7582;
  assign n7586 = n7585 ^ n7582;
  assign n7587 = ~n7261 & n7586;
  assign n7588 = n7587 ^ n7582;
  assign n7589 = n7279 & n7588;
  assign n7590 = n7589 ^ n7582;
  assign n7591 = ~n7581 & ~n7590;
  assign n7592 = n7268 ^ n7245;
  assign n7593 = n7592 ^ n7241;
  assign n7594 = ~n7260 & n7593;
  assign n7595 = n7594 ^ n7241;
  assign n7596 = n7261 & n7595;
  assign n7597 = n7591 & ~n7596;
  assign n7598 = ~n7580 & n7597;
  assign n7599 = ~n7294 & n7598;
  assign n7600 = n7576 & n7599;
  assign n7601 = ~n7276 & n7600;
  assign n7602 = ~n7307 & n7601;
  assign n7603 = ~n7265 & n7602;
  assign n7604 = n7603 ^ n5172;
  assign n7605 = n7604 ^ x307;
  assign n5667 = ~n5585 & n5666;
  assign n5668 = n5667 ^ n5665;
  assign n5669 = n5584 & n5668;
  assign n5671 = n5670 ^ n5642;
  assign n5675 = n5674 ^ n5671;
  assign n5676 = n5584 & n5675;
  assign n5677 = n5676 ^ n5671;
  assign n5678 = ~n5585 & n5677;
  assign n5679 = ~n5669 & ~n5678;
  assign n5680 = ~n5663 & n5679;
  assign n5681 = n5658 & ~n5660;
  assign n5691 = n5690 ^ n5681;
  assign n5697 = n5696 ^ n5662;
  assign n5700 = n5699 ^ n5660;
  assign n5701 = ~n5696 & n5700;
  assign n5702 = n5701 ^ n5660;
  assign n5703 = ~n5697 & ~n5702;
  assign n5704 = n5703 ^ n5662;
  assign n5710 = ~n5659 & ~n5672;
  assign n5711 = n5674 & ~n5710;
  assign n5709 = n5705 ^ n5641;
  assign n5712 = n5711 ^ n5709;
  assign n5708 = n5707 ^ n5665;
  assign n5713 = n5712 ^ n5708;
  assign n5714 = n5713 ^ n5708;
  assign n5715 = n5662 & n5714;
  assign n5716 = n5715 ^ n5708;
  assign n5717 = n5660 & n5716;
  assign n5718 = n5717 ^ n5708;
  assign n5719 = n5704 & ~n5718;
  assign n5720 = ~n5695 & n5719;
  assign n5721 = ~n5691 & n5720;
  assign n5722 = n5680 & n5721;
  assign n5723 = ~n5656 & n5722;
  assign n5724 = n5723 ^ n3966;
  assign n5725 = n5724 ^ x275;
  assign n5766 = n5765 ^ x278;
  assign n5770 = ~n4708 & n4868;
  assign n5771 = n5770 ^ n4863;
  assign n5772 = n4728 & n5771;
  assign n5777 = n4883 ^ n4873;
  assign n5778 = n4895 & n5777;
  assign n5784 = n4855 ^ n4846;
  assign n5785 = n5784 ^ n4864;
  assign n5786 = n5785 ^ n4852;
  assign n5787 = n5786 ^ n4898;
  assign n5788 = n4708 & ~n5787;
  assign n5789 = n5788 ^ n4898;
  assign n5781 = n4871 ^ n4861;
  assign n5782 = ~n4708 & n5781;
  assign n5783 = n5782 ^ n4861;
  assign n5790 = n5789 ^ n5783;
  assign n5791 = n4728 & n5790;
  assign n5792 = n5791 ^ n5789;
  assign n5793 = ~n4878 & ~n5792;
  assign n5794 = ~n5780 & n5793;
  assign n5795 = ~n5778 & n5794;
  assign n5796 = n5784 ^ n4882;
  assign n5797 = n4708 & n5796;
  assign n5798 = n5797 ^ n5784;
  assign n5799 = n4889 & n5798;
  assign n5800 = n5795 & ~n5799;
  assign n5803 = n4842 & ~n4889;
  assign n5801 = n4874 ^ n4857;
  assign n5802 = ~n4901 & n5801;
  assign n5804 = n5803 ^ n5802;
  assign n5805 = n5800 & ~n5804;
  assign n5806 = ~n5776 & n5805;
  assign n5807 = ~n5772 & n5806;
  assign n5808 = n5807 ^ n3994;
  assign n5809 = n5808 ^ x277;
  assign n4310 = n4309 ^ x232;
  assign n4457 = n4456 ^ x237;
  assign n4654 = n4310 & ~n4457;
  assign n4655 = n4654 ^ n4457;
  assign n4556 = n4555 ^ x236;
  assign n4564 = n4563 ^ n3209;
  assign n4565 = ~n3199 & ~n4564;
  assign n4566 = n3254 ^ n3194;
  assign n4567 = n3221 & n4566;
  assign n4578 = n3229 ^ n3201;
  assign n4577 = n3243 ^ n3231;
  assign n4579 = n4578 ^ n4577;
  assign n4580 = ~n2846 & ~n4579;
  assign n4581 = n4580 ^ n4577;
  assign n4572 = n3250 ^ n3223;
  assign n4573 = n4572 ^ n3216;
  assign n4574 = n4573 ^ n3227;
  assign n4575 = ~n2846 & n4574;
  assign n4576 = n4575 ^ n3227;
  assign n4582 = n4581 ^ n4576;
  assign n4583 = n2809 & n4582;
  assign n4584 = n4583 ^ n4576;
  assign n4585 = ~n3232 & ~n4584;
  assign n4586 = ~n3234 & n4585;
  assign n4587 = ~n4571 & n4586;
  assign n4588 = ~n4567 & n4587;
  assign n4589 = ~n4565 & n4588;
  assign n4590 = n3229 ^ n3195;
  assign n4591 = n2846 & ~n4590;
  assign n4592 = n4591 ^ n3195;
  assign n4593 = n2809 & n4592;
  assign n4594 = n4589 & ~n4593;
  assign n4595 = ~n4562 & n4594;
  assign n4596 = ~n4560 & n4595;
  assign n4597 = ~n3225 & n4596;
  assign n4598 = n4597 ^ n3088;
  assign n4599 = n4598 ^ x234;
  assign n4600 = ~n4556 & n4599;
  assign n4601 = n4600 ^ n4599;
  assign n4602 = n4601 ^ n4556;
  assign n4480 = n4479 ^ n3666;
  assign n4478 = n3688 ^ n3661;
  assign n4481 = n4480 ^ n4478;
  assign n4482 = n3542 & ~n4481;
  assign n4483 = n4482 ^ n4478;
  assign n4474 = n4473 ^ n3674;
  assign n4472 = n4471 ^ n3644;
  assign n4475 = n4474 ^ n4472;
  assign n4476 = n3542 & n4475;
  assign n4477 = n4476 ^ n4472;
  assign n4484 = n4483 ^ n4477;
  assign n4485 = ~n3679 & n4484;
  assign n4486 = n4485 ^ n4483;
  assign n4487 = ~n3687 & ~n4486;
  assign n4488 = ~n4468 & n4487;
  assign n4489 = ~n4463 & n4488;
  assign n4490 = ~n3678 & n4489;
  assign n4491 = ~n3639 & n4490;
  assign n4492 = n4491 ^ n3067;
  assign n4493 = n4492 ^ x235;
  assign n4544 = n4543 ^ x233;
  assign n4545 = n4493 & n4544;
  assign n4604 = n4545 ^ n4493;
  assign n4605 = n4604 ^ n4544;
  assign n4606 = n4605 ^ n4493;
  assign n4656 = n4602 & n4606;
  assign n4620 = n4601 & n4606;
  assign n4669 = n4656 ^ n4620;
  assign n4670 = n4669 ^ n4606;
  assign n4607 = n4600 & n4606;
  assign n4671 = n4670 ^ n4607;
  assign n4675 = ~n4655 & n4671;
  assign n4617 = n4600 & ~n4605;
  assign n4616 = n4602 & ~n4605;
  assign n4618 = n4617 ^ n4616;
  assign n5812 = n4618 & n4654;
  assign n4458 = n4457 ^ n4310;
  assign n4628 = n4617 ^ n4600;
  assign n4603 = n4545 & n4602;
  assign n4625 = n4603 ^ n4545;
  assign n4609 = n4601 & n4604;
  assign n4621 = n4620 ^ n4609;
  assign n4622 = n4621 ^ n4601;
  assign n4612 = n4600 ^ n4556;
  assign n4614 = ~n4605 & ~n4612;
  assign n4615 = n4614 ^ n4605;
  assign n4619 = n4618 ^ n4615;
  assign n4623 = n4622 ^ n4619;
  assign n4613 = n4545 & ~n4612;
  assign n4624 = n4623 ^ n4613;
  assign n4626 = n4625 ^ n4624;
  assign n4627 = n4626 ^ n4607;
  assign n4629 = n4628 ^ n4627;
  assign n4611 = n4602 & n4604;
  assign n4630 = n4629 ^ n4611;
  assign n4642 = n4630 ^ n4614;
  assign n4643 = n4310 & ~n4642;
  assign n4644 = n4643 ^ n4614;
  assign n4645 = ~n4458 & n4644;
  assign n5813 = n5812 ^ n4645;
  assign n4610 = n4609 ^ n4604;
  assign n4631 = n4630 ^ n4610;
  assign n4637 = n4631 ^ n4616;
  assign n4638 = n4637 ^ n4624;
  assign n4639 = n4457 & n4638;
  assign n4640 = n4639 ^ n4624;
  assign n4641 = ~n4310 & ~n4640;
  assign n5814 = ~n4457 & n4620;
  assign n4667 = n4629 ^ n4619;
  assign n5815 = n4667 ^ n4611;
  assign n5816 = ~n4655 & n5815;
  assign n5817 = ~n5814 & ~n5816;
  assign n4672 = n4671 ^ n4656;
  assign n5825 = n4672 ^ n4607;
  assign n5826 = n5825 ^ n4623;
  assign n4632 = n4631 ^ n4617;
  assign n5827 = n5826 ^ n4632;
  assign n4657 = n4656 ^ n4609;
  assign n4658 = n4657 ^ n4617;
  assign n5820 = n4658 ^ n4619;
  assign n4666 = n4626 ^ n4603;
  assign n5821 = n5820 ^ n4666;
  assign n5818 = n4666 ^ n4613;
  assign n5819 = n5818 ^ n4657;
  assign n5822 = n5821 ^ n5819;
  assign n5823 = ~n4310 & ~n5822;
  assign n5824 = n5823 ^ n5819;
  assign n5828 = n5827 ^ n5824;
  assign n5829 = n5828 ^ n5824;
  assign n5830 = n4310 & n5829;
  assign n5831 = n5830 ^ n5824;
  assign n5832 = ~n4458 & ~n5831;
  assign n5833 = n5832 ^ n5824;
  assign n5834 = n5817 & n5833;
  assign n5835 = ~n4641 & n5834;
  assign n5836 = ~n5813 & n5835;
  assign n5837 = ~n4675 & n5836;
  assign n5838 = n5837 ^ n4016;
  assign n5839 = n5838 ^ x276;
  assign n5841 = ~n5809 & ~n5839;
  assign n5842 = ~n5766 & n5841;
  assign n5840 = n5839 ^ n5809;
  assign n5843 = n5842 ^ n5840;
  assign n5844 = ~n5725 & ~n5843;
  assign n5866 = n5766 & n5839;
  assign n5870 = n5866 ^ n5841;
  assign n5871 = n5870 ^ n5809;
  assign n5768 = n5766 ^ n5725;
  assign n5848 = n5839 ^ n5766;
  assign n5849 = n5848 ^ n5725;
  assign n5850 = ~n5768 & ~n5849;
  assign n5851 = n5850 ^ n5766;
  assign n5858 = ~n5809 & ~n5851;
  assign n5859 = n5725 & n5858;
  assign n5860 = n5859 ^ n5858;
  assign n5872 = n5871 ^ n5860;
  assign n5873 = ~n5844 & n5872;
  assign n5845 = n5844 ^ n5725;
  assign n5881 = n5873 ^ n5845;
  assign n5882 = n5881 ^ n5725;
  assign n5767 = ~n5725 & ~n5766;
  assign n5853 = n5767 & n5809;
  assign n5854 = n5853 ^ n5809;
  assign n5810 = n5725 & n5809;
  assign n5855 = n5854 ^ n5810;
  assign n5883 = n5882 ^ n5855;
  assign n5875 = n5810 ^ n5725;
  assign n5876 = n5875 ^ n5859;
  assign n5867 = n5866 ^ n5809;
  assign n5868 = n5867 ^ n5843;
  assign n5869 = n5868 ^ n5766;
  assign n5874 = n5873 ^ n5869;
  assign n5877 = n5876 ^ n5874;
  assign n5865 = n5858 ^ n5849;
  assign n5878 = n5877 ^ n5865;
  assign n5879 = n5878 ^ n5855;
  assign n5884 = n5883 ^ n5879;
  assign n5769 = n5768 ^ n5767;
  assign n5811 = n5810 ^ n5769;
  assign n5846 = n5845 ^ n5811;
  assign n5847 = n5846 ^ n5843;
  assign n5852 = n5851 ^ n5847;
  assign n5856 = n5855 ^ n5852;
  assign n5862 = n5859 ^ n5856;
  assign n5861 = n5860 ^ n5846;
  assign n5863 = n5862 ^ n5861;
  assign n5864 = n5863 ^ n5766;
  assign n5880 = n5879 ^ n5864;
  assign n5885 = n5884 ^ n5880;
  assign n5857 = n5856 ^ n5839;
  assign n5886 = n5885 ^ n5857;
  assign n5887 = n5886 ^ n5860;
  assign n5954 = n5953 ^ x279;
  assign n4926 = n4838 ^ x249;
  assign n4962 = n4961 ^ x244;
  assign n4963 = ~n4926 & n4962;
  assign n4964 = n4963 ^ n4926;
  assign n4965 = n4964 ^ n4962;
  assign n4966 = n4965 ^ n4963;
  assign n4967 = n4717 ^ n4713;
  assign n4968 = n4967 ^ n4714;
  assign n4969 = n4968 ^ n4547;
  assign n4970 = ~n3918 & ~n4969;
  assign n4971 = n4970 ^ n4547;
  assign n4972 = n4971 ^ n2886;
  assign n4973 = n4972 ^ x246;
  assign n4974 = n4707 ^ x248;
  assign n4975 = ~n4973 & n4974;
  assign n4976 = n4975 ^ n4974;
  assign n5019 = n5018 ^ x245;
  assign n5025 = n4411 ^ n4379;
  assign n5026 = n5025 ^ n4387;
  assign n5027 = ~n4426 & ~n5026;
  assign n5033 = n4414 ^ n4311;
  assign n5034 = ~n5032 & n5033;
  assign n5035 = n5034 ^ n5031;
  assign n5036 = n5035 ^ n4311;
  assign n5037 = n5036 ^ n5029;
  assign n5038 = ~n4313 & ~n5037;
  assign n5039 = ~n5027 & ~n5038;
  assign n5040 = n4405 ^ n4388;
  assign n5041 = n4425 & n5040;
  assign n5042 = n4372 ^ n4367;
  assign n5043 = n5042 ^ n4420;
  assign n5044 = n4311 & n5043;
  assign n5045 = n5044 ^ n4420;
  assign n5046 = n4313 & n5045;
  assign n5047 = n5046 ^ n4420;
  assign n5048 = ~n5041 & ~n5047;
  assign n5049 = n5039 & n5048;
  assign n5050 = ~n5024 & n5049;
  assign n5051 = ~n4432 & n5050;
  assign n5052 = ~n4399 & n5051;
  assign n5053 = n5052 ^ n2916;
  assign n5054 = n5053 ^ x247;
  assign n5055 = n5019 & ~n5054;
  assign n5088 = n4976 & n5055;
  assign n5093 = n5088 ^ n5055;
  assign n4977 = n4976 ^ n4973;
  assign n5056 = n5055 ^ n5019;
  assign n5068 = n4977 & n5056;
  assign n5089 = n5088 ^ n5068;
  assign n5081 = n5019 ^ n4974;
  assign n5082 = n4973 & n5081;
  assign n5083 = n5082 ^ n5019;
  assign n5079 = n5054 ^ n5019;
  assign n5084 = n5079 ^ n4973;
  assign n5085 = ~n5083 & ~n5084;
  assign n5067 = n4977 & n5055;
  assign n5069 = n5068 ^ n5067;
  assign n5086 = n5085 ^ n5069;
  assign n5080 = n5079 ^ n4974;
  assign n5087 = n5086 ^ n5080;
  assign n5090 = n5089 ^ n5087;
  assign n4978 = n4977 ^ n4974;
  assign n5076 = ~n4978 & n5056;
  assign n5059 = n4974 ^ n4973;
  assign n5062 = ~n5019 & n5059;
  assign n5077 = n5076 ^ n5062;
  assign n5057 = n5056 ^ n5054;
  assign n5060 = n5057 ^ n5019;
  assign n5064 = n4975 & ~n5060;
  assign n5061 = n5059 & ~n5060;
  assign n5065 = n5064 ^ n5061;
  assign n5066 = n5065 ^ n4977;
  assign n5070 = n5069 ^ n5066;
  assign n5073 = n5070 ^ n5057;
  assign n5063 = n5062 ^ n5061;
  assign n5071 = n5070 ^ n5063;
  assign n5058 = ~n4978 & n5057;
  assign n5072 = n5071 ^ n5058;
  assign n5074 = n5073 ^ n5072;
  assign n5075 = n5074 ^ n5068;
  assign n5078 = n5077 ^ n5075;
  assign n5091 = n5090 ^ n5078;
  assign n5092 = n5091 ^ n5067;
  assign n5094 = n5093 ^ n5092;
  assign n5095 = ~n4966 & ~n5094;
  assign n5890 = n5092 ^ n5089;
  assign n5891 = ~n4962 & ~n5890;
  assign n5892 = n5891 ^ n5089;
  assign n5893 = n4926 & n5892;
  assign n5888 = n5070 ^ n5064;
  assign n5889 = n4965 & n5888;
  assign n5894 = n5893 ^ n5889;
  assign n5895 = n5082 ^ n5067;
  assign n5896 = n5895 ^ n5075;
  assign n5897 = n5896 ^ n5058;
  assign n5898 = ~n4962 & n5897;
  assign n5901 = n5888 ^ n5088;
  assign n5101 = n5056 & ~n5059;
  assign n5902 = n5901 ^ n5101;
  assign n5903 = n5902 ^ n5087;
  assign n5904 = n4962 & n5903;
  assign n5905 = n5904 ^ n5902;
  assign n5899 = n4962 & n5078;
  assign n5900 = n5899 ^ n5075;
  assign n5906 = n5905 ^ n5900;
  assign n5907 = ~n4926 & n5906;
  assign n5908 = n5907 ^ n5900;
  assign n5909 = ~n5898 & ~n5908;
  assign n5910 = ~n5894 & n5909;
  assign n5911 = ~n5095 & n5910;
  assign n5912 = n5911 ^ n3936;
  assign n5913 = n5912 ^ x274;
  assign n5955 = n5954 ^ n5913;
  assign n5961 = n5860 ^ n5844;
  assign n5962 = n5961 ^ n5768;
  assign n5963 = n5962 ^ n5878;
  assign n5958 = n5868 ^ n5839;
  assign n5959 = ~n5725 & n5958;
  assign n5960 = n5884 & ~n5959;
  assign n5964 = n5963 ^ n5960;
  assign n5965 = n5954 & ~n5964;
  assign n5966 = n5965 ^ n5963;
  assign n5956 = ~n5885 & ~n5954;
  assign n5957 = n5956 ^ n5884;
  assign n5967 = n5966 ^ n5957;
  assign n5968 = ~n5955 & n5967;
  assign n5969 = n5968 ^ n5966;
  assign n5970 = ~n5887 & n5969;
  assign n5971 = n5970 ^ n4727;
  assign n7606 = n5971 ^ x305;
  assign n7607 = n7605 & ~n7606;
  assign n7608 = n7607 ^ n7605;
  assign n7609 = n7608 ^ n7606;
  assign n6739 = n6738 ^ x286;
  assign n6258 = ~n4457 & n4611;
  assign n6259 = n4656 ^ n4631;
  assign n6260 = ~n4655 & ~n6259;
  assign n6261 = ~n6258 & ~n6260;
  assign n4661 = n4654 ^ n4310;
  assign n6262 = n4619 ^ n4614;
  assign n6263 = n4661 & ~n6262;
  assign n6264 = ~n4457 & n4621;
  assign n6265 = n6264 ^ n4609;
  assign n6266 = ~n4310 & n6265;
  assign n6270 = n4671 ^ n4624;
  assign n6271 = n6270 ^ n4603;
  assign n6269 = n4667 ^ n4631;
  assign n6272 = n6271 ^ n6269;
  assign n6273 = ~n4457 & n6272;
  assign n6274 = n6273 ^ n6269;
  assign n6267 = n4310 & n4545;
  assign n6268 = n6267 ^ n4627;
  assign n6275 = n6274 ^ n6268;
  assign n6276 = n4458 & n6275;
  assign n6277 = n6276 ^ n6268;
  assign n6278 = ~n6266 & n6277;
  assign n6279 = ~n4675 & n6278;
  assign n6280 = ~n6263 & n6279;
  assign n6281 = n6261 & n6280;
  assign n6282 = n5826 ^ n4629;
  assign n6283 = ~n4310 & n6282;
  assign n6284 = n6283 ^ n4629;
  assign n6285 = n4458 & ~n6284;
  assign n6286 = n6281 & ~n6285;
  assign n6287 = ~n5813 & n6286;
  assign n6288 = n6287 ^ n3540;
  assign n6740 = n6288 ^ x291;
  assign n6778 = n4965 & n5072;
  assign n6779 = ~n4964 & n5061;
  assign n5109 = ~n4966 & n5056;
  assign n5110 = n4975 & n5109;
  assign n6780 = n6779 ^ n5110;
  assign n6781 = n5897 ^ n5070;
  assign n6782 = n6781 ^ n5085;
  assign n6783 = n4926 & n6782;
  assign n6784 = n6783 ^ n6781;
  assign n6785 = n4962 & n6784;
  assign n6788 = ~n4963 & ~n4976;
  assign n5096 = n4965 & n5088;
  assign n6790 = n5101 ^ n5096;
  assign n6789 = n5094 ^ n5091;
  assign n6791 = n6790 ^ n6789;
  assign n6792 = ~n6788 & n6791;
  assign n6786 = n5089 ^ n5072;
  assign n6787 = ~n4962 & n6786;
  assign n6793 = n6792 ^ n6787;
  assign n6794 = ~n4966 & n6793;
  assign n6795 = n6794 ^ n6792;
  assign n6796 = ~n6785 & ~n6795;
  assign n6797 = ~n5893 & n6796;
  assign n6798 = ~n6780 & n6797;
  assign n6799 = ~n6778 & n6798;
  assign n6801 = n4964 & n5074;
  assign n6800 = ~n4962 & ~n5094;
  assign n6802 = n6801 ^ n6800;
  assign n6803 = n6799 & ~n6802;
  assign n6804 = n6803 ^ n3606;
  assign n6805 = n6804 ^ x288;
  assign n6831 = n6830 ^ x287;
  assign n6832 = ~n6805 & ~n6831;
  assign n6833 = n6832 ^ n6831;
  assign n6834 = n6833 ^ n6805;
  assign n6746 = n5256 ^ n5254;
  assign n5324 = n5323 ^ n5258;
  assign n6747 = n6746 ^ n5324;
  assign n6748 = ~n5298 & ~n6747;
  assign n6749 = n6748 ^ n6746;
  assign n6742 = n5238 ^ n5234;
  assign n6743 = n6742 ^ n5256;
  assign n6744 = ~n5298 & ~n6743;
  assign n6745 = n6744 ^ n5256;
  assign n6750 = n6749 ^ n6745;
  assign n6751 = ~n5297 & n6750;
  assign n6752 = n6751 ^ n6745;
  assign n6763 = n5298 & ~n5334;
  assign n6755 = n5927 ^ n5268;
  assign n6753 = n5264 ^ n5243;
  assign n6754 = n6753 ^ n5242;
  assign n6756 = n6755 ^ n6754;
  assign n6757 = n6755 ^ n5298;
  assign n6758 = n5303 & n6757;
  assign n6759 = n6758 ^ n5298;
  assign n6760 = ~n6756 & ~n6759;
  assign n6761 = n6760 ^ n6754;
  assign n6762 = ~n5254 & n6761;
  assign n6764 = n6763 ^ n6762;
  assign n6765 = n6764 ^ n6762;
  assign n6766 = ~n5252 & ~n6765;
  assign n6767 = n6766 ^ n6762;
  assign n6768 = n5303 & n6767;
  assign n6769 = n6768 ^ n6762;
  assign n6770 = n6752 & n6769;
  assign n6771 = n5922 & n6770;
  assign n6772 = ~n5314 & n6771;
  assign n6773 = n6772 ^ n3576;
  assign n6774 = n6773 ^ x289;
  assign n4136 = n4135 ^ n4108;
  assign n4137 = ~n2772 & n4136;
  assign n4138 = n4137 ^ n4108;
  assign n4139 = n3274 & n4138;
  assign n4133 = n3275 & n4132;
  assign n4140 = n4139 ^ n4133;
  assign n6016 = ~n2772 & n4143;
  assign n6017 = n6016 ^ n4104;
  assign n6013 = n4172 ^ n4106;
  assign n6014 = ~n2772 & n6013;
  assign n6015 = n6014 ^ n4172;
  assign n6018 = n6017 ^ n6015;
  assign n6019 = n3274 & n6018;
  assign n6020 = n6019 ^ n6017;
  assign n6036 = n4132 ^ n4121;
  assign n6037 = ~n3274 & n6036;
  assign n6034 = n3276 & n4135;
  assign n4118 = n4110 & ~n4117;
  assign n4130 = n4129 ^ n4118;
  assign n6035 = n6034 ^ n4130;
  assign n6038 = n6037 ^ n6035;
  assign n6026 = n4143 ^ n4123;
  assign n6027 = ~n3274 & n6026;
  assign n6028 = n6027 ^ n4143;
  assign n6029 = n6028 ^ n4117;
  assign n6030 = n4141 & ~n6029;
  assign n6031 = n6030 ^ n4117;
  assign n6023 = n5739 ^ n4115;
  assign n6024 = ~n4141 & n6023;
  assign n6025 = n6024 ^ n4115;
  assign n6032 = n6031 ^ n6025;
  assign n6021 = n4106 & ~n4141;
  assign n6022 = n6021 ^ n5726;
  assign n6033 = n6032 ^ n6022;
  assign n6039 = n6038 ^ n6033;
  assign n6040 = ~n6020 & n6039;
  assign n6041 = ~n4140 & n6040;
  assign n6042 = n6041 ^ n3635;
  assign n6775 = n6042 ^ x290;
  assign n6776 = ~n6774 & ~n6775;
  assign n6777 = n6776 ^ n6775;
  assign n6836 = n6777 ^ n6774;
  assign n6840 = ~n6834 & ~n6836;
  assign n6837 = n6836 ^ n6775;
  assign n6838 = ~n6834 & ~n6837;
  assign n6835 = ~n6777 & ~n6834;
  assign n6839 = n6838 ^ n6835;
  assign n6841 = n6840 ^ n6839;
  assign n6842 = n6841 ^ n6834;
  assign n6892 = n6740 & ~n6842;
  assign n6843 = n6832 ^ n6805;
  assign n6844 = ~n6837 & ~n6843;
  assign n6870 = n6844 ^ n6843;
  assign n6868 = ~n6836 & ~n6843;
  assign n6849 = n6776 & ~n6843;
  assign n6869 = n6868 ^ n6849;
  assign n6871 = n6870 ^ n6869;
  assign n6888 = n6871 ^ n6838;
  assign n6854 = ~n6833 & ~n6837;
  assign n6852 = n6844 ^ n6838;
  assign n6853 = n6852 ^ n6837;
  assign n6855 = n6854 ^ n6853;
  assign n6846 = n6805 ^ n6775;
  assign n6847 = ~n6774 & n6846;
  assign n6845 = n6844 ^ n6842;
  assign n6848 = n6847 ^ n6845;
  assign n6872 = n6855 ^ n6848;
  assign n6851 = ~n6777 & ~n6833;
  assign n6856 = n6855 ^ n6851;
  assign n6857 = n6856 ^ n6849;
  assign n6858 = n6857 ^ n6854;
  assign n6859 = n6858 ^ n6833;
  assign n6850 = n6849 ^ n6848;
  assign n6860 = n6859 ^ n6850;
  assign n6873 = n6872 ^ n6860;
  assign n6874 = n6873 ^ n6844;
  assign n6889 = n6888 ^ n6874;
  assign n6890 = ~n6740 & n6889;
  assign n6891 = n6890 ^ n6888;
  assign n6893 = n6892 ^ n6891;
  assign n6894 = n6739 & ~n6893;
  assign n6895 = n6894 ^ n6891;
  assign n7610 = n6873 ^ n6839;
  assign n7611 = ~n6740 & ~n7610;
  assign n7612 = n7611 ^ n6873;
  assign n7613 = n6739 & ~n7612;
  assign n6877 = n6848 ^ n6844;
  assign n6875 = n6776 & n6832;
  assign n6861 = ~n6777 & n6832;
  assign n6862 = n6861 ^ n6860;
  assign n6876 = n6875 ^ n6862;
  assign n6878 = n6877 ^ n6876;
  assign n6879 = n6878 ^ n6832;
  assign n6880 = n6879 ^ n6874;
  assign n6881 = n6880 ^ n6871;
  assign n6882 = n6740 & n6881;
  assign n6883 = n6882 ^ n6871;
  assign n6884 = n6739 & ~n6883;
  assign n7614 = ~n6739 & ~n6842;
  assign n6885 = n6739 & n6740;
  assign n7615 = n6885 ^ n6740;
  assign n7616 = n7615 ^ n6739;
  assign n7617 = n6870 ^ n6836;
  assign n7618 = n7617 ^ n6860;
  assign n7619 = ~n7616 & ~n7618;
  assign n7620 = ~n7614 & ~n7619;
  assign n6741 = n6740 ^ n6739;
  assign n7629 = n6831 ^ n6805;
  assign n7630 = n7629 ^ n6774;
  assign n7631 = n6847 ^ n6775;
  assign n7632 = n7630 & ~n7631;
  assign n7633 = n6740 & n7632;
  assign n7621 = n6858 & ~n7615;
  assign n6863 = n6861 ^ n6854;
  assign n7622 = n6885 ^ n6739;
  assign n7623 = n6855 & ~n7622;
  assign n7624 = ~n6857 & ~n7623;
  assign n7625 = ~n6863 & ~n7624;
  assign n7626 = ~n6875 & n7625;
  assign n7627 = ~n7621 & ~n7626;
  assign n7628 = ~n6868 & ~n7627;
  assign n7634 = n7633 ^ n7628;
  assign n7635 = ~n6741 & ~n7634;
  assign n7636 = n7635 ^ n7628;
  assign n7637 = n7620 & n7636;
  assign n7638 = ~n6884 & n7637;
  assign n7639 = ~n7613 & n7638;
  assign n7640 = n6895 & n7639;
  assign n7641 = n7640 ^ n5230;
  assign n7642 = n7641 ^ x308;
  assign n5435 = n5354 ^ n5353;
  assign n5442 = n5441 ^ n5439;
  assign n5438 = n5437 ^ n5428;
  assign n5443 = n5442 ^ n5438;
  assign n5444 = ~n5354 & n5443;
  assign n5445 = n5444 ^ n5438;
  assign n5446 = n5435 & n5445;
  assign n5451 = ~n5353 & ~n5450;
  assign n5458 = n5457 ^ n5452;
  assign n5459 = ~n5435 & ~n5458;
  assign n5460 = ~n5451 & ~n5459;
  assign n5465 = n5464 ^ n5441;
  assign n5466 = n5461 & ~n5465;
  assign n5481 = n5471 ^ n5430;
  assign n5484 = n5483 ^ n5481;
  assign n5472 = n5471 ^ n5470;
  assign n5473 = n5472 ^ n5354;
  assign n5474 = ~n5435 & ~n5473;
  assign n5475 = n5474 ^ n5354;
  assign n5476 = n5463 & ~n5475;
  assign n5479 = n5478 ^ n5476;
  assign n5480 = ~n5467 & n5479;
  assign n5485 = n5484 ^ n5480;
  assign n5486 = n5485 ^ n5480;
  assign n5487 = ~n5354 & ~n5486;
  assign n5488 = n5487 ^ n5480;
  assign n5489 = ~n5435 & ~n5488;
  assign n5490 = n5489 ^ n5480;
  assign n5491 = ~n5466 & n5490;
  assign n5492 = n5460 & n5491;
  assign n5493 = n5354 & n5449;
  assign n5494 = n5493 ^ n5448;
  assign n5495 = n5435 & n5494;
  assign n5496 = n5492 & ~n5495;
  assign n5497 = ~n5446 & n5496;
  assign n5498 = ~n5434 & n5497;
  assign n5499 = n5498 ^ n2845;
  assign n5500 = n5499 ^ x262;
  assign n5313 = n5309 & n5312;
  assign n5315 = n5314 ^ n5313;
  assign n5317 = n5312 ^ n5242;
  assign n5318 = n5316 & n5317;
  assign n5319 = ~n5255 & n5303;
  assign n5320 = n5319 ^ n5256;
  assign n5338 = n5322 ^ n5242;
  assign n5337 = n5336 ^ n5243;
  assign n5339 = n5338 ^ n5337;
  assign n5340 = n5297 & ~n5339;
  assign n5341 = n5340 ^ n5337;
  assign n5328 = n5267 ^ n5247;
  assign n5329 = n5328 ^ n5254;
  assign n5327 = n5326 ^ n5324;
  assign n5330 = n5329 ^ n5327;
  assign n5331 = ~n5297 & ~n5330;
  assign n5332 = n5331 ^ n5327;
  assign n5342 = n5341 ^ n5332;
  assign n5343 = ~n5298 & ~n5342;
  assign n5344 = n5343 ^ n5341;
  assign n5345 = n5320 & ~n5344;
  assign n5346 = ~n5318 & n5345;
  assign n5347 = ~n5315 & n5346;
  assign n5348 = ~n5307 & n5347;
  assign n5349 = ~n5302 & n5348;
  assign n5350 = ~n5270 & n5349;
  assign n5351 = n5350 ^ n2808;
  assign n5352 = n5351 ^ x267;
  assign n5540 = n5500 ^ n5352;
  assign n4608 = n4607 ^ n4603;
  assign n4633 = n4632 ^ n4608;
  assign n4634 = n4310 & ~n4633;
  assign n4635 = n4634 ^ n4608;
  assign n4636 = n4458 & n4635;
  assign n4646 = n4624 ^ n4614;
  assign n4647 = n4646 ^ n4609;
  assign n4648 = n4647 ^ n4620;
  assign n4649 = n4648 ^ n4620;
  assign n4650 = n4457 & ~n4649;
  assign n4651 = n4650 ^ n4620;
  assign n4652 = n4458 & n4651;
  assign n4653 = n4652 ^ n4620;
  assign n4677 = ~n4458 & n4671;
  assign n4668 = n4667 ^ n4666;
  assign n4673 = n4672 ^ n4668;
  assign n4674 = n4654 & ~n4673;
  assign n4676 = n4675 ^ n4674;
  assign n4678 = n4677 ^ n4676;
  assign n4662 = n4618 ^ n4613;
  assign n4663 = n4662 ^ n4614;
  assign n4664 = n4661 & n4663;
  assign n4659 = n4658 ^ n4626;
  assign n4660 = ~n4655 & ~n4659;
  assign n4665 = n4664 ^ n4660;
  assign n4679 = n4678 ^ n4665;
  assign n4680 = ~n4653 & ~n4679;
  assign n4681 = ~n4645 & n4680;
  assign n4682 = ~n4641 & n4681;
  assign n4683 = ~n4636 & n4682;
  assign n4684 = n4683 ^ n3183;
  assign n4685 = n4684 ^ x266;
  assign n4890 = n4865 ^ n4863;
  assign n4891 = n4708 & n4890;
  assign n4892 = n4891 ^ n4863;
  assign n4893 = n4889 & n4892;
  assign n4900 = n4894 & n4899;
  assign n4902 = n4865 & ~n4901;
  assign n4910 = n4728 & ~n4854;
  assign n4905 = n4870 ^ n4854;
  assign n4906 = n4905 ^ n4883;
  assign n4903 = n4860 ^ n4852;
  assign n4904 = n4903 ^ n4856;
  assign n4907 = n4906 ^ n4904;
  assign n4908 = ~n4728 & n4907;
  assign n4909 = n4908 ^ n4904;
  assign n4911 = n4910 ^ n4909;
  assign n4912 = ~n4708 & ~n4911;
  assign n4913 = n4912 ^ n4909;
  assign n4915 = n4874 & ~n4901;
  assign n4914 = n4881 & ~n4889;
  assign n4916 = n4915 ^ n4914;
  assign n4917 = n4913 & ~n4916;
  assign n4918 = ~n4902 & n4917;
  assign n4919 = ~n4900 & n4918;
  assign n4920 = ~n4897 & n4919;
  assign n4921 = ~n4893 & n4920;
  assign n4922 = ~n4888 & n4921;
  assign n4923 = ~n4878 & n4922;
  assign n4924 = n4923 ^ n2880;
  assign n4925 = n4924 ^ x263;
  assign n5098 = n4965 & n5076;
  assign n5097 = n4964 & ~n5091;
  assign n5099 = n5098 ^ n5097;
  assign n5119 = n4965 ^ n4926;
  assign n5120 = n5068 & n5119;
  assign n5118 = n4966 & n5071;
  assign n5121 = n5120 ^ n5118;
  assign n5114 = n5061 ^ n5060;
  assign n5111 = n5110 ^ n5061;
  assign n5112 = n5111 ^ n5070;
  assign n5113 = n5112 ^ n5110;
  assign n5115 = n5114 ^ n5113;
  assign n5116 = n4966 & ~n5115;
  assign n5117 = n5116 ^ n5111;
  assign n5122 = n5121 ^ n5117;
  assign n5106 = n4963 & n5089;
  assign n5105 = ~n4966 & n5074;
  assign n5107 = n5106 ^ n5105;
  assign n5100 = n5067 ^ n5058;
  assign n5102 = n5101 ^ n5100;
  assign n5103 = ~n4964 & n5102;
  assign n5104 = n5103 ^ n5058;
  assign n5108 = n5107 ^ n5104;
  assign n5123 = n5122 ^ n5108;
  assign n5124 = ~n5099 & ~n5123;
  assign n5125 = ~n5096 & n5124;
  assign n5126 = ~n5095 & n5125;
  assign n5127 = n5126 ^ n3001;
  assign n5128 = n5127 ^ x265;
  assign n5129 = ~n4925 & ~n5128;
  assign n5130 = n5129 ^ n5128;
  assign n5507 = ~n4685 & ~n5130;
  assign n5560 = n5507 ^ n5130;
  assign n4145 = n3274 & n4144;
  assign n4146 = n4145 ^ n4132;
  assign n4147 = ~n4141 & n4146;
  assign n4155 = ~n4141 & n4154;
  assign n4157 = n4113 ^ n4104;
  assign n4158 = ~n4156 & n4157;
  assign n4159 = ~n4155 & ~n4158;
  assign n4162 = n4125 ^ n4112;
  assign n4161 = n4160 ^ n4106;
  assign n4163 = n4162 ^ n4161;
  assign n4164 = n4163 ^ n4161;
  assign n4165 = ~n2772 & n4164;
  assign n4166 = n4165 ^ n4161;
  assign n4167 = n3274 & n4166;
  assign n4168 = n4167 ^ n4161;
  assign n4169 = n4159 & ~n4168;
  assign n4173 = n4141 & n4172;
  assign n4170 = n2772 & n4123;
  assign n4174 = n4173 ^ n4170;
  assign n4175 = n4169 & ~n4174;
  assign n4176 = ~n4152 & n4175;
  assign n4177 = ~n4151 & n4176;
  assign n4178 = ~n4147 & n4177;
  assign n4179 = ~n4140 & n4178;
  assign n4180 = ~n4130 & n4179;
  assign n4181 = ~n4109 & n4180;
  assign n4182 = n4181 ^ n3042;
  assign n4183 = n4182 ^ x264;
  assign n5531 = n4685 & n5129;
  assign n5534 = ~n4183 & n5531;
  assign n5542 = n5534 ^ n5531;
  assign n5508 = ~n4183 & ~n4685;
  assign n5509 = n5508 ^ n4685;
  assign n5510 = ~n5130 & ~n5509;
  assign n5527 = n5510 ^ n4925;
  assign n5520 = n5128 ^ n4925;
  assign n5521 = n5520 ^ n4685;
  assign n5515 = n4685 ^ n4183;
  assign n5522 = ~n5128 & ~n5515;
  assign n5523 = n5522 ^ n4183;
  assign n5524 = n5521 & n5523;
  assign n5525 = n5524 ^ n4925;
  assign n5131 = n5130 ^ n4925;
  assign n5516 = ~n5131 & n5515;
  assign n5517 = n5516 ^ n5131;
  assign n5512 = ~n4925 & n5508;
  assign n5513 = n5512 ^ n5508;
  assign n5511 = n5510 ^ n5507;
  assign n5514 = n5513 ^ n5511;
  assign n5518 = n5517 ^ n5514;
  assign n5519 = n5518 ^ n5511;
  assign n5526 = n5525 ^ n5519;
  assign n5528 = n5527 ^ n5526;
  assign n5132 = n5131 ^ n5128;
  assign n5133 = n4685 & ~n5132;
  assign n5506 = n5133 ^ n5132;
  assign n5529 = n5528 ^ n5506;
  assign n5530 = n5529 ^ n5512;
  assign n5543 = n5542 ^ n5530;
  assign n5541 = n5522 ^ n5511;
  assign n5544 = n5543 ^ n5541;
  assign n5561 = n5560 ^ n5544;
  assign n7332 = n5561 ^ n5514;
  assign n7643 = n7332 ^ n5528;
  assign n7644 = n5500 & n7643;
  assign n7645 = n7644 ^ n5528;
  assign n7646 = n5540 & ~n7645;
  assign n5501 = ~n5352 & n5500;
  assign n5502 = n5501 ^ n5352;
  assign n7647 = ~n5502 & n5516;
  assign n7328 = n5543 ^ n5528;
  assign n7329 = n5352 & ~n7328;
  assign n7330 = n7329 ^ n5543;
  assign n7331 = n5500 & n7330;
  assign n5134 = n4183 & n5133;
  assign n7333 = n7332 ^ n5134;
  assign n7334 = ~n5352 & ~n7333;
  assign n7335 = n7334 ^ n7332;
  assign n7336 = n5540 & ~n7335;
  assign n7648 = n5544 ^ n5518;
  assign n5562 = n4685 & ~n5131;
  assign n7649 = n7648 ^ n5562;
  assign n7650 = ~n5500 & ~n7649;
  assign n7651 = n7650 ^ n5562;
  assign n7652 = n5352 & n7651;
  assign n7660 = ~n5352 & ~n5528;
  assign n5554 = n5134 ^ n5133;
  assign n5559 = n5554 ^ n5530;
  assign n7653 = n5559 ^ n5534;
  assign n7654 = n5502 & ~n7653;
  assign n7340 = n5529 ^ n5511;
  assign n7655 = n7340 ^ n5534;
  assign n5503 = n5502 ^ n5500;
  assign n5504 = n5503 ^ n5352;
  assign n7656 = n5504 ^ n5134;
  assign n5505 = n5134 & n5504;
  assign n7657 = n7656 ^ n5505;
  assign n7658 = ~n7655 & ~n7657;
  assign n7659 = ~n7654 & ~n7658;
  assign n7661 = n7660 ^ n7659;
  assign n7662 = n5540 & n7661;
  assign n7663 = n7662 ^ n7659;
  assign n7664 = ~n7652 & ~n7663;
  assign n7665 = ~n7336 & n7664;
  assign n7666 = ~n7331 & n7665;
  assign n5567 = n5544 ^ n5510;
  assign n7667 = ~n5540 & n5567;
  assign n7668 = n7666 & ~n7667;
  assign n7669 = ~n7647 & n7668;
  assign n7670 = n7655 ^ n5507;
  assign n7671 = n5352 & n7670;
  assign n7672 = n7671 ^ n5507;
  assign n7673 = n5540 & n7672;
  assign n7674 = n7669 & ~n7673;
  assign n7675 = ~n7646 & n7674;
  assign n7676 = n7675 ^ n5204;
  assign n7677 = n7676 ^ x306;
  assign n7678 = n7642 & n7677;
  assign n7725 = n7678 ^ n7677;
  assign n7726 = n7609 & n7725;
  assign n7688 = n7642 ^ n7605;
  assign n7689 = n7677 ^ n7605;
  assign n7690 = n7688 & n7689;
  assign n7703 = n7690 ^ n7678;
  assign n7680 = n7678 ^ n7642;
  assign n7681 = n7680 ^ n7677;
  assign n7684 = n7607 & ~n7681;
  assign n7683 = n7607 & n7678;
  assign n7685 = n7684 ^ n7683;
  assign n7682 = n7608 & ~n7681;
  assign n7686 = n7685 ^ n7682;
  assign n7704 = n7703 ^ n7686;
  assign n6167 = n6044 & ~n6076;
  assign n6168 = ~n6166 & n6167;
  assign n6171 = n6170 ^ n6168;
  assign n6048 = n6047 ^ n6044;
  assign n6131 = n6130 ^ n6119;
  assign n6132 = n6131 ^ n6049;
  assign n6163 = n6162 ^ n6132;
  assign n6164 = n6163 ^ n6156;
  assign n6165 = ~n6048 & n6164;
  assign n6172 = n6171 ^ n6165;
  assign n6435 = n6157 ^ n6045;
  assign n6433 = ~n6045 & n6160;
  assign n6434 = n6433 ^ n6159;
  assign n6436 = n6435 ^ n6434;
  assign n6437 = n6436 ^ n6159;
  assign n6438 = n6044 & n6437;
  assign n6448 = n6123 & ~n6137;
  assign n6449 = ~n6048 & n6448;
  assign n6440 = n6076 ^ n6049;
  assign n6441 = n6440 ^ n6109;
  assign n6442 = n6441 ^ n6136;
  assign n6446 = ~n6048 & ~n6442;
  assign n6447 = n6077 & n6446;
  assign n6450 = n6449 ^ n6447;
  assign n6439 = n6164 ^ n6131;
  assign n6443 = n6442 ^ n6439;
  assign n6444 = ~n6047 & n6443;
  assign n6445 = n6444 ^ n6442;
  assign n6451 = n6450 ^ n6445;
  assign n6452 = ~n6438 & ~n6451;
  assign n6453 = ~n6172 & n6452;
  assign n6454 = n6453 ^ n3306;
  assign n7479 = n6454 ^ x303;
  assign n6199 = n5687 ^ n5657;
  assign n6197 = n6196 ^ n5642;
  assign n6198 = n6197 ^ n5672;
  assign n6200 = n6199 ^ n6198;
  assign n6201 = ~n5661 & n6200;
  assign n6209 = n6208 ^ n5648;
  assign n6203 = n6202 ^ n5644;
  assign n6204 = n6203 ^ n5698;
  assign n6205 = n6204 ^ n6198;
  assign n6206 = n5585 & n6205;
  assign n6207 = n6206 ^ n6204;
  assign n6210 = n6209 ^ n6207;
  assign n6211 = n6210 ^ n6207;
  assign n6212 = ~n5585 & n6211;
  assign n6213 = n6212 ^ n6207;
  assign n6214 = n5584 & n6213;
  assign n6215 = n6214 ^ n6207;
  assign n6216 = ~n6201 & ~n6215;
  assign n6217 = ~n6193 & n6216;
  assign n6218 = ~n5691 & n6217;
  assign n6219 = n5680 & n6218;
  assign n6220 = n6219 ^ n3827;
  assign n7478 = n6220 ^ x298;
  assign n7483 = n7479 ^ n7478;
  assign n5974 = n5385 & n5424;
  assign n5975 = n5354 & n5974;
  assign n5976 = n5975 ^ n5441;
  assign n5977 = ~n5435 & n5976;
  assign n5978 = n5977 ^ n5441;
  assign n5982 = ~n5353 & n5428;
  assign n5981 = n5979 & ~n5980;
  assign n5983 = n5982 ^ n5981;
  assign n5984 = ~n5978 & ~n5983;
  assign n5988 = ~n5985 & n5987;
  assign n5989 = n5457 ^ n5448;
  assign n5990 = ~n5986 & ~n5989;
  assign n5991 = n5483 ^ n5456;
  assign n5992 = n5991 ^ n5450;
  assign n5993 = n5979 & n5992;
  assign n6000 = n5452 ^ n5448;
  assign n6001 = n6000 ^ n5430;
  assign n6002 = n6001 ^ n5437;
  assign n6003 = n5353 & n6002;
  assign n5995 = n5478 ^ n5450;
  assign n5994 = n5974 ^ n5426;
  assign n5996 = n5995 ^ n5994;
  assign n5997 = n5986 & ~n5996;
  assign n5998 = n5997 ^ n5994;
  assign n5999 = n5998 ^ n5353;
  assign n6004 = n6003 ^ n5999;
  assign n6005 = n5354 & n6004;
  assign n6006 = n6005 ^ n5999;
  assign n6007 = ~n5993 & ~n6006;
  assign n6008 = ~n5990 & n6007;
  assign n6009 = ~n5988 & n6008;
  assign n6010 = n5984 & n6009;
  assign n6011 = n6010 ^ n3760;
  assign n7419 = n6011 ^ x299;
  assign n7420 = n3276 & ~n4117;
  assign n7421 = n4121 & ~n4156;
  assign n7428 = n4125 ^ n4115;
  assign n7427 = n4135 ^ n4122;
  assign n7429 = n7428 ^ n7427;
  assign n7430 = n3274 & n7429;
  assign n7431 = n7430 ^ n7427;
  assign n7423 = n4172 ^ n4123;
  assign n7422 = n4154 ^ n4132;
  assign n7424 = n7423 ^ n7422;
  assign n7425 = n3274 & n7424;
  assign n7426 = n7425 ^ n7422;
  assign n7432 = n7431 ^ n7426;
  assign n7433 = n7432 ^ n7431;
  assign n7434 = ~n6028 & ~n7433;
  assign n7435 = n7434 ^ n7431;
  assign n7436 = n4141 & ~n7435;
  assign n7437 = n7436 ^ n7431;
  assign n7438 = ~n5726 & ~n7437;
  assign n7439 = ~n7421 & n7438;
  assign n7440 = ~n7420 & n7439;
  assign n7441 = n2772 & n4172;
  assign n7442 = n7441 ^ n6021;
  assign n7443 = n7440 & ~n7442;
  assign n7444 = ~n4139 & n7443;
  assign n7445 = ~n5728 & n7444;
  assign n7446 = ~n4147 & n7445;
  assign n7447 = ~n4109 & n7446;
  assign n7448 = ~n4104 & n7447;
  assign n7449 = n7448 ^ n4343;
  assign n7450 = n7449 ^ x300;
  assign n7451 = n7419 & ~n7450;
  assign n7452 = n7451 ^ n7419;
  assign n7453 = ~n5297 & ~n6749;
  assign n7459 = n5927 ^ n5322;
  assign n7458 = n5323 ^ n5261;
  assign n7460 = n7459 ^ n7458;
  assign n7461 = ~n5297 & ~n7460;
  assign n7462 = n7461 ^ n7458;
  assign n7454 = n5333 ^ n5265;
  assign n7455 = n7454 ^ n5310;
  assign n7456 = n5298 & n7455;
  assign n7457 = n7456 ^ n5310;
  assign n7463 = n7462 ^ n7457;
  assign n7464 = ~n5303 & n7463;
  assign n7465 = n7464 ^ n7462;
  assign n7466 = ~n5318 & ~n7465;
  assign n7467 = ~n5929 & n7466;
  assign n7468 = ~n5926 & n7467;
  assign n7469 = ~n5315 & n7468;
  assign n7470 = ~n7453 & n7469;
  assign n7471 = ~n5302 & n7470;
  assign n7472 = n7471 ^ n4364;
  assign n7473 = n7472 ^ x301;
  assign n6372 = ~n4964 & n5087;
  assign n6373 = n5114 ^ n5074;
  assign n6374 = n5119 & ~n6373;
  assign n6376 = n5076 ^ n4965;
  assign n6377 = n6376 ^ n5098;
  assign n6375 = n4965 & ~n5101;
  assign n6378 = n6377 ^ n6375;
  assign n6379 = n6378 ^ n5065;
  assign n6380 = n6379 ^ n5091;
  assign n6381 = n4926 & ~n6380;
  assign n6382 = ~n6374 & ~n6381;
  assign n6383 = ~n6372 & n6382;
  assign n6384 = n5902 ^ n5067;
  assign n6385 = n6384 ^ n5114;
  assign n6386 = n6385 ^ n5071;
  assign n6387 = n4962 & ~n6386;
  assign n6388 = n6387 ^ n5071;
  assign n6389 = n4966 & n6388;
  assign n6390 = n6383 & ~n6389;
  assign n6391 = ~n5894 & n6390;
  assign n6392 = n6391 ^ n3436;
  assign n7474 = n6392 ^ x302;
  assign n7475 = n7473 & ~n7474;
  assign n7476 = n7475 ^ n7474;
  assign n7486 = n7476 ^ n7473;
  assign n7498 = n7452 & n7486;
  assign n7477 = n7452 & ~n7476;
  assign n7499 = n7498 ^ n7477;
  assign n7496 = n7452 & n7475;
  assign n7497 = n7496 ^ n7452;
  assign n7500 = n7499 ^ n7497;
  assign n7492 = n7474 ^ n7450;
  assign n7493 = n7419 & ~n7492;
  assign n7494 = n7493 ^ n7492;
  assign n7484 = n7451 ^ n7450;
  assign n7489 = ~n7476 & ~n7484;
  assign n7487 = n7484 ^ n7419;
  assign n7488 = n7486 & n7487;
  assign n7490 = n7489 ^ n7488;
  assign n7485 = n7475 & ~n7484;
  assign n7491 = n7490 ^ n7485;
  assign n7495 = n7494 ^ n7491;
  assign n7501 = n7500 ^ n7495;
  assign n7502 = ~n7478 & ~n7501;
  assign n7503 = n7502 ^ n7495;
  assign n7504 = n7483 & ~n7503;
  assign n7480 = n7478 & n7479;
  assign n7481 = n7480 ^ n7479;
  assign n7482 = n7477 & n7481;
  assign n7505 = n7504 ^ n7482;
  assign n7506 = n7480 ^ n7478;
  assign n7507 = n7506 ^ n7479;
  assign n7526 = n7475 & n7487;
  assign n7527 = n7526 ^ n7488;
  assign n7525 = n7495 ^ n7487;
  assign n7528 = n7527 ^ n7525;
  assign n7520 = n7486 ^ n7474;
  assign n7510 = n7451 & n7475;
  assign n7511 = n7510 ^ n7500;
  assign n7517 = n7511 ^ n7477;
  assign n7518 = n7517 ^ n7419;
  assign n7513 = n7451 & n7486;
  assign n7509 = n7498 ^ n7493;
  assign n7512 = n7511 ^ n7509;
  assign n7514 = n7513 ^ n7512;
  assign n7515 = n7514 ^ n7498;
  assign n7516 = n7515 ^ n7496;
  assign n7519 = n7518 ^ n7516;
  assign n7521 = n7520 ^ n7519;
  assign n7522 = n7521 ^ n7501;
  assign n7523 = n7522 ^ n7491;
  assign n7508 = n7488 ^ n7484;
  assign n7524 = n7523 ^ n7508;
  assign n7529 = n7528 ^ n7524;
  assign n7530 = ~n7507 & ~n7529;
  assign n7531 = n7529 ^ n7495;
  assign n7532 = n7478 & n7531;
  assign n7533 = n7532 ^ n7495;
  assign n7534 = ~n7483 & ~n7533;
  assign n7536 = n7485 & n7506;
  assign n7535 = n7478 & n7489;
  assign n7537 = n7536 ^ n7535;
  assign n7538 = ~n7534 & ~n7537;
  assign n7539 = n7513 ^ n7510;
  assign n7540 = n7539 ^ n7522;
  assign n7541 = n7481 & ~n7540;
  assign n7542 = n7541 ^ n7522;
  assign n7543 = n7495 ^ n7489;
  assign n7544 = n7543 ^ n7499;
  assign n7545 = n7544 ^ n7499;
  assign n7546 = ~n7478 & ~n7545;
  assign n7547 = n7546 ^ n7499;
  assign n7548 = n7483 & n7547;
  assign n7549 = n7548 ^ n7499;
  assign n7554 = n7527 ^ n7511;
  assign n7555 = n7479 & n7554;
  assign n7556 = n7555 ^ n7511;
  assign n7550 = n7519 ^ n7496;
  assign n7551 = n7550 ^ n7516;
  assign n7552 = ~n7479 & n7551;
  assign n7553 = n7552 ^ n7550;
  assign n7557 = n7556 ^ n7553;
  assign n7558 = ~n7478 & n7557;
  assign n7559 = n7558 ^ n7553;
  assign n7560 = ~n7549 & ~n7559;
  assign n7561 = n7542 & n7560;
  assign n7562 = n7538 & n7561;
  assign n7563 = ~n7530 & n7562;
  assign n7564 = ~n7505 & n7563;
  assign n7565 = n7564 ^ n5296;
  assign n7566 = n7565 ^ x309;
  assign n6012 = n6011 ^ x297;
  assign n6043 = n6042 ^ x292;
  assign n6179 = n6163 ^ n6148;
  assign n6180 = ~n6045 & n6179;
  assign n6181 = n6180 ^ n6148;
  assign n6176 = n6175 ^ n6045;
  assign n6177 = n6176 ^ n6161;
  assign n6178 = n6177 ^ n6144;
  assign n6182 = n6181 ^ n6178;
  assign n6183 = n6173 & n6182;
  assign n6184 = n6183 ^ n6181;
  assign n6185 = ~n6172 & ~n6184;
  assign n6186 = n6185 ^ n3763;
  assign n6187 = n6186 ^ x294;
  assign n6221 = n6220 ^ x296;
  assign n6222 = n6187 & ~n6221;
  assign n6223 = n6222 ^ n6187;
  assign n6226 = n4895 & n5784;
  assign n6227 = n5785 ^ n4850;
  assign n6228 = ~n4901 & n6227;
  assign n6236 = n4903 ^ n4848;
  assign n6235 = n4862 ^ n4853;
  assign n6237 = n6236 ^ n6235;
  assign n6238 = n4728 & ~n6237;
  assign n6239 = n6238 ^ n6235;
  assign n6232 = n5801 ^ n4870;
  assign n6233 = n4728 & n6232;
  assign n6234 = n6233 ^ n4870;
  assign n6240 = n6239 ^ n6234;
  assign n6241 = n4708 & n6240;
  assign n6242 = n6241 ^ n6239;
  assign n6243 = ~n6231 & ~n6242;
  assign n6244 = ~n5772 & n6243;
  assign n6245 = ~n6230 & n6244;
  assign n6246 = ~n6228 & n6245;
  assign n6247 = ~n6226 & n6246;
  assign n6248 = n4884 ^ n4873;
  assign n6249 = n6248 ^ n4856;
  assign n6250 = n4708 & n6249;
  assign n6251 = n6250 ^ n6248;
  assign n6252 = n4889 & n6251;
  assign n6253 = n6247 & ~n6252;
  assign n6254 = ~n4893 & n6253;
  assign n6255 = ~n5780 & n6254;
  assign n6256 = n6255 ^ n3796;
  assign n6257 = n6256 ^ x295;
  assign n6289 = n6288 ^ x293;
  assign n6290 = ~n6257 & ~n6289;
  assign n6306 = n6290 ^ n6257;
  assign n6312 = n6223 & ~n6306;
  assign n6224 = n6223 ^ n6221;
  assign n6225 = n6224 ^ n6187;
  assign n6307 = ~n6225 & ~n6306;
  assign n6313 = n6312 ^ n6307;
  assign n6310 = n6222 & ~n6306;
  assign n6311 = n6310 ^ n6306;
  assign n6314 = n6313 ^ n6311;
  assign n6308 = n6307 ^ n6225;
  assign n6300 = n6187 & ~n6289;
  assign n6298 = n6222 & n6290;
  assign n6295 = n6224 & n6290;
  assign n6299 = n6298 ^ n6295;
  assign n6301 = n6300 ^ n6299;
  assign n6291 = n6290 ^ n6289;
  assign n6294 = n6222 & ~n6291;
  assign n6296 = n6295 ^ n6294;
  assign n6293 = n6223 & ~n6291;
  assign n6297 = n6296 ^ n6293;
  assign n6302 = n6301 ^ n6297;
  assign n6303 = n6302 ^ n6290;
  assign n6304 = n6303 ^ n6299;
  assign n6292 = ~n6225 & ~n6291;
  assign n6305 = n6304 ^ n6292;
  assign n6309 = n6308 ^ n6305;
  assign n6315 = n6314 ^ n6309;
  assign n6316 = n6315 ^ n6313;
  assign n6317 = ~n6043 & n6316;
  assign n6318 = n6317 ^ n6315;
  assign n6319 = n6012 & n6318;
  assign n6320 = n6043 & n6305;
  assign n6321 = n6320 ^ n6292;
  assign n6322 = n6012 & n6321;
  assign n6324 = n6294 ^ n6291;
  assign n6323 = n6293 ^ n6292;
  assign n6325 = n6324 ^ n6323;
  assign n6326 = n6043 ^ n6012;
  assign n6327 = n6012 & n6326;
  assign n6328 = n6327 ^ n6326;
  assign n6329 = n6328 ^ n6043;
  assign n6330 = ~n6325 & n6329;
  assign n6338 = n6314 ^ n6292;
  assign n6336 = n6304 ^ n6302;
  assign n6337 = n6336 ^ n6293;
  assign n6339 = n6338 ^ n6337;
  assign n6331 = n6310 ^ n6296;
  assign n6332 = n6331 ^ n6222;
  assign n6333 = n6332 ^ n6299;
  assign n6334 = n6333 ^ n6312;
  assign n6335 = n6334 ^ n6325;
  assign n6340 = n6339 ^ n6335;
  assign n6341 = n6327 ^ n6043;
  assign n6342 = ~n6340 & ~n6341;
  assign n6344 = n6292 ^ n6291;
  assign n6345 = n6344 ^ n6224;
  assign n6343 = n6314 ^ n6297;
  assign n6346 = n6345 ^ n6343;
  assign n6347 = n6346 ^ n6333;
  assign n6348 = n6347 ^ n6337;
  assign n6349 = n6348 ^ n6299;
  assign n6350 = n6349 ^ n6299;
  assign n6351 = n6012 & n6350;
  assign n6352 = n6351 ^ n6299;
  assign n6353 = ~n6043 & n6352;
  assign n6354 = n6353 ^ n6299;
  assign n6355 = ~n6342 & ~n6354;
  assign n6358 = n6300 ^ n6221;
  assign n6359 = n6257 ^ n6221;
  assign n6360 = n6358 & ~n6359;
  assign n6356 = n6289 ^ n6257;
  assign n6357 = n6356 ^ n6187;
  assign n6361 = n6360 ^ n6357;
  assign n6362 = n6361 ^ n6334;
  assign n6363 = ~n6012 & n6362;
  assign n6364 = n6363 ^ n6334;
  assign n6365 = n6043 & n6364;
  assign n6366 = n6355 & ~n6365;
  assign n6367 = ~n6330 & n6366;
  assign n6368 = ~n6322 & n6367;
  assign n6369 = ~n6319 & n6368;
  assign n6370 = n6369 ^ n4812;
  assign n7567 = n6370 ^ x304;
  assign n7568 = ~n7566 & n7567;
  assign n7569 = n7568 ^ n7567;
  assign n7746 = n7569 ^ n7566;
  assign n8783 = n7704 & n7746;
  assign n7693 = n7607 ^ n7606;
  assign n7696 = ~n7681 & ~n7693;
  assign n7695 = n7680 & ~n7693;
  assign n7697 = n7696 ^ n7695;
  assign n7713 = n7697 ^ n7685;
  assign n7714 = n7713 ^ n7606;
  assign n7701 = n7642 ^ n7606;
  assign n7708 = n7690 ^ n7605;
  assign n7709 = ~n7701 & n7708;
  assign n7702 = ~n7688 & ~n7701;
  assign n7705 = n7704 ^ n7702;
  assign n7691 = n7690 ^ n7683;
  assign n7679 = n7609 & n7678;
  assign n7687 = n7686 ^ n7679;
  assign n7692 = n7691 ^ n7687;
  assign n7694 = n7693 ^ n7692;
  assign n7698 = n7697 ^ n7694;
  assign n7700 = n7698 ^ n7696;
  assign n7706 = n7705 ^ n7700;
  assign n7707 = n7706 ^ n7679;
  assign n7710 = n7709 ^ n7707;
  assign n7711 = n7710 ^ n7704;
  assign n7699 = n7698 ^ n7692;
  assign n7712 = n7711 ^ n7699;
  assign n7715 = n7714 ^ n7712;
  assign n7742 = n7715 ^ n7695;
  assign n7743 = n7567 & ~n7742;
  assign n7744 = n7743 ^ n7695;
  assign n7745 = ~n7566 & n7744;
  assign n8784 = n8783 ^ n7745;
  assign n8785 = n7569 & n7682;
  assign n7718 = n7715 ^ n7696;
  assign n7719 = n7718 ^ n7704;
  assign n7720 = n7719 ^ n7684;
  assign n7717 = n7704 ^ n7682;
  assign n7721 = n7720 ^ n7717;
  assign n7716 = n7715 ^ n7681;
  assign n7722 = n7721 ^ n7716;
  assign n7723 = n7569 & ~n7722;
  assign n7738 = n7704 ^ n7692;
  assign n7739 = ~n7567 & n7738;
  assign n7740 = n7739 ^ n7704;
  assign n7741 = n7566 & n7740;
  assign n7767 = n7699 ^ n7695;
  assign n8786 = n7569 & ~n7767;
  assign n8792 = n7606 ^ n7605;
  assign n8793 = n8792 ^ n7642;
  assign n8794 = n8793 ^ n7721;
  assign n7730 = n7706 ^ n7608;
  assign n7731 = n7730 ^ n7717;
  assign n7764 = n7731 ^ n7679;
  assign n7765 = n7764 ^ n7722;
  assign n8787 = n7765 ^ n7715;
  assign n8788 = n8787 ^ n7682;
  assign n8789 = n8788 ^ n7713;
  assign n8790 = ~n7566 & ~n8789;
  assign n8791 = n8790 ^ n7713;
  assign n8795 = n8794 ^ n8791;
  assign n8796 = n8795 ^ n8791;
  assign n8797 = ~n7566 & n8796;
  assign n8798 = n8797 ^ n8791;
  assign n8799 = n7567 & n8798;
  assign n8800 = n8799 ^ n8791;
  assign n8801 = ~n8786 & ~n8800;
  assign n7763 = n7567 ^ n7566;
  assign n8802 = n7566 & ~n7706;
  assign n8803 = n8802 ^ n7711;
  assign n8804 = n7763 & ~n8803;
  assign n8805 = n8804 ^ n7711;
  assign n8806 = n8801 & n8805;
  assign n8807 = ~n7741 & n8806;
  assign n8808 = ~n7723 & n8807;
  assign n8809 = ~n8785 & n8808;
  assign n8810 = ~n8784 & n8809;
  assign n8811 = ~n7726 & n8810;
  assign n8812 = n8811 ^ n5351;
  assign n9064 = n8812 ^ x363;
  assign n7783 = ~n5863 & ~n5913;
  assign n7784 = n7783 ^ n5861;
  assign n7780 = ~n5878 & ~n5913;
  assign n7781 = n7780 ^ n5865;
  assign n7785 = n7784 ^ n7781;
  assign n7786 = ~n5954 & n7785;
  assign n7787 = n7786 ^ n7784;
  assign n7782 = n7781 ^ n5954;
  assign n7788 = n7787 ^ n7782;
  assign n7789 = n7788 ^ n7784;
  assign n7790 = n7789 ^ n4555;
  assign n7791 = n7790 ^ x334;
  assign n7280 = n7278 & ~n7279;
  assign n7281 = n7255 ^ n7246;
  assign n7282 = ~n7260 & ~n7281;
  assign n7283 = n7282 ^ n7255;
  assign n7284 = ~n7261 & ~n7283;
  assign n7285 = ~n7280 & ~n7284;
  assign n7792 = n7255 ^ n7248;
  assign n7793 = n7792 ^ n7269;
  assign n7311 = n7251 ^ n7238;
  assign n7794 = n7793 ^ n7311;
  assign n7795 = n7794 ^ n7235;
  assign n7796 = n7260 & n7795;
  assign n7797 = n7796 ^ n7235;
  assign n7798 = n7261 & n7797;
  assign n7805 = ~n7261 & n7272;
  assign n7800 = n7244 ^ n7242;
  assign n7801 = n7800 ^ n7251;
  assign n7799 = n7792 ^ n7245;
  assign n7802 = n7801 ^ n7799;
  assign n7803 = ~n7261 & n7802;
  assign n7804 = n7803 ^ n7799;
  assign n7806 = n7805 ^ n7804;
  assign n7807 = n7260 & n7806;
  assign n7808 = n7807 ^ n7804;
  assign n7809 = ~n7798 & ~n7808;
  assign n7811 = n7236 & ~n7261;
  assign n7810 = n7227 & ~n7279;
  assign n7812 = n7811 ^ n7810;
  assign n7813 = n7809 & ~n7812;
  assign n7814 = ~n7580 & n7813;
  assign n7815 = n7285 & n7814;
  assign n7816 = ~n7275 & n7815;
  assign n7817 = n7816 ^ n5018;
  assign n7818 = n7817 ^ x339;
  assign n7819 = n7791 & ~n7818;
  assign n7974 = n7819 ^ n7818;
  assign n7820 = n7819 ^ n7791;
  assign n7975 = n7974 ^ n7820;
  assign n6633 = n5912 ^ x272;
  assign n6638 = n6045 & n6439;
  assign n6639 = n6448 ^ n6150;
  assign n6640 = n6047 & n6639;
  assign n6641 = ~n6638 & ~n6640;
  assign n6642 = ~n6446 & n6641;
  assign n6643 = n6044 & n6434;
  assign n6644 = n6642 & ~n6643;
  assign n6645 = ~n6637 & n6644;
  assign n6646 = n6645 ^ n4222;
  assign n6647 = n6646 ^ x270;
  assign n6595 = n6000 ^ n5468;
  assign n6596 = n6595 ^ n5980;
  assign n6597 = n6596 ^ n5441;
  assign n6598 = n6597 ^ n5441;
  assign n6599 = n5354 & ~n6598;
  assign n6600 = n6599 ^ n5441;
  assign n6601 = n5353 & n6600;
  assign n6602 = n6601 ^ n5441;
  assign n6605 = n6604 ^ n5477;
  assign n6603 = n5456 ^ n5437;
  assign n6606 = n6605 ^ n6603;
  assign n6607 = n6606 ^ n6603;
  assign n6608 = ~n5979 & ~n6607;
  assign n6609 = n6608 ^ n6603;
  assign n6610 = ~n5987 & n6609;
  assign n6611 = n6610 ^ n6603;
  assign n6612 = ~n6602 & ~n6611;
  assign n6613 = n5452 & n5979;
  assign n6621 = n5985 ^ n5482;
  assign n6614 = n5482 ^ n5472;
  assign n6615 = ~n5987 & n6614;
  assign n6618 = n6604 ^ n5481;
  assign n6616 = n5482 ^ n5470;
  assign n6617 = n5979 & ~n6616;
  assign n6619 = n6618 ^ n6617;
  assign n6620 = ~n6615 & ~n6619;
  assign n6622 = n6621 ^ n6620;
  assign n6623 = n6622 ^ n6620;
  assign n6624 = ~n5354 & ~n6623;
  assign n6625 = n6624 ^ n6620;
  assign n6626 = ~n5435 & n6625;
  assign n6627 = n6626 ^ n6620;
  assign n6628 = ~n6613 & ~n6627;
  assign n6629 = n6612 & n6628;
  assign n6630 = ~n5446 & n6629;
  assign n6631 = n6630 ^ n4217;
  assign n6632 = n6631 ^ x271;
  assign n6665 = n6647 ^ n6632;
  assign n6666 = ~n6633 & n6665;
  assign n6648 = n5351 ^ x269;
  assign n6657 = ~n6633 & n6648;
  assign n6660 = ~n6632 & n6647;
  assign n6662 = n6657 & n6660;
  assign n6667 = n6666 ^ n6662;
  assign n6653 = n6633 & n6647;
  assign n6654 = n6632 & n6653;
  assign n6659 = n6654 ^ n6653;
  assign n6661 = n6660 ^ n6659;
  assign n6663 = n6662 ^ n6661;
  assign n6649 = n6632 & ~n6648;
  assign n6650 = ~n6647 & n6649;
  assign n6651 = ~n6633 & n6650;
  assign n6664 = n6663 ^ n6651;
  assign n6668 = n6667 ^ n6664;
  assign n6658 = n6632 & n6657;
  assign n6669 = n6668 ^ n6658;
  assign n6652 = n6651 ^ n6650;
  assign n6655 = n6654 ^ n6652;
  assign n6634 = n6633 ^ n6632;
  assign n6635 = n6632 & ~n6634;
  assign n6656 = n6655 ^ n6635;
  assign n6670 = n6669 ^ n6656;
  assign n6671 = n4684 ^ x268;
  assign n6672 = n5724 ^ x273;
  assign n6673 = n6671 & ~n6672;
  assign n6674 = n6673 ^ n6671;
  assign n6675 = n6674 ^ n6672;
  assign n6676 = n6670 & n6675;
  assign n6677 = n6672 ^ n6671;
  assign n6680 = n6648 & n6654;
  assign n6681 = n6680 ^ n6654;
  assign n6682 = n6681 ^ n6663;
  assign n6678 = n6648 & n6659;
  assign n6679 = n6678 ^ n6659;
  assign n6683 = n6682 ^ n6679;
  assign n6684 = n6671 & n6683;
  assign n6685 = n6684 ^ n6679;
  assign n6686 = ~n6677 & n6685;
  assign n6701 = n6658 ^ n6657;
  assign n6702 = n6701 ^ n6662;
  assign n7826 = n6673 & n6702;
  assign n7822 = n6679 ^ n6656;
  assign n7823 = ~n6671 & n7822;
  assign n7824 = n7823 ^ n6656;
  assign n7825 = n6677 & n7824;
  assign n7827 = n7826 ^ n7825;
  assign n6690 = n6661 ^ n6634;
  assign n6691 = n6690 ^ n6635;
  assign n6689 = n6660 ^ n6632;
  assign n6692 = n6691 ^ n6689;
  assign n6693 = n6648 & n6692;
  assign n6694 = n6693 ^ n6692;
  assign n6687 = n6681 ^ n6649;
  assign n6688 = n6687 ^ n6650;
  assign n6695 = n6694 ^ n6688;
  assign n6696 = ~n6671 & n6695;
  assign n6697 = n6696 ^ n6693;
  assign n6698 = n6677 & n6697;
  assign n6699 = n6698 ^ n6693;
  assign n7828 = n6702 ^ n6691;
  assign n7829 = n6675 & ~n7828;
  assign n7830 = n6673 ^ n6672;
  assign n7831 = n6694 & ~n7830;
  assign n6706 = n6662 ^ n6651;
  assign n7832 = n6675 & n6706;
  assign n6709 = n6688 ^ n6652;
  assign n6710 = n6709 ^ n6662;
  assign n6708 = n6678 ^ n6669;
  assign n6711 = n6710 ^ n6708;
  assign n6707 = n6706 ^ n6695;
  assign n6712 = n6711 ^ n6707;
  assign n7838 = n6712 ^ n6634;
  assign n7837 = n6695 ^ n6679;
  assign n7839 = n7838 ^ n7837;
  assign n7840 = n7839 ^ n6634;
  assign n7834 = n6680 ^ n6668;
  assign n7835 = n7834 ^ n6652;
  assign n7833 = n7828 ^ n6662;
  assign n7836 = n7835 ^ n7833;
  assign n7841 = n7840 ^ n7836;
  assign n7842 = n7841 ^ n7836;
  assign n7843 = n6671 & n7842;
  assign n7844 = n7843 ^ n7836;
  assign n7845 = n6677 & ~n7844;
  assign n7846 = n7845 ^ n7836;
  assign n7847 = ~n7832 & n7846;
  assign n7848 = ~n7831 & n7847;
  assign n7849 = ~n7829 & n7848;
  assign n7850 = ~n6699 & n7849;
  assign n7851 = ~n7827 & n7850;
  assign n7852 = ~n6686 & n7851;
  assign n7853 = ~n6676 & n7852;
  assign n7854 = n7853 ^ n4961;
  assign n7855 = n7854 ^ x338;
  assign n6393 = n6392 ^ x256;
  assign n6394 = n4924 ^ x261;
  assign n6395 = n4611 & n4654;
  assign n6396 = n4631 ^ n4619;
  assign n6397 = ~n4458 & n6396;
  assign n6398 = n5825 ^ n4613;
  assign n6399 = n4654 & n6398;
  assign n6401 = n6270 ^ n4626;
  assign n6400 = n4629 ^ n4616;
  assign n6402 = n6401 ^ n6400;
  assign n6403 = n6400 ^ n4661;
  assign n6404 = n6400 & n6403;
  assign n6405 = n6404 ^ n6400;
  assign n6406 = ~n6402 & n6405;
  assign n6407 = n6406 ^ n6404;
  assign n6408 = n6407 ^ n6400;
  assign n6409 = n6408 ^ n4661;
  assign n6410 = ~n6399 & n6409;
  assign n6411 = n6410 ^ n6399;
  assign n6412 = n4617 ^ n4614;
  assign n6413 = n6412 ^ n4629;
  assign n6414 = n6413 ^ n5818;
  assign n6415 = n4457 & n6414;
  assign n6416 = n6415 ^ n5818;
  assign n6417 = ~n4310 & ~n6416;
  assign n6418 = ~n6411 & ~n6417;
  assign n6419 = ~n6266 & n6418;
  assign n6420 = ~n6397 & n6419;
  assign n6421 = ~n6395 & n6420;
  assign n6422 = ~n4310 & n4669;
  assign n6423 = n6422 ^ n4609;
  assign n6424 = n4457 & n6423;
  assign n6425 = n6424 ^ n4609;
  assign n6426 = n6421 & ~n6425;
  assign n6427 = ~n4636 & n6426;
  assign n6428 = ~n4675 & n6427;
  assign n6429 = n6428 ^ n3347;
  assign n6430 = n6429 ^ x259;
  assign n6431 = n5499 ^ x260;
  assign n6432 = ~n6430 & ~n6431;
  assign n6495 = n6432 ^ n6430;
  assign n6455 = n6454 ^ x257;
  assign n6457 = n5659 & n6456;
  assign n6464 = n6463 ^ n5670;
  assign n6462 = n5705 ^ n5686;
  assign n6465 = n6464 ^ n6462;
  assign n6466 = n5660 & ~n5698;
  assign n6467 = n6466 ^ n5662;
  assign n6468 = ~n6464 & ~n6467;
  assign n6469 = n6468 ^ n6466;
  assign n6470 = n6465 & ~n6469;
  assign n6471 = n6470 ^ n6462;
  assign n6460 = ~n5661 & n5684;
  assign n6458 = n5711 ^ n5686;
  assign n6459 = n6458 ^ n5682;
  assign n6461 = n6460 ^ n6459;
  assign n6472 = n6471 ^ n6461;
  assign n6473 = ~n6189 & n6472;
  assign n6474 = n6473 ^ n6471;
  assign n6475 = ~n6457 & ~n6474;
  assign n6476 = n5660 & n5670;
  assign n6477 = n6476 ^ n5642;
  assign n6478 = n5662 & n6477;
  assign n6479 = n6478 ^ n5642;
  assign n6480 = n6475 & ~n6479;
  assign n6481 = n6202 ^ n5658;
  assign n6482 = ~n5584 & n6481;
  assign n6483 = n6482 ^ n5658;
  assign n6484 = n5585 & n6483;
  assign n6485 = n6480 & ~n6484;
  assign n6486 = ~n5669 & n6485;
  assign n6487 = ~n5663 & n6486;
  assign n6488 = ~n5656 & n6487;
  assign n6489 = n6488 ^ n3392;
  assign n6490 = n6489 ^ x258;
  assign n6491 = ~n6455 & n6490;
  assign n6492 = n6491 ^ n6455;
  assign n6504 = n6492 ^ n6490;
  assign n6508 = n6504 ^ n6455;
  assign n6518 = ~n6495 & n6508;
  assign n6498 = n6495 ^ n6431;
  assign n6515 = ~n6498 & n6504;
  assign n6499 = n6498 ^ n6430;
  assign n6511 = ~n6492 & ~n6499;
  assign n6516 = n6515 ^ n6511;
  assign n6510 = ~n6492 & ~n6498;
  assign n6512 = n6511 ^ n6510;
  assign n6501 = n6491 & ~n6498;
  assign n6513 = n6512 ^ n6501;
  assign n6514 = n6513 ^ n6498;
  assign n6517 = n6516 ^ n6514;
  assign n6519 = n6518 ^ n6517;
  assign n7039 = ~n6394 & ~n6519;
  assign n7040 = n7039 ^ n6518;
  assign n7041 = n6393 & n7040;
  assign n6500 = n6491 & ~n6499;
  assign n6502 = n6501 ^ n6500;
  assign n6523 = n6510 ^ n6502;
  assign n6505 = n6432 & n6504;
  assign n6496 = n6491 & ~n6495;
  assign n6497 = n6496 ^ n6491;
  assign n6503 = n6502 ^ n6497;
  assign n6506 = n6505 ^ n6503;
  assign n6493 = n6432 & ~n6492;
  assign n6494 = n6493 ^ n6432;
  assign n6507 = n6506 ^ n6494;
  assign n6509 = n6508 ^ n6507;
  assign n6520 = n6519 ^ n6509;
  assign n6524 = n6523 ^ n6520;
  assign n6525 = n6524 ^ n6430;
  assign n6526 = n6525 ^ n6514;
  assign n6527 = n6526 ^ n6518;
  assign n6528 = n6393 & n6527;
  assign n6529 = n6528 ^ n6518;
  assign n6530 = ~n6394 & n6529;
  assign n6521 = ~n6394 & ~n6520;
  assign n6522 = n6393 & n6521;
  assign n6531 = n6530 ^ n6522;
  assign n6538 = n6520 ^ n6507;
  assign n6539 = n6538 ^ n6515;
  assign n6548 = ~n6393 & ~n6394;
  assign n7856 = ~n6539 & n6548;
  assign n6532 = n6493 ^ n6492;
  assign n6533 = n6532 ^ n6512;
  assign n7857 = ~n6393 & ~n6513;
  assign n6544 = n6394 ^ n6393;
  assign n7858 = ~n6493 & n6544;
  assign n7859 = ~n6510 & n7858;
  assign n6577 = n6511 ^ n6496;
  assign n7860 = n6394 & ~n6577;
  assign n7861 = ~n7859 & ~n7860;
  assign n7862 = ~n6503 & ~n7861;
  assign n7863 = ~n7857 & ~n7862;
  assign n7864 = n6533 & ~n7863;
  assign n7865 = n7864 ^ n6393;
  assign n7866 = n6517 ^ n6505;
  assign n7867 = n7866 ^ n6500;
  assign n7868 = n7867 ^ n7864;
  assign n7869 = n7864 ^ n6394;
  assign n7870 = n7864 & n7869;
  assign n7871 = n7870 ^ n7864;
  assign n7872 = n7868 & n7871;
  assign n7873 = n7872 ^ n7870;
  assign n7874 = n7873 ^ n7864;
  assign n7875 = n7874 ^ n6394;
  assign n7876 = ~n7865 & n7875;
  assign n7877 = n7876 ^ n7864;
  assign n7878 = ~n7856 & n7877;
  assign n7880 = n6523 ^ n6518;
  assign n7045 = n6526 ^ n6507;
  assign n7046 = n7045 ^ n6517;
  assign n7879 = n7046 ^ n6493;
  assign n7881 = n7880 ^ n7879;
  assign n6575 = ~n6495 & n6504;
  assign n7882 = n7881 ^ n6575;
  assign n7883 = n6394 & ~n7882;
  assign n7884 = n7883 ^ n6575;
  assign n7885 = n6544 & n7884;
  assign n7886 = n7878 & ~n7885;
  assign n7887 = ~n6531 & n7886;
  assign n7888 = ~n7041 & n7887;
  assign n7889 = n7888 ^ n5420;
  assign n7890 = n7889 ^ x337;
  assign n7891 = ~n7855 & ~n7890;
  assign n7892 = n7891 ^ n7855;
  assign n7893 = n7892 ^ n7890;
  assign n7894 = n6302 & n6329;
  assign n7895 = n6291 ^ n6257;
  assign n7896 = n7895 ^ n6309;
  assign n7897 = n7896 ^ n6347;
  assign n7898 = n7897 ^ n6315;
  assign n7899 = n7898 ^ n6344;
  assign n7900 = n6344 ^ n6012;
  assign n7901 = n6043 & n7900;
  assign n7902 = n7901 ^ n6012;
  assign n7903 = ~n7899 & n7902;
  assign n7904 = n7903 ^ n7898;
  assign n7905 = ~n6310 & ~n7904;
  assign n7906 = n7905 ^ n6292;
  assign n7907 = ~n6043 & ~n7906;
  assign n7908 = n7907 ^ n6292;
  assign n7909 = n6326 & n6346;
  assign n7910 = ~n7908 & ~n7909;
  assign n7917 = n6337 ^ n6294;
  assign n7915 = n7897 ^ n6307;
  assign n7916 = n7915 ^ n6298;
  assign n7918 = n7917 ^ n7916;
  assign n7919 = ~n6043 & n7918;
  assign n7920 = n7919 ^ n7916;
  assign n7911 = n6335 ^ n6331;
  assign n7912 = n7911 ^ n6314;
  assign n7913 = ~n6012 & n7912;
  assign n7914 = n7913 ^ n6314;
  assign n7921 = n7920 ^ n7914;
  assign n7922 = ~n6326 & ~n7921;
  assign n7923 = n7922 ^ n7914;
  assign n7924 = n7910 & n7923;
  assign n7925 = ~n7894 & n7924;
  assign n7926 = ~n6330 & n7925;
  assign n7927 = ~n6319 & n7926;
  assign n7928 = n7927 ^ n5384;
  assign n7929 = n7928 ^ x336;
  assign n7930 = n7528 ^ n7522;
  assign n7931 = n7930 ^ n7490;
  assign n7932 = ~n7478 & n7931;
  assign n7933 = n7932 ^ n7490;
  assign n7934 = n7479 & n7933;
  assign n7935 = ~n7481 & n7485;
  assign n7937 = n7550 ^ n7498;
  assign n7936 = n7522 ^ n7512;
  assign n7938 = n7937 ^ n7936;
  assign n7939 = ~n7507 & ~n7938;
  assign n7946 = n7510 ^ n7498;
  assign n7947 = n7946 ^ n7495;
  assign n7948 = n7947 ^ n7512;
  assign n7949 = n7479 & ~n7948;
  assign n7940 = n7550 ^ n7526;
  assign n7941 = n7480 & n7940;
  assign n7942 = ~n7506 & ~n7513;
  assign n7943 = n7514 ^ n7511;
  assign n7944 = ~n7942 & n7943;
  assign n7945 = ~n7941 & ~n7944;
  assign n7950 = n7949 ^ n7945;
  assign n7951 = ~n7478 & ~n7950;
  assign n7952 = n7951 ^ n7945;
  assign n7953 = ~n7939 & n7952;
  assign n7954 = ~n7935 & n7953;
  assign n7955 = ~n7479 & ~n7525;
  assign n7956 = n7955 ^ n7528;
  assign n7957 = n7478 & ~n7956;
  assign n7958 = n7954 & ~n7957;
  assign n7959 = ~n7934 & n7958;
  assign n7960 = ~n7530 & n7959;
  assign n7961 = ~n7505 & n7960;
  assign n7962 = n7961 ^ n4456;
  assign n7963 = n7962 ^ x335;
  assign n7964 = ~n7929 & ~n7963;
  assign n8014 = ~n7893 & n7964;
  assign n7990 = n7891 & n7964;
  assign n8024 = n8014 ^ n7990;
  assign n7991 = n7990 ^ n7891;
  assign n7965 = n7964 ^ n7963;
  assign n7966 = n7965 ^ n7929;
  assign n7970 = ~n7892 & ~n7966;
  assign n7986 = n7970 ^ n7892;
  assign n7987 = n7986 ^ n7964;
  assign n7980 = n7963 ^ n7855;
  assign n7981 = n7929 ^ n7890;
  assign n7982 = ~n7855 & ~n7981;
  assign n7983 = n7982 ^ n7929;
  assign n7984 = ~n7980 & ~n7983;
  assign n7985 = n7984 ^ n7929;
  assign n7988 = n7987 ^ n7985;
  assign n7968 = n7891 & ~n7966;
  assign n7989 = n7988 ^ n7968;
  assign n7992 = n7991 ^ n7989;
  assign n7978 = ~n7892 & ~n7965;
  assign n7976 = n7893 ^ n7855;
  assign n7977 = ~n7965 & ~n7976;
  assign n7979 = n7978 ^ n7977;
  assign n7993 = n7992 ^ n7979;
  assign n7994 = n7993 ^ n7965;
  assign n8816 = n8024 ^ n7994;
  assign n8817 = n7791 & ~n8816;
  assign n8818 = n8817 ^ n7994;
  assign n8819 = n7975 & ~n8818;
  assign n7821 = n7820 ^ n7818;
  assign n7971 = n7970 ^ n7966;
  assign n7967 = ~n7893 & ~n7966;
  assign n7969 = n7968 ^ n7967;
  assign n7972 = n7971 ^ n7969;
  assign n7973 = n7821 & ~n7972;
  assign n7995 = n7994 ^ n7977;
  assign n7996 = n7791 & ~n7995;
  assign n7999 = n7996 ^ n7977;
  assign n8000 = ~n7818 & n7999;
  assign n9065 = n7988 ^ n7972;
  assign n9066 = n7819 & ~n9065;
  assign n8001 = n7964 ^ n7929;
  assign n8002 = ~n7893 & ~n8001;
  assign n8022 = n8002 ^ n7970;
  assign n8004 = ~n7892 & n7964;
  assign n9067 = n8022 ^ n8004;
  assign n9068 = n7791 & n9067;
  assign n9069 = n9068 ^ n8004;
  assign n9070 = ~n7818 & n9069;
  assign n8023 = n8004 ^ n7964;
  assign n8025 = n8024 ^ n8023;
  assign n9071 = n8025 ^ n7985;
  assign n9072 = ~n7791 & ~n9071;
  assign n9073 = n9072 ^ n8025;
  assign n9074 = n7975 & n9073;
  assign n9075 = n9074 ^ n8025;
  assign n9076 = ~n9070 & ~n9075;
  assign n8005 = n8004 ^ n7978;
  assign n8006 = n8005 ^ n7986;
  assign n8007 = n8006 ^ n8001;
  assign n8003 = n8002 ^ n7988;
  assign n8008 = n8007 ^ n8003;
  assign n8009 = n8008 ^ n8006;
  assign n9078 = ~n7974 & ~n8009;
  assign n9079 = ~n8008 & ~n9078;
  assign n9080 = n9079 ^ n7967;
  assign n8822 = n7820 & n7988;
  assign n9077 = n8822 ^ n7970;
  assign n9081 = n9080 ^ n9077;
  assign n9082 = ~n7975 & ~n9081;
  assign n9083 = n7993 ^ n7968;
  assign n9084 = n7820 & n9083;
  assign n9085 = n9084 ^ n7968;
  assign n9086 = ~n9082 & ~n9085;
  assign n9087 = n9076 & n9086;
  assign n9088 = ~n9066 & n9087;
  assign n9089 = ~n8000 & n9088;
  assign n9090 = ~n7973 & n9089;
  assign n9091 = ~n8819 & n9090;
  assign n9092 = n9091 ^ n5499;
  assign n9093 = n9092 ^ x358;
  assign n9095 = n9064 & ~n9093;
  assign n9094 = n9093 ^ n9064;
  assign n9096 = n9095 ^ n9094;
  assign n8664 = ~n7483 & n7526;
  assign n8665 = n7947 ^ n7485;
  assign n8666 = n8665 ^ n7514;
  assign n8667 = ~n7507 & ~n8666;
  assign n8668 = ~n8664 & ~n8667;
  assign n8673 = n7550 ^ n7490;
  assign n8669 = n7519 ^ n7517;
  assign n8670 = n8669 ^ n7493;
  assign n8671 = n7479 & n8670;
  assign n8672 = n8671 ^ n7493;
  assign n8674 = n8673 ^ n8672;
  assign n8675 = n8674 ^ n8672;
  assign n8676 = n7479 & n8675;
  assign n8677 = n8676 ^ n8672;
  assign n8678 = ~n7478 & n8677;
  assign n8679 = n8678 ^ n8672;
  assign n8680 = n8668 & ~n8679;
  assign n8682 = ~n7481 & n7524;
  assign n8681 = n7506 & n7930;
  assign n8683 = n8682 ^ n8681;
  assign n8684 = n8680 & ~n8683;
  assign n8685 = ~n7934 & n8684;
  assign n8686 = ~n7505 & n8685;
  assign n8687 = n8686 ^ n5053;
  assign n8688 = n8687 ^ x343;
  assign n5535 = n5534 ^ n5529;
  assign n5532 = n5531 ^ n5129;
  assign n5533 = n5532 ^ n5530;
  assign n5536 = n5535 ^ n5533;
  assign n5537 = n5352 & n5536;
  assign n5538 = n5537 ^ n5533;
  assign n5539 = n5500 & n5538;
  assign n5550 = n5503 & n5543;
  assign n5545 = n5544 ^ n5514;
  assign n5546 = n5545 ^ n5510;
  assign n5547 = ~n5500 & n5546;
  assign n5548 = n5547 ^ n5510;
  assign n5549 = ~n5540 & n5548;
  assign n5551 = n5550 ^ n5549;
  assign n5552 = n5534 ^ n5528;
  assign n5553 = ~n5502 & ~n5552;
  assign n5555 = n5554 ^ n5533;
  assign n5556 = n5504 & n5555;
  assign n5557 = n5542 ^ n5529;
  assign n5558 = ~n5502 & n5557;
  assign n5568 = n5567 ^ n5134;
  assign n5563 = n5514 ^ n5131;
  assign n5564 = n5563 ^ n5562;
  assign n5565 = n5564 ^ n5561;
  assign n5566 = n5565 ^ n5559;
  assign n5569 = n5568 ^ n5566;
  assign n5570 = n5501 & n5569;
  assign n5571 = ~n5500 & n5525;
  assign n5572 = n5571 ^ n5519;
  assign n5573 = n5540 & ~n5572;
  assign n5574 = n5573 ^ n5519;
  assign n5575 = ~n5570 & n5574;
  assign n5576 = ~n5558 & n5575;
  assign n5577 = ~n5556 & n5576;
  assign n5578 = ~n5553 & n5577;
  assign n5579 = ~n5551 & n5578;
  assign n5580 = ~n5539 & n5579;
  assign n5581 = ~n5505 & n5580;
  assign n5582 = n5581 ^ n4707;
  assign n8689 = n5582 ^ x344;
  assign n8690 = n8688 & ~n8689;
  assign n8691 = n8690 ^ n8689;
  assign n8693 = n7817 ^ x341;
  assign n8694 = n7787 ^ n4972;
  assign n8695 = n8694 ^ x342;
  assign n8696 = n8693 & n8695;
  assign n8706 = ~n8691 & n8696;
  assign n6864 = n6863 ^ n6862;
  assign n6865 = ~n6740 & ~n6864;
  assign n6866 = n6865 ^ n6862;
  assign n6867 = n6741 & ~n6866;
  assign n6886 = n6875 & n6885;
  assign n6887 = n6886 ^ n6884;
  assign n6896 = ~n6740 & ~n6845;
  assign n6897 = n6896 ^ n6844;
  assign n6898 = ~n6741 & n6897;
  assign n6899 = ~n6740 & n6841;
  assign n6900 = n6899 ^ n6839;
  assign n6901 = n6739 & n6900;
  assign n6902 = n6851 ^ n6840;
  assign n6903 = n6885 & n6902;
  assign n6904 = n6868 ^ n6854;
  assign n6905 = n6904 ^ n6875;
  assign n6906 = n6905 ^ n6850;
  assign n6907 = n6906 ^ n6850;
  assign n6908 = ~n6740 & n6907;
  assign n6909 = n6908 ^ n6850;
  assign n6910 = ~n6741 & ~n6909;
  assign n6911 = n6910 ^ n6850;
  assign n6912 = ~n6903 & n6911;
  assign n6913 = ~n6740 & ~n6860;
  assign n6914 = n6913 ^ n6835;
  assign n6915 = n6739 & n6914;
  assign n6916 = n6915 ^ n6835;
  assign n6917 = n6912 & ~n6916;
  assign n6918 = ~n6901 & n6917;
  assign n6919 = ~n6898 & n6918;
  assign n6920 = n6895 & n6919;
  assign n6921 = ~n6887 & n6920;
  assign n6922 = ~n6867 & n6921;
  assign n6923 = n6922 ^ n4838;
  assign n8724 = n6923 ^ x345;
  assign n8723 = n7854 ^ x340;
  assign n8735 = n8724 ^ n8723;
  assign n8744 = n8706 & ~n8735;
  assign n8697 = n8696 ^ n8693;
  assign n8712 = n8690 & n8697;
  assign n8725 = n8723 & ~n8724;
  assign n8726 = n8725 ^ n8724;
  assign n8727 = n8726 ^ n8723;
  assign n8728 = n8727 ^ n8724;
  assign n8739 = n8712 & n8728;
  assign n8708 = n8690 ^ n8688;
  assign n8709 = n8696 & n8708;
  assign n8710 = n8709 ^ n8696;
  assign n8692 = n8691 ^ n8688;
  assign n8702 = n8692 & n8696;
  assign n8707 = n8706 ^ n8702;
  assign n8711 = n8710 ^ n8707;
  assign n8713 = n8712 ^ n8711;
  assign n8736 = n8713 & ~n8723;
  assign n8737 = n8736 ^ n8712;
  assign n8740 = n8739 ^ n8737;
  assign n8738 = n8735 & n8737;
  assign n8741 = n8740 ^ n8738;
  assign n8731 = ~n8691 & n8697;
  assign n8732 = n8731 ^ n8697;
  assign n8698 = n8697 ^ n8695;
  assign n8716 = ~n8698 & n8708;
  assign n8715 = ~n8691 & ~n8698;
  assign n8717 = n8716 ^ n8715;
  assign n8718 = n8717 ^ n8698;
  assign n8699 = n8698 ^ n8693;
  assign n8701 = n8690 & n8699;
  assign n8705 = n8701 ^ n8690;
  assign n8714 = n8713 ^ n8705;
  assign n8719 = n8718 ^ n8714;
  assign n8720 = n8719 ^ n8701;
  assign n8721 = n8720 ^ n8692;
  assign n8703 = n8702 ^ n8701;
  assign n8700 = n8692 & n8699;
  assign n8704 = n8703 ^ n8700;
  assign n8722 = n8721 ^ n8704;
  assign n8730 = n8722 ^ n8712;
  assign n8733 = n8732 ^ n8730;
  assign n8734 = ~n8726 & ~n8733;
  assign n8742 = n8741 ^ n8734;
  assign n8743 = n8742 ^ n8739;
  assign n8745 = n8744 ^ n8743;
  assign n8764 = n8709 ^ n8700;
  assign n8936 = n8723 & n8764;
  assign n8937 = n8936 ^ n8700;
  assign n8938 = ~n8735 & n8937;
  assign n8939 = n8709 & ~n8726;
  assign n8944 = ~n8723 & n8731;
  assign n8941 = n8722 ^ n8702;
  assign n8754 = n8714 ^ n8700;
  assign n8753 = ~n8691 & n8699;
  assign n8755 = n8754 ^ n8753;
  assign n8752 = n8720 ^ n8714;
  assign n8756 = n8755 ^ n8752;
  assign n8751 = n8719 ^ n8699;
  assign n8757 = n8756 ^ n8751;
  assign n8942 = n8941 ^ n8757;
  assign n8940 = n8753 ^ n8752;
  assign n8943 = n8942 ^ n8940;
  assign n8945 = n8944 ^ n8943;
  assign n8946 = ~n8735 & n8945;
  assign n8947 = n8946 ^ n8943;
  assign n8950 = n8704 & n8728;
  assign n8948 = n8717 & ~n8735;
  assign n8949 = n8948 ^ n8738;
  assign n8951 = n8950 ^ n8949;
  assign n8952 = ~n8947 & ~n8951;
  assign n8953 = ~n8939 & n8952;
  assign n8954 = ~n8938 & n8953;
  assign n8955 = ~n8745 & n8954;
  assign n8956 = n8955 ^ n5127;
  assign n8957 = n8956 ^ x361;
  assign n8077 = n6680 ^ n6657;
  assign n8078 = n8077 ^ n6662;
  assign n8079 = ~n6671 & n8078;
  assign n8076 = n6708 ^ n6693;
  assign n8080 = n8079 ^ n8076;
  assign n8081 = n6677 & n8080;
  assign n8082 = n8081 ^ n8076;
  assign n8084 = n7837 ^ n6663;
  assign n8083 = n7828 ^ n6710;
  assign n8085 = n8084 ^ n8083;
  assign n8086 = ~n6672 & ~n8085;
  assign n8087 = n8086 ^ n8083;
  assign n8088 = n6671 & ~n8087;
  assign n8089 = ~n8082 & ~n8088;
  assign n8096 = n7834 ^ n6656;
  assign n8097 = ~n6672 & n8096;
  assign n8098 = n8097 ^ n6656;
  assign n8091 = n6649 ^ n6635;
  assign n8092 = n8091 ^ n7822;
  assign n8093 = n8092 ^ n6648;
  assign n8094 = ~n6672 & ~n8093;
  assign n8090 = n6694 ^ n6664;
  assign n8095 = n8094 ^ n8090;
  assign n8099 = n8098 ^ n8095;
  assign n8100 = n6671 & n8099;
  assign n8101 = n8100 ^ n8095;
  assign n8102 = n8089 & ~n8101;
  assign n8103 = ~n7827 & n8102;
  assign n8104 = n8103 ^ n4309;
  assign n8451 = n8104 ^ x328;
  assign n8452 = n7962 ^ x333;
  assign n6540 = n6394 & ~n6539;
  assign n6534 = n6533 ^ n6507;
  assign n6535 = n6534 ^ n6526;
  assign n6536 = ~n6394 & ~n6535;
  assign n6537 = n6536 ^ n6526;
  assign n6541 = n6540 ^ n6537;
  assign n6542 = ~n6393 & n6541;
  assign n6543 = n6542 ^ n6537;
  assign n6553 = ~n6393 & n6505;
  assign n6551 = n6393 & n6502;
  assign n6552 = n6551 ^ n6501;
  assign n6554 = n6553 ^ n6552;
  assign n6555 = ~n6394 & n6554;
  assign n6556 = n6555 ^ n6552;
  assign n6549 = n6548 ^ n6544;
  assign n8053 = n6575 ^ n6549;
  assign n6578 = n6577 ^ n6510;
  assign n6579 = n6578 ^ n6507;
  assign n8054 = n6579 ^ n6548;
  assign n8055 = ~n6575 & ~n8054;
  assign n8056 = n8055 ^ n6548;
  assign n8057 = ~n8053 & n8056;
  assign n8058 = n8057 ^ n6549;
  assign n8064 = ~n6394 & n7880;
  assign n8060 = n6524 ^ n6503;
  assign n6574 = n6496 ^ n6493;
  assign n8059 = n7866 ^ n6574;
  assign n8061 = n8060 ^ n8059;
  assign n8062 = ~n6394 & n8061;
  assign n8063 = n8062 ^ n8059;
  assign n8065 = n8064 ^ n8063;
  assign n8066 = n6393 & ~n8065;
  assign n8067 = n8066 ^ n8063;
  assign n8068 = n8058 & n8067;
  assign n8069 = ~n6530 & n8068;
  assign n8070 = ~n6556 & n8069;
  assign n8071 = ~n6543 & n8070;
  assign n8072 = ~n7041 & n8071;
  assign n8073 = n8072 ^ n4543;
  assign n8483 = n8073 ^ x329;
  assign n7337 = n5533 ^ n5134;
  assign n7338 = ~n5502 & n7337;
  assign n8490 = n5569 ^ n5130;
  assign n8491 = n8490 ^ n5554;
  assign n8489 = n5515 ^ n4925;
  assign n8492 = n8491 ^ n8489;
  assign n8493 = ~n5134 & ~n8492;
  assign n7339 = n5518 ^ n5510;
  assign n7326 = n5554 ^ n5529;
  assign n8488 = n7339 ^ n7326;
  assign n8494 = n8493 ^ n8488;
  assign n8495 = n5352 & n8494;
  assign n8496 = n8495 ^ n8488;
  assign n8484 = n5561 ^ n5534;
  assign n8485 = ~n5352 & ~n8484;
  assign n8486 = n8485 ^ n5561;
  assign n8487 = ~n5516 & n8486;
  assign n8497 = n8496 ^ n8487;
  assign n8498 = n5500 & n8497;
  assign n8499 = n8498 ^ n8496;
  assign n8500 = ~n5549 & n8499;
  assign n8501 = ~n7338 & n8500;
  assign n8502 = ~n7646 & n8501;
  assign n8503 = ~n5539 & n8502;
  assign n8504 = ~n5505 & n8503;
  assign n8505 = ~n7331 & n8504;
  assign n8506 = n8505 ^ n4598;
  assign n8507 = n8506 ^ x330;
  assign n8508 = ~n8483 & n8507;
  assign n8537 = n8508 ^ n8483;
  assign n8453 = ~n6739 & n6849;
  assign n8454 = n6904 ^ n6902;
  assign n8455 = n8454 ^ n6848;
  assign n8456 = n7615 & ~n8455;
  assign n8457 = ~n8453 & ~n8456;
  assign n8458 = n6839 & ~n7616;
  assign n8459 = n6880 ^ n6740;
  assign n8460 = n6739 & n6878;
  assign n8461 = n8460 ^ n6876;
  assign n8462 = n8461 ^ n6880;
  assign n8463 = ~n8459 & n8462;
  assign n8464 = n8463 ^ n8460;
  assign n8465 = n8464 ^ n6876;
  assign n8466 = n8465 ^ n6740;
  assign n8467 = n6880 & ~n8466;
  assign n8468 = n8467 ^ n6880;
  assign n8469 = n8468 ^ n6740;
  assign n8470 = ~n8458 & n8469;
  assign n8471 = n8457 & n8470;
  assign n8473 = ~n6871 & n7616;
  assign n8472 = ~n6856 & n6885;
  assign n8474 = n8473 ^ n8472;
  assign n8475 = n8471 & ~n8474;
  assign n8476 = ~n6901 & n8475;
  assign n8477 = ~n7613 & n8476;
  assign n8478 = ~n6898 & n8477;
  assign n8479 = n8478 ^ n4492;
  assign n8480 = n8479 ^ x331;
  assign n8536 = n8480 & n8508;
  assign n8538 = n8537 ^ n8536;
  assign n8481 = n7790 ^ x332;
  assign n8524 = n8507 ^ n8481;
  assign n8525 = n8524 ^ n8480;
  assign n8526 = ~n8483 & ~n8525;
  assign n8482 = n8480 & n8481;
  assign n8518 = n8482 ^ n8480;
  assign n8519 = n8518 ^ n8481;
  assign n8520 = n8508 & ~n8519;
  assign n8521 = n8520 ^ n8508;
  assign n8516 = n8481 ^ n8480;
  assign n8517 = n8508 & n8516;
  assign n8522 = n8521 ^ n8517;
  assign n8514 = n8482 ^ n8481;
  assign n8515 = ~n8483 & n8514;
  assign n8523 = n8522 ^ n8515;
  assign n8527 = n8526 ^ n8523;
  assign n8539 = n8538 ^ n8527;
  assign n8533 = n8483 ^ n8480;
  assign n8534 = n8507 ^ n8483;
  assign n8535 = n8533 & ~n8534;
  assign n8540 = n8539 ^ n8535;
  assign n8531 = n8515 ^ n8514;
  assign n8509 = n8508 ^ n8507;
  assign n8529 = n8509 ^ n8483;
  assign n8530 = n8514 & n8529;
  assign n8532 = n8531 ^ n8530;
  assign n8541 = n8540 ^ n8532;
  assign n8511 = n8507 ^ n8480;
  assign n8512 = ~n8483 & n8511;
  assign n8513 = n8512 ^ n8483;
  assign n8528 = n8527 ^ n8513;
  assign n8542 = n8541 ^ n8528;
  assign n8554 = n8542 ^ n8519;
  assign n8550 = n8482 & n8529;
  assign n8551 = n8550 ^ n8529;
  assign n8545 = n8516 ^ n8483;
  assign n8546 = n8545 ^ n8507;
  assign n8547 = n8546 ^ n8526;
  assign n8543 = n8542 ^ n8530;
  assign n8510 = n8482 & n8509;
  assign n8544 = n8543 ^ n8510;
  assign n8548 = n8547 ^ n8544;
  assign n8549 = n8548 ^ n8530;
  assign n8552 = n8551 ^ n8549;
  assign n8553 = n8552 ^ n8520;
  assign n8555 = n8554 ^ n8553;
  assign n8556 = n8555 ^ n8552;
  assign n8557 = n8452 & ~n8556;
  assign n8558 = n8557 ^ n8552;
  assign n8559 = ~n8451 & ~n8558;
  assign n8560 = n8451 & ~n8452;
  assign n8561 = n8548 ^ n8528;
  assign n8562 = n8560 & n8561;
  assign n8564 = n8560 ^ n8452;
  assign n8563 = n8560 ^ n8451;
  assign n8565 = n8564 ^ n8563;
  assign n8568 = n8526 ^ n8483;
  assign n8566 = n8522 ^ n8520;
  assign n8567 = n8566 ^ n8539;
  assign n8569 = n8568 ^ n8567;
  assign n8570 = n8569 ^ n8539;
  assign n8571 = n8570 ^ n8532;
  assign n8572 = n8452 & ~n8571;
  assign n8573 = n8572 ^ n8532;
  assign n8574 = ~n8565 & n8573;
  assign n8582 = n8520 & n8563;
  assign n8575 = n8531 ^ n8509;
  assign n8576 = n8575 ^ n8544;
  assign n8577 = n8576 ^ n8532;
  assign n8578 = n8577 ^ n8550;
  assign n8579 = n8451 & n8578;
  assign n8580 = n8579 ^ n8550;
  assign n8581 = ~n8452 & n8580;
  assign n8583 = n8582 ^ n8581;
  assign n8584 = ~n8452 & ~n8549;
  assign n8585 = n8584 ^ n8530;
  assign n8586 = ~n8451 & n8585;
  assign n8597 = n8566 ^ n8543;
  assign n8595 = n8569 ^ n8517;
  assign n8596 = n8595 ^ n8522;
  assign n8598 = n8597 ^ n8596;
  assign n8599 = n8451 & n8598;
  assign n8600 = n8599 ^ n8596;
  assign n8589 = n8548 ^ n8510;
  assign n8590 = n8589 ^ n8517;
  assign n8591 = n8590 ^ n8480;
  assign n8587 = n8552 ^ n8528;
  assign n8588 = n8587 ^ n8544;
  assign n8592 = n8591 ^ n8588;
  assign n8593 = ~n8451 & ~n8592;
  assign n8594 = n8593 ^ n8588;
  assign n8601 = n8600 ^ n8594;
  assign n8602 = n8452 & n8601;
  assign n8603 = n8602 ^ n8600;
  assign n8604 = ~n8586 & ~n8603;
  assign n8605 = ~n8583 & n8604;
  assign n8606 = ~n8574 & n8605;
  assign n8607 = ~n8562 & n8606;
  assign n8608 = ~n8559 & n8607;
  assign n8609 = n8608 ^ n4684;
  assign n8958 = n8609 ^ x362;
  assign n9032 = n8957 & n8958;
  assign n5583 = n5582 ^ x346;
  assign n5972 = n5971 ^ x351;
  assign n6948 = ~n5583 & n5972;
  assign n6700 = n6656 & ~n6677;
  assign n6703 = n6702 ^ n6678;
  assign n6704 = n6703 ^ n6682;
  assign n6705 = n6675 & n6704;
  assign n6715 = n6711 ^ n6652;
  assign n6716 = n6715 ^ n6670;
  assign n6717 = n6716 ^ n6634;
  assign n6713 = n6671 & n6712;
  assign n6714 = n6713 ^ n6711;
  assign n6718 = n6717 ^ n6714;
  assign n6719 = n6718 ^ n6714;
  assign n6720 = n6671 & ~n6719;
  assign n6721 = n6720 ^ n6714;
  assign n6722 = n6677 & n6721;
  assign n6723 = n6722 ^ n6714;
  assign n6724 = ~n6705 & ~n6723;
  assign n6725 = ~n6700 & n6724;
  assign n6726 = ~n6699 & n6725;
  assign n6727 = ~n6686 & n6726;
  assign n6728 = ~n6676 & n6727;
  assign n6729 = n6728 ^ n4761;
  assign n6730 = n6729 ^ x348;
  assign n6924 = n6923 ^ x347;
  assign n6925 = ~n6730 & ~n6924;
  assign n6933 = n6925 ^ n6924;
  assign n6371 = n6370 ^ x350;
  assign n6545 = ~n6393 & n6516;
  assign n6546 = n6545 ^ n6515;
  assign n6547 = n6544 & n6546;
  assign n6550 = n6505 & ~n6549;
  assign n6557 = n6556 ^ n6550;
  assign n6558 = n6518 ^ n6501;
  assign n6559 = n6393 & n6558;
  assign n6560 = n6559 ^ n6518;
  assign n6561 = n6394 & n6560;
  assign n6562 = n6506 ^ n6501;
  assign n6563 = n6562 ^ n6500;
  assign n6564 = n6563 ^ n6500;
  assign n6565 = ~n6394 & n6564;
  assign n6566 = n6565 ^ n6500;
  assign n6567 = n6393 & n6566;
  assign n6568 = n6567 ^ n6500;
  assign n6569 = ~n6393 & ~n6533;
  assign n6570 = n6569 ^ n6517;
  assign n6571 = n6544 & ~n6570;
  assign n6572 = n6571 ^ n6517;
  assign n6573 = ~n6568 & n6572;
  assign n6576 = n6575 ^ n6574;
  assign n6580 = n6579 ^ n6576;
  assign n6581 = ~n6393 & n6580;
  assign n6582 = n6581 ^ n6576;
  assign n6583 = ~n6544 & n6582;
  assign n6584 = n6573 & ~n6583;
  assign n6585 = ~n6561 & n6584;
  assign n6586 = ~n6557 & n6585;
  assign n6587 = ~n6547 & n6586;
  assign n6588 = ~n6543 & n6587;
  assign n6589 = ~n6531 & n6588;
  assign n6590 = n6589 ^ n4788;
  assign n6591 = n6590 ^ x349;
  assign n6592 = ~n6371 & n6591;
  assign n6593 = n6592 ^ n6371;
  assign n6594 = n6593 ^ n6591;
  assign n6944 = n6594 ^ n6371;
  assign n6945 = ~n6933 & n6944;
  assign n6974 = n6945 ^ n6944;
  assign n6934 = ~n6371 & ~n6933;
  assign n6935 = n6591 & n6934;
  assign n6964 = n6935 ^ n6934;
  assign n6969 = n6964 ^ n6593;
  assign n6952 = ~n6593 & n6925;
  assign n6926 = n6925 ^ n6730;
  assign n6937 = ~n6593 & ~n6926;
  assign n6953 = n6952 ^ n6937;
  assign n6970 = n6969 ^ n6953;
  assign n6957 = n6926 ^ n6924;
  assign n6971 = n6970 ^ n6957;
  assign n6958 = n6592 & ~n6957;
  assign n6928 = n6924 ^ n6594;
  assign n6929 = n6730 & ~n6928;
  assign n6943 = n6934 ^ n6929;
  assign n6946 = n6945 ^ n6943;
  assign n6959 = n6958 ^ n6946;
  assign n6972 = n6971 ^ n6959;
  assign n6968 = ~n6926 & n6944;
  assign n6973 = n6972 ^ n6968;
  assign n6975 = n6974 ^ n6973;
  assign n6976 = n6975 ^ n6925;
  assign n6931 = n6928 ^ n6925;
  assign n6927 = n6594 & ~n6926;
  assign n6930 = n6929 ^ n6927;
  assign n6932 = n6931 ^ n6930;
  assign n6967 = n6952 ^ n6932;
  assign n6977 = n6976 ^ n6967;
  assign n6978 = n6977 ^ n6945;
  assign n8961 = n6948 & ~n6978;
  assign n8959 = n6948 ^ n5583;
  assign n8960 = n6937 & ~n8959;
  assign n8962 = n8961 ^ n8960;
  assign n5973 = n5972 ^ n5583;
  assign n6954 = n5583 & n6953;
  assign n6955 = n6954 ^ n6937;
  assign n6956 = n5973 & n6955;
  assign n6960 = n6959 ^ n6927;
  assign n6961 = ~n5583 & n6960;
  assign n6962 = n6961 ^ n6927;
  assign n6963 = n5972 & n6962;
  assign n6942 = n6592 & ~n6926;
  assign n6982 = n6970 ^ n6942;
  assign n6993 = n6982 ^ n6925;
  assign n6990 = n6973 ^ n6937;
  assign n6991 = n6990 ^ n6958;
  assign n6992 = n6991 ^ n6930;
  assign n6994 = n6993 ^ n6992;
  assign n8963 = ~n5972 & n6994;
  assign n8965 = n6959 & ~n8959;
  assign n6936 = n6935 ^ n6932;
  assign n6980 = n6975 ^ n6936;
  assign n8964 = ~n5973 & ~n6980;
  assign n8966 = n8965 ^ n8964;
  assign n6949 = n6948 ^ n5972;
  assign n8967 = n6977 ^ n6949;
  assign n8968 = n6977 & n8967;
  assign n8969 = n8968 ^ n6977;
  assign n8970 = n6972 ^ n6958;
  assign n8971 = n8970 ^ n6977;
  assign n8972 = n8969 & ~n8971;
  assign n8973 = n8972 ^ n8968;
  assign n8974 = n8973 ^ n6977;
  assign n8975 = n8974 ^ n6949;
  assign n8976 = ~n8966 & n8975;
  assign n8977 = n8976 ^ n8966;
  assign n8978 = ~n8963 & ~n8977;
  assign n8981 = n6982 ^ n6932;
  assign n8980 = n6977 ^ n6973;
  assign n8982 = n8981 ^ n8980;
  assign n7007 = n6994 ^ n6964;
  assign n8979 = n7007 ^ n6968;
  assign n8983 = n8982 ^ n8979;
  assign n8984 = n5583 & ~n8983;
  assign n8985 = n8984 ^ n8979;
  assign n7011 = n6972 ^ n6970;
  assign n7012 = n5583 & ~n7011;
  assign n7013 = n7012 ^ n6972;
  assign n8986 = n8985 ^ n7013;
  assign n8987 = n5973 & n8986;
  assign n8988 = n8987 ^ n7013;
  assign n8989 = n8978 & ~n8988;
  assign n8990 = ~n6963 & n8989;
  assign n8991 = ~n6956 & n8990;
  assign n8992 = ~n8962 & n8991;
  assign n8993 = n8992 ^ n4924;
  assign n8994 = n8993 ^ x359;
  assign n7029 = n5809 ^ n5766;
  assign n7030 = n7029 ^ n5961;
  assign n7028 = n5963 ^ n5887;
  assign n7031 = n7030 ^ n7028;
  assign n7032 = ~n5913 & ~n7031;
  assign n7033 = n7032 ^ n7028;
  assign n7024 = n5887 ^ n5884;
  assign n7025 = n7024 ^ n5960;
  assign n7026 = n5913 & ~n7025;
  assign n7027 = n7026 ^ n5960;
  assign n7034 = n7033 ^ n7027;
  assign n7035 = n5954 & n7034;
  assign n7036 = n7035 ^ n7027;
  assign n7037 = n7036 ^ n4099;
  assign n7038 = n7037 ^ x318;
  assign n7042 = n6393 & n6537;
  assign n7043 = n6510 ^ n6503;
  assign n7044 = n7043 ^ n6548;
  assign n7047 = n7046 ^ n6533;
  assign n7048 = n7047 ^ n6549;
  assign n7049 = ~n7043 & n7048;
  assign n7050 = n7049 ^ n6549;
  assign n7051 = n7044 & ~n7050;
  assign n7052 = n7051 ^ n6548;
  assign n7054 = n6576 ^ n6510;
  assign n7053 = n6574 ^ n6500;
  assign n7055 = n7054 ^ n7053;
  assign n7056 = ~n6393 & n7055;
  assign n7057 = n7056 ^ n7053;
  assign n7058 = n6544 & n7057;
  assign n7059 = ~n7052 & ~n7058;
  assign n7060 = ~n7042 & n7059;
  assign n7061 = ~n6561 & n7060;
  assign n7062 = ~n6557 & n7061;
  assign n7063 = ~n6547 & n7062;
  assign n7064 = ~n7041 & n7063;
  assign n7065 = n6520 & n7064;
  assign n7066 = n7065 ^ n3514;
  assign n7067 = n7066 ^ x317;
  assign n7068 = ~n7038 & ~n7067;
  assign n7089 = ~n6326 & n6338;
  assign n7086 = n6326 ^ n6296;
  assign n7087 = ~n6043 & ~n7086;
  assign n7084 = n6325 ^ n6309;
  assign n7085 = n6327 & n7084;
  assign n7088 = n7087 ^ n7085;
  assign n7090 = n7089 ^ n7088;
  assign n7070 = n6333 ^ n6323;
  assign n7071 = n7070 ^ n6338;
  assign n7081 = n6043 & n7071;
  assign n7075 = n6341 ^ n6310;
  assign n7076 = n6347 ^ n6329;
  assign n7077 = ~n6341 & ~n7076;
  assign n7078 = n7077 ^ n6329;
  assign n7079 = ~n7075 & ~n7078;
  assign n7080 = n7079 ^ n6310;
  assign n7082 = n7081 ^ n7080;
  assign n7069 = n6340 ^ n6302;
  assign n7072 = n7071 ^ n7069;
  assign n7073 = n6328 & ~n7072;
  assign n7074 = n7073 ^ n6302;
  assign n7083 = n7082 ^ n7074;
  assign n7091 = n7090 ^ n7083;
  assign n7092 = ~n6322 & ~n7091;
  assign n7093 = ~n6319 & n7092;
  assign n7094 = n7093 ^ n3916;
  assign n7095 = n7094 ^ x320;
  assign n7096 = ~n6739 & n6869;
  assign n7102 = n6862 ^ n6848;
  assign n7103 = n7102 ^ n6856;
  assign n7104 = ~n6740 & ~n7103;
  assign n7105 = n7104 ^ n6856;
  assign n7098 = n6869 ^ n6839;
  assign n7097 = n6880 ^ n6851;
  assign n7099 = n7098 ^ n7097;
  assign n7100 = n6740 & ~n7099;
  assign n7101 = n7100 ^ n7097;
  assign n7106 = n7105 ^ n7101;
  assign n7107 = n6739 & n7106;
  assign n7108 = n7107 ^ n7105;
  assign n7109 = ~n6867 & n7108;
  assign n7110 = ~n7096 & n7109;
  assign n7111 = n6740 & n6852;
  assign n7112 = n7111 ^ n6838;
  assign n7113 = n6741 & n7112;
  assign n7114 = n7110 & ~n7113;
  assign n7115 = ~n6740 & n6840;
  assign n7116 = n6848 ^ n6835;
  assign n7117 = n6740 & ~n7116;
  assign n7118 = n7117 ^ n6835;
  assign n7119 = n7118 ^ n6842;
  assign n7120 = ~n6741 & ~n7119;
  assign n7121 = n7120 ^ n6842;
  assign n7122 = ~n7115 & n7121;
  assign n7123 = n7114 & n7122;
  assign n7124 = ~n6887 & n7123;
  assign n7125 = n7124 ^ n3717;
  assign n7126 = n7125 ^ x319;
  assign n7127 = ~n7095 & n7126;
  assign n7129 = n7127 ^ n7095;
  assign n7138 = n7129 ^ n7126;
  assign n7141 = n7068 & n7138;
  assign n7286 = n7239 & n7260;
  assign n7287 = n7286 ^ n7238;
  assign n7288 = ~n7261 & n7287;
  assign n7295 = n7274 ^ n7227;
  assign n7296 = n7295 ^ n7234;
  assign n7297 = n7263 & ~n7296;
  assign n7299 = n7246 ^ n7241;
  assign n7298 = n7271 ^ n7248;
  assign n7300 = n7299 ^ n7298;
  assign n7301 = n7300 ^ n7274;
  assign n7302 = n7261 & n7301;
  assign n7303 = n7302 ^ n7274;
  assign n7304 = ~n7260 & ~n7303;
  assign n7312 = ~n7261 & n7311;
  assign n7305 = n7245 ^ n7230;
  assign n7306 = n7266 & ~n7305;
  assign n7308 = n7307 ^ n7242;
  assign n7309 = n7308 ^ n7255;
  assign n7310 = ~n7306 & ~n7309;
  assign n7313 = n7312 ^ n7310;
  assign n7314 = n7279 & n7313;
  assign n7315 = n7314 ^ n7310;
  assign n7316 = ~n7304 & ~n7315;
  assign n7317 = ~n7297 & n7316;
  assign n7318 = ~n7294 & n7317;
  assign n7319 = ~n7288 & n7318;
  assign n7320 = n7285 & n7319;
  assign n7321 = ~n7276 & n7320;
  assign n7322 = ~n7265 & n7321;
  assign n7323 = n7322 ^ n2771;
  assign n7324 = n7323 ^ x316;
  assign n7325 = ~n5502 & n5565;
  assign n7327 = n5503 & n7326;
  assign n7341 = n7340 ^ n5516;
  assign n7342 = n7341 ^ n7339;
  assign n7343 = n5500 & ~n7342;
  assign n7344 = n7343 ^ n7339;
  assign n7345 = n5540 & ~n7344;
  assign n7346 = ~n7338 & ~n7345;
  assign n7347 = ~n5556 & n7346;
  assign n7348 = ~n5553 & n7347;
  assign n7349 = ~n7336 & n7348;
  assign n7350 = ~n5505 & n7349;
  assign n7351 = ~n7331 & n7350;
  assign n7352 = ~n7327 & n7351;
  assign n7353 = ~n7325 & n7352;
  assign n7355 = n5500 & n5544;
  assign n7354 = n5504 & ~n7332;
  assign n7356 = n7355 ^ n7354;
  assign n7357 = n7353 & ~n7356;
  assign n7358 = ~n5551 & n7357;
  assign n7359 = n7358 ^ n3273;
  assign n7360 = n7359 ^ x321;
  assign n7361 = n7324 & n7360;
  assign n7368 = n7361 ^ n7360;
  assign n7383 = n7141 & n7368;
  assign n7161 = n7068 ^ n7038;
  assign n7364 = ~n7129 & ~n7161;
  assign n7162 = n7127 & ~n7161;
  assign n7365 = n7364 ^ n7162;
  assign n7366 = n7365 ^ n7161;
  assign n7139 = n7138 ^ n7095;
  assign n7159 = n7141 ^ n7139;
  assign n7133 = n7126 ^ n7038;
  assign n7134 = n7133 ^ n7067;
  assign n7155 = n7134 ^ n7038;
  assign n7156 = n7133 & n7155;
  assign n7157 = n7156 ^ n7134;
  assign n7158 = n7095 & ~n7157;
  assign n7160 = n7159 ^ n7158;
  assign n7163 = n7162 ^ n7160;
  assign n7164 = n7163 ^ n7126;
  assign n7130 = n7068 ^ n7067;
  assign n7147 = ~n7130 & n7138;
  assign n7146 = n7127 & ~n7130;
  assign n7148 = n7147 ^ n7146;
  assign n7131 = ~n7129 & ~n7130;
  assign n7145 = n7131 ^ n7130;
  assign n7149 = n7148 ^ n7145;
  assign n7140 = n7068 & n7139;
  assign n7144 = n7140 ^ n7131;
  assign n7150 = n7149 ^ n7144;
  assign n7153 = n7150 ^ n7146;
  assign n7142 = n7141 ^ n7140;
  assign n7135 = n7134 ^ n7095;
  assign n7136 = n7133 ^ n7129;
  assign n7137 = n7135 & n7136;
  assign n7143 = n7142 ^ n7137;
  assign n7151 = n7150 ^ n7143;
  assign n7128 = n7068 & n7127;
  assign n7132 = n7131 ^ n7128;
  assign n7152 = n7151 ^ n7132;
  assign n7154 = n7153 ^ n7152;
  assign n7165 = n7164 ^ n7154;
  assign n7367 = n7366 ^ n7165;
  assign n7369 = n7368 ^ n7324;
  assign n7370 = ~n7367 & ~n7369;
  assign n7380 = n7360 ^ n7324;
  assign n8995 = n7163 ^ n7148;
  assign n8996 = n7360 & n8995;
  assign n8997 = n8996 ^ n7163;
  assign n8998 = ~n7380 & n8997;
  assign n7372 = n7165 & n7368;
  assign n7371 = n7160 & n7368;
  assign n7373 = n7372 ^ n7371;
  assign n7378 = n7130 ^ n7038;
  assign n7379 = ~n7129 & ~n7378;
  assign n8999 = n7379 ^ n7367;
  assign n9000 = n7361 & ~n8999;
  assign n7374 = n7160 ^ n7149;
  assign n7375 = n7360 & ~n7374;
  assign n7376 = n7375 ^ n7160;
  assign n7377 = n7324 & n7376;
  assign n7391 = n7147 ^ n7138;
  assign n7392 = n7391 ^ n7367;
  assign n7393 = n7392 ^ n7141;
  assign n9001 = n7393 ^ n7162;
  assign n9002 = n7380 & ~n9001;
  assign n9003 = n7146 ^ n7144;
  assign n9004 = n7368 & n9003;
  assign n7384 = n7128 ^ n7068;
  assign n7385 = n7384 ^ n7142;
  assign n7386 = n7385 ^ n7141;
  assign n7387 = n7386 ^ n7364;
  assign n7388 = ~n7360 & n7387;
  assign n7389 = n7388 ^ n7364;
  assign n7390 = n7324 & n7389;
  assign n9007 = n7150 ^ n7128;
  assign n9006 = n7142 ^ n7067;
  assign n9008 = n9007 ^ n9006;
  assign n9005 = n7165 ^ n7128;
  assign n9009 = n9008 ^ n9005;
  assign n9010 = ~n7360 & n9009;
  assign n9011 = n9010 ^ n9005;
  assign n9012 = ~n7380 & n9011;
  assign n9014 = ~n7151 & ~n7360;
  assign n7362 = n7361 ^ n7324;
  assign n9013 = n7144 & n7362;
  assign n9015 = n9014 ^ n9013;
  assign n9016 = ~n9012 & ~n9015;
  assign n9017 = ~n7390 & n9016;
  assign n9018 = ~n9004 & n9017;
  assign n9019 = ~n9002 & n9018;
  assign n9020 = ~n7377 & n9019;
  assign n9021 = ~n9000 & n9020;
  assign n9022 = ~n7373 & n9021;
  assign n9023 = ~n8998 & n9022;
  assign n9024 = ~n7370 & n9023;
  assign n9025 = ~n7383 & n9024;
  assign n9026 = n9025 ^ n4182;
  assign n9027 = n9026 ^ x360;
  assign n9028 = ~n8994 & n9027;
  assign n9039 = n9028 ^ n9027;
  assign n9045 = n9032 & n9039;
  assign n9110 = n9045 ^ n9032;
  assign n9040 = n9039 ^ n8994;
  assign n9042 = n9032 & n9040;
  assign n9033 = n9032 ^ n8957;
  assign n9034 = n9033 ^ n8958;
  assign n9035 = n9034 ^ n8957;
  assign n9036 = n9028 & n9035;
  assign n9029 = ~n8958 & n9028;
  assign n9031 = n9029 ^ n9028;
  assign n9037 = n9036 ^ n9031;
  assign n9101 = n9042 ^ n9037;
  assign n9111 = n9110 ^ n9101;
  assign n9060 = n9028 ^ n8994;
  assign n9112 = n9111 ^ n9060;
  assign n9108 = n9035 & ~n9060;
  assign n9048 = n9035 & n9040;
  assign n9054 = n9048 ^ n9040;
  assign n9041 = ~n9034 & n9040;
  assign n9043 = n9042 ^ n9041;
  assign n9055 = n9054 ^ n9043;
  assign n9056 = n9055 ^ n9033;
  assign n9030 = ~n8957 & n9029;
  assign n9052 = n9030 ^ n9029;
  assign n9051 = n9033 & n9039;
  assign n9053 = n9052 ^ n9051;
  assign n9057 = n9056 ^ n9053;
  assign n9109 = n9108 ^ n9057;
  assign n9113 = n9112 ^ n9109;
  assign n9114 = n9096 & ~n9113;
  assign n9104 = n9051 & n9064;
  assign n9102 = n9064 & n9101;
  assign n9103 = n9102 ^ n9037;
  assign n9105 = n9104 ^ n9103;
  assign n9106 = ~n9093 & n9105;
  assign n9107 = n9106 ^ n9103;
  assign n9115 = n9114 ^ n9107;
  assign n10763 = n9051 & n9096;
  assign n10764 = ~n9115 & ~n10763;
  assign n9061 = n9060 ^ n9033;
  assign n9047 = ~n9034 & n9039;
  assign n9049 = n9048 ^ n9047;
  assign n9046 = n9045 ^ n9036;
  assign n9050 = n9049 ^ n9046;
  assign n9058 = n9057 ^ n9050;
  assign n9038 = n9037 ^ n9030;
  assign n9044 = n9043 ^ n9038;
  assign n9059 = n9058 ^ n9044;
  assign n9062 = n9061 ^ n9059;
  assign n9063 = n9062 ^ n9055;
  assign n10765 = n9063 & ~n9093;
  assign n10766 = n10765 ^ n9052;
  assign n10767 = n9094 & n10766;
  assign n10768 = n10767 ^ n9052;
  assign n10374 = n9113 ^ n9057;
  assign n10375 = n9093 & ~n10374;
  assign n10376 = n10375 ^ n9113;
  assign n10377 = ~n9064 & ~n10376;
  assign n11470 = n9108 ^ n9095;
  assign n11471 = n9052 ^ n9046;
  assign n11472 = n11471 ^ n9093;
  assign n11473 = ~n9095 & ~n11472;
  assign n11474 = n11473 ^ n11471;
  assign n11475 = n11470 & n11474;
  assign n11476 = n11475 ^ n9108;
  assign n11482 = n9055 ^ n9038;
  assign n11483 = n11482 ^ n9047;
  assign n11484 = n9093 & n11483;
  assign n10775 = n9055 ^ n9042;
  assign n11478 = n10775 ^ n9050;
  assign n10387 = n9045 ^ n9042;
  assign n11477 = n10387 ^ n9062;
  assign n11479 = n11478 ^ n11477;
  assign n11480 = ~n9093 & n11479;
  assign n11481 = n11480 ^ n11477;
  assign n11485 = n11484 ^ n11481;
  assign n11486 = n11485 ^ n11481;
  assign n11487 = ~n9041 & ~n11486;
  assign n11488 = n11487 ^ n11481;
  assign n11489 = n9064 & ~n11488;
  assign n11490 = n11489 ^ n11481;
  assign n11491 = ~n11476 & ~n11490;
  assign n11492 = ~n10377 & n11491;
  assign n11493 = ~n10768 & n11492;
  assign n11494 = n10764 & n11493;
  assign n11495 = n11494 ^ n7676;
  assign n11496 = n11495 ^ x402;
  assign n6938 = n6937 ^ n6936;
  assign n6939 = ~n5583 & ~n6938;
  assign n6940 = n6939 ^ n6937;
  assign n6941 = n5973 & n6940;
  assign n6947 = n6946 ^ n6942;
  assign n6950 = n6949 ^ n5583;
  assign n6951 = n6947 & n6950;
  assign n6965 = n6949 & n6964;
  assign n6966 = n6965 ^ n6963;
  assign n6979 = n6949 & ~n6978;
  assign n6981 = n6980 ^ n6927;
  assign n6983 = n6982 ^ n6981;
  assign n6984 = n6983 ^ n6968;
  assign n6985 = n6984 ^ n6968;
  assign n6986 = ~n5972 & n6985;
  assign n6987 = n6986 ^ n6968;
  assign n6988 = ~n5583 & n6987;
  assign n6989 = n6988 ^ n6968;
  assign n6995 = n6994 ^ n6942;
  assign n6996 = n6995 ^ n6945;
  assign n6997 = ~n5583 & n6996;
  assign n6998 = n6997 ^ n6945;
  assign n6999 = n5973 & n6998;
  assign n7000 = ~n6989 & ~n6999;
  assign n7003 = ~n5973 & n6952;
  assign n7001 = n6949 & ~n6980;
  assign n7002 = n6934 & n7001;
  assign n7004 = n7003 ^ n7002;
  assign n7005 = n7000 & ~n7004;
  assign n7006 = ~n6979 & n7005;
  assign n7008 = n7007 ^ n6972;
  assign n7009 = n5583 & n7008;
  assign n7010 = n7009 ^ n6972;
  assign n7014 = n7013 ^ n7010;
  assign n7015 = ~n5973 & n7014;
  assign n7016 = n7015 ^ n7010;
  assign n7017 = n7006 & ~n7016;
  assign n7018 = ~n6966 & n7017;
  assign n7019 = ~n6956 & n7018;
  assign n7020 = ~n6951 & n7019;
  assign n7021 = ~n6941 & n7020;
  assign n7022 = n7021 ^ n6830;
  assign n9816 = n7022 ^ x383;
  assign n9817 = n7746 & n7765;
  assign n9818 = n7569 & n7683;
  assign n7728 = n7707 ^ n7609;
  assign n7724 = n7722 ^ n7706;
  assign n7727 = n7726 ^ n7724;
  assign n7729 = n7728 ^ n7727;
  assign n7732 = n7731 ^ n7729;
  assign n7733 = n7732 ^ n7726;
  assign n7747 = n7746 ^ n7567;
  assign n9819 = n7733 & ~n7747;
  assign n9820 = n7679 ^ n7567;
  assign n9821 = n7727 ^ n7698;
  assign n9822 = ~n7566 & ~n9821;
  assign n9823 = n9822 ^ n7698;
  assign n9824 = n9823 ^ n7679;
  assign n9825 = ~n9820 & ~n9824;
  assign n9826 = n9825 ^ n9822;
  assign n9827 = n9826 ^ n7698;
  assign n9828 = n9827 ^ n7567;
  assign n9829 = ~n7679 & n9828;
  assign n9830 = n9829 ^ n7679;
  assign n9831 = n9830 ^ n7567;
  assign n9832 = ~n9819 & n9831;
  assign n9835 = n7720 ^ n7695;
  assign n9836 = ~n7763 & n9835;
  assign n9837 = n9836 ^ n7695;
  assign n9838 = n9837 ^ n7568;
  assign n9833 = n7699 & n7746;
  assign n9834 = n9833 ^ n7684;
  assign n9839 = n9838 ^ n9834;
  assign n9840 = n9832 & n9839;
  assign n9841 = ~n8785 & n9840;
  assign n9842 = ~n9818 & n9841;
  assign n9843 = ~n9817 & n9842;
  assign n9844 = ~n7566 & n7692;
  assign n9845 = n9844 ^ n7711;
  assign n9846 = ~n7567 & ~n9845;
  assign n9847 = n9846 ^ n7711;
  assign n9848 = n9843 & n9847;
  assign n9849 = ~n8784 & n9848;
  assign n9850 = n9849 ^ n6773;
  assign n9851 = n9850 ^ x385;
  assign n9852 = n9816 & n9851;
  assign n9853 = n9852 ^ n9851;
  assign n9222 = n7148 & n7368;
  assign n9223 = n9222 ^ n9000;
  assign n9232 = n7385 ^ n7151;
  assign n9401 = n7361 & ~n9232;
  assign n9402 = n7386 ^ n7131;
  assign n9403 = ~n7369 & n9402;
  assign n7363 = n7165 & n7362;
  assign n9405 = n7364 ^ n7151;
  assign n9406 = n9405 ^ n7393;
  assign n9404 = n7360 & ~n9007;
  assign n9407 = n9406 ^ n9404;
  assign n9408 = ~n7380 & n9407;
  assign n9409 = n9408 ^ n9406;
  assign n9410 = n7379 ^ n7163;
  assign n9411 = n9410 ^ n7142;
  assign n9412 = ~n7324 & n9411;
  assign n9413 = n9412 ^ n7142;
  assign n9414 = ~n7360 & n9413;
  assign n9415 = ~n9409 & ~n9414;
  assign n9416 = ~n7363 & n9415;
  assign n9417 = ~n7372 & n9416;
  assign n9418 = ~n7370 & n9417;
  assign n9419 = ~n9403 & n9418;
  assign n9420 = ~n9401 & n9419;
  assign n9422 = n7128 & n7380;
  assign n9421 = ~n7149 & ~n7360;
  assign n9423 = n9422 ^ n9421;
  assign n9424 = n9420 & ~n9423;
  assign n9425 = ~n9223 & n9424;
  assign n9426 = ~n7383 & n9425;
  assign n9427 = n9426 ^ n6042;
  assign n9780 = n9427 ^ x386;
  assign n8729 = ~n8722 & n8728;
  assign n9282 = n8733 ^ n8725;
  assign n9283 = n8727 ^ n8711;
  assign n9284 = n8733 & ~n9283;
  assign n9285 = n9284 ^ n8727;
  assign n9286 = ~n9282 & n9285;
  assign n9287 = n9286 ^ n8725;
  assign n9288 = ~n8739 & ~n9287;
  assign n9781 = n8724 & n8731;
  assign n9782 = n8707 & n8725;
  assign n9791 = n8755 ^ n8724;
  assign n9792 = ~n8723 & ~n9791;
  assign n9793 = n9792 ^ n8724;
  assign n9794 = ~n8756 & n9793;
  assign n9795 = n9794 ^ n8752;
  assign n9796 = ~n8716 & n9795;
  assign n9296 = n8757 ^ n8716;
  assign n9783 = n9296 ^ n8701;
  assign n9784 = n9783 ^ n8730;
  assign n9785 = n9783 ^ n8724;
  assign n9786 = n8723 & ~n9785;
  assign n9787 = n9786 ^ n8724;
  assign n9788 = ~n9784 & n9787;
  assign n9789 = n9788 ^ n8730;
  assign n9790 = ~n8706 & n9789;
  assign n9797 = n9796 ^ n9790;
  assign n9798 = n8723 & n9797;
  assign n9799 = n9798 ^ n9790;
  assign n9800 = ~n8939 & n9799;
  assign n9801 = ~n9782 & n9800;
  assign n9802 = ~n9781 & n9801;
  assign n8758 = n8757 ^ n8715;
  assign n9803 = n8758 ^ n8701;
  assign n9804 = n9803 ^ n8941;
  assign n9805 = ~n8724 & ~n9804;
  assign n9806 = n9805 ^ n8941;
  assign n9807 = ~n8723 & ~n9806;
  assign n9808 = n9802 & ~n9807;
  assign n9809 = ~n8938 & n9808;
  assign n9810 = n9288 & n9809;
  assign n9811 = ~n8729 & n9810;
  assign n9812 = n9811 ^ n6804;
  assign n9813 = n9812 ^ x384;
  assign n9814 = n9780 & n9813;
  assign n9864 = n9814 ^ n9813;
  assign n9868 = n9864 ^ n9780;
  assign n9886 = n9853 & ~n9868;
  assign n9887 = n9886 ^ n9853;
  assign n9857 = n9852 ^ n9816;
  assign n9858 = n9814 & n9857;
  assign n9879 = n9858 ^ n9857;
  assign n9870 = ~n9813 & n9857;
  assign n9880 = n9879 ^ n9870;
  assign n9856 = n9814 & n9852;
  assign n9875 = n9856 ^ n9852;
  assign n9873 = n9852 & n9864;
  assign n9815 = n9814 ^ n9780;
  assign n9872 = n9815 & n9852;
  assign n9874 = n9873 ^ n9872;
  assign n9876 = n9875 ^ n9874;
  assign n9869 = n9857 & ~n9868;
  assign n9871 = n9870 ^ n9869;
  assign n9877 = n9876 ^ n9871;
  assign n9881 = n9880 ^ n9877;
  assign n9882 = n9881 ^ n9873;
  assign n9883 = n9882 ^ n9864;
  assign n9854 = n9853 ^ n9816;
  assign n9865 = ~n9854 & n9864;
  assign n9878 = n9877 ^ n9865;
  assign n9884 = n9883 ^ n9878;
  assign n9860 = n9814 & n9853;
  assign n9885 = n9884 ^ n9860;
  assign n9888 = n9887 ^ n9885;
  assign n9866 = n9865 ^ n9854;
  assign n9861 = n9860 ^ n9814;
  assign n9859 = n9858 ^ n9856;
  assign n9862 = n9861 ^ n9859;
  assign n9855 = n9815 & ~n9854;
  assign n9863 = n9862 ^ n9855;
  assign n9867 = n9866 ^ n9863;
  assign n9889 = n9888 ^ n9867;
  assign n9462 = n8563 & ~n8589;
  assign n9471 = n8588 ^ n8517;
  assign n9469 = n8550 ^ n8542;
  assign n9470 = n9469 ^ n8595;
  assign n9472 = n9471 ^ n9470;
  assign n9473 = ~n8451 & n9472;
  assign n9474 = n9473 ^ n9470;
  assign n9466 = n8535 ^ n8481;
  assign n9467 = ~n8451 & n9466;
  assign n9463 = n8555 ^ n8510;
  assign n9464 = n9463 ^ n8569;
  assign n9465 = n9464 ^ n8550;
  assign n9468 = n9467 ^ n9465;
  assign n9475 = n9474 ^ n9468;
  assign n9476 = ~n8452 & n9475;
  assign n9477 = n9476 ^ n9474;
  assign n9478 = ~n8583 & ~n9477;
  assign n9479 = ~n8562 & n9478;
  assign n9480 = ~n9462 & n9479;
  assign n9481 = ~n8559 & n9480;
  assign n9482 = n9481 ^ n6288;
  assign n9890 = n9482 ^ x387;
  assign n8074 = n8073 ^ x327;
  assign n8075 = n7094 ^ x322;
  assign n8141 = n7258 ^ n7231;
  assign n8142 = n7262 & n8141;
  assign n8143 = ~n7299 & ~n8142;
  assign n8144 = n7279 & ~n8143;
  assign n8145 = n7583 ^ n7278;
  assign n8146 = n8145 ^ n7256;
  assign n8147 = n8146 ^ n7250;
  assign n8148 = ~n7261 & n8147;
  assign n8149 = n8148 ^ n7250;
  assign n8150 = ~n7260 & ~n8149;
  assign n8151 = ~n8144 & ~n8150;
  assign n8152 = n7253 ^ n7236;
  assign n8153 = n8152 ^ n7269;
  assign n8154 = n8153 ^ n7269;
  assign n8155 = n7260 & n8154;
  assign n8156 = n8155 ^ n7269;
  assign n8157 = n7261 & n8156;
  assign n8158 = n8157 ^ n7269;
  assign n8159 = n8151 & ~n8158;
  assign n8160 = ~n7297 & n8159;
  assign n8161 = ~n7288 & n8160;
  assign n8162 = n7576 & n8161;
  assign n8163 = ~n7275 & n8162;
  assign n8164 = ~n7265 & n8163;
  assign n8165 = n8164 ^ n6108;
  assign n8166 = n8165 ^ x324;
  assign n8106 = ~n7478 & n7556;
  assign n8107 = n7479 & ~n7529;
  assign n8108 = n8107 ^ n7477;
  assign n8109 = ~n7478 & n8108;
  assign n8110 = n8109 ^ n7477;
  assign n8111 = n7946 ^ n7513;
  assign n8112 = n8111 ^ n7519;
  assign n8113 = n7478 & n8112;
  assign n8114 = n8113 ^ n7519;
  assign n8115 = ~n7479 & n8114;
  assign n8116 = ~n8110 & ~n8115;
  assign n8117 = ~n7483 & n7512;
  assign n8118 = n7500 ^ n7496;
  assign n8119 = n7480 & n8118;
  assign n8124 = n7526 ^ n7524;
  assign n8125 = n8124 ^ n7489;
  assign n8126 = n8125 ^ n7527;
  assign n8127 = n7478 & n8126;
  assign n8128 = n8127 ^ n7527;
  assign n8120 = n7946 ^ n7519;
  assign n8121 = n8120 ^ n7523;
  assign n8122 = n7478 & ~n8121;
  assign n8123 = n8122 ^ n8120;
  assign n8129 = n8128 ^ n8123;
  assign n8130 = n7479 & n8129;
  assign n8131 = n8130 ^ n8128;
  assign n8132 = ~n7504 & ~n8131;
  assign n8133 = ~n7530 & n8132;
  assign n8134 = ~n8119 & n8133;
  assign n8135 = ~n8117 & n8134;
  assign n8136 = n8116 & n8135;
  assign n8137 = ~n8106 & n8136;
  assign n8138 = n8137 ^ n6073;
  assign n8139 = n8138 ^ x325;
  assign n8182 = n8166 ^ n8139;
  assign n8167 = n7359 ^ x323;
  assign n8168 = n8167 ^ n8166;
  assign n8105 = n8104 ^ x326;
  assign n8140 = n8139 ^ n8105;
  assign n8196 = n8167 ^ n8140;
  assign n8197 = n8168 & ~n8196;
  assign n8198 = n8197 ^ n8167;
  assign n8208 = ~n8182 & ~n8198;
  assign n8209 = n8208 ^ n8140;
  assign n8170 = ~n8166 & ~n8167;
  assign n8171 = n8170 ^ n8167;
  assign n8172 = ~n8105 & n8171;
  assign n8173 = n8172 ^ n8167;
  assign n8169 = n8139 & n8168;
  assign n8174 = n8173 ^ n8169;
  assign n8175 = n8140 & ~n8174;
  assign n8176 = n8175 ^ n8173;
  assign n8210 = n8209 ^ n8176;
  assign n8177 = n8167 ^ n8139;
  assign n8178 = n8105 & n8177;
  assign n8179 = ~n8166 & n8178;
  assign n8180 = n8167 & n8179;
  assign n8211 = n8210 ^ n8180;
  assign n8212 = n8211 ^ n8177;
  assign n8213 = n8075 & n8212;
  assign n8191 = n8166 ^ n8105;
  assign n8192 = n8191 ^ n8139;
  assign n8183 = n8167 & ~n8182;
  assign n8184 = n8183 ^ n8166;
  assign n8187 = n8167 ^ n8105;
  assign n8189 = n8184 & ~n8187;
  assign n8188 = n8187 ^ n8184;
  assign n8190 = n8189 ^ n8188;
  assign n8193 = n8192 ^ n8190;
  assign n8214 = n8213 ^ n8193;
  assign n8195 = n8173 ^ n8168;
  assign n8199 = n8198 ^ n8195;
  assign n8181 = n8180 ^ n8176;
  assign n8200 = n8199 ^ n8181;
  assign n8201 = n8193 & n8200;
  assign n8202 = n8201 ^ n8187;
  assign n8185 = n8184 ^ n8181;
  assign n8186 = n8185 ^ n8177;
  assign n8194 = n8193 ^ n8186;
  assign n8203 = n8202 ^ n8194;
  assign n8204 = n8203 ^ n8140;
  assign n8205 = n8204 ^ n8186;
  assign n8206 = n8075 & ~n8205;
  assign n8207 = n8206 ^ n8186;
  assign n8215 = n8214 ^ n8207;
  assign n8216 = n8074 & ~n8215;
  assign n8217 = n8216 ^ n8207;
  assign n8218 = n8217 ^ n6738;
  assign n9891 = n8218 ^ x382;
  assign n9892 = ~n9890 & ~n9891;
  assign n9893 = n9892 ^ n9890;
  assign n9894 = ~n9889 & ~n9893;
  assign n9899 = ~n9889 & ~n9891;
  assign n9895 = n9880 ^ n9860;
  assign n9896 = n9895 ^ n9877;
  assign n9897 = n9891 & n9896;
  assign n9898 = n9897 ^ n9877;
  assign n9900 = n9899 ^ n9898;
  assign n9901 = n9890 & n9900;
  assign n9902 = n9901 ^ n9898;
  assign n9903 = ~n9890 & n9895;
  assign n9904 = n9903 ^ n9860;
  assign n9905 = ~n9891 & n9904;
  assign n9906 = n9886 & n9892;
  assign n9907 = n9891 ^ n9890;
  assign n9908 = n9863 ^ n9856;
  assign n9909 = n9908 ^ n9873;
  assign n9910 = ~n9907 & n9909;
  assign n9911 = ~n9906 & ~n9910;
  assign n9912 = n9892 ^ n9891;
  assign n9913 = n9884 & ~n9912;
  assign n9920 = n9870 ^ n9865;
  assign n9921 = n9920 ^ n9884;
  assign n9914 = n9869 ^ n9858;
  assign n9915 = n9880 ^ n9876;
  assign n9916 = n9915 ^ n9874;
  assign n9917 = ~n9890 & n9916;
  assign n9918 = n9917 ^ n9915;
  assign n9919 = ~n9914 & ~n9918;
  assign n9922 = n9921 ^ n9919;
  assign n9923 = n9922 ^ n9919;
  assign n9924 = n9890 & n9923;
  assign n9925 = n9924 ^ n9919;
  assign n9926 = ~n9907 & ~n9925;
  assign n9927 = n9926 ^ n9919;
  assign n9928 = ~n9913 & n9927;
  assign n9929 = n9911 & n9928;
  assign n9930 = ~n9905 & n9929;
  assign n9931 = ~n9902 & n9930;
  assign n9932 = ~n9894 & n9931;
  assign n9933 = n9932 ^ n7641;
  assign n11497 = n9933 ^ x404;
  assign n11498 = ~n11496 & ~n11497;
  assign n11499 = n11498 ^ n11497;
  assign n11500 = n11499 ^ n11496;
  assign n8221 = n7641 ^ x310;
  assign n8220 = n7066 ^ x315;
  assign n8222 = n8221 ^ n8220;
  assign n8223 = n7323 ^ x314;
  assign n8234 = n7899 ^ n7071;
  assign n8235 = n8234 ^ n6335;
  assign n8232 = n7915 ^ n6325;
  assign n8233 = n8232 ^ n6336;
  assign n8236 = n8235 ^ n8233;
  assign n8237 = ~n6012 & n8236;
  assign n8238 = n8237 ^ n8235;
  assign n8227 = n6338 ^ n6309;
  assign n8228 = n8227 ^ n6314;
  assign n8229 = n6328 & ~n8228;
  assign n8230 = n8229 ^ n6343;
  assign n8224 = n6327 & n6333;
  assign n8225 = n8224 ^ n6312;
  assign n8226 = n8225 ^ n6298;
  assign n8231 = n8230 ^ n8226;
  assign n8239 = n8238 ^ n8231;
  assign n8240 = ~n6326 & n8239;
  assign n8241 = n8240 ^ n8231;
  assign n8242 = ~n7080 & n8241;
  assign n8243 = ~n7894 & n8242;
  assign n8244 = ~n6330 & n8243;
  assign n8245 = ~n6322 & n8244;
  assign n8246 = n8245 ^ n5637;
  assign n8247 = n8246 ^ x313;
  assign n8248 = ~n8223 & n8247;
  assign n8249 = n7565 ^ x311;
  assign n8250 = n6663 & n6671;
  assign n8251 = n8250 ^ n6651;
  assign n8252 = n6672 & n8251;
  assign n8253 = n8252 ^ n6651;
  assign n8254 = n7828 ^ n6682;
  assign n8255 = n6675 & ~n8254;
  assign n8256 = n6703 ^ n6680;
  assign n8257 = n8256 ^ n6693;
  assign n8258 = n6673 & n6703;
  assign n8259 = n8258 ^ n6674;
  assign n8260 = n8257 & n8259;
  assign n8261 = ~n8255 & ~n8260;
  assign n8262 = n7830 ^ n6662;
  assign n8263 = n8256 ^ n6673;
  assign n8264 = ~n7830 & ~n8263;
  assign n8265 = n8264 ^ n6673;
  assign n8266 = ~n8262 & ~n8265;
  assign n8267 = n8266 ^ n6662;
  assign n8268 = n8261 & ~n8267;
  assign n8269 = ~n7825 & n8268;
  assign n8275 = n6695 ^ n6652;
  assign n8271 = n6694 ^ n6682;
  assign n8270 = n6693 ^ n6668;
  assign n8272 = n8271 ^ n8270;
  assign n8273 = n6671 & n8272;
  assign n8274 = n8273 ^ n8270;
  assign n8276 = n8275 ^ n8274;
  assign n8277 = n6677 & n8276;
  assign n8278 = n8277 ^ n8275;
  assign n8279 = n8269 & ~n8278;
  assign n8280 = ~n8253 & n8279;
  assign n8281 = ~n6676 & n8280;
  assign n8282 = n8281 ^ n5605;
  assign n8283 = n8282 ^ x312;
  assign n8284 = n8249 & n8283;
  assign n8299 = n8284 ^ n8283;
  assign n8300 = n8248 & n8299;
  assign n8321 = n8300 ^ n8299;
  assign n8287 = n8248 ^ n8223;
  assign n8290 = n8287 ^ n8247;
  assign n8297 = n8290 ^ n8223;
  assign n8319 = n8297 & n8299;
  assign n8313 = n8284 & n8297;
  assign n8311 = n8284 & n8290;
  assign n8302 = n8248 & n8284;
  assign n8312 = n8311 ^ n8302;
  assign n8314 = n8313 ^ n8312;
  assign n8315 = n8314 ^ n8284;
  assign n8285 = n8284 ^ n8249;
  assign n8288 = n8285 & ~n8287;
  assign n8316 = n8315 ^ n8288;
  assign n8317 = n8316 ^ n8287;
  assign n8294 = n8285 ^ n8283;
  assign n8295 = n8290 & ~n8294;
  assign n8306 = n8295 ^ n8294;
  assign n8303 = n8302 ^ n8248;
  assign n8286 = n8248 & n8285;
  assign n8301 = n8300 ^ n8286;
  assign n8304 = n8303 ^ n8301;
  assign n8298 = ~n8294 & n8297;
  assign n8305 = n8304 ^ n8298;
  assign n8307 = n8306 ^ n8305;
  assign n8318 = n8317 ^ n8307;
  assign n8320 = n8319 ^ n8318;
  assign n8322 = n8321 ^ n8320;
  assign n8323 = ~n8221 & n8322;
  assign n8291 = n8285 & n8290;
  assign n8292 = n8291 ^ n8285;
  assign n8289 = n8288 ^ n8286;
  assign n8293 = n8292 ^ n8289;
  assign n8296 = n8295 ^ n8293;
  assign n8308 = n8307 ^ n8296;
  assign n8309 = n8221 & ~n8308;
  assign n8310 = n8309 ^ n8307;
  assign n8324 = n8323 ^ n8310;
  assign n8325 = n8222 & ~n8324;
  assign n8326 = n8325 ^ n8310;
  assign n8327 = n8307 ^ n8304;
  assign n8328 = n8221 & ~n8327;
  assign n8329 = n8328 ^ n8304;
  assign n8330 = n8220 & n8329;
  assign n8331 = n8220 & ~n8221;
  assign n8333 = n8331 ^ n8221;
  assign n8335 = n8286 & ~n8333;
  assign n8611 = n8327 ^ n8319;
  assign n8612 = n8611 ^ n8312;
  assign n8613 = ~n8220 & ~n8612;
  assign n8614 = n8613 ^ n8312;
  assign n8615 = n8222 & n8614;
  assign n8340 = n8315 ^ n8291;
  assign n8341 = n8340 ^ n8293;
  assign n8342 = n8221 & n8341;
  assign n8343 = n8342 ^ n8293;
  assign n8344 = n8222 & n8343;
  assign n8618 = n8221 & n8313;
  assign n8616 = ~n8221 & n8289;
  assign n8617 = n8616 ^ n8286;
  assign n8619 = n8618 ^ n8617;
  assign n8620 = ~n8220 & n8619;
  assign n8621 = n8620 ^ n8617;
  assign n8622 = n8300 ^ n8291;
  assign n8623 = n8622 ^ n8320;
  assign n8624 = ~n8220 & n8623;
  assign n8625 = n8624 ^ n8320;
  assign n8626 = ~n8221 & n8625;
  assign n8632 = n8322 ^ n8286;
  assign n8628 = n8331 ^ n8220;
  assign n8629 = n8318 & n8628;
  assign n8630 = n8629 ^ n8295;
  assign n8627 = n8312 ^ n8298;
  assign n8631 = n8630 ^ n8627;
  assign n8633 = n8632 ^ n8631;
  assign n8634 = n8633 ^ n8631;
  assign n8635 = ~n8220 & n8634;
  assign n8636 = n8635 ^ n8631;
  assign n8637 = n8222 & n8636;
  assign n8638 = n8637 ^ n8631;
  assign n8639 = ~n8626 & ~n8638;
  assign n8640 = ~n8621 & n8639;
  assign n8641 = ~n8344 & n8640;
  assign n8642 = ~n8615 & n8641;
  assign n8643 = ~n8335 & n8642;
  assign n8644 = ~n8330 & n8643;
  assign n8645 = n8326 & n8644;
  assign n8646 = n8645 ^ n5724;
  assign n10257 = n8646 ^ x371;
  assign n9575 = ~n8451 & n9469;
  assign n9576 = n9575 ^ n8530;
  assign n9577 = n8452 & n9576;
  assign n9578 = n9577 ^ n8530;
  assign n10258 = ~n8452 & n8576;
  assign n10259 = n8553 ^ n8532;
  assign n10260 = n10259 ^ n8567;
  assign n10261 = n10259 ^ n8452;
  assign n10262 = n8565 & n10261;
  assign n10263 = n10262 ^ n8452;
  assign n10264 = n10260 & n10263;
  assign n10265 = n10264 ^ n8567;
  assign n10266 = n8548 & n10265;
  assign n10267 = ~n8565 & ~n10266;
  assign n10268 = ~n10258 & ~n10267;
  assign n10272 = n8452 & ~n8536;
  assign n10269 = ~n8527 & n8560;
  assign n10270 = n10269 ^ n8523;
  assign n10273 = n10272 ^ n10270;
  assign n10274 = ~n8565 & n10273;
  assign n10271 = n10270 ^ n8451;
  assign n10275 = n10274 ^ n10271;
  assign n10276 = n10268 & ~n10275;
  assign n10277 = n9469 ^ n8589;
  assign n10278 = ~n8452 & ~n10277;
  assign n10279 = n10278 ^ n8589;
  assign n10280 = n8565 & ~n10279;
  assign n10281 = n10276 & ~n10280;
  assign n10282 = ~n9578 & n10281;
  assign n10283 = ~n8574 & n10282;
  assign n10284 = ~n8559 & n10283;
  assign n10285 = n10284 ^ n5838;
  assign n10286 = n10285 ^ x372;
  assign n10287 = ~n10257 & ~n10286;
  assign n10288 = n10287 ^ n10257;
  assign n9435 = n6927 & n6948;
  assign n9436 = n9435 ^ n6979;
  assign n10289 = n5973 & n7010;
  assign n10290 = n6950 & ~n6977;
  assign n10291 = n6949 & ~n6967;
  assign n9431 = n6959 ^ n6942;
  assign n9432 = n5583 & n9431;
  assign n9433 = n9432 ^ n6942;
  assign n9434 = ~n5973 & n9433;
  assign n10294 = n5583 & ~n6982;
  assign n10292 = ~n5583 & n6992;
  assign n10293 = n10292 ^ n6991;
  assign n10295 = n10294 ^ n10293;
  assign n10296 = n5972 & n10295;
  assign n10297 = n10296 ^ n10293;
  assign n10298 = ~n9434 & ~n10297;
  assign n10299 = ~n10291 & n10298;
  assign n10300 = ~n10290 & n10299;
  assign n10301 = n6975 ^ n6937;
  assign n10302 = n10301 ^ n6929;
  assign n10303 = n10302 ^ n6975;
  assign n10304 = n10303 ^ n6975;
  assign n10305 = ~n5583 & n10304;
  assign n10306 = n10305 ^ n6975;
  assign n10307 = n5972 & n10306;
  assign n10308 = n10307 ^ n6975;
  assign n10309 = n10300 & ~n10308;
  assign n10310 = ~n8960 & n10309;
  assign n10311 = ~n10289 & n10310;
  assign n10312 = ~n9436 & n10311;
  assign n10313 = n10312 ^ n5808;
  assign n10314 = n10313 ^ x373;
  assign n7381 = n7379 & n7380;
  assign n7382 = ~n7367 & n7368;
  assign n7394 = ~n7360 & ~n7393;
  assign n7397 = n7154 & ~n7360;
  assign n7398 = n7397 ^ n7152;
  assign n7395 = n7147 ^ n7128;
  assign n7396 = ~n7360 & n7395;
  assign n7399 = n7398 ^ n7396;
  assign n7400 = n7324 & ~n7399;
  assign n7401 = n7400 ^ n7398;
  assign n7402 = ~n7394 & n7401;
  assign n7403 = n7158 ^ n7134;
  assign n7404 = n7403 ^ n7365;
  assign n7405 = n7360 & ~n7404;
  assign n7406 = n7405 ^ n7365;
  assign n7407 = ~n7380 & n7406;
  assign n7408 = n7402 & ~n7407;
  assign n7409 = ~n7390 & n7408;
  assign n7410 = ~n7383 & n7409;
  assign n7411 = ~n7382 & n7410;
  assign n7412 = ~n7381 & n7411;
  assign n7413 = ~n7377 & n7412;
  assign n7414 = ~n7373 & n7413;
  assign n7415 = ~n7370 & n7414;
  assign n7416 = ~n7363 & n7415;
  assign n7417 = n7416 ^ n5765;
  assign n10315 = n7417 ^ x374;
  assign n10316 = n10315 ^ n10314;
  assign n10317 = ~n10314 & n10316;
  assign n10331 = ~n10288 & n10317;
  assign n10320 = n10288 ^ n10286;
  assign n10321 = n10320 ^ n10287;
  assign n10322 = n10317 & n10321;
  assign n10346 = n10331 ^ n10322;
  assign n7734 = n7733 ^ n7698;
  assign n7735 = ~n7567 & ~n7734;
  assign n7736 = n7735 ^ n7698;
  assign n7737 = n7566 & ~n7736;
  assign n7748 = n7712 & ~n7747;
  assign n7749 = ~n7569 & ~n7717;
  assign n7752 = ~n7731 & ~n7749;
  assign n7753 = n7752 ^ n7706;
  assign n7750 = n7749 ^ n7726;
  assign n7751 = ~n7747 & ~n7750;
  assign n7754 = n7753 ^ n7751;
  assign n7755 = n7754 ^ n7569;
  assign n7756 = n7697 ^ n7683;
  assign n7757 = n7756 ^ n7747;
  assign n7758 = n7754 & n7757;
  assign n7759 = n7758 ^ n7747;
  assign n7760 = ~n7755 & ~n7759;
  assign n7761 = n7760 ^ n7569;
  assign n7762 = ~n7748 & ~n7761;
  assign n7766 = n7765 ^ n7704;
  assign n7768 = n7767 ^ n7766;
  assign n7769 = n7768 ^ n7687;
  assign n7770 = ~n7566 & ~n7769;
  assign n7771 = n7770 ^ n7687;
  assign n7772 = n7763 & n7771;
  assign n7773 = n7762 & ~n7772;
  assign n7774 = ~n7745 & n7773;
  assign n7775 = ~n7741 & n7774;
  assign n7776 = ~n7737 & n7775;
  assign n7777 = ~n7723 & n7776;
  assign n7778 = n7777 ^ n5953;
  assign n10255 = n7778 ^ x375;
  assign n8759 = n8758 ^ n8711;
  assign n8748 = n8733 ^ n8716;
  assign n8749 = n8748 ^ n8707;
  assign n8746 = n8695 ^ n8693;
  assign n8747 = n8746 ^ n8689;
  assign n8750 = n8749 ^ n8747;
  assign n8760 = n8759 ^ n8750;
  assign n8761 = ~n8724 & ~n8760;
  assign n8762 = n8761 ^ n8759;
  assign n8763 = n8723 & n8762;
  assign n8770 = ~n8722 & ~n8726;
  assign n8768 = ~n8720 & ~n8723;
  assign n8765 = n8764 ^ n8747;
  assign n8766 = n8765 ^ n8756;
  assign n8767 = n8727 & ~n8766;
  assign n8769 = n8768 ^ n8767;
  assign n8771 = n8770 ^ n8769;
  assign n8772 = n8767 ^ n8754;
  assign n8773 = n8771 ^ n8725;
  assign n8774 = ~n8772 & ~n8773;
  assign n8775 = n8774 ^ n8725;
  assign n8776 = ~n8771 & n8775;
  assign n8777 = ~n8763 & n8776;
  assign n8778 = ~n8745 & n8777;
  assign n8779 = ~n8729 & n8778;
  assign n8780 = n8779 ^ n5912;
  assign n10256 = n8780 ^ x370;
  assign n10333 = n10315 ^ n10257;
  assign n10358 = n10314 ^ n10286;
  assign n10359 = ~n10315 & ~n10358;
  assign n10360 = n10359 ^ n10314;
  assign n10361 = ~n10333 & n10360;
  assign n10341 = n10314 ^ n10257;
  assign n10357 = n10341 ^ n10286;
  assign n10362 = n10361 ^ n10357;
  assign n10334 = n10333 ^ n10286;
  assign n10335 = ~n10286 & ~n10334;
  assign n10336 = n10335 ^ n10315;
  assign n10337 = ~n10314 & ~n10336;
  assign n10338 = n10337 ^ n10334;
  assign n10797 = n10362 ^ n10338;
  assign n10798 = ~n10256 & n10797;
  assign n10799 = n10798 ^ n10362;
  assign n10325 = n10317 ^ n10314;
  assign n10326 = n10325 ^ n10315;
  assign n10327 = n10257 & n10326;
  assign n10328 = n10322 ^ n10317;
  assign n10329 = n10328 ^ n10287;
  assign n10330 = ~n10327 & ~n10329;
  assign n10791 = n10330 ^ n10322;
  assign n10347 = n10317 ^ n10315;
  assign n10348 = ~n10257 & n10347;
  assign n10339 = ~n10321 & ~n10338;
  assign n10349 = n10339 ^ n10315;
  assign n10350 = ~n10348 & n10349;
  assign n10351 = n10350 ^ n10346;
  assign n10792 = n10791 ^ n10351;
  assign n10793 = n10256 & n10792;
  assign n10794 = n10793 ^ n10791;
  assign n10795 = n10794 ^ n10351;
  assign n10796 = n10795 ^ n10350;
  assign n10800 = n10799 ^ n10796;
  assign n10801 = ~n10255 & ~n10800;
  assign n10802 = n10801 ^ n10799;
  assign n10803 = ~n10346 & ~n10802;
  assign n10804 = n10803 ^ n5971;
  assign n11501 = n10804 ^ x401;
  assign n7023 = n7022 ^ x381;
  assign n7418 = n7417 ^ x376;
  assign n8389 = n7023 & n7418;
  assign n8390 = n8389 ^ n7023;
  assign n8391 = n8390 ^ n7418;
  assign n8392 = n8391 ^ n7023;
  assign n7779 = n7778 ^ x377;
  assign n7997 = n7996 ^ n7994;
  assign n7998 = ~n7975 & ~n7997;
  assign n8010 = n7821 & ~n8009;
  assign n8011 = ~n7972 & ~n7974;
  assign n8012 = n7821 & n7970;
  assign n8013 = n7992 ^ n7978;
  assign n8015 = n8014 ^ n8013;
  assign n8016 = n8015 ^ n7990;
  assign n8017 = n8016 ^ n7990;
  assign n8018 = n7791 & n8017;
  assign n8019 = n8018 ^ n7990;
  assign n8020 = n7975 & n8019;
  assign n8021 = n8020 ^ n7990;
  assign n8034 = n8022 ^ n7989;
  assign n8035 = n7791 & n8034;
  assign n8036 = n8035 ^ n8022;
  assign n8029 = n8024 ^ n7977;
  assign n8030 = n8029 ^ n8004;
  assign n8026 = n8025 ^ n8022;
  assign n8027 = n8026 ^ n8004;
  assign n8028 = n8027 ^ n7969;
  assign n8031 = n8030 ^ n8028;
  assign n8032 = ~n7791 & n8031;
  assign n8033 = n8032 ^ n8028;
  assign n8037 = n8036 ^ n8033;
  assign n8038 = n8037 ^ n8033;
  assign n8039 = n8009 & ~n8038;
  assign n8040 = n8039 ^ n8033;
  assign n8041 = ~n7818 & ~n8040;
  assign n8042 = n8041 ^ n8033;
  assign n8043 = ~n8021 & ~n8042;
  assign n8044 = ~n8012 & n8043;
  assign n8045 = ~n8011 & n8044;
  assign n8046 = ~n8010 & n8045;
  assign n8047 = ~n8000 & n8046;
  assign n8048 = ~n7998 & n8047;
  assign n8049 = ~n7973 & n8048;
  assign n8050 = n8049 ^ n7223;
  assign n8051 = n8050 ^ x379;
  assign n8052 = n7779 & n8051;
  assign n8219 = n8218 ^ x380;
  assign n8332 = n8295 & n8331;
  assign n8334 = n8293 & ~n8333;
  assign n8336 = n8335 ^ n8334;
  assign n8337 = n8221 & n8314;
  assign n8338 = n8337 ^ n8313;
  assign n8339 = n8222 & n8338;
  assign n8345 = ~n8220 & n8319;
  assign n8346 = n8345 ^ n8322;
  assign n8347 = n8222 & n8346;
  assign n8348 = n8347 ^ n8322;
  assign n8349 = n8311 ^ n8288;
  assign n8350 = ~n8333 & n8349;
  assign n8359 = n8318 ^ n8298;
  assign n8358 = n8305 ^ n8300;
  assign n8360 = n8359 ^ n8358;
  assign n8361 = n8221 & n8360;
  assign n8362 = n8361 ^ n8359;
  assign n8353 = n8340 ^ n8300;
  assign n8354 = n8353 ^ n8302;
  assign n8351 = n8307 ^ n8302;
  assign n8352 = n8351 ^ n8315;
  assign n8355 = n8354 ^ n8352;
  assign n8356 = n8221 & ~n8355;
  assign n8357 = n8356 ^ n8352;
  assign n8363 = n8362 ^ n8357;
  assign n8364 = n8220 & ~n8363;
  assign n8365 = n8364 ^ n8362;
  assign n8366 = ~n8350 & ~n8365;
  assign n8367 = ~n8348 & n8366;
  assign n8368 = ~n8344 & n8367;
  assign n8369 = ~n8339 & n8368;
  assign n8370 = ~n8336 & n8369;
  assign n8371 = ~n8332 & n8370;
  assign n8372 = ~n8330 & n8371;
  assign n8373 = n8326 & n8372;
  assign n8374 = n8373 ^ n7185;
  assign n8375 = n8374 ^ x378;
  assign n8376 = ~n8219 & n8375;
  assign n8443 = n8052 & n8376;
  assign n8377 = n8376 ^ n8375;
  assign n8419 = ~n7779 & n8377;
  assign n8430 = n8419 ^ n8377;
  assign n8378 = n8052 & n8377;
  assign n8431 = n8430 ^ n8378;
  assign n10103 = n8443 ^ n8431;
  assign n10104 = n8392 & n10103;
  assign n8379 = n8052 ^ n7779;
  assign n8382 = n8379 ^ n8051;
  assign n8383 = n8377 ^ n8219;
  assign n8384 = ~n8382 & n8383;
  assign n8406 = n8384 ^ n8383;
  assign n8396 = n8052 & n8383;
  assign n8393 = n8379 & n8383;
  assign n8405 = n8396 ^ n8393;
  assign n8407 = n8406 ^ n8405;
  assign n10102 = n8389 & n8407;
  assign n10105 = n10104 ^ n10102;
  assign n8397 = n8376 ^ n8219;
  assign n8398 = n8052 & ~n8397;
  assign n11502 = n8398 ^ n8378;
  assign n11503 = ~n8391 & n11502;
  assign n8428 = n8376 & ~n8382;
  assign n10107 = n8428 ^ n8384;
  assign n8401 = n8382 ^ n7779;
  assign n8402 = n8376 & n8401;
  assign n11504 = n10107 ^ n8402;
  assign n11505 = n11504 ^ n8396;
  assign n11506 = n8392 & n11505;
  assign n8404 = n7418 ^ n7023;
  assign n8420 = n8051 & n8419;
  assign n8421 = n8420 ^ n8419;
  assign n8422 = n8421 ^ n8402;
  assign n10126 = n8422 ^ n8384;
  assign n8410 = ~n8397 & n8401;
  assign n10654 = ~n8392 & ~n8410;
  assign n11514 = ~n10126 & n10654;
  assign n8408 = n8379 & ~n8397;
  assign n8409 = n8408 ^ n8398;
  assign n11509 = n8443 ^ n8409;
  assign n11510 = n11509 ^ n8378;
  assign n8429 = n8428 ^ n8420;
  assign n8411 = n8410 ^ n8409;
  assign n8412 = n8411 ^ n8397;
  assign n11507 = n8429 ^ n8412;
  assign n11508 = n11507 ^ n8384;
  assign n11511 = n11510 ^ n11508;
  assign n11512 = n7418 & ~n11511;
  assign n11513 = n11512 ^ n11508;
  assign n11515 = n11514 ^ n11513;
  assign n11516 = n11515 ^ n11513;
  assign n11517 = n7023 & ~n11516;
  assign n11518 = n11517 ^ n11513;
  assign n11519 = n8404 & ~n11518;
  assign n11520 = n11519 ^ n11513;
  assign n11521 = ~n11506 & n11520;
  assign n11522 = ~n11503 & n11521;
  assign n11524 = n8429 ^ n8421;
  assign n8380 = n8376 & n8379;
  assign n11523 = n8431 ^ n8380;
  assign n11525 = n11524 ^ n11523;
  assign n11526 = n7418 & n11525;
  assign n11527 = n11526 ^ n11523;
  assign n11528 = n7023 & n11527;
  assign n11529 = n11522 & ~n11528;
  assign n8417 = n8408 ^ n8393;
  assign n11530 = ~n7023 & n8417;
  assign n11531 = n11530 ^ n8405;
  assign n11532 = n7418 & n11531;
  assign n11533 = n11532 ^ n8405;
  assign n11534 = n11529 & ~n11533;
  assign n11535 = ~n10105 & n11534;
  assign n11536 = n11535 ^ n7604;
  assign n11537 = n11536 ^ x403;
  assign n11538 = n11501 & n11537;
  assign n11539 = n11538 ^ n11501;
  assign n11540 = ~n11500 & n11539;
  assign n9144 = ~n8221 & n8286;
  assign n9145 = n9144 ^ n8300;
  assign n9146 = n8222 & n9145;
  assign n9147 = n9146 ^ n8300;
  assign n9148 = n8298 & n8628;
  assign n9149 = n8304 ^ n8295;
  assign n9150 = ~n8333 & n9149;
  assign n9155 = n8293 ^ n8291;
  assign n9156 = n9155 ^ n8286;
  assign n9157 = n9156 ^ n8319;
  assign n9158 = ~n8220 & n9157;
  assign n9159 = n9158 ^ n8319;
  assign n9151 = n8293 ^ n8288;
  assign n9152 = n8628 & n9151;
  assign n9153 = n9152 ^ n8335;
  assign n9154 = n9153 ^ n8313;
  assign n9160 = n9159 ^ n9154;
  assign n9161 = n9160 ^ n9154;
  assign n9162 = ~n8302 & ~n9161;
  assign n9163 = n9162 ^ n9154;
  assign n9164 = n8222 & ~n9163;
  assign n9165 = n9164 ^ n9154;
  assign n9166 = ~n9150 & ~n9165;
  assign n9167 = ~n9148 & n9166;
  assign n9169 = n8359 ^ n8307;
  assign n9168 = n8340 ^ n8311;
  assign n9170 = n9169 ^ n9168;
  assign n9171 = n8221 & ~n9170;
  assign n9172 = n9171 ^ n9168;
  assign n9173 = n8222 & n9172;
  assign n9174 = n9167 & ~n9173;
  assign n9175 = ~n8350 & n9174;
  assign n9176 = ~n8348 & n9175;
  assign n9177 = ~n9147 & n9176;
  assign n9178 = ~n8629 & n9177;
  assign n9179 = ~n8332 & n9178;
  assign n9180 = ~n8330 & n9179;
  assign n9181 = n9180 ^ n6220;
  assign n9182 = n9181 ^ x394;
  assign n8649 = n8192 ^ n8189;
  assign n9185 = n8649 ^ n8200;
  assign n9186 = ~n8075 & ~n9185;
  assign n9187 = n9186 ^ n8649;
  assign n9183 = n8075 & ~n8210;
  assign n9184 = n9183 ^ n8209;
  assign n9188 = n9187 ^ n9184;
  assign n9189 = ~n8074 & ~n9188;
  assign n9190 = n9189 ^ n9187;
  assign n9191 = ~n8179 & n9190;
  assign n9192 = n9191 ^ n6454;
  assign n9193 = n9192 ^ x399;
  assign n9330 = ~n9182 & n9193;
  assign n9331 = n9330 ^ n9193;
  assign n9355 = n9331 ^ n9182;
  assign n9356 = n9355 ^ n9193;
  assign n9195 = n7820 & ~n8009;
  assign n9196 = n7975 & n7992;
  assign n8820 = n7819 & ~n8006;
  assign n8821 = n8820 ^ n8010;
  assign n9202 = n8025 ^ n7967;
  assign n9203 = n9202 ^ n8003;
  assign n9204 = ~n7791 & n9203;
  assign n9205 = n9204 ^ n9202;
  assign n9199 = ~n7974 & n8025;
  assign n9200 = n9199 ^ n7968;
  assign n9197 = n7979 ^ n7970;
  assign n9198 = n9197 ^ n8024;
  assign n9201 = n9200 ^ n9198;
  assign n9206 = n9205 ^ n9201;
  assign n9207 = n7975 & n9206;
  assign n9208 = n9207 ^ n9201;
  assign n9209 = ~n8821 & ~n9208;
  assign n9210 = ~n9196 & n9209;
  assign n9211 = ~n9195 & n9210;
  assign n9212 = n8004 ^ n8002;
  assign n9213 = n7818 & n9212;
  assign n9214 = n9213 ^ n8002;
  assign n9215 = ~n7791 & n9214;
  assign n9216 = n9211 & ~n9215;
  assign n9217 = ~n9066 & n9216;
  assign n9218 = ~n8819 & n9217;
  assign n9219 = ~n7973 & n9218;
  assign n9220 = n9219 ^ n6011;
  assign n9221 = n9220 ^ x395;
  assign n9252 = ~n7700 & ~n7747;
  assign n9256 = n7718 ^ n7699;
  assign n9253 = n7707 & n7747;
  assign n9254 = n7749 & n7764;
  assign n9255 = ~n9253 & ~n9254;
  assign n9257 = n9256 ^ n9255;
  assign n9258 = n9257 ^ n9255;
  assign n9259 = n7566 & n9258;
  assign n9260 = n9259 ^ n9255;
  assign n9261 = n7763 & n9260;
  assign n9262 = n9261 ^ n9255;
  assign n9263 = ~n9252 & ~n9262;
  assign n9264 = n7709 ^ n7606;
  assign n9265 = n9264 ^ n7683;
  assign n9266 = n9265 ^ n7683;
  assign n9267 = ~n7566 & n9266;
  assign n9268 = n9267 ^ n7683;
  assign n9269 = n7763 & n9268;
  assign n9270 = n9269 ^ n7683;
  assign n9271 = n9263 & ~n9270;
  assign n9273 = n7567 & n7692;
  assign n9272 = n7569 & n7684;
  assign n9274 = n9273 ^ n9272;
  assign n9275 = n9271 & ~n9274;
  assign n9276 = ~n7737 & n9275;
  assign n9277 = ~n7723 & n9276;
  assign n9278 = ~n8785 & n9277;
  assign n9279 = ~n8784 & n9278;
  assign n9280 = n9279 ^ n7472;
  assign n9281 = n9280 ^ x397;
  assign n9224 = ~n7360 & ~n7392;
  assign n9225 = n9224 ^ n7367;
  assign n9226 = ~n7380 & ~n9225;
  assign n9227 = n9226 ^ n7367;
  assign n9229 = n7163 & n7361;
  assign n9228 = n7144 & n7360;
  assign n9230 = n9229 ^ n9228;
  assign n9231 = n9227 & ~n9230;
  assign n9233 = n7368 & ~n9232;
  assign n9234 = ~n7137 & n7369;
  assign n9235 = n9234 ^ n7362;
  assign n9237 = n7148 ^ n7132;
  assign n9236 = n7379 ^ n7160;
  assign n9238 = n9237 ^ n9236;
  assign n9239 = ~n9234 & ~n9238;
  assign n9240 = n9239 ^ n9236;
  assign n9241 = ~n9235 & ~n9240;
  assign n9242 = n9241 ^ n7362;
  assign n9243 = ~n9233 & ~n9242;
  assign n9244 = n9231 & n9243;
  assign n9245 = ~n9223 & n9244;
  assign n9246 = ~n8998 & n9245;
  assign n9247 = ~n7363 & n9246;
  assign n9248 = ~n7372 & n9247;
  assign n9249 = n9248 ^ n7449;
  assign n9250 = n9249 ^ x396;
  assign n9332 = n9281 ^ n9250;
  assign n9333 = ~n9221 & n9332;
  assign n9251 = ~n9221 & ~n9250;
  assign n9318 = n9251 ^ n9221;
  assign n9361 = n9333 ^ n9318;
  assign n9289 = n8754 ^ n8731;
  assign n9290 = n9289 ^ n8725;
  assign n9291 = n8727 ^ n8722;
  assign n9292 = ~n9289 & n9291;
  assign n9293 = n9292 ^ n8727;
  assign n9294 = n9290 & n9293;
  assign n9295 = n9294 ^ n8725;
  assign n9297 = n8723 & n9296;
  assign n9298 = n9297 ^ n8758;
  assign n9299 = n8724 & n9298;
  assign n9300 = ~n9295 & ~n9299;
  assign n9301 = n8753 ^ n8719;
  assign n9302 = n8723 & ~n9301;
  assign n9303 = n8711 ^ n8702;
  assign n9304 = n8724 & n9303;
  assign n9305 = ~n9302 & ~n9304;
  assign n9306 = ~n8726 & ~n8750;
  assign n9307 = n9305 & ~n9306;
  assign n9308 = n9300 & n9307;
  assign n9309 = n9288 & n9308;
  assign n9310 = ~n8729 & n9309;
  assign n9311 = n9310 ^ n6392;
  assign n9312 = n9311 ^ x398;
  assign n9313 = n9281 & n9312;
  assign n9322 = n9251 & n9313;
  assign n9323 = n9322 ^ n9313;
  assign n9319 = n9318 ^ n9250;
  assign n9320 = n9313 & ~n9319;
  assign n9316 = n9251 ^ n9250;
  assign n9317 = n9313 & ~n9316;
  assign n9321 = n9320 ^ n9317;
  assign n9324 = n9323 ^ n9321;
  assign n9314 = n9313 ^ n9281;
  assign n9315 = n9251 & n9314;
  assign n9325 = n9324 ^ n9315;
  assign n9326 = n9325 ^ n9322;
  assign n9362 = n9361 ^ n9326;
  assign n9363 = ~n9356 & ~n9362;
  assign n9194 = n9193 ^ n9182;
  assign n9338 = n9312 ^ n9281;
  assign n9339 = ~n9250 & ~n9338;
  assign n9340 = n9339 ^ n9322;
  assign n9341 = n9340 ^ n9317;
  assign n9336 = n9314 ^ n9312;
  assign n9364 = n9341 ^ n9336;
  assign n9352 = n9320 ^ n9319;
  assign n9348 = n9332 ^ n9221;
  assign n9334 = n9313 ^ n9312;
  assign n9343 = ~n9319 & n9334;
  assign n9349 = n9348 ^ n9343;
  assign n9337 = n9251 & ~n9336;
  assign n9342 = n9341 ^ n9337;
  assign n9344 = n9343 ^ n9342;
  assign n9345 = n9344 ^ n9320;
  assign n9335 = ~n9316 & n9334;
  assign n9346 = n9345 ^ n9335;
  assign n9347 = n9346 ^ n9333;
  assign n9350 = n9349 ^ n9347;
  assign n9351 = n9350 ^ n9343;
  assign n9353 = n9352 ^ n9351;
  assign n9365 = n9364 ^ n9353;
  assign n9366 = n9365 ^ n9324;
  assign n10011 = n9366 ^ n9318;
  assign n10012 = n10011 ^ n9362;
  assign n10014 = n10012 ^ n9351;
  assign n10015 = ~n9182 & n10014;
  assign n10016 = n10015 ^ n10012;
  assign n10017 = n9194 & n10016;
  assign n10013 = ~n9356 & n10012;
  assign n10018 = n10017 ^ n10013;
  assign n10019 = n9362 ^ n9342;
  assign n10020 = ~n9182 & ~n10019;
  assign n10021 = n10020 ^ n9362;
  assign n10022 = n9193 & ~n10021;
  assign n10023 = n9337 & n9355;
  assign n10024 = n9317 & n9330;
  assign n9354 = n9331 & ~n9353;
  assign n9367 = n9366 ^ n9321;
  assign n9368 = ~n9182 & n9367;
  assign n9369 = n9368 ^ n9321;
  assign n9370 = n9194 & n9369;
  assign n9357 = n9221 & ~n9312;
  assign n9358 = n9357 ^ n9319;
  assign n9359 = n9358 ^ n9345;
  assign n10026 = n9355 & ~n9359;
  assign n10025 = n9331 & n9335;
  assign n10027 = n10026 ^ n10025;
  assign n10028 = n9356 ^ n9320;
  assign n10029 = n9344 ^ n9331;
  assign n10030 = ~n9320 & ~n10029;
  assign n10031 = n10030 ^ n9331;
  assign n10032 = ~n10028 & n10031;
  assign n10033 = n10032 ^ n9356;
  assign n10034 = n9353 ^ n9315;
  assign n10035 = n9182 & ~n10034;
  assign n10036 = n10035 ^ n9354;
  assign n10037 = n10033 & ~n10036;
  assign n10038 = n9350 ^ n9322;
  assign n10039 = ~n9194 & n10038;
  assign n10041 = n9251 & n9334;
  assign n10040 = n10012 ^ n9315;
  assign n10042 = n10041 ^ n10040;
  assign n10043 = n9330 & n10042;
  assign n10044 = n10043 ^ n10041;
  assign n10045 = ~n10039 & ~n10044;
  assign n10046 = n10037 & n10045;
  assign n10047 = ~n10027 & n10046;
  assign n10048 = ~n9370 & n10047;
  assign n10049 = ~n9354 & n10048;
  assign n10050 = ~n10024 & n10049;
  assign n10051 = ~n10023 & n10050;
  assign n10052 = ~n10022 & n10051;
  assign n10053 = ~n10018 & n10052;
  assign n10054 = ~n9363 & n10053;
  assign n10055 = n10054 ^ n7565;
  assign n11541 = n10055 ^ x405;
  assign n9429 = n9220 ^ x393;
  assign n9428 = n9427 ^ x388;
  assign n9514 = n9429 ^ n9428;
  assign n9430 = n9181 ^ x392;
  assign n9437 = ~n5583 & ~n6970;
  assign n9438 = n9437 ^ n6975;
  assign n9439 = n5973 & n9438;
  assign n9440 = n9439 ^ n6975;
  assign n9448 = n5583 & n6937;
  assign n9443 = n6980 ^ n6972;
  assign n9444 = n9443 ^ n6994;
  assign n9441 = n6973 ^ n6952;
  assign n9442 = n9441 ^ n7007;
  assign n9445 = n9444 ^ n9442;
  assign n9446 = n5583 & ~n9445;
  assign n9447 = n9446 ^ n9442;
  assign n9449 = n9448 ^ n9447;
  assign n9450 = n5972 & n9449;
  assign n9451 = n9450 ^ n9447;
  assign n9452 = ~n9440 & ~n9451;
  assign n9453 = ~n6966 & n9452;
  assign n9454 = ~n6951 & n9453;
  assign n9455 = ~n9436 & n9454;
  assign n9456 = ~n9434 & n9455;
  assign n9457 = ~n6941 & n9456;
  assign n9458 = ~n8962 & n9457;
  assign n9459 = n9458 ^ n6256;
  assign n9460 = n9459 ^ x391;
  assign n9461 = ~n9430 & ~n9460;
  assign n9483 = n9482 ^ x389;
  assign n9484 = n8214 ^ n8074;
  assign n9485 = n9484 ^ n8216;
  assign n9486 = n9485 ^ n6186;
  assign n9487 = n9486 ^ x390;
  assign n9488 = ~n9483 & n9487;
  assign n9492 = n9488 ^ n9483;
  assign n9493 = n9492 ^ n9487;
  assign n9539 = n9461 & n9493;
  assign n9489 = n9488 ^ n9487;
  assign n9491 = n9461 ^ n9460;
  assign n9505 = n9491 ^ n9430;
  assign n9508 = n9489 & ~n9505;
  assign n9506 = n9505 ^ n9460;
  assign n9507 = n9493 & ~n9506;
  assign n9509 = n9508 ^ n9507;
  assign n9540 = n9539 ^ n9509;
  assign n9494 = ~n9491 & n9493;
  assign n9541 = n9540 ^ n9494;
  assign n9529 = n9487 ^ n9483;
  assign n9530 = n9529 ^ n9430;
  assign n9531 = n9530 ^ n9460;
  assign n9532 = n9531 ^ n9483;
  assign n9533 = n9532 ^ n9430;
  assign n9534 = n9483 ^ n9430;
  assign n9535 = n9460 & n9534;
  assign n9536 = n9535 ^ n9483;
  assign n9537 = ~n9533 & n9536;
  assign n9538 = n9537 ^ n9507;
  assign n9542 = n9541 ^ n9538;
  assign n9528 = n9461 & n9488;
  assign n9543 = n9542 ^ n9528;
  assign n9972 = n9429 & n9543;
  assign n9496 = ~n9491 & ~n9492;
  assign n9490 = n9461 & n9489;
  assign n9495 = n9494 ^ n9490;
  assign n9497 = n9496 ^ n9495;
  assign n9503 = n9497 ^ n9491;
  assign n9501 = n9489 & ~n9491;
  assign n9502 = n9501 ^ n9490;
  assign n9504 = n9503 ^ n9502;
  assign n9527 = n9504 ^ n9488;
  assign n9544 = n9543 ^ n9527;
  assign n9973 = n9972 ^ n9544;
  assign n9974 = ~n9514 & ~n9973;
  assign n9975 = n9974 ^ n9544;
  assign n9515 = n9429 & n9514;
  assign n9516 = n9515 ^ n9429;
  assign n9518 = n9508 ^ n9489;
  assign n9519 = n9518 ^ n9502;
  assign n9517 = n9507 ^ n9501;
  assign n9520 = n9519 ^ n9517;
  assign n9521 = n9516 & n9520;
  assign n10809 = n9495 & n9515;
  assign n10810 = n9509 ^ n9496;
  assign n9969 = n9516 ^ n9428;
  assign n10811 = n10810 ^ n9969;
  assign n10812 = n9515 ^ n9502;
  assign n10813 = ~n10810 & ~n10812;
  assign n10814 = n10813 ^ n9515;
  assign n10815 = n10811 & n10814;
  assign n10816 = n10815 ^ n9969;
  assign n10817 = n9494 ^ n9429;
  assign n10818 = n9516 & n10817;
  assign n10819 = n10818 ^ n9515;
  assign n10820 = n10819 ^ n9429;
  assign n10821 = n10820 ^ n9428;
  assign n9522 = ~n9492 & ~n9506;
  assign n9523 = n9522 ^ n9496;
  assign n9976 = n9523 ^ n9492;
  assign n9547 = n9505 ^ n9493;
  assign n9548 = n9547 ^ n9538;
  assign n9977 = n9976 ^ n9548;
  assign n10822 = n9977 ^ n9504;
  assign n10823 = n10821 & n10822;
  assign n10824 = n10823 ^ n9428;
  assign n10825 = ~n10816 & ~n10824;
  assign n9560 = n9537 ^ n9530;
  assign n9549 = n9548 ^ n9528;
  assign n10826 = n9560 ^ n9549;
  assign n10827 = ~n9429 & n10826;
  assign n10828 = n10827 ^ n9549;
  assign n10829 = ~n9428 & ~n10828;
  assign n10830 = n10825 & ~n10829;
  assign n10831 = ~n10809 & n10830;
  assign n10832 = ~n9521 & n10831;
  assign n10833 = n9975 & n10832;
  assign n10834 = n10833 ^ n6370;
  assign n11542 = n10834 ^ x400;
  assign n11543 = n11541 & n11542;
  assign n11544 = n11543 ^ n11541;
  assign n11545 = n11540 & n11544;
  assign n11737 = n11542 ^ n11541;
  assign n11548 = n11539 ^ n11537;
  assign n11563 = n11498 & ~n11548;
  assign n11555 = ~n11500 & ~n11548;
  assign n11564 = n11563 ^ n11555;
  assign n11550 = n11548 ^ n11501;
  assign n11556 = n11498 & n11550;
  assign n11565 = n11564 ^ n11556;
  assign n11566 = n11565 ^ n11501;
  assign n11559 = n11555 ^ n11550;
  assign n11557 = n11556 ^ n11555;
  assign n11552 = n11498 ^ n11496;
  assign n11553 = n11550 & ~n11552;
  assign n11551 = ~n11499 & n11550;
  assign n11554 = n11553 ^ n11551;
  assign n11558 = n11557 ^ n11554;
  assign n11560 = n11559 ^ n11558;
  assign n11561 = n11560 ^ n11554;
  assign n11549 = ~n11499 & ~n11548;
  assign n11562 = n11561 ^ n11549;
  assign n11567 = n11566 ^ n11562;
  assign n12110 = n11567 ^ n11560;
  assign n12111 = ~n11541 & ~n12110;
  assign n12112 = n12111 ^ n11560;
  assign n12113 = n11737 & n12112;
  assign n11578 = n11539 & ~n11552;
  assign n12114 = n11544 & n11578;
  assign n11546 = n11543 ^ n11542;
  assign n11547 = n11546 ^ n11541;
  assign n11588 = n11567 ^ n11549;
  assign n11569 = n11501 ^ n11497;
  assign n11570 = n11569 ^ n11537;
  assign n11571 = n11570 ^ n11501;
  assign n11572 = ~n11569 & ~n11571;
  assign n11573 = n11572 ^ n11570;
  assign n11574 = ~n11496 & n11573;
  assign n11575 = n11574 ^ n11563;
  assign n11568 = n11567 ^ n11556;
  assign n11576 = n11575 ^ n11568;
  assign n11597 = n11588 ^ n11576;
  assign n12115 = n11597 ^ n11553;
  assign n12116 = ~n11547 & n12115;
  assign n11601 = n11574 ^ n11570;
  assign n11590 = n11497 ^ n11496;
  assign n11591 = n11538 & n11590;
  assign n11592 = n11591 ^ n11538;
  assign n11602 = n11601 ^ n11592;
  assign n11600 = n11564 ^ n11551;
  assign n11603 = n11602 ^ n11600;
  assign n11595 = n11548 ^ n11498;
  assign n11596 = n11595 ^ n11557;
  assign n11598 = n11597 ^ n11596;
  assign n11579 = n11578 ^ n11539;
  assign n11577 = n11576 ^ n11540;
  assign n11580 = n11579 ^ n11577;
  assign n11594 = n11591 ^ n11580;
  assign n11599 = n11598 ^ n11594;
  assign n11604 = n11603 ^ n11599;
  assign n11581 = ~n11547 & ~n11580;
  assign n12117 = n11565 ^ n11553;
  assign n12118 = n11544 & n12117;
  assign n12119 = n11598 ^ n11577;
  assign n12120 = n12119 ^ n11562;
  assign n12121 = n11562 ^ n11543;
  assign n12122 = ~n11562 & ~n12121;
  assign n12123 = n12122 ^ n11562;
  assign n12124 = n12120 & ~n12123;
  assign n12125 = n12124 ^ n12122;
  assign n12126 = n12125 ^ n11562;
  assign n12127 = n12126 ^ n11543;
  assign n12128 = ~n12118 & ~n12127;
  assign n12129 = n12128 ^ n12118;
  assign n12130 = n11542 & n11602;
  assign n12131 = n12130 ^ n11592;
  assign n12132 = ~n11541 & n12131;
  assign n12133 = ~n12129 & ~n12132;
  assign n12134 = ~n11581 & n12133;
  assign n12135 = ~n11604 & n12134;
  assign n12136 = ~n12116 & n12135;
  assign n12137 = ~n12114 & n12136;
  assign n12138 = ~n12113 & n12137;
  assign n12139 = ~n11545 & n12138;
  assign n12140 = n12139 ^ n8812;
  assign n12934 = n12140 ^ x459;
  assign n8781 = n8780 ^ x368;
  assign n8813 = n8812 ^ x365;
  assign n8859 = n8781 & ~n8813;
  assign n8863 = n8859 ^ n8781;
  assign n8864 = n8863 ^ n8813;
  assign n8650 = ~n8074 & ~n8075;
  assign n8651 = n8650 ^ n8074;
  assign n8652 = n8649 & ~n8651;
  assign n8653 = ~n8200 & n8650;
  assign n8654 = ~n8179 & n8653;
  assign n8655 = ~n8652 & ~n8654;
  assign n8656 = n8209 ^ n8179;
  assign n8657 = n8656 ^ n8181;
  assign n8658 = n8075 & ~n8657;
  assign n8659 = n8658 ^ n8656;
  assign n8660 = n8074 & n8659;
  assign n8661 = n8655 & ~n8660;
  assign n8662 = n8661 ^ n6646;
  assign n8663 = n8662 ^ x366;
  assign n8823 = n8014 ^ n7971;
  assign n8824 = n7820 & ~n8823;
  assign n8831 = n8008 ^ n7988;
  assign n8832 = n8831 ^ n8026;
  assign n8826 = n7992 ^ n7969;
  assign n8825 = n7990 ^ n7977;
  assign n8827 = n8826 ^ n8825;
  assign n8828 = n8827 ^ n7979;
  assign n8829 = ~n7791 & n8828;
  assign n8830 = n8829 ^ n7979;
  assign n8833 = n8832 ^ n8830;
  assign n8834 = n8833 ^ n8830;
  assign n8835 = ~n7791 & n8834;
  assign n8836 = n8835 ^ n8830;
  assign n8837 = ~n7975 & n8836;
  assign n8838 = n8837 ^ n8830;
  assign n8839 = ~n8824 & ~n8838;
  assign n8840 = n8002 ^ n7969;
  assign n8841 = n8840 ^ n8005;
  assign n8842 = n8841 ^ n8005;
  assign n8843 = n7791 & n8842;
  assign n8844 = n8843 ^ n8005;
  assign n8845 = n7975 & n8844;
  assign n8846 = n8845 ^ n8005;
  assign n8847 = n8839 & ~n8846;
  assign n8848 = ~n7998 & n8847;
  assign n8849 = ~n8822 & n8848;
  assign n8850 = ~n8821 & n8849;
  assign n8851 = ~n8819 & n8850;
  assign n8852 = n8851 ^ n6631;
  assign n8853 = n8852 ^ x367;
  assign n8860 = n8663 & n8853;
  assign n8861 = n8860 ^ n8663;
  assign n8869 = n8861 ^ n8853;
  assign n8874 = n8869 ^ n8663;
  assign n8875 = n8864 & n8874;
  assign n8873 = n8853 & n8864;
  assign n8876 = n8875 ^ n8873;
  assign n8872 = n8663 & n8864;
  assign n8877 = n8876 ^ n8872;
  assign n8782 = n8781 ^ n8663;
  assign n8814 = n8813 ^ n8782;
  assign n8815 = n8813 ^ n8663;
  assign n8854 = n8853 ^ n8813;
  assign n8855 = ~n8815 & n8854;
  assign n8856 = ~n8814 & n8855;
  assign n8878 = n8877 ^ n8856;
  assign n8610 = n8609 ^ x364;
  assign n8647 = n8646 ^ x369;
  assign n10059 = n8610 & ~n8647;
  assign n10060 = n10059 ^ n8610;
  assign n10061 = n10060 ^ n8647;
  assign n10062 = n8878 & n10061;
  assign n8884 = n8853 ^ n8782;
  assign n8885 = ~n8815 & n8884;
  assign n8883 = n8860 & n8863;
  assign n8886 = n8885 ^ n8883;
  assign n8887 = n8886 ^ n8856;
  assign n8865 = n8864 ^ n8781;
  assign n8870 = ~n8865 & ~n8869;
  assign n8867 = n8859 & n8860;
  assign n8871 = n8870 ^ n8867;
  assign n8879 = n8878 ^ n8871;
  assign n8880 = n8879 ^ n8865;
  assign n8866 = n8861 & ~n8865;
  assign n8868 = n8867 ^ n8866;
  assign n8881 = n8880 ^ n8868;
  assign n8862 = n8859 & n8861;
  assign n8882 = n8881 ^ n8862;
  assign n8888 = n8887 ^ n8882;
  assign n8889 = n8888 ^ n8866;
  assign n8890 = n8889 ^ n8813;
  assign n8891 = n8890 ^ n8879;
  assign n10530 = n8891 & n10059;
  assign n10527 = n10059 ^ n8647;
  assign n10528 = n8862 & ~n10527;
  assign n8648 = n8647 ^ n8610;
  assign n10526 = n8648 & n8883;
  assign n10529 = n10528 ^ n10526;
  assign n10531 = n10530 ^ n10529;
  assign n10532 = n8870 & ~n10527;
  assign n8896 = n8863 & n8874;
  assign n10063 = n8896 ^ n8876;
  assign n8857 = n8856 ^ n8855;
  assign n8900 = n8891 ^ n8857;
  assign n8894 = n8872 ^ n8864;
  assign n8895 = n8894 ^ n8875;
  assign n8901 = n8900 ^ n8895;
  assign n10064 = n10063 ^ n8901;
  assign n10065 = n8610 & n10064;
  assign n10066 = n10065 ^ n10063;
  assign n10067 = ~n8648 & n10066;
  assign n10533 = n10532 ^ n10067;
  assign n8858 = ~n8610 & n8857;
  assign n8892 = n8891 ^ n8858;
  assign n8893 = ~n8648 & n8892;
  assign n10068 = ~n8881 & n10060;
  assign n10069 = ~n8893 & ~n10068;
  assign n10535 = n8891 ^ n8866;
  assign n10536 = n10535 ^ n8895;
  assign n8897 = n8896 ^ n8895;
  assign n8898 = n8897 ^ n8883;
  assign n8899 = n8898 ^ n8863;
  assign n8902 = n8901 ^ n8899;
  assign n8916 = n8902 ^ n8872;
  assign n10534 = n8916 ^ n8873;
  assign n10537 = n10536 ^ n10534;
  assign n10538 = n10537 ^ n10534;
  assign n10539 = ~n8610 & n10538;
  assign n10540 = n10539 ^ n10534;
  assign n10541 = ~n8648 & n10540;
  assign n10542 = n10541 ^ n10534;
  assign n10548 = n8647 & ~n8888;
  assign n10544 = n8882 ^ n8867;
  assign n10075 = n8875 ^ n8866;
  assign n10543 = n10075 ^ n8871;
  assign n10545 = n10544 ^ n10543;
  assign n10546 = ~n8647 & ~n10545;
  assign n10547 = n10546 ^ n10543;
  assign n10549 = n10548 ^ n10547;
  assign n10550 = ~n8610 & n10549;
  assign n10551 = n10550 ^ n10547;
  assign n10552 = ~n10542 & ~n10551;
  assign n10553 = n10069 & n10552;
  assign n10554 = ~n10533 & n10553;
  assign n10555 = ~n10531 & n10554;
  assign n10556 = ~n10062 & n10555;
  assign n10557 = n10556 ^ n7854;
  assign n10558 = n10557 ^ x434;
  assign n9498 = ~n9429 & n9497;
  assign n9499 = n9498 ^ n9495;
  assign n9500 = ~n9428 & n9499;
  assign n9985 = n9541 ^ n9483;
  assign n10559 = n9516 & n9985;
  assign n9552 = n9522 ^ n9504;
  assign n9970 = ~n9552 & n9969;
  assign n9524 = ~n9428 & n9523;
  assign n9525 = n9524 ^ n9496;
  assign n9526 = n9429 & n9525;
  assign n9971 = n9970 ^ n9526;
  assign n10560 = n9516 & n9977;
  assign n9993 = ~n9516 & ~n9539;
  assign n10562 = ~n9501 & n9993;
  assign n10563 = n9993 ^ n9505;
  assign n10564 = n10562 ^ n9493;
  assign n10565 = ~n10563 & n10564;
  assign n10566 = n10565 ^ n9493;
  assign n10567 = n10562 & n10566;
  assign n9986 = n9985 ^ n9518;
  assign n9996 = n9986 ^ n9539;
  assign n9980 = n9519 ^ n9501;
  assign n10561 = n9996 ^ n9980;
  assign n10568 = n10567 ^ n10561;
  assign n10569 = n9429 & ~n10568;
  assign n10570 = n10569 ^ n10561;
  assign n9555 = n9544 ^ n9542;
  assign n10571 = n10570 ^ n9555;
  assign n10572 = ~n9428 & ~n10571;
  assign n10573 = n10572 ^ n9555;
  assign n10574 = ~n10560 & n10573;
  assign n10575 = ~n9971 & n10574;
  assign n10576 = ~n10559 & n10575;
  assign n10577 = n9549 ^ n9522;
  assign n10578 = n10577 ^ n9541;
  assign n10579 = n9428 & ~n10578;
  assign n10580 = n10579 ^ n10577;
  assign n10581 = ~n9429 & ~n10580;
  assign n10582 = n10576 & ~n10581;
  assign n10583 = ~n9500 & n10582;
  assign n10584 = n10583 ^ n7928;
  assign n10585 = n10584 ^ x432;
  assign n10586 = n10558 & n10585;
  assign n9573 = n8993 ^ x357;
  assign n9572 = n9311 ^ x352;
  assign n9574 = n9573 ^ n9572;
  assign n9579 = ~n8564 & n9464;
  assign n9586 = n8483 ^ n8481;
  assign n9587 = n8533 ^ n8507;
  assign n9588 = n9586 & n9587;
  assign n9589 = n8452 & ~n9588;
  assign n9581 = n8541 ^ n8524;
  assign n9580 = n8595 ^ n8539;
  assign n9582 = n9581 ^ n9580;
  assign n9583 = n8560 & ~n9582;
  assign n9584 = n9583 ^ n9580;
  assign n9590 = n9589 ^ n9584;
  assign n9591 = ~n8565 & ~n9590;
  assign n9585 = n9584 ^ n8451;
  assign n9592 = n9591 ^ n9585;
  assign n9593 = n8552 ^ n8532;
  assign n9594 = n8452 & ~n9593;
  assign n9595 = n9594 ^ n8552;
  assign n9596 = n9595 ^ n8566;
  assign n9597 = ~n8565 & ~n9596;
  assign n9598 = n9597 ^ n9595;
  assign n9599 = n9592 & n9598;
  assign n9600 = ~n9579 & n9599;
  assign n9601 = ~n9578 & n9600;
  assign n9602 = ~n8581 & n9601;
  assign n9603 = ~n8586 & n9602;
  assign n9604 = ~n9462 & n9603;
  assign n9605 = n9604 ^ n6429;
  assign n9606 = n9605 ^ x355;
  assign n9632 = n9192 ^ x353;
  assign n9611 = n8340 ^ n8322;
  assign n9612 = n9611 ^ n8313;
  assign n9610 = n8319 ^ n8316;
  assign n9613 = n9612 ^ n9610;
  assign n9614 = ~n8221 & n9613;
  assign n9615 = n9614 ^ n9610;
  assign n9607 = n8300 ^ n8296;
  assign n9608 = ~n8221 & n9607;
  assign n9609 = n9608 ^ n8296;
  assign n9616 = n9615 ^ n9609;
  assign n9617 = n8222 & n9616;
  assign n9618 = n9617 ^ n9615;
  assign n9619 = ~n8621 & ~n9618;
  assign n9620 = ~n9147 & n9619;
  assign n9621 = ~n8615 & n9620;
  assign n9622 = ~n8339 & n9621;
  assign n9623 = ~n8336 & n9622;
  assign n9624 = ~n8629 & n9623;
  assign n9625 = ~n8332 & n9624;
  assign n9626 = n8326 & n9625;
  assign n9627 = n9626 ^ n6489;
  assign n9628 = n9627 ^ x354;
  assign n9643 = n9632 ^ n9628;
  assign n9633 = n9092 ^ x356;
  assign n9644 = n9643 ^ n9633;
  assign n9645 = ~n9606 & ~n9644;
  assign n9646 = n9645 ^ n9606;
  assign n9634 = n9632 & n9633;
  assign n9635 = n9634 ^ n9632;
  assign n9629 = n9606 & ~n9628;
  assign n9639 = n9629 ^ n9628;
  assign n9640 = n9635 & ~n9639;
  assign n9630 = n9629 ^ n9606;
  assign n9631 = n9630 ^ n9628;
  assign n9638 = n9631 & n9634;
  assign n9641 = n9640 ^ n9638;
  assign n9636 = n9635 ^ n9633;
  assign n9637 = n9631 & ~n9636;
  assign n9642 = n9641 ^ n9637;
  assign n9647 = n9646 ^ n9642;
  assign n9648 = n9647 ^ n9637;
  assign n9649 = n9573 & ~n9648;
  assign n9650 = n9649 ^ n9647;
  assign n9651 = ~n9574 & ~n9650;
  assign n9658 = n9630 & n9635;
  assign n10587 = n9658 ^ n9638;
  assign n10588 = n9572 & n10587;
  assign n10589 = n10588 ^ n9658;
  assign n10590 = ~n9574 & n10589;
  assign n9652 = n9572 & ~n9573;
  assign n9653 = n9652 ^ n9572;
  assign n9938 = n9653 ^ n9573;
  assign n9675 = ~n9636 & ~n9639;
  assign n9700 = n9675 ^ n9636;
  assign n9666 = n9630 & ~n9636;
  assign n9697 = n9666 ^ n9637;
  assign n9701 = n9700 ^ n9697;
  assign n9939 = n9701 ^ n9647;
  assign n9940 = n9938 & n9939;
  assign n9678 = n9630 & n9634;
  assign n9693 = n9653 & n9678;
  assign n9941 = n9940 ^ n9693;
  assign n10591 = n9632 & n9938;
  assign n10592 = n9630 & n10591;
  assign n9667 = n9666 ^ n9647;
  assign n9663 = n9633 ^ n9606;
  assign n9664 = n9644 & n9663;
  assign n9665 = n9664 ^ n9638;
  assign n9668 = n9667 ^ n9665;
  assign n9942 = n9653 & ~n9668;
  assign n10593 = n10592 ^ n9942;
  assign n9684 = n9667 ^ n9630;
  assign n9682 = n9658 ^ n9647;
  assign n9683 = n9682 ^ n9678;
  assign n9685 = n9684 ^ n9683;
  assign n9686 = n9685 ^ n9675;
  assign n9687 = n9686 ^ n9641;
  assign n9688 = ~n9573 & n9687;
  assign n9689 = n9688 ^ n9686;
  assign n9676 = n9675 ^ n9645;
  assign n9656 = n9634 & ~n9639;
  assign n9655 = n9631 & n9635;
  assign n9657 = n9656 ^ n9655;
  assign n9677 = n9676 ^ n9657;
  assign n9679 = n9678 ^ n9677;
  assign n9680 = ~n9573 & n9679;
  assign n9681 = n9680 ^ n9677;
  assign n9690 = n9689 ^ n9681;
  assign n9691 = ~n9572 & n9690;
  assign n9692 = n9691 ^ n9689;
  assign n9662 = n9629 & n9634;
  assign n9669 = n9668 ^ n9662;
  assign n9699 = n9669 ^ n9629;
  assign n9702 = n9701 ^ n9699;
  assign n10599 = n9702 ^ n9645;
  assign n9959 = n9702 ^ n9666;
  assign n10600 = n10599 ^ n9959;
  assign n10601 = ~n9572 & n10600;
  assign n10602 = n10601 ^ n9959;
  assign n9694 = n9662 ^ n9655;
  assign n10594 = n9939 ^ n9694;
  assign n10595 = n10594 ^ n9959;
  assign n10596 = n10595 ^ n9642;
  assign n10597 = n9572 & n10596;
  assign n10598 = n10597 ^ n9642;
  assign n10603 = n10602 ^ n10598;
  assign n10604 = ~n9574 & n10603;
  assign n10605 = n10604 ^ n10598;
  assign n10606 = ~n9692 & ~n10605;
  assign n10607 = ~n10593 & n10606;
  assign n10608 = ~n9941 & n10607;
  assign n10609 = ~n10590 & n10608;
  assign n10610 = ~n9651 & n10609;
  assign n10611 = n10610 ^ n7889;
  assign n10612 = n10611 ^ x433;
  assign n9327 = n9182 & n9326;
  assign n9328 = n9327 ^ n9322;
  assign n9329 = ~n9194 & n9328;
  assign n9360 = ~n9356 & ~n9359;
  assign n10215 = n10041 ^ n9362;
  assign n10216 = n10215 ^ n9320;
  assign n10217 = n9193 & ~n10216;
  assign n10218 = n10217 ^ n9320;
  assign n10219 = ~n9182 & n10218;
  assign n10220 = n9182 & n9317;
  assign n10221 = n10041 ^ n9353;
  assign n10222 = ~n9356 & ~n10221;
  assign n10223 = n9337 ^ n9194;
  assign n10224 = n9335 ^ n9182;
  assign n10225 = ~n9337 & ~n10224;
  assign n10226 = n10225 ^ n9182;
  assign n10227 = ~n10223 & ~n10226;
  assign n10228 = n10227 ^ n9337;
  assign n9379 = n9366 ^ n9344;
  assign n10229 = n9379 ^ n9320;
  assign n10230 = n9182 & n10229;
  assign n10231 = n10230 ^ n9320;
  assign n10232 = n9194 & n10231;
  assign n10233 = ~n10228 & ~n10232;
  assign n10234 = ~n10222 & n10233;
  assign n10235 = ~n10220 & n10234;
  assign n10236 = n10012 ^ n9359;
  assign n10237 = n10236 ^ n9365;
  assign n10238 = ~n9182 & ~n10237;
  assign n10239 = n10238 ^ n9365;
  assign n10240 = n9193 & n10239;
  assign n10241 = n10235 & ~n10240;
  assign n10242 = ~n10026 & n10241;
  assign n10243 = ~n10017 & n10242;
  assign n10244 = ~n10022 & n10243;
  assign n10245 = ~n10219 & n10244;
  assign n10246 = ~n9363 & n10245;
  assign n10247 = ~n9360 & n10246;
  assign n10248 = ~n9354 & n10247;
  assign n10249 = ~n9329 & n10248;
  assign n10250 = n10249 ^ n7962;
  assign n10613 = n10250 ^ x431;
  assign n10614 = n10612 & n10613;
  assign n10636 = n10614 ^ n10612;
  assign n10644 = n10586 & n10636;
  assign n10645 = n10644 ^ n10636;
  assign n10616 = n10586 ^ n10585;
  assign n10642 = n10616 & n10636;
  assign n10637 = n10586 ^ n10558;
  assign n10638 = n10636 & n10637;
  assign n10643 = n10642 ^ n10638;
  assign n10646 = n10645 ^ n10643;
  assign n10625 = n10585 & n10613;
  assign n10626 = n10625 ^ n10614;
  assign n10620 = n10614 ^ n10613;
  assign n10623 = n10616 & n10620;
  assign n10621 = n10586 & n10620;
  assign n10617 = n10616 ^ n10558;
  assign n10618 = n10614 & ~n10617;
  assign n10622 = n10621 ^ n10618;
  assign n10624 = n10623 ^ n10622;
  assign n10627 = n10626 ^ n10624;
  assign n10640 = n10637 ^ n10627;
  assign n10632 = n10585 ^ n10558;
  assign n10633 = n10613 & n10632;
  assign n10634 = n10633 ^ n10627;
  assign n10628 = n10627 ^ n10614;
  assign n10615 = n10586 & n10614;
  assign n10619 = n10618 ^ n10615;
  assign n10629 = n10628 ^ n10619;
  assign n10630 = n10629 ^ n10622;
  assign n10631 = n10630 ^ n10624;
  assign n10635 = n10634 ^ n10631;
  assign n10639 = n10638 ^ n10635;
  assign n10641 = n10640 ^ n10639;
  assign n10647 = n10646 ^ n10641;
  assign n10352 = n10317 ^ n10287;
  assign n10318 = ~n10286 & n10317;
  assign n10353 = n10352 ^ n10318;
  assign n10363 = n10362 ^ n10353;
  assign n10354 = n10353 ^ n10351;
  assign n10355 = n10354 ^ n10334;
  assign n10332 = n10331 ^ n10330;
  assign n10340 = n10339 ^ n10332;
  assign n10342 = n10341 ^ n10340;
  assign n10356 = n10355 ^ n10342;
  assign n10364 = n10363 ^ n10356;
  assign n10365 = n10364 ^ n10357;
  assign n10366 = n10365 ^ n10355;
  assign n10367 = ~n10256 & ~n10366;
  assign n10368 = n10367 ^ n10355;
  assign n10319 = n10318 ^ n10288;
  assign n10323 = n10322 ^ n10319;
  assign n10324 = n10323 ^ n10316;
  assign n10343 = n10342 ^ n10324;
  assign n10344 = ~n10256 & ~n10343;
  assign n10345 = n10344 ^ n10324;
  assign n10369 = n10368 ^ n10345;
  assign n10370 = ~n10255 & n10369;
  assign n10371 = n10370 ^ n10368;
  assign n10372 = n10371 ^ n7790;
  assign n10648 = n10372 ^ x430;
  assign n8413 = n8412 ^ n8407;
  assign n8414 = ~n7418 & ~n8413;
  assign n8415 = n8414 ^ n8407;
  assign n8416 = n8404 & n8415;
  assign n8381 = n8380 ^ n8378;
  assign n10096 = n8407 ^ n8381;
  assign n10097 = n7418 & n10096;
  assign n10098 = n10097 ^ n8407;
  assign n10099 = n7023 & n10098;
  assign n8385 = n8384 ^ n8381;
  assign n8386 = ~n7418 & n8385;
  assign n8387 = n8386 ^ n8384;
  assign n8388 = n7023 & n8387;
  assign n10649 = n8422 ^ n8380;
  assign n10650 = n7023 & n10649;
  assign n10651 = n10650 ^ n8380;
  assign n10652 = ~n7418 & n10651;
  assign n8399 = n8398 ^ n8396;
  assign n10661 = n8428 ^ n8399;
  assign n10662 = n10661 ^ n8422;
  assign n10658 = ~n8391 & n8419;
  assign n10655 = n8398 ^ n8391;
  assign n10656 = n10655 ^ n8384;
  assign n10657 = ~n10654 & ~n10656;
  assign n10659 = n10658 ^ n10657;
  assign n10653 = n8412 ^ n8396;
  assign n10660 = n10659 ^ n10653;
  assign n10663 = n10662 ^ n10660;
  assign n10664 = n10663 ^ n10660;
  assign n10665 = n7418 & n10664;
  assign n10666 = n10665 ^ n10660;
  assign n10667 = n7023 & ~n10666;
  assign n10668 = n10667 ^ n10660;
  assign n10669 = ~n10652 & n10668;
  assign n10670 = ~n7023 & n8378;
  assign n10671 = n10670 ^ n8417;
  assign n10672 = n7418 & n10671;
  assign n10673 = n10672 ^ n8417;
  assign n10674 = n10669 & ~n10673;
  assign n10675 = ~n10104 & n10674;
  assign n10676 = ~n8388 & n10675;
  assign n10677 = ~n10099 & n10676;
  assign n10678 = ~n8416 & n10677;
  assign n10679 = n10678 ^ n7817;
  assign n10680 = n10679 ^ x435;
  assign n10681 = ~n10648 & ~n10680;
  assign n10682 = n10681 ^ n10680;
  assign n10683 = n10682 ^ n10648;
  assign n10684 = n10647 & ~n10683;
  assign n10685 = n10642 ^ n10616;
  assign n10686 = n10685 ^ n10631;
  assign n10687 = n10686 ^ n10644;
  assign n10688 = n10687 ^ n10641;
  assign n10689 = n10648 & n10688;
  assign n10690 = n10689 ^ n10641;
  assign n10691 = ~n10680 & n10690;
  assign n10692 = n10681 ^ n10648;
  assign n10693 = n10692 ^ n10682;
  assign n10694 = n10644 ^ n10619;
  assign n10695 = n10694 ^ n10586;
  assign n10696 = n10695 ^ n10622;
  assign n10697 = ~n10693 & n10696;
  assign n10703 = n10687 ^ n10646;
  assign n10699 = n10621 ^ n10620;
  assign n10698 = n10635 ^ n10623;
  assign n10700 = n10699 ^ n10698;
  assign n10701 = n10700 ^ n10629;
  assign n10702 = n10701 ^ n10638;
  assign n10704 = n10703 ^ n10702;
  assign n10705 = ~n10692 & n10704;
  assign n10706 = n10680 ^ n10630;
  assign n10707 = n10693 & n10706;
  assign n10708 = n10707 ^ n10680;
  assign n10709 = n10631 & ~n10708;
  assign n10710 = n10709 ^ n10624;
  assign n10711 = ~n10627 & ~n10710;
  assign n10712 = n10711 ^ n10698;
  assign n10713 = ~n10693 & ~n10712;
  assign n10714 = n10713 ^ n10698;
  assign n10715 = ~n10705 & ~n10714;
  assign n10717 = n10620 ^ n10612;
  assign n10718 = n10717 ^ n10696;
  assign n10716 = n10686 ^ n10641;
  assign n10719 = n10718 ^ n10716;
  assign n10720 = n10719 ^ n10619;
  assign n10721 = ~n10680 & ~n10720;
  assign n10722 = n10721 ^ n10719;
  assign n10723 = n10648 & ~n10722;
  assign n10724 = n10715 & ~n10723;
  assign n10725 = ~n10697 & n10724;
  assign n10726 = n10643 & ~n10648;
  assign n10727 = n10726 ^ n10638;
  assign n10728 = n10727 ^ n10700;
  assign n10729 = n10727 ^ n10680;
  assign n10730 = ~n10727 & n10729;
  assign n10731 = n10730 ^ n10727;
  assign n10732 = n10728 & ~n10731;
  assign n10733 = n10732 ^ n10730;
  assign n10734 = n10733 ^ n10727;
  assign n10735 = n10734 ^ n10680;
  assign n10736 = n10725 & n10735;
  assign n10737 = n10736 ^ n10725;
  assign n10738 = ~n10691 & n10737;
  assign n10739 = ~n10684 & n10738;
  assign n10740 = n10739 ^ n9092;
  assign n12933 = n10740 ^ x454;
  assign n13013 = n12934 ^ n12933;
  assign n10885 = n9878 & ~n9912;
  assign n10886 = n9888 ^ n9862;
  assign n10887 = n10886 ^ n9890;
  assign n10888 = n10886 ^ n9907;
  assign n10889 = n10886 & ~n10888;
  assign n10890 = n10889 ^ n10886;
  assign n10891 = n10887 & n10890;
  assign n10892 = n10891 ^ n10889;
  assign n10893 = n10892 ^ n10886;
  assign n10894 = n10893 ^ n9907;
  assign n10895 = ~n9884 & ~n10894;
  assign n10896 = n10895 ^ n9907;
  assign n10412 = n9886 & ~n9912;
  assign n10413 = n9869 ^ n9865;
  assign n10414 = n10413 ^ n9867;
  assign n10415 = n10414 ^ n9867;
  assign n10416 = ~n9890 & n10415;
  assign n10417 = n10416 ^ n9867;
  assign n10418 = n9907 & ~n10417;
  assign n10419 = n10418 ^ n9867;
  assign n10420 = ~n10412 & n10419;
  assign n10897 = n9855 & ~n9893;
  assign n10422 = n9874 ^ n9863;
  assign n10898 = n10422 ^ n9888;
  assign n10899 = n9892 & n10898;
  assign n10904 = n9876 ^ n9859;
  assign n10900 = n9914 ^ n9872;
  assign n10901 = n10900 ^ n9882;
  assign n10902 = n9891 & n10901;
  assign n10903 = n10902 ^ n10900;
  assign n10905 = n10904 ^ n10903;
  assign n10906 = n10905 ^ n10903;
  assign n10907 = n9891 & n10906;
  assign n10908 = n10907 ^ n10903;
  assign n10909 = ~n9890 & n10908;
  assign n10910 = n10909 ^ n10903;
  assign n10911 = ~n10899 & ~n10910;
  assign n10912 = ~n10897 & n10911;
  assign n10913 = n10420 & n10912;
  assign n10914 = ~n9905 & n10913;
  assign n10915 = n10896 & n10914;
  assign n10916 = ~n10885 & n10915;
  assign n10917 = ~n9894 & n10916;
  assign n10918 = n10917 ^ n6923;
  assign n11050 = n10918 ^ x441;
  assign n11051 = n10557 ^ x436;
  assign n11010 = ~n9194 & n9250;
  assign n11011 = ~n9221 & n11010;
  assign n11012 = ~n9336 & n11011;
  assign n11013 = n9353 ^ n9335;
  assign n11014 = n9330 & ~n11013;
  assign n11015 = ~n9193 & n9340;
  assign n11016 = n11015 ^ n9322;
  assign n11017 = ~n9182 & n11016;
  assign n11018 = n11017 ^ n9322;
  assign n11024 = n9193 & n9325;
  assign n11020 = n10215 ^ n9345;
  assign n11019 = n9350 ^ n9344;
  assign n11021 = n11020 ^ n11019;
  assign n11022 = ~n9193 & ~n11021;
  assign n11023 = n11022 ^ n11019;
  assign n11025 = n11024 ^ n11023;
  assign n11026 = ~n9182 & n11025;
  assign n11027 = n11026 ^ n11023;
  assign n11028 = ~n11018 & ~n11027;
  assign n11029 = ~n10027 & n11028;
  assign n11030 = ~n10219 & n11029;
  assign n11031 = ~n9360 & n11030;
  assign n11032 = ~n11014 & n11031;
  assign n11033 = ~n11012 & n11032;
  assign n11034 = ~n10018 & n11033;
  assign n11035 = ~n9329 & n11034;
  assign n11036 = n11035 ^ n8687;
  assign n11037 = n11036 ^ x439;
  assign n9097 = n9096 ^ n9064;
  assign n9098 = n9063 & ~n9097;
  assign n10769 = n9064 & ~n9113;
  assign n10770 = n10769 ^ n9109;
  assign n10771 = n9093 & n10770;
  assign n10772 = n10771 ^ n9109;
  assign n9116 = n9111 ^ n9030;
  assign n10773 = n9093 & n9116;
  assign n10777 = n9049 ^ n9037;
  assign n10776 = n10775 ^ n9048;
  assign n10778 = n10777 ^ n10776;
  assign n10779 = ~n9093 & n10778;
  assign n10780 = n10779 ^ n10776;
  assign n10774 = n9046 ^ n9041;
  assign n10781 = n10780 ^ n10774;
  assign n10782 = n9094 & n10781;
  assign n10783 = n10782 ^ n10774;
  assign n10784 = ~n10773 & ~n10783;
  assign n10785 = ~n10772 & n10784;
  assign n10786 = ~n10768 & n10785;
  assign n10787 = n10764 & n10786;
  assign n10788 = ~n9098 & n10787;
  assign n10789 = n10788 ^ n5582;
  assign n11038 = n10789 ^ x440;
  assign n11039 = ~n11037 & ~n11038;
  assign n11040 = n11039 ^ n11038;
  assign n11042 = n10679 ^ x437;
  assign n11043 = n10345 ^ n10255;
  assign n11044 = n11043 ^ n10370;
  assign n11045 = n11044 ^ n8694;
  assign n11046 = n11045 ^ x438;
  assign n11047 = n11042 & ~n11046;
  assign n11048 = n11047 ^ n11042;
  assign n11049 = n11048 ^ n11046;
  assign n11069 = ~n11040 & n11049;
  assign n11041 = n11040 ^ n11037;
  assign n11064 = n11041 ^ n11038;
  assign n11065 = n11047 & ~n11064;
  assign n11070 = n11069 ^ n11065;
  assign n11084 = ~n11051 & n11070;
  assign n11085 = n11084 ^ n11065;
  assign n11086 = n11050 & n11085;
  assign n11117 = n11051 ^ n11050;
  assign n11299 = n11039 & n11047;
  assign n11103 = ~n11041 & n11049;
  assign n11101 = n11039 & n11049;
  assign n11055 = n11047 ^ n11046;
  assign n11057 = n11039 & ~n11055;
  assign n11056 = ~n11041 & ~n11055;
  assign n11058 = n11057 ^ n11056;
  assign n11096 = n11058 ^ n11055;
  assign n11090 = ~n11040 & n11047;
  assign n11072 = n11042 ^ n11037;
  assign n11073 = n11049 ^ n11038;
  assign n11074 = n11072 & n11073;
  assign n11071 = n11070 ^ n11056;
  assign n11075 = n11074 ^ n11071;
  assign n11091 = n11090 ^ n11075;
  assign n11092 = n11091 ^ n11056;
  assign n11093 = n11092 ^ n11065;
  assign n11094 = n11093 ^ n11040;
  assign n11077 = ~n11041 & n11048;
  assign n11078 = n11077 ^ n11048;
  assign n11063 = n11039 & n11048;
  assign n11076 = n11075 ^ n11063;
  assign n11079 = n11078 ^ n11076;
  assign n11089 = n11079 ^ n11074;
  assign n11095 = n11094 ^ n11089;
  assign n11097 = n11096 ^ n11095;
  assign n11102 = n11101 ^ n11097;
  assign n11104 = n11103 ^ n11102;
  assign n12936 = n11299 ^ n11104;
  assign n11098 = n11097 ^ n11069;
  assign n11100 = n11098 ^ n11049;
  assign n11105 = n11104 ^ n11100;
  assign n11106 = n11105 ^ n11057;
  assign n12935 = n11106 ^ n11095;
  assign n12937 = n12936 ^ n12935;
  assign n12938 = ~n11117 & ~n12937;
  assign n12939 = n12938 ^ n12935;
  assign n11301 = n11078 ^ n11042;
  assign n11119 = n11090 ^ n11077;
  assign n11298 = n11119 ^ n11065;
  assign n11300 = n11299 ^ n11298;
  assign n11302 = n11301 ^ n11300;
  assign n11303 = n11302 ^ n11079;
  assign n12945 = n11303 ^ n11095;
  assign n12946 = n12945 ^ n11089;
  assign n12947 = ~n11050 & ~n12946;
  assign n12948 = n12947 ^ n12945;
  assign n12940 = n11119 ^ n11063;
  assign n12941 = n12940 ^ n11302;
  assign n12942 = n12941 ^ n11093;
  assign n12943 = n11050 & n12942;
  assign n12944 = n12943 ^ n12941;
  assign n12949 = n12948 ^ n12944;
  assign n12950 = n11051 & ~n12949;
  assign n12951 = n12950 ^ n12944;
  assign n12952 = n12939 & ~n12951;
  assign n12953 = ~n11086 & n12952;
  assign n12954 = n12953 ^ n8956;
  assign n12955 = n12954 ^ x457;
  assign n10790 = n10789 ^ x442;
  assign n10805 = n10804 ^ x447;
  assign n10806 = ~n10790 & ~n10805;
  assign n10807 = n10806 ^ n10805;
  assign n10808 = n10807 ^ n10790;
  assign n10835 = n10834 ^ x446;
  assign n8903 = n8902 ^ n8878;
  assign n8904 = ~n8610 & n8903;
  assign n8905 = n8904 ^ n8878;
  assign n8906 = ~n8648 & n8905;
  assign n10073 = n8887 ^ n8878;
  assign n10837 = n10073 ^ n8881;
  assign n10836 = n8887 ^ n8871;
  assign n10838 = n10837 ^ n10836;
  assign n10839 = n10838 ^ n10836;
  assign n10840 = ~n8610 & ~n10839;
  assign n10841 = n10840 ^ n10836;
  assign n10842 = ~n8647 & n10841;
  assign n10843 = n10842 ^ n10836;
  assign n8921 = n8875 ^ n8870;
  assign n10844 = n8921 ^ n8862;
  assign n10845 = n10844 ^ n8897;
  assign n10846 = n10845 ^ n10075;
  assign n10847 = n8610 & n10846;
  assign n10848 = n10847 ^ n10075;
  assign n10849 = n8648 & n10848;
  assign n10850 = ~n10843 & ~n10849;
  assign n10851 = n8610 & n10063;
  assign n10852 = n10851 ^ n8900;
  assign n10853 = ~n8648 & n10852;
  assign n10854 = n10853 ^ n8900;
  assign n10855 = n10850 & ~n10854;
  assign n10856 = ~n8906 & n10855;
  assign n10857 = ~n10533 & n10856;
  assign n10858 = ~n10531 & n10857;
  assign n10859 = ~n10062 & n10858;
  assign n10860 = n10859 ^ n6729;
  assign n10861 = n10860 ^ x444;
  assign n9654 = n9640 & n9653;
  assign n9670 = ~n9573 & ~n9669;
  assign n9671 = n9670 ^ n9662;
  assign n9659 = n9658 ^ n9657;
  assign n9660 = n9573 & n9659;
  assign n9661 = n9660 ^ n9658;
  assign n9672 = n9671 ^ n9661;
  assign n9673 = n9574 & n9672;
  assign n9674 = n9673 ^ n9671;
  assign n9935 = n9653 & n9677;
  assign n9936 = n9935 ^ n9651;
  assign n10862 = ~n9572 & n9681;
  assign n10869 = n9664 ^ n9606;
  assign n10870 = n9572 & ~n10869;
  assign n9703 = n9702 ^ n9637;
  assign n10868 = n9703 ^ n9675;
  assign n10871 = n10870 ^ n10868;
  assign n10863 = n9686 ^ n9637;
  assign n10864 = n10863 ^ n9638;
  assign n9708 = n9701 ^ n9685;
  assign n10865 = n10864 ^ n9708;
  assign n10866 = ~n9572 & ~n10865;
  assign n10867 = n10866 ^ n9708;
  assign n10872 = n10871 ^ n10867;
  assign n10873 = ~n9574 & ~n10872;
  assign n10874 = n10873 ^ n10871;
  assign n10875 = ~n10862 & ~n10874;
  assign n10876 = ~n9936 & n10875;
  assign n10877 = ~n10593 & n10876;
  assign n10878 = ~n10590 & n10877;
  assign n10879 = ~n9674 & n10878;
  assign n10880 = ~n9654 & n10879;
  assign n10881 = n10880 ^ n6590;
  assign n10882 = n10881 ^ x445;
  assign n10919 = n10918 ^ x443;
  assign n10920 = ~n10882 & ~n10919;
  assign n10921 = ~n10861 & n10920;
  assign n10922 = n10921 ^ n10920;
  assign n10883 = n10861 & n10882;
  assign n10884 = n10883 ^ n10861;
  assign n10923 = n10922 ^ n10884;
  assign n10924 = ~n10835 & n10923;
  assign n10925 = ~n10808 & n10924;
  assign n10931 = n10883 & n10919;
  assign n10929 = n10924 ^ n10923;
  assign n10926 = n10835 & n10919;
  assign n10927 = ~n10861 & n10926;
  assign n10928 = n10927 ^ n10926;
  assign n10930 = n10929 ^ n10928;
  assign n10932 = n10931 ^ n10930;
  assign n10933 = ~n10808 & n10932;
  assign n10934 = n10805 ^ n10790;
  assign n10936 = ~n10835 & ~n10861;
  assign n10937 = ~n10919 & n10936;
  assign n10938 = n10937 ^ n10936;
  assign n10939 = n10882 & n10938;
  assign n10940 = n10939 ^ n10938;
  assign n10935 = n10930 ^ n10924;
  assign n10941 = n10940 ^ n10935;
  assign n10942 = n10805 & n10941;
  assign n10943 = n10942 ^ n10940;
  assign n10944 = n10934 & n10943;
  assign n10945 = ~n10807 & n10929;
  assign n10953 = n10931 ^ n10883;
  assign n10955 = n10953 ^ n10919;
  assign n10956 = n10955 ^ n10920;
  assign n10958 = n10835 & ~n10956;
  assign n10950 = n10835 & n10922;
  assign n10951 = n10950 ^ n10922;
  assign n10968 = n10958 ^ n10951;
  assign n10969 = n10968 ^ n10921;
  assign n10966 = n10939 ^ n10930;
  assign n10967 = n10966 ^ n10924;
  assign n10970 = n10969 ^ n10967;
  assign n10946 = n10861 ^ n10835;
  assign n10964 = n10946 ^ n10882;
  assign n10965 = n10964 ^ n10919;
  assign n10971 = n10970 ^ n10965;
  assign n10957 = n10956 ^ n10937;
  assign n10959 = n10958 ^ n10957;
  assign n10960 = n10959 ^ n10921;
  assign n10961 = n10960 ^ n10951;
  assign n10962 = n10961 ^ n10950;
  assign n10947 = n10919 ^ n10861;
  assign n10948 = n10946 & n10947;
  assign n10949 = n10948 ^ n10927;
  assign n10952 = n10951 ^ n10949;
  assign n10963 = n10962 ^ n10952;
  assign n10972 = n10971 ^ n10963;
  assign n10973 = n10972 ^ n10927;
  assign n10974 = n10790 & n10973;
  assign n10954 = n10953 ^ n10952;
  assign n10975 = n10974 ^ n10954;
  assign n10976 = n10805 & n10975;
  assign n10977 = n10976 ^ n10954;
  assign n10978 = ~n10945 & ~n10977;
  assign n10979 = n10972 ^ n10961;
  assign n10980 = ~n10790 & ~n10979;
  assign n10981 = n10980 ^ n10972;
  assign n10982 = ~n10805 & n10981;
  assign n10983 = n10929 & ~n10934;
  assign n10984 = ~n10807 & n10932;
  assign n10989 = ~n10807 & n10937;
  assign n10990 = n10989 ^ n10958;
  assign n10986 = n10953 ^ n10950;
  assign n10987 = n10986 ^ n10959;
  assign n10985 = n10972 ^ n10939;
  assign n10988 = n10987 ^ n10985;
  assign n10991 = n10990 ^ n10988;
  assign n10992 = n10991 ^ n10990;
  assign n10993 = ~n10790 & ~n10992;
  assign n10994 = n10993 ^ n10990;
  assign n10995 = n10805 & n10994;
  assign n10996 = n10995 ^ n10990;
  assign n10997 = n10805 & n10970;
  assign n10998 = n10997 ^ n10967;
  assign n10999 = ~n10934 & n10998;
  assign n11000 = ~n10996 & ~n10999;
  assign n11001 = ~n10984 & n11000;
  assign n11002 = ~n10983 & n11001;
  assign n11003 = ~n10982 & n11002;
  assign n11004 = n10978 & n11003;
  assign n11005 = ~n10944 & n11004;
  assign n11006 = ~n10933 & n11005;
  assign n11007 = ~n10925 & n11006;
  assign n11008 = n11007 ^ n8993;
  assign n12956 = n11008 ^ x455;
  assign n12957 = n12955 & ~n12956;
  assign n12958 = n12957 ^ n12955;
  assign n12959 = n12958 ^ n12956;
  assign n10100 = n8390 & n8410;
  assign n10101 = ~n7418 & n8420;
  assign n8394 = n8393 ^ n8380;
  assign n8395 = n8392 & n8394;
  assign n10114 = n8443 ^ n8405;
  assign n10115 = n10114 ^ n8421;
  assign n10112 = n8431 ^ n8399;
  assign n10113 = n10112 ^ n8408;
  assign n10116 = n10115 ^ n10113;
  assign n10117 = n7023 & n10116;
  assign n10118 = n10117 ^ n10113;
  assign n10108 = n10107 ^ n8410;
  assign n10106 = n8429 ^ n8398;
  assign n10109 = n10108 ^ n10106;
  assign n10110 = n7023 & n10109;
  assign n10111 = n10110 ^ n10106;
  assign n10119 = n10118 ^ n10111;
  assign n10120 = ~n7418 & n10119;
  assign n10121 = n10120 ^ n10111;
  assign n10122 = ~n10105 & ~n10121;
  assign n10123 = ~n8395 & n10122;
  assign n10124 = ~n10101 & n10123;
  assign n10125 = ~n10100 & n10124;
  assign n10127 = n10126 ^ n8417;
  assign n10128 = n7418 & n10127;
  assign n10129 = n10128 ^ n10126;
  assign n10130 = ~n8404 & n10129;
  assign n10131 = n10125 & ~n10130;
  assign n10132 = ~n10099 & n10131;
  assign n10133 = ~n8416 & n10132;
  assign n10134 = n10133 ^ n7323;
  assign n11382 = n10134 ^ x412;
  assign n9099 = n9057 ^ n9036;
  assign n9100 = n9095 & n9099;
  assign n9126 = n9059 & n9093;
  assign n9127 = n9126 ^ n9044;
  assign n9117 = n9052 ^ n9048;
  assign n9118 = n9117 ^ n9111;
  assign n9119 = n9118 ^ n9116;
  assign n9120 = ~n9093 & n9119;
  assign n9121 = n9120 ^ n9116;
  assign n9122 = n9113 ^ n9108;
  assign n9123 = n9122 ^ n9051;
  assign n9124 = n9123 ^ n9121;
  assign n9125 = ~n9121 & n9124;
  assign n9128 = n9127 ^ n9125;
  assign n9129 = n9094 & ~n9128;
  assign n9130 = n9129 ^ n9125;
  assign n9132 = n9062 & n9064;
  assign n9131 = n9055 & n9093;
  assign n9133 = n9132 ^ n9131;
  assign n9134 = n9130 & ~n9133;
  assign n9135 = ~n9115 & n9134;
  assign n9136 = ~n9100 & n9135;
  assign n9137 = ~n9098 & n9136;
  assign n9138 = n9137 ^ n7359;
  assign n11381 = n9138 ^ x417;
  assign n11385 = n11382 ^ n11381;
  assign n10404 = n9880 ^ n9856;
  assign n10405 = n10404 ^ n9874;
  assign n10406 = ~n9890 & n10405;
  assign n10407 = n10406 ^ n10404;
  assign n10408 = ~n9907 & n10407;
  assign n10409 = n9885 & n9891;
  assign n10410 = n10409 ^ n9860;
  assign n10411 = ~n9890 & n10410;
  assign n11339 = n9867 ^ n9860;
  assign n11340 = n11339 ^ n9886;
  assign n11341 = n11340 ^ n9886;
  assign n11342 = n9890 & ~n11341;
  assign n11343 = n11342 ^ n9886;
  assign n11344 = n9907 & n11343;
  assign n11345 = n11344 ^ n9886;
  assign n11347 = n9876 ^ n9872;
  assign n11346 = n9870 ^ n9855;
  assign n11348 = n11347 ^ n11346;
  assign n11349 = n9891 & n11348;
  assign n11350 = n11349 ^ n11346;
  assign n11351 = ~n9890 & n11350;
  assign n11352 = ~n11345 & ~n11351;
  assign n11354 = n9890 & n9914;
  assign n11353 = n10404 ^ n9862;
  assign n11355 = n11354 ^ n11353;
  assign n11356 = ~n9907 & n11355;
  assign n11357 = n11356 ^ n11353;
  assign n11358 = n11352 & ~n11357;
  assign n11359 = n10896 & n11358;
  assign n11360 = ~n10411 & n11359;
  assign n11361 = ~n10885 & n11360;
  assign n11362 = ~n10408 & n11361;
  assign n11363 = ~n9894 & n11362;
  assign n11364 = n11363 ^ n7125;
  assign n11365 = n11364 ^ x415;
  assign n9510 = n9509 ^ n9504;
  assign n9511 = ~n9429 & ~n9510;
  assign n9512 = n9511 ^ n9504;
  assign n9513 = ~n9428 & ~n9512;
  assign n9545 = n9544 ^ n9539;
  assign n9546 = ~n9514 & ~n9545;
  assign n9550 = n9516 & ~n9549;
  assign n9551 = ~n9546 & ~n9550;
  assign n9561 = ~n9429 & ~n9560;
  assign n9554 = n9519 ^ n9496;
  assign n9556 = n9555 ^ n9554;
  assign n9553 = n9552 ^ n9501;
  assign n9557 = n9556 ^ n9553;
  assign n9558 = n9429 & n9557;
  assign n9559 = n9558 ^ n9553;
  assign n9562 = n9561 ^ n9559;
  assign n9563 = n9428 & ~n9562;
  assign n9564 = n9563 ^ n9559;
  assign n9565 = n9551 & n9564;
  assign n9566 = ~n9526 & n9565;
  assign n9567 = ~n9521 & n9566;
  assign n9568 = ~n9513 & n9567;
  assign n9569 = ~n9500 & n9568;
  assign n9570 = n9569 ^ n7094;
  assign n11366 = n9570 ^ x416;
  assign n11367 = n11365 & n11366;
  assign n11368 = n11367 ^ n11365;
  assign n11369 = n11368 ^ n11366;
  assign n11370 = n11369 ^ n11365;
  assign n11371 = n10799 ^ n10794;
  assign n11372 = n10255 & n11371;
  assign n11373 = n11372 ^ n10799;
  assign n11374 = n11373 ^ n7037;
  assign n11375 = n11374 ^ x414;
  assign n9937 = n9653 & ~n9667;
  assign n9949 = ~n9572 & n9686;
  assign n9709 = n9708 ^ n9658;
  assign n9710 = n9709 ^ n9638;
  assign n9944 = n9710 ^ n9656;
  assign n9945 = n9944 ^ n9703;
  assign n9943 = n9658 ^ n9641;
  assign n9946 = n9945 ^ n9943;
  assign n9947 = n9572 & ~n9946;
  assign n9948 = n9947 ^ n9943;
  assign n9950 = n9949 ^ n9948;
  assign n9951 = n9573 & n9950;
  assign n9952 = n9951 ^ n9948;
  assign n9953 = ~n9942 & ~n9952;
  assign n9954 = ~n9941 & n9953;
  assign n9955 = ~n9654 & n9954;
  assign n9956 = ~n9655 & n9955;
  assign n9957 = ~n9937 & n9956;
  assign n9960 = n9959 ^ n9668;
  assign n9958 = n9679 ^ n9662;
  assign n9961 = n9960 ^ n9958;
  assign n9962 = ~n9573 & ~n9961;
  assign n9963 = n9962 ^ n9958;
  assign n9964 = ~n9572 & n9963;
  assign n9965 = n9957 & ~n9964;
  assign n9966 = ~n9936 & n9965;
  assign n9967 = n9966 ^ n7066;
  assign n11376 = n9967 ^ x413;
  assign n11377 = ~n11375 & ~n11376;
  assign n11434 = n11370 & n11377;
  assign n11435 = n11434 ^ n11377;
  assign n11418 = ~n11369 & n11377;
  assign n11405 = n11367 & n11377;
  assign n11419 = n11418 ^ n11405;
  assign n11436 = n11435 ^ n11419;
  assign n11378 = n11377 ^ n11376;
  assign n11401 = n11368 & ~n11378;
  assign n11400 = n11370 & ~n11378;
  assign n11402 = n11401 ^ n11400;
  assign n11398 = ~n11369 & ~n11378;
  assign n11399 = n11398 ^ n11378;
  assign n11403 = n11402 ^ n11399;
  assign n11777 = n11436 ^ n11403;
  assign n11778 = n11382 & ~n11777;
  assign n11779 = n11778 ^ n11403;
  assign n11780 = ~n11385 & ~n11779;
  assign n11383 = ~n11381 & n11382;
  assign n11384 = n11383 ^ n11381;
  assign n11386 = n11385 ^ n11384;
  assign n11415 = n11386 ^ n11381;
  assign n11416 = n11398 & n11415;
  assign n11406 = n11405 ^ n11367;
  assign n11379 = n11378 ^ n11375;
  assign n11395 = n11368 & ~n11379;
  assign n11380 = n11370 & ~n11379;
  assign n11396 = n11395 ^ n11380;
  assign n11393 = ~n11369 & ~n11379;
  assign n11394 = n11393 ^ n11379;
  assign n11397 = n11396 ^ n11394;
  assign n11404 = n11403 ^ n11397;
  assign n11407 = n11406 ^ n11404;
  assign n11414 = ~n11384 & n11407;
  assign n11417 = n11416 ^ n11414;
  assign n11446 = n11397 ^ n11393;
  assign n12232 = n11446 ^ n11434;
  assign n12233 = n11382 & ~n12232;
  assign n12234 = n12233 ^ n11434;
  assign n12235 = n11385 & n12234;
  assign n11420 = ~n11386 & n11419;
  assign n11388 = n11377 ^ n11375;
  assign n11390 = n11368 & ~n11388;
  assign n11389 = n11370 & ~n11388;
  assign n11391 = n11390 ^ n11389;
  assign n11392 = n11391 ^ n11388;
  assign n11408 = n11407 ^ n11392;
  assign n11781 = n11420 ^ n11408;
  assign n11782 = n11384 & ~n11781;
  assign n11783 = n11782 ^ n11408;
  assign n11423 = n11390 & n11415;
  assign n11422 = ~n11397 & n11415;
  assign n11424 = n11423 ^ n11422;
  assign n12961 = n11408 ^ n11402;
  assign n12962 = n12961 ^ n11389;
  assign n12960 = n11407 ^ n11380;
  assign n12963 = n12962 ^ n12960;
  assign n12964 = ~n11381 & ~n12963;
  assign n12965 = n12964 ^ n12960;
  assign n12966 = n11382 & n12965;
  assign n11784 = n11393 ^ n11389;
  assign n12969 = n11436 ^ n11402;
  assign n12237 = n11418 ^ n11400;
  assign n12968 = n12237 ^ n11403;
  assign n12970 = n12969 ^ n12968;
  assign n12971 = n12969 ^ n11382;
  assign n12972 = n11385 & n12971;
  assign n12973 = n12972 ^ n11382;
  assign n12974 = ~n12970 & ~n12973;
  assign n12975 = n12974 ^ n12968;
  assign n12976 = ~n11784 & n12975;
  assign n12967 = n11381 & n11396;
  assign n12977 = n12976 ^ n12967;
  assign n12978 = n11385 & ~n12977;
  assign n12979 = n12978 ^ n12976;
  assign n12980 = ~n12966 & n12979;
  assign n12981 = ~n11424 & n12980;
  assign n12982 = n11783 & n12981;
  assign n12983 = ~n12235 & n12982;
  assign n12984 = ~n11417 & n12983;
  assign n12985 = ~n11780 & n12984;
  assign n12986 = n12985 ^ n9026;
  assign n12987 = n12986 ^ x456;
  assign n8910 = n8900 ^ n8872;
  assign n8911 = n8647 & n8910;
  assign n8912 = n8911 ^ n8872;
  assign n8907 = n8902 ^ n8868;
  assign n8908 = n8647 & n8907;
  assign n8909 = n8908 ^ n8902;
  assign n8913 = n8912 ^ n8909;
  assign n8914 = ~n8610 & n8913;
  assign n8915 = n8914 ^ n8909;
  assign n8922 = n8921 ^ n8882;
  assign n8923 = n8922 ^ n8889;
  assign n8924 = n8610 & n8923;
  assign n8925 = n8924 ^ n8922;
  assign n8926 = n8925 ^ n8898;
  assign n8927 = n8925 & n8926;
  assign n8917 = n8916 ^ n8895;
  assign n8918 = n8917 ^ n8890;
  assign n8919 = ~n8610 & n8918;
  assign n8920 = n8919 ^ n8917;
  assign n8928 = n8927 ^ n8920;
  assign n8929 = ~n8648 & ~n8928;
  assign n8930 = n8929 ^ n8927;
  assign n8931 = ~n8915 & n8930;
  assign n8932 = ~n8906 & n8931;
  assign n8933 = ~n8893 & n8932;
  assign n8934 = n8933 ^ n8104;
  assign n10214 = n8934 ^ x424;
  assign n10251 = n10250 ^ x429;
  assign n10252 = ~n10214 & ~n10251;
  assign n10253 = n10252 ^ n10214;
  assign n10254 = n10253 ^ n10251;
  assign n10373 = n10372 ^ x428;
  assign n10378 = n9093 & n9111;
  assign n10379 = n10378 ^ n9036;
  assign n10380 = n9094 & n10379;
  assign n10381 = n10380 ^ n9036;
  assign n10382 = n9064 & ~n9122;
  assign n10388 = n10387 ^ n9047;
  assign n10386 = n9116 ^ n9043;
  assign n10389 = n10388 ^ n10386;
  assign n10390 = n9064 & n10389;
  assign n10391 = n10390 ^ n10386;
  assign n10383 = n9062 & n9096;
  assign n10384 = n10383 ^ n9049;
  assign n10385 = n10384 ^ n9053;
  assign n10392 = n10391 ^ n10385;
  assign n10393 = ~n9093 & n10392;
  assign n10394 = n10393 ^ n10385;
  assign n10395 = ~n10382 & ~n10394;
  assign n10396 = ~n10381 & n10395;
  assign n10397 = ~n9107 & n10396;
  assign n10398 = ~n10377 & n10397;
  assign n10399 = ~n9100 & n10398;
  assign n10400 = ~n9098 & n10399;
  assign n10401 = n10400 ^ n8506;
  assign n10402 = n10401 ^ x426;
  assign n10403 = n10373 & n10402;
  assign n10423 = n10422 ^ n9886;
  assign n10421 = n9862 ^ n9858;
  assign n10424 = n10423 ^ n10421;
  assign n10425 = n10424 ^ n10421;
  assign n10426 = n9890 & n10425;
  assign n10427 = n10426 ^ n10421;
  assign n10428 = n9891 & n10427;
  assign n10429 = n10428 ^ n10421;
  assign n10430 = n9888 ^ n9873;
  assign n10431 = n9890 & n10430;
  assign n10432 = n10431 ^ n9888;
  assign n10433 = n10432 ^ n9877;
  assign n10434 = n10432 ^ n9907;
  assign n10435 = ~n10432 & ~n10434;
  assign n10436 = n10435 ^ n10432;
  assign n10437 = n10433 & ~n10436;
  assign n10438 = n10437 ^ n10435;
  assign n10439 = n10438 ^ n10432;
  assign n10440 = n10439 ^ n9907;
  assign n10441 = ~n10429 & ~n10440;
  assign n10442 = n10441 ^ n10429;
  assign n10443 = n10420 & ~n10442;
  assign n10444 = ~n10411 & n10443;
  assign n10445 = ~n9902 & n10444;
  assign n10446 = ~n10408 & n10445;
  assign n10447 = n10446 ^ n8479;
  assign n10448 = n10447 ^ x427;
  assign n9695 = n9652 ^ n9573;
  assign n9696 = n9694 & ~n9695;
  assign n9711 = n9710 ^ n9668;
  assign n9698 = ~n9652 & ~n9697;
  assign n9704 = n9695 & ~n9703;
  assign n9705 = n9647 & n9704;
  assign n9706 = ~n9698 & ~n9705;
  assign n9707 = ~n9677 & ~n9706;
  assign n9712 = n9711 ^ n9707;
  assign n9713 = n9712 ^ n9707;
  assign n9714 = ~n9572 & n9713;
  assign n9715 = n9714 ^ n9707;
  assign n9716 = n9573 & ~n9715;
  assign n9717 = n9716 ^ n9707;
  assign n9718 = ~n9696 & n9717;
  assign n9719 = n9573 & ~n9683;
  assign n9720 = n9719 ^ n9678;
  assign n9721 = n9572 & n9720;
  assign n9722 = n9718 & ~n9721;
  assign n9723 = ~n9693 & n9722;
  assign n9724 = ~n9692 & n9723;
  assign n9725 = ~n9674 & n9724;
  assign n9726 = ~n9654 & n9725;
  assign n9727 = ~n9651 & n9726;
  assign n9728 = n9727 ^ n8073;
  assign n10449 = n9728 ^ x425;
  assign n10450 = ~n10448 & ~n10449;
  assign n10451 = n10450 ^ n10449;
  assign n10452 = n10403 & ~n10451;
  assign n10453 = ~n10254 & n10452;
  assign n10454 = n10254 ^ n10252;
  assign n10455 = n10403 ^ n10373;
  assign n10456 = n10455 ^ n10402;
  assign n10468 = n10456 ^ n10373;
  assign n10475 = n10451 ^ n10448;
  assign n10501 = n10468 & ~n10475;
  assign n11959 = ~n10251 & n10501;
  assign n10485 = n10403 & ~n10475;
  assign n10484 = ~n10456 & ~n10475;
  assign n10486 = n10485 ^ n10484;
  assign n10473 = n10450 & ~n10456;
  assign n11956 = n10486 ^ n10473;
  assign n11957 = ~n10251 & n11956;
  assign n11958 = n11957 ^ n10473;
  assign n11960 = n11959 ^ n11958;
  assign n11961 = ~n10454 & n11960;
  assign n11962 = n11961 ^ n11958;
  assign n11963 = n10252 & n10485;
  assign n10496 = ~n10451 & n10468;
  assign n10478 = n10450 & n10455;
  assign n10470 = ~n10451 & n10455;
  assign n10479 = n10478 ^ n10470;
  assign n11964 = n10496 ^ n10479;
  assign n11965 = ~n10253 & n11964;
  assign n10476 = n10455 & ~n10475;
  assign n10477 = n10476 ^ n10455;
  assign n10480 = n10479 ^ n10477;
  assign n11966 = n10214 & n10480;
  assign n10494 = n10254 ^ n10214;
  assign n10469 = n10450 & n10468;
  assign n10471 = n10470 ^ n10469;
  assign n11967 = n10471 ^ n10452;
  assign n10462 = n10403 & n10450;
  assign n11968 = n11967 ^ n10462;
  assign n11969 = ~n10494 & n11968;
  assign n11970 = ~n11966 & ~n11969;
  assign n11212 = n10484 ^ n10476;
  assign n11213 = n11212 ^ n10501;
  assign n10457 = n10450 ^ n10448;
  assign n10459 = n10403 & ~n10457;
  assign n11981 = n11213 ^ n10459;
  assign n10461 = ~n10451 & ~n10456;
  assign n10463 = n10462 ^ n10461;
  assign n11973 = n10473 ^ n10463;
  assign n11971 = n10496 ^ n10462;
  assign n10458 = ~n10456 & ~n10457;
  assign n11972 = n11971 ^ n10458;
  assign n11974 = n11973 ^ n11972;
  assign n11975 = n11973 ^ n10251;
  assign n11976 = n10454 & ~n11975;
  assign n11977 = n11976 ^ n10251;
  assign n11978 = n11974 & n11977;
  assign n11979 = n11978 ^ n11972;
  assign n11980 = ~n10478 & ~n11979;
  assign n11982 = n11981 ^ n11980;
  assign n11983 = n11982 ^ n11980;
  assign n11984 = n10251 & n11983;
  assign n11985 = n11984 ^ n11980;
  assign n11986 = n10454 & ~n11985;
  assign n11987 = n11986 ^ n11980;
  assign n11988 = n11970 & n11987;
  assign n11989 = ~n11965 & n11988;
  assign n11990 = ~n11963 & n11989;
  assign n11991 = ~n10251 & n10458;
  assign n10482 = ~n10457 & n10468;
  assign n10483 = n10482 ^ n10476;
  assign n11992 = n11991 ^ n10483;
  assign n11993 = n10454 & n11992;
  assign n11994 = n11993 ^ n10483;
  assign n11995 = n11990 & ~n11994;
  assign n11996 = ~n11962 & n11995;
  assign n11997 = ~n10453 & n11996;
  assign n11998 = n11997 ^ n8609;
  assign n12988 = n11998 ^ x458;
  assign n12989 = ~n12987 & ~n12988;
  assign n13009 = n12989 ^ n12987;
  assign n13010 = n12959 & ~n13009;
  assign n12990 = n12989 ^ n12988;
  assign n12991 = n12990 ^ n12987;
  assign n12995 = n12959 ^ n12955;
  assign n12997 = ~n12991 & ~n12995;
  assign n12996 = n12989 & ~n12995;
  assign n12998 = n12997 ^ n12996;
  assign n13271 = n13010 ^ n12998;
  assign n13272 = n12933 & n13271;
  assign n13273 = n13272 ^ n13010;
  assign n13274 = n13013 & n13273;
  assign n12993 = n12958 & n12989;
  assign n12992 = n12959 & ~n12991;
  assign n12994 = n12993 ^ n12992;
  assign n12999 = n12998 ^ n12994;
  assign n13000 = ~n12934 & n12999;
  assign n13001 = n13000 ^ n12998;
  assign n13002 = ~n12933 & n13001;
  assign n13004 = n12933 & ~n12934;
  assign n13036 = n12957 & ~n13009;
  assign n13037 = n13036 ^ n12957;
  assign n13008 = n12957 & ~n12990;
  assign n13003 = n12957 & ~n12991;
  assign n13035 = n13008 ^ n13003;
  assign n13038 = n13037 ^ n13035;
  assign n13268 = n13038 ^ n13003;
  assign n13465 = n13004 & n13268;
  assign n13032 = ~n12990 & ~n12995;
  assign n13466 = n13035 ^ n13032;
  assign n13467 = ~n13013 & n13466;
  assign n13015 = n12959 & ~n12990;
  assign n13020 = n13015 ^ n12994;
  assign n13019 = n12958 & ~n12991;
  assign n13021 = n13020 ^ n13019;
  assign n13014 = n12958 & ~n13009;
  assign n13016 = n13015 ^ n13014;
  assign n13017 = n13016 ^ n12992;
  assign n13018 = n13017 ^ n12958;
  assign n13022 = n13021 ^ n13018;
  assign n13065 = n13004 & n13022;
  assign n13474 = n13065 ^ n12933;
  assign n13026 = n13015 ^ n12956;
  assign n13023 = n13022 ^ n13010;
  assign n13024 = n13023 ^ n13016;
  assign n13025 = n13024 ^ n13021;
  assign n13027 = n13026 ^ n13025;
  assign n13472 = n13004 & n13027;
  assign n13068 = n12992 & n13004;
  assign n13473 = n13472 ^ n13068;
  assign n13475 = n13474 ^ n13473;
  assign n13470 = n13004 & ~n13014;
  assign n13005 = n13004 ^ n12933;
  assign n13468 = n13020 ^ n13010;
  assign n13469 = n13005 & ~n13468;
  assign n13471 = n13470 ^ n13469;
  assign n13476 = n13475 ^ n13471;
  assign n13477 = ~n13467 & ~n13476;
  assign n13478 = ~n13465 & n13477;
  assign n13480 = n13015 ^ n12993;
  assign n13481 = n13480 ^ n13038;
  assign n13482 = n13481 ^ n13036;
  assign n13033 = n13032 ^ n12995;
  assign n13034 = n13033 ^ n12998;
  assign n13479 = n13034 ^ n13023;
  assign n13483 = n13482 ^ n13479;
  assign n13484 = n12934 & ~n13483;
  assign n13485 = n13484 ^ n13479;
  assign n13486 = ~n12933 & ~n13485;
  assign n13487 = n13478 & ~n13486;
  assign n13283 = n13036 ^ n13019;
  assign n13488 = n12933 & n13283;
  assign n13489 = n13488 ^ n13019;
  assign n13490 = n12934 & n13489;
  assign n13491 = n13487 & ~n13490;
  assign n13492 = ~n13002 & n13491;
  assign n13493 = ~n13274 & n13492;
  assign n13494 = n13493 ^ n9138;
  assign n13645 = n13494 ^ x513;
  assign n11255 = ~n10807 & n10966;
  assign n11253 = n10959 ^ n10950;
  assign n11254 = ~n10808 & ~n11253;
  assign n11256 = n11255 ^ n11254;
  assign n11257 = n10940 ^ n10929;
  assign n11258 = n11257 ^ n10968;
  assign n11259 = ~n10805 & n11258;
  assign n11260 = n11259 ^ n10968;
  assign n11261 = ~n10790 & n11260;
  assign n11262 = ~n10944 & ~n11261;
  assign n11269 = n10986 ^ n10948;
  assign n11270 = n10805 & n11269;
  assign n11271 = n11270 ^ n10986;
  assign n11264 = n10973 ^ n10932;
  assign n11265 = n11264 ^ n10958;
  assign n11263 = n10954 ^ n10938;
  assign n11266 = n11265 ^ n11263;
  assign n11267 = ~n10805 & n11266;
  assign n11268 = n11267 ^ n11263;
  assign n11272 = n11271 ^ n11268;
  assign n11273 = n10790 & n11272;
  assign n11274 = n11273 ^ n11268;
  assign n11275 = n10959 ^ n10937;
  assign n11276 = n11275 ^ n10929;
  assign n11277 = n10790 & ~n11276;
  assign n11278 = n11277 ^ n10929;
  assign n11279 = n11278 ^ n11275;
  assign n11280 = n10805 & ~n11279;
  assign n11281 = n11280 ^ n11275;
  assign n11282 = ~n11274 & n11281;
  assign n11283 = n11262 & n11282;
  assign n11284 = ~n11256 & n11283;
  assign n11285 = ~n10982 & n11284;
  assign n11286 = ~n10933 & n11285;
  assign n11287 = n11286 ^ n7022;
  assign n12231 = n11287 ^ x477;
  assign n11387 = n11386 ^ n11380;
  assign n11409 = n11408 ^ n11384;
  assign n11410 = ~n11380 & ~n11409;
  assign n11411 = n11410 ^ n11384;
  assign n11412 = n11387 & ~n11411;
  assign n11413 = n11412 ^ n11386;
  assign n11428 = n11407 ^ n11395;
  assign n12236 = n11383 & n11428;
  assign n12250 = n11398 ^ n11391;
  assign n12239 = n11376 ^ n11365;
  assign n12240 = n11375 ^ n11365;
  assign n12241 = n12240 ^ n11366;
  assign n12242 = n12241 ^ n11376;
  assign n12243 = ~n11366 & ~n12242;
  assign n12244 = n12243 ^ n12241;
  assign n12245 = n12239 & ~n12244;
  assign n12246 = n12245 ^ n12241;
  assign n11437 = n11436 ^ n11434;
  assign n12238 = n12237 ^ n11437;
  assign n12247 = n12246 ^ n12238;
  assign n12248 = ~n11382 & ~n12247;
  assign n12249 = n12248 ^ n12238;
  assign n12251 = n12250 ^ n12249;
  assign n12252 = n11385 & n12251;
  assign n12253 = n12252 ^ n12250;
  assign n12254 = ~n11423 & ~n12253;
  assign n12255 = ~n12236 & n12254;
  assign n12256 = n11405 ^ n11401;
  assign n12257 = n12256 ^ n11404;
  assign n12258 = ~n11382 & n12257;
  assign n12259 = n12258 ^ n11404;
  assign n12260 = ~n11385 & n12259;
  assign n12261 = n12255 & ~n12260;
  assign n12262 = ~n11414 & n12261;
  assign n12263 = ~n12235 & n12262;
  assign n12264 = ~n11413 & n12263;
  assign n12265 = ~n11780 & n12264;
  assign n12266 = n12265 ^ n7417;
  assign n12267 = n12266 ^ x472;
  assign n12268 = n12231 & ~n12267;
  assign n12269 = n12268 ^ n12231;
  assign n12075 = n10680 & n10716;
  assign n12071 = n10646 ^ n10644;
  assign n12070 = n10700 ^ n10627;
  assign n12072 = n12071 ^ n12070;
  assign n12073 = ~n10680 & n12072;
  assign n12074 = n12073 ^ n12070;
  assign n12076 = n12075 ^ n12074;
  assign n12077 = ~n10648 & n12076;
  assign n12078 = n12077 ^ n12074;
  assign n12270 = n10629 ^ n10621;
  assign n12271 = ~n10680 & n12270;
  assign n11753 = n10719 ^ n10638;
  assign n12272 = n11753 ^ n10700;
  assign n12273 = n12272 ^ n10623;
  assign n12274 = ~n10682 & ~n12273;
  assign n12275 = ~n12271 & ~n12274;
  assign n12277 = n10644 ^ n10642;
  assign n12276 = n10635 ^ n10630;
  assign n12278 = n12277 ^ n12276;
  assign n12279 = ~n10692 & n12278;
  assign n12089 = n10696 ^ n10642;
  assign n12280 = n12089 ^ n10639;
  assign n12281 = n12089 ^ n10680;
  assign n12282 = n10693 & ~n12281;
  assign n12283 = n12282 ^ n10680;
  assign n12284 = n12280 & n12283;
  assign n12285 = n12284 ^ n10639;
  assign n12286 = ~n10716 & ~n12285;
  assign n12287 = n12286 ^ n10619;
  assign n12288 = n12286 ^ n10693;
  assign n12289 = n12286 & ~n12288;
  assign n12290 = n12289 ^ n12286;
  assign n12291 = ~n12287 & n12290;
  assign n12292 = n12291 ^ n12289;
  assign n12293 = n12292 ^ n12286;
  assign n12294 = n12293 ^ n10693;
  assign n12295 = ~n12279 & ~n12294;
  assign n12296 = n12295 ^ n12279;
  assign n12297 = n12275 & ~n12296;
  assign n12298 = ~n12078 & n12297;
  assign n12299 = n12298 ^ n8050;
  assign n12300 = n12299 ^ x475;
  assign n11582 = n11560 ^ n11553;
  assign n11583 = ~n11547 & n11582;
  assign n11584 = n11580 ^ n11557;
  assign n11585 = n11542 & ~n11584;
  assign n11586 = n11585 ^ n11580;
  assign n11587 = n11541 & ~n11586;
  assign n12301 = n11546 & n11560;
  assign n12311 = n11537 ^ n11501;
  assign n12312 = n12311 ^ n11596;
  assign n12313 = n11541 & n12312;
  assign n12302 = n11598 ^ n11578;
  assign n12303 = n12302 ^ n11592;
  assign n12304 = n12302 ^ n11541;
  assign n12305 = ~n11542 & n12304;
  assign n12306 = n12305 ^ n11541;
  assign n12307 = ~n12303 & n12306;
  assign n12308 = n12307 ^ n11592;
  assign n12309 = ~n11540 & ~n12308;
  assign n12310 = n11580 & n12309;
  assign n12314 = n12313 ^ n12310;
  assign n12315 = ~n11542 & ~n12314;
  assign n12316 = n12315 ^ n12310;
  assign n12317 = ~n12301 & n12316;
  assign n12318 = n11539 ^ n11499;
  assign n12319 = n12318 ^ n11554;
  assign n12320 = n12319 ^ n11554;
  assign n12321 = ~n11541 & ~n12320;
  assign n12322 = n12321 ^ n11554;
  assign n12323 = ~n11542 & n12322;
  assign n12324 = n12323 ^ n11554;
  assign n12325 = n12317 & ~n12324;
  assign n12326 = ~n11587 & n12325;
  assign n12327 = ~n11583 & n12326;
  assign n12328 = ~n12113 & n12327;
  assign n12329 = n12328 ^ n7778;
  assign n12330 = n12329 ^ x473;
  assign n12331 = n12300 & n12330;
  assign n12332 = n12331 ^ n12300;
  assign n9571 = n9570 ^ x418;
  assign n9729 = n9728 ^ x423;
  assign n8400 = n8390 & n8399;
  assign n8403 = n8389 & n8402;
  assign n8418 = ~n8391 & n8417;
  assign n8432 = n8431 ^ n8429;
  assign n8433 = n8432 ^ n8411;
  assign n8434 = n8433 ^ n7418;
  assign n8424 = n8419 ^ n8384;
  assign n8423 = n8422 ^ n8412;
  assign n8425 = n8424 ^ n8423;
  assign n8426 = n8390 & n8425;
  assign n8427 = n8426 ^ n8423;
  assign n8435 = n8434 ^ n8427;
  assign n8436 = n8404 & n8435;
  assign n8437 = n8436 ^ n8433;
  assign n8438 = ~n8418 & ~n8437;
  assign n8439 = ~n8416 & n8438;
  assign n8440 = ~n8403 & n8439;
  assign n8441 = ~n8400 & n8440;
  assign n8444 = ~n7023 & n8443;
  assign n8442 = n8392 & n8396;
  assign n8445 = n8444 ^ n8442;
  assign n8446 = n8441 & ~n8445;
  assign n8447 = ~n8395 & n8446;
  assign n8448 = ~n8388 & n8447;
  assign n8449 = n8448 ^ n8165;
  assign n8450 = n8449 ^ x420;
  assign n9139 = n9138 ^ x419;
  assign n9140 = n9139 ^ n8450;
  assign n8935 = n8934 ^ x422;
  assign n9141 = n9140 ^ n8935;
  assign n9142 = n8450 & ~n9141;
  assign n9143 = n9142 ^ n8935;
  assign n11196 = n9143 ^ n9140;
  assign n11197 = n11196 ^ n8935;
  assign n9372 = n9314 ^ n9251;
  assign n9373 = n9372 ^ n9351;
  assign n9374 = n9182 & n9373;
  assign n9371 = n9362 ^ n9322;
  assign n9375 = n9374 ^ n9371;
  assign n9376 = n9193 & ~n9375;
  assign n9380 = n9379 ^ n9335;
  assign n9377 = n9182 & n9347;
  assign n9378 = n9377 ^ n9346;
  assign n9381 = n9380 ^ n9378;
  assign n9382 = n9381 ^ n9378;
  assign n9383 = ~n9182 & n9382;
  assign n9384 = n9383 ^ n9378;
  assign n9385 = ~n9194 & n9384;
  assign n9386 = n9385 ^ n9378;
  assign n9387 = ~n9376 & ~n9386;
  assign n9389 = n9342 & n9355;
  assign n9388 = n9182 & n9350;
  assign n9390 = n9389 ^ n9388;
  assign n9391 = n9387 & ~n9390;
  assign n9392 = ~n9370 & n9391;
  assign n9393 = ~n9363 & n9392;
  assign n9394 = ~n9360 & n9393;
  assign n9395 = ~n9354 & n9394;
  assign n9396 = ~n9329 & n9395;
  assign n9397 = n9396 ^ n8138;
  assign n9398 = n9397 ^ x421;
  assign n9399 = n9143 & n9398;
  assign n11198 = n11197 ^ n9399;
  assign n9737 = n9398 ^ n8450;
  assign n9738 = ~n8450 & n8935;
  assign n9739 = n9738 ^ n8935;
  assign n9740 = ~n9737 & n9739;
  assign n11199 = n11198 ^ n9740;
  assign n9735 = n9398 ^ n9139;
  assign n9734 = n9398 ^ n8935;
  assign n9736 = n9735 ^ n9734;
  assign n9748 = ~n8935 & n9398;
  assign n9756 = n9748 ^ n9398;
  assign n9757 = n9756 ^ n9738;
  assign n9758 = n9757 ^ n8450;
  assign n9759 = ~n9736 & ~n9758;
  assign n9755 = n9735 ^ n8450;
  assign n9760 = n9759 ^ n9755;
  assign n11200 = n11199 ^ n9760;
  assign n11201 = n9729 & ~n11200;
  assign n11202 = n11201 ^ n11199;
  assign n9749 = n9748 ^ n8935;
  assign n9750 = ~n8450 & ~n9749;
  assign n9751 = n9750 ^ n8450;
  assign n9753 = n9751 ^ n9398;
  assign n9754 = ~n9139 & ~n9753;
  assign n9761 = n9760 ^ n9754;
  assign n9741 = n9740 ^ n9398;
  assign n9742 = ~n9736 & n9741;
  assign n9743 = n9742 ^ n9738;
  assign n11192 = n9761 ^ n9743;
  assign n9765 = n9748 ^ n8450;
  assign n11190 = ~n9139 & ~n9765;
  assign n11191 = n11190 ^ n9734;
  assign n11193 = n11192 ^ n11191;
  assign n11194 = ~n9729 & n11193;
  assign n11195 = n11194 ^ n11192;
  assign n11203 = n11202 ^ n11195;
  assign n11204 = ~n9571 & n11203;
  assign n11205 = n11204 ^ n11195;
  assign n11206 = n11205 ^ n8218;
  assign n12334 = n11206 ^ x476;
  assign n9934 = n9933 ^ x406;
  assign n9968 = n9967 ^ x411;
  assign n10070 = n8866 & n10059;
  assign n10071 = n8885 & n10060;
  assign n10072 = n8856 ^ n8814;
  assign n10080 = n8883 ^ n8875;
  assign n10081 = n8610 & n10080;
  assign n10082 = n10081 ^ n8883;
  assign n10074 = n10073 ^ n8867;
  assign n10076 = n10075 ^ n10074;
  assign n10077 = n10076 ^ n10072;
  assign n10078 = n10077 ^ n10072;
  assign n10079 = ~n8610 & n10078;
  assign n10083 = n10082 ^ n10079;
  assign n10084 = n10083 ^ n10079;
  assign n10085 = n10072 & ~n10084;
  assign n10086 = n10085 ^ n10079;
  assign n10087 = n8648 & ~n10086;
  assign n10088 = n10087 ^ n10079;
  assign n10089 = ~n10071 & ~n10088;
  assign n10090 = ~n10070 & n10089;
  assign n10091 = n10069 & n10090;
  assign n10092 = ~n10067 & n10091;
  assign n10093 = ~n10062 & n10092;
  assign n10094 = n10093 ^ n8282;
  assign n10095 = n10094 ^ x408;
  assign n10135 = n10134 ^ x410;
  assign n10136 = ~n10095 & n10135;
  assign n10137 = n10136 ^ n10095;
  assign n10138 = n10137 ^ n10135;
  assign n10150 = n10138 ^ n10095;
  assign n9987 = n9986 ^ n9490;
  assign n9988 = n9987 ^ n9522;
  assign n9989 = ~n9429 & n9988;
  assign n9990 = n9989 ^ n9522;
  assign n9981 = n9969 & n9980;
  assign n9979 = n9515 & n9517;
  assign n9982 = n9981 ^ n9979;
  assign n9983 = n9982 ^ n9548;
  assign n9978 = n9977 ^ n9494;
  assign n9984 = n9983 ^ n9978;
  assign n9991 = n9990 ^ n9984;
  assign n9992 = n9991 ^ n9984;
  assign n9994 = ~n9496 & n9993;
  assign n9995 = n9554 ^ n9494;
  assign n9997 = n9996 ^ n9995;
  assign n9998 = ~n9994 & n9997;
  assign n9999 = ~n9543 & ~n9998;
  assign n10000 = n9999 ^ n9984;
  assign n10001 = n10000 ^ n9984;
  assign n10002 = ~n9992 & n10001;
  assign n10003 = n10002 ^ n9984;
  assign n10004 = ~n9514 & n10003;
  assign n10005 = n10004 ^ n9984;
  assign n10006 = n9975 & n10005;
  assign n10007 = ~n9513 & n10006;
  assign n10008 = ~n9971 & n10007;
  assign n10009 = n10008 ^ n8246;
  assign n10010 = n10009 ^ x409;
  assign n10056 = n10055 ^ x407;
  assign n10057 = ~n10010 & ~n10056;
  assign n10058 = n10057 ^ n10056;
  assign n10153 = n10058 ^ n10010;
  assign n10154 = n10150 & ~n10153;
  assign n10155 = n10154 ^ n10150;
  assign n10151 = ~n10058 & n10150;
  assign n10143 = n10057 ^ n10010;
  assign n10147 = ~n10137 & ~n10143;
  assign n10148 = n10147 ^ n10143;
  assign n10145 = n10136 & ~n10143;
  assign n10144 = n10138 & ~n10143;
  assign n10146 = n10145 ^ n10144;
  assign n10149 = n10148 ^ n10146;
  assign n10152 = n10151 ^ n10149;
  assign n10156 = n10155 ^ n10152;
  assign n10157 = n10156 ^ n10057;
  assign n10141 = n10057 & n10136;
  assign n10140 = n10057 & n10138;
  assign n10142 = n10141 ^ n10140;
  assign n10158 = n10157 ^ n10142;
  assign n10159 = n10158 ^ n10156;
  assign n10139 = ~n10058 & n10138;
  assign n10160 = n10159 ^ n10139;
  assign n10161 = ~n9968 & n10160;
  assign n10162 = n10161 ^ n10139;
  assign n10163 = n9934 & n10162;
  assign n10176 = n9934 & n9968;
  assign n10180 = n10176 ^ n9968;
  assign n10181 = n10180 ^ n9934;
  assign n10183 = ~n10149 & ~n10181;
  assign n10166 = n10136 & ~n10153;
  assign n10165 = n10138 & ~n10153;
  assign n10167 = n10166 ^ n10165;
  assign n10168 = n10167 ^ n10153;
  assign n10169 = n10168 ^ n10154;
  assign n11832 = ~n10169 & ~n10181;
  assign n11829 = n9934 & n10146;
  assign n11830 = n11829 ^ n10145;
  assign n11831 = n9968 & n11830;
  assign n11833 = n11832 ^ n11831;
  assign n12000 = n10167 ^ n10151;
  assign n12001 = n9934 & n12000;
  assign n12002 = n12001 ^ n10151;
  assign n12003 = ~n9968 & n12002;
  assign n10164 = n9968 ^ n9934;
  assign n10187 = ~n10058 & ~n10137;
  assign n11845 = ~n10164 & n10187;
  assign n11844 = n10141 & n10176;
  assign n11846 = n11845 ^ n11844;
  assign n12004 = n10187 ^ n10156;
  assign n12005 = n10180 & ~n12004;
  assign n10177 = n10176 ^ n9934;
  assign n10178 = n10169 ^ n10145;
  assign n10179 = n10177 & ~n10178;
  assign n12335 = n12000 ^ n10145;
  assign n12336 = n10176 & n12335;
  assign n10192 = n10147 ^ n10139;
  assign n10193 = n10192 ^ n10151;
  assign n12340 = n10193 ^ n10144;
  assign n12341 = n12340 ^ n10166;
  assign n12017 = n10154 ^ n10144;
  assign n10188 = n10187 ^ n10147;
  assign n11834 = n10188 ^ n10058;
  assign n11835 = n11834 ^ n10193;
  assign n12018 = n12017 ^ n11835;
  assign n12019 = n12018 ^ n10140;
  assign n12337 = n12019 ^ n10142;
  assign n12338 = ~n9934 & ~n12337;
  assign n12339 = n12338 ^ n10142;
  assign n12342 = n12341 ^ n12339;
  assign n12343 = n12342 ^ n12339;
  assign n12344 = ~n9934 & n12343;
  assign n12345 = n12344 ^ n12339;
  assign n12346 = n9968 & n12345;
  assign n12347 = n12346 ^ n12339;
  assign n12348 = ~n12336 & ~n12347;
  assign n12349 = ~n10179 & n12348;
  assign n12350 = ~n12005 & n12349;
  assign n12351 = ~n11846 & n12350;
  assign n12352 = ~n12003 & n12351;
  assign n12353 = ~n11833 & n12352;
  assign n12354 = ~n10183 & n12353;
  assign n12355 = ~n10163 & n12354;
  assign n12356 = n12355 ^ n8374;
  assign n12357 = n12356 ^ x474;
  assign n12358 = n12334 & n12357;
  assign n12399 = n12332 & n12358;
  assign n12333 = n12332 ^ n12330;
  assign n12359 = n12358 ^ n12334;
  assign n12363 = n12359 ^ n12357;
  assign n12385 = ~n12333 & ~n12363;
  assign n12400 = n12399 ^ n12385;
  assign n12386 = n12385 ^ n12363;
  assign n12373 = n12357 ^ n12300;
  assign n12374 = n12330 & n12373;
  assign n12369 = n12331 & n12358;
  assign n12375 = n12374 ^ n12369;
  assign n12368 = n12331 & ~n12363;
  assign n12370 = n12369 ^ n12368;
  assign n12367 = n12331 & n12359;
  assign n12371 = n12370 ^ n12367;
  assign n12361 = n12333 ^ n12300;
  assign n12364 = n12363 ^ n12334;
  assign n12365 = n12361 & n12364;
  assign n12372 = n12371 ^ n12365;
  assign n12376 = n12375 ^ n12372;
  assign n12377 = n12376 ^ n12361;
  assign n12362 = n12359 & n12361;
  assign n12366 = n12365 ^ n12362;
  assign n12378 = n12377 ^ n12366;
  assign n12384 = n12378 ^ n12368;
  assign n12387 = n12386 ^ n12384;
  assign n12401 = n12400 ^ n12387;
  assign n12402 = n12401 ^ n12332;
  assign n12389 = n12334 ^ n12330;
  assign n12390 = n12389 ^ n12300;
  assign n12391 = n12390 ^ n12330;
  assign n12392 = n12391 ^ n12357;
  assign n12393 = n12374 ^ n12300;
  assign n12394 = n12392 & n12393;
  assign n12395 = n12394 ^ n12389;
  assign n12383 = ~n12333 & n12358;
  assign n12388 = n12387 ^ n12383;
  assign n12396 = n12395 ^ n12388;
  assign n12380 = n12371 ^ n12331;
  assign n12381 = n12380 ^ n12370;
  assign n12360 = ~n12333 & n12359;
  assign n12379 = n12378 ^ n12360;
  assign n12382 = n12381 ^ n12379;
  assign n12397 = n12396 ^ n12382;
  assign n12398 = n12397 ^ n12385;
  assign n12403 = n12402 ^ n12398;
  assign n12404 = n12269 & n12403;
  assign n12405 = n12380 ^ n12376;
  assign n12406 = n12405 ^ n12378;
  assign n12407 = ~n12267 & n12406;
  assign n12408 = n12407 ^ n12378;
  assign n12409 = ~n12231 & n12408;
  assign n12410 = n12269 ^ n12267;
  assign n12411 = n12367 ^ n12362;
  assign n12412 = n12411 ^ n12380;
  assign n12413 = n12410 & n12412;
  assign n12414 = n12401 ^ n12360;
  assign n12415 = n12268 & ~n12414;
  assign n12420 = ~n12267 & n12370;
  assign n12416 = n12384 ^ n12376;
  assign n12417 = n12416 ^ n12372;
  assign n12418 = ~n12267 & n12417;
  assign n12419 = n12418 ^ n12416;
  assign n12421 = n12420 ^ n12419;
  assign n12422 = ~n12231 & n12421;
  assign n12423 = n12422 ^ n12419;
  assign n12424 = n12267 ^ n12231;
  assign n12437 = n12403 ^ n12388;
  assign n12427 = n12414 ^ n12333;
  assign n12426 = n12399 ^ n12388;
  assign n12428 = n12427 ^ n12426;
  assign n12438 = n12437 ^ n12428;
  assign n12425 = n12410 ^ n12231;
  assign n12429 = n12428 ^ n12360;
  assign n12430 = n12429 ^ n12397;
  assign n12431 = n12425 & ~n12430;
  assign n12432 = ~n12385 & n12431;
  assign n12433 = n12428 ^ n12400;
  assign n12434 = n12433 ^ n12362;
  assign n12435 = ~n12269 & n12434;
  assign n12436 = ~n12432 & ~n12435;
  assign n12439 = n12438 ^ n12436;
  assign n12440 = n12439 ^ n12436;
  assign n12441 = n12267 & n12440;
  assign n12442 = n12441 ^ n12436;
  assign n12443 = n12424 & n12442;
  assign n12444 = n12443 ^ n12436;
  assign n12445 = ~n12423 & ~n12444;
  assign n12446 = ~n12415 & n12445;
  assign n12447 = ~n12413 & n12446;
  assign n12448 = ~n12409 & n12447;
  assign n12449 = ~n12404 & n12448;
  assign n12450 = n12449 ^ n10134;
  assign n13646 = n12450 ^ x508;
  assign n13647 = ~n13645 & ~n13646;
  assign n9400 = n9399 ^ n9141;
  assign n9731 = n9729 ^ n9571;
  assign n9730 = n9571 & ~n9729;
  assign n9732 = n9731 ^ n9730;
  assign n9733 = n9400 & n9732;
  assign n9744 = n9743 ^ n9398;
  assign n9745 = n9744 ^ n8935;
  assign n9746 = n9745 ^ n9735;
  assign n9747 = n9730 & ~n9746;
  assign n9752 = n9751 ^ n9143;
  assign n9762 = n9761 ^ n9752;
  assign n9763 = ~n9747 & ~n9762;
  assign n9764 = ~n9733 & n9763;
  assign n9769 = n9141 ^ n8450;
  assign n9770 = n9757 ^ n9398;
  assign n9771 = n9769 & ~n9770;
  assign n9772 = n9771 ^ n9755;
  assign n9766 = n9765 ^ n9734;
  assign n9767 = n9139 & n9766;
  assign n9768 = n9767 ^ n9765;
  assign n9773 = n9772 ^ n9768;
  assign n9774 = n9729 & n9773;
  assign n9775 = n9774 ^ n9768;
  assign n9776 = ~n9731 & n9775;
  assign n9777 = n9764 & ~n9776;
  assign n9778 = n9777 ^ n9192;
  assign n9779 = n9778 ^ x449;
  assign n10170 = n10169 ^ n10149;
  assign n10171 = n10170 ^ n10139;
  assign n10172 = n10171 ^ n10144;
  assign n10173 = n9968 & n10172;
  assign n10174 = n10173 ^ n10144;
  assign n10175 = n10164 & n10174;
  assign n10182 = n10165 & ~n10181;
  assign n10184 = n10183 ^ n10182;
  assign n10185 = n10151 ^ n10144;
  assign n10186 = ~n10181 & n10185;
  assign n10189 = n10188 ^ n10141;
  assign n10190 = ~n9934 & n10189;
  assign n10191 = ~n10186 & ~n10190;
  assign n10194 = n10177 & n10193;
  assign n10195 = n10154 ^ n10145;
  assign n10196 = n10180 & n10195;
  assign n10197 = ~n10164 & n10166;
  assign n10199 = n10187 ^ n10165;
  assign n10198 = n10095 ^ n10056;
  assign n10200 = n10199 ^ n10198;
  assign n10201 = n10176 & ~n10200;
  assign n10202 = ~n10197 & ~n10201;
  assign n10203 = ~n10196 & n10202;
  assign n10204 = ~n10194 & n10203;
  assign n10205 = n10191 & n10204;
  assign n10206 = ~n10184 & n10205;
  assign n10207 = ~n10179 & n10206;
  assign n10208 = ~n10175 & n10207;
  assign n10209 = ~n10163 & n10208;
  assign n10210 = n10209 ^ n9627;
  assign n10211 = n10210 ^ x450;
  assign n10212 = n9779 & ~n10211;
  assign n10213 = n10212 ^ n9779;
  assign n10460 = n10459 ^ n10458;
  assign n10464 = n10463 ^ n10460;
  assign n10465 = ~n10251 & n10464;
  assign n10466 = n10465 ^ n10460;
  assign n10467 = n10454 & n10466;
  assign n10472 = ~n10454 & n10471;
  assign n10474 = ~n10254 & n10473;
  assign n10487 = n10486 ^ n10483;
  assign n10481 = n10480 ^ n10476;
  assign n10488 = n10487 ^ n10481;
  assign n10489 = n10488 ^ n10481;
  assign n10490 = ~n10251 & n10489;
  assign n10491 = n10490 ^ n10481;
  assign n10492 = ~n10214 & n10491;
  assign n10493 = n10492 ^ n10481;
  assign n10497 = ~n10251 & n10496;
  assign n10495 = n10460 & ~n10494;
  assign n10498 = n10497 ^ n10495;
  assign n10499 = ~n10493 & ~n10498;
  assign n10500 = ~n10254 & n10485;
  assign n10503 = n10496 ^ n10452;
  assign n10502 = ~n10254 & n10501;
  assign n10504 = n10503 ^ n10502;
  assign n10505 = n10504 ^ n10478;
  assign n10506 = n10505 ^ n10462;
  assign n10507 = n10506 ^ n10253;
  assign n10508 = n10484 ^ n10482;
  assign n10509 = n10508 ^ n10506;
  assign n10510 = n10509 ^ n10502;
  assign n10511 = ~n10507 & ~n10510;
  assign n10512 = n10511 ^ n10253;
  assign n10513 = ~n10500 & n10512;
  assign n10514 = n10499 & n10513;
  assign n10515 = ~n10474 & n10514;
  assign n10516 = ~n10472 & n10515;
  assign n10517 = n10480 ^ n10470;
  assign n10518 = n10214 & n10517;
  assign n10519 = n10518 ^ n10480;
  assign n10520 = ~n10251 & n10519;
  assign n10521 = n10516 & ~n10520;
  assign n10522 = ~n10467 & n10521;
  assign n10523 = ~n10453 & n10522;
  assign n10524 = n10523 ^ n9605;
  assign n10525 = n10524 ^ x451;
  assign n10741 = n10740 ^ x452;
  assign n10742 = ~n10525 & ~n10741;
  assign n10750 = n10742 ^ n10525;
  assign n10751 = n10750 ^ n10741;
  assign n10754 = n10213 & ~n10751;
  assign n10761 = n10754 ^ n10213;
  assign n10756 = n10212 & ~n10751;
  assign n10757 = n10756 ^ n10751;
  assign n10752 = n10751 ^ n10525;
  assign n10753 = n10212 & ~n10752;
  assign n10755 = n10754 ^ n10753;
  assign n10758 = n10757 ^ n10755;
  assign n10744 = n10525 ^ n9779;
  assign n10745 = n10744 ^ n10741;
  assign n10746 = n10741 ^ n10525;
  assign n10747 = n10211 & n10746;
  assign n10748 = n10747 ^ n10525;
  assign n10749 = ~n10745 & n10748;
  assign n10759 = n10758 ^ n10749;
  assign n10743 = n10213 & n10742;
  assign n10760 = n10759 ^ n10743;
  assign n10762 = n10761 ^ n10760;
  assign n11009 = n11008 ^ x453;
  assign n11052 = n11050 & n11051;
  assign n11053 = n11049 & n11052;
  assign n11054 = ~n11041 & n11053;
  assign n11059 = n11051 & n11058;
  assign n11060 = n11059 ^ n11056;
  assign n11061 = n11050 & n11060;
  assign n11062 = ~n11054 & ~n11061;
  assign n11082 = n11039 & n11053;
  assign n11080 = n11052 & n11079;
  assign n11066 = n11065 ^ n11063;
  assign n11067 = n11052 ^ n11050;
  assign n11068 = n11066 & n11067;
  assign n11081 = n11080 ^ n11068;
  assign n11083 = n11082 ^ n11081;
  assign n11087 = n11053 & ~n11064;
  assign n11088 = n11052 ^ n11051;
  assign n11099 = n11098 ^ n11076;
  assign n11107 = n11106 ^ n11099;
  assign n11108 = n11088 & n11107;
  assign n11109 = ~n11087 & ~n11108;
  assign n11110 = n11104 ^ n11090;
  assign n11111 = n11110 ^ n11074;
  assign n11112 = n11111 ^ n11102;
  assign n11113 = ~n11050 & ~n11112;
  assign n11114 = n11113 ^ n11102;
  assign n11115 = ~n11051 & n11114;
  assign n11116 = n11109 & ~n11115;
  assign n11118 = n11050 & n11091;
  assign n11120 = n11119 ^ n11118;
  assign n11121 = ~n11117 & n11120;
  assign n11122 = n11121 ^ n11119;
  assign n11123 = n11116 & ~n11122;
  assign n11124 = ~n11086 & n11123;
  assign n11125 = ~n11083 & n11124;
  assign n11126 = n11062 & n11125;
  assign n11127 = n11126 ^ n9311;
  assign n11128 = n11127 ^ x448;
  assign n11132 = n10213 ^ n10211;
  assign n11142 = n11132 ^ n9779;
  assign n11143 = n10742 & ~n11142;
  assign n11144 = n11143 ^ n11142;
  assign n11133 = ~n10750 & n11132;
  assign n11139 = n11133 ^ n10750;
  assign n11137 = n10212 & ~n10750;
  assign n11138 = n11137 ^ n10759;
  assign n11140 = n11139 ^ n11138;
  assign n11134 = n11133 ^ n10743;
  assign n11135 = n11134 ^ n10748;
  assign n11129 = n10756 ^ n10743;
  assign n11130 = n11129 ^ n10754;
  assign n11131 = n11130 ^ n10749;
  assign n11136 = n11135 ^ n11131;
  assign n11141 = n11140 ^ n11136;
  assign n11145 = n11144 ^ n11141;
  assign n11146 = n11145 ^ n11140;
  assign n11147 = ~n11128 & ~n11146;
  assign n11148 = n11147 ^ n11140;
  assign n11149 = ~n11009 & n11148;
  assign n11150 = n11145 ^ n10754;
  assign n11151 = n11150 ^ n10757;
  assign n11153 = ~n11009 & n11128;
  assign n11152 = n11128 ^ n11009;
  assign n11154 = n11153 ^ n11152;
  assign n11155 = n11151 & n11154;
  assign n11156 = ~n11138 & n11154;
  assign n11158 = n11143 ^ n11133;
  assign n11157 = n10212 & n10742;
  assign n11159 = n11158 ^ n11157;
  assign n11160 = n11159 ^ n10742;
  assign n11161 = n11160 ^ n11134;
  assign n11162 = n11161 ^ n11157;
  assign n11163 = ~n11152 & n11162;
  assign n11172 = n11009 & n11131;
  assign n11173 = n11172 ^ n11130;
  assign n11167 = n11145 ^ n11143;
  assign n11166 = n11136 ^ n11133;
  assign n11168 = n11167 ^ n11166;
  assign n11164 = n11140 ^ n10743;
  assign n11165 = n11164 ^ n10755;
  assign n11169 = n11168 ^ n11165;
  assign n11170 = n11009 & ~n11169;
  assign n11171 = n11170 ^ n11165;
  assign n11174 = n11173 ^ n11171;
  assign n11175 = ~n11128 & n11174;
  assign n11176 = n11175 ^ n11173;
  assign n11177 = ~n11163 & ~n11176;
  assign n11178 = ~n11156 & n11177;
  assign n11180 = n11135 ^ n10525;
  assign n11181 = n11180 ^ n10761;
  assign n11182 = n11128 & n11181;
  assign n11179 = n11153 & n11158;
  assign n11183 = n11182 ^ n11179;
  assign n11184 = n11178 & ~n11183;
  assign n11185 = ~n11155 & n11184;
  assign n11186 = ~n11149 & n11185;
  assign n11187 = n10762 & n11186;
  assign n11188 = n11187 ^ n9967;
  assign n13648 = n11188 ^ x509;
  assign n12915 = n12329 ^ x471;
  assign n11292 = ~n11051 & n11075;
  assign n11289 = n11098 ^ n11095;
  assign n11290 = n11051 & ~n11289;
  assign n11291 = n11290 ^ n11095;
  assign n11293 = n11292 ^ n11291;
  assign n11294 = ~n11050 & ~n11293;
  assign n11295 = n11294 ^ n11291;
  assign n12053 = n11111 ^ n11092;
  assign n12054 = ~n11050 & ~n12053;
  assign n12055 = n12054 ^ n11092;
  assign n12048 = n11105 ^ n11103;
  assign n12049 = n12048 ^ n11079;
  assign n11296 = n11105 ^ n11095;
  assign n12047 = n11296 ^ n11119;
  assign n12050 = n12049 ^ n12047;
  assign n12051 = ~n11050 & ~n12050;
  assign n12052 = n12051 ^ n12049;
  assign n12056 = n12055 ^ n12052;
  assign n12057 = n11051 & n12056;
  assign n12058 = n12057 ^ n12052;
  assign n12060 = ~n11117 & n11299;
  assign n12059 = ~n11051 & n11098;
  assign n12061 = n12060 ^ n12059;
  assign n12062 = ~n12058 & ~n12061;
  assign n12063 = ~n11083 & n12062;
  assign n12064 = n11295 & n12063;
  assign n12065 = n12064 ^ n8780;
  assign n12916 = n12065 ^ x466;
  assign n12818 = n10805 & n11278;
  assign n12819 = ~n10805 & n10952;
  assign n12820 = n10973 ^ n10966;
  assign n12821 = n10806 ^ n10790;
  assign n12822 = n12820 & ~n12821;
  assign n12823 = n10922 ^ n10882;
  assign n12824 = n12823 ^ n11263;
  assign n12825 = ~n10807 & ~n12824;
  assign n12832 = n10805 & ~n10963;
  assign n12826 = n12820 ^ n10933;
  assign n12827 = n12826 ^ n10931;
  assign n12828 = n10806 & n12827;
  assign n12829 = n12828 ^ n10931;
  assign n12830 = n12826 & n12829;
  assign n12831 = ~n10940 & ~n12830;
  assign n12833 = n12832 ^ n12831;
  assign n12834 = n10934 & ~n12833;
  assign n12835 = n12834 ^ n12831;
  assign n12836 = ~n12825 & n12835;
  assign n12837 = ~n10925 & n12836;
  assign n12838 = ~n12822 & n12837;
  assign n12839 = ~n12819 & n12838;
  assign n12840 = n10962 ^ n10958;
  assign n12841 = ~n10805 & ~n12840;
  assign n12842 = n12841 ^ n10958;
  assign n12843 = ~n10934 & n12842;
  assign n12844 = n12839 & ~n12843;
  assign n12845 = ~n12818 & n12844;
  assign n12846 = ~n11254 & n12845;
  assign n12847 = n12846 ^ n10313;
  assign n12848 = n12847 ^ x469;
  assign n11208 = n10473 & ~n10494;
  assign n11209 = n11208 ^ n10453;
  assign n11240 = n10469 ^ n10452;
  assign n11221 = n10478 ^ n10461;
  assign n12852 = n11240 ^ n11221;
  assign n12850 = n10470 ^ n10463;
  assign n12851 = n12850 ^ n10460;
  assign n12853 = n12852 ^ n12851;
  assign n12854 = ~n10251 & n12853;
  assign n12855 = n12854 ^ n12851;
  assign n12856 = ~n10454 & n12855;
  assign n12862 = n10486 ^ n10471;
  assign n12863 = ~n10253 & n12862;
  assign n12858 = n11972 ^ n10480;
  assign n12859 = n10454 & n12858;
  assign n12860 = n12859 ^ n10480;
  assign n12857 = ~n10251 & n10483;
  assign n12861 = n12860 ^ n12857;
  assign n12864 = n12863 ^ n12861;
  assign n12865 = ~n12856 & ~n12864;
  assign n12866 = ~n11962 & n12865;
  assign n12867 = ~n11209 & n12866;
  assign n12868 = ~n10502 & n12867;
  assign n12869 = n12868 ^ n10285;
  assign n12870 = n12869 ^ x468;
  assign n11828 = ~n10152 & n10177;
  assign n11840 = ~n9934 & n10139;
  assign n11836 = n11835 ^ n10140;
  assign n11837 = n11836 ^ n10158;
  assign n11838 = n9934 & n11837;
  assign n11839 = n11838 ^ n10158;
  assign n11841 = n11840 ^ n11839;
  assign n11842 = ~n9968 & ~n11841;
  assign n11843 = n11842 ^ n11839;
  assign n11847 = n10151 ^ n10141;
  assign n11848 = ~n9968 & n11847;
  assign n11849 = n11848 ^ n10151;
  assign n11850 = ~n10164 & n11849;
  assign n12006 = ~n9968 & n10188;
  assign n12007 = n12006 ^ n10145;
  assign n12008 = n10164 & n12007;
  assign n12009 = n12008 ^ n10145;
  assign n12010 = n10176 ^ n10169;
  assign n12011 = n10149 ^ n9934;
  assign n12012 = ~n10169 & ~n12011;
  assign n12013 = n12012 ^ n10149;
  assign n12014 = ~n12010 & n12013;
  assign n12015 = n12014 ^ n10176;
  assign n12016 = ~n12009 & ~n12015;
  assign n12020 = n9968 & ~n12019;
  assign n12021 = n12020 ^ n10140;
  assign n12022 = ~n9934 & n12021;
  assign n12023 = n12016 & ~n12022;
  assign n12024 = ~n10184 & n12023;
  assign n12025 = ~n12005 & n12024;
  assign n12026 = ~n11850 & n12025;
  assign n12027 = ~n11831 & n12026;
  assign n12028 = n11843 & n12027;
  assign n12029 = ~n12003 & n12028;
  assign n12030 = ~n11828 & n12029;
  assign n12031 = ~n10163 & n12030;
  assign n12032 = n12031 ^ n8646;
  assign n12849 = n12032 ^ x467;
  assign n12878 = n12870 ^ n12849;
  assign n12872 = n12266 ^ x470;
  assign n12873 = ~n12870 & ~n12872;
  assign n12874 = n12873 ^ n12849;
  assign n12871 = n12849 & n12870;
  assign n12875 = n12874 ^ n12871;
  assign n12876 = n12875 ^ n12872;
  assign n12894 = n12878 ^ n12876;
  assign n12895 = n12894 ^ n12872;
  assign n12922 = n12848 & ~n12895;
  assign n12879 = n12878 ^ n12872;
  assign n12923 = n12922 ^ n12879;
  assign n13686 = ~n12916 & ~n12923;
  assign n12906 = n12848 & n12849;
  assign n12891 = n12849 ^ n12848;
  assign n12899 = ~n12870 & n12891;
  assign n12900 = n12899 ^ n12849;
  assign n12901 = ~n12879 & ~n12900;
  assign n12902 = n12901 ^ n12872;
  assign n12882 = n12870 ^ n12848;
  assign n12883 = ~n12849 & ~n12872;
  assign n12884 = n12883 ^ n12873;
  assign n12885 = n12884 ^ n12879;
  assign n12886 = n12885 ^ n12870;
  assign n12887 = ~n12882 & n12886;
  assign n12897 = n12887 ^ n12872;
  assign n12898 = n12897 ^ n12848;
  assign n12903 = n12902 ^ n12898;
  assign n12905 = n12903 ^ n12891;
  assign n12907 = n12906 ^ n12905;
  assign n12896 = n12895 ^ n12884;
  assign n12904 = n12903 ^ n12896;
  assign n12908 = n12907 ^ n12904;
  assign n12909 = n12908 ^ n12848;
  assign n12910 = n12909 ^ n12883;
  assign n12889 = n12872 ^ n12871;
  assign n12890 = n12882 & ~n12889;
  assign n12892 = n12891 ^ n12890;
  assign n12877 = ~n12848 & ~n12876;
  assign n12888 = n12887 ^ n12877;
  assign n12893 = n12892 ^ n12888;
  assign n12911 = n12910 ^ n12893;
  assign n12881 = n12878 ^ n12848;
  assign n12912 = n12911 ^ n12881;
  assign n12880 = n12879 ^ n12877;
  assign n12913 = n12912 ^ n12880;
  assign n12914 = n12913 ^ n12905;
  assign n13687 = n13686 ^ n12914;
  assign n13688 = ~n12915 & ~n13687;
  assign n13689 = n13688 ^ n12914;
  assign n13693 = n12898 & n12915;
  assign n12919 = n12872 ^ n12870;
  assign n12920 = n12919 ^ n12848;
  assign n12921 = n12920 ^ n12893;
  assign n13690 = n12921 ^ n12902;
  assign n13691 = n12915 & ~n13690;
  assign n13692 = n13691 ^ n12921;
  assign n13694 = n13693 ^ n13692;
  assign n13695 = ~n12916 & ~n13694;
  assign n13696 = n13695 ^ n13692;
  assign n13697 = n13689 & n13696;
  assign n13698 = n13697 ^ n11374;
  assign n13699 = n13698 ^ x510;
  assign n13706 = n13648 & n13699;
  assign n13707 = n13706 ^ n13699;
  assign n13708 = n13707 ^ n13648;
  assign n11207 = n11206 ^ x478;
  assign n11210 = n10501 ^ n10480;
  assign n11211 = ~n10253 & n11210;
  assign n11214 = n11213 ^ n10480;
  assign n11215 = ~n10494 & n11214;
  assign n11216 = n10502 ^ n10253;
  assign n11217 = n10504 ^ n10471;
  assign n11218 = ~n11216 & n11217;
  assign n11219 = ~n11215 & ~n11218;
  assign n11220 = ~n11211 & n11219;
  assign n11222 = n10482 ^ n10480;
  assign n11223 = n11222 ^ n10485;
  assign n11224 = n11223 ^ n11212;
  assign n11225 = n11223 ^ n10251;
  assign n11226 = n10454 & n11225;
  assign n11227 = n11226 ^ n10251;
  assign n11228 = n11224 & ~n11227;
  assign n11229 = n11228 ^ n11212;
  assign n11230 = ~n11221 & ~n11229;
  assign n11231 = ~n10459 & n11230;
  assign n11232 = n11231 ^ n10252;
  assign n11233 = n10470 ^ n10458;
  assign n11234 = n11233 ^ n10254;
  assign n11235 = n11231 & n11234;
  assign n11236 = n11235 ^ n10254;
  assign n11237 = ~n11232 & ~n11236;
  assign n11238 = n11237 ^ n10252;
  assign n11239 = n11220 & ~n11238;
  assign n11241 = n10251 & n11240;
  assign n11242 = n11241 ^ n10452;
  assign n11243 = n10214 & n11242;
  assign n11244 = n11239 & ~n11243;
  assign n11245 = ~n10467 & n11244;
  assign n11246 = ~n11209 & n11245;
  assign n11247 = n11246 ^ n9482;
  assign n11248 = n11247 ^ x483;
  assign n11421 = n11420 ^ n11419;
  assign n11425 = n11424 ^ n11421;
  assign n11426 = n11403 ^ n11398;
  assign n11427 = n11426 ^ n11386;
  assign n11429 = n11428 ^ n11384;
  assign n11430 = n11426 & n11429;
  assign n11431 = n11430 ^ n11384;
  assign n11432 = ~n11427 & ~n11431;
  assign n11433 = n11432 ^ n11386;
  assign n11439 = n11408 ^ n11400;
  assign n11440 = n11439 ^ n11434;
  assign n11441 = n11440 ^ n11395;
  assign n11438 = n11437 ^ n11403;
  assign n11442 = n11441 ^ n11438;
  assign n11443 = ~n11382 & n11442;
  assign n11444 = n11443 ^ n11438;
  assign n11445 = ~n11381 & ~n11444;
  assign n11448 = n11439 ^ n11437;
  assign n11447 = n11446 ^ n11391;
  assign n11449 = n11448 ^ n11447;
  assign n11450 = ~n11382 & n11449;
  assign n11451 = n11450 ^ n11447;
  assign n11452 = n11451 ^ n11401;
  assign n11453 = n11451 ^ n11385;
  assign n11454 = n11451 & n11453;
  assign n11455 = n11454 ^ n11451;
  assign n11456 = ~n11452 & n11455;
  assign n11457 = n11456 ^ n11454;
  assign n11458 = n11457 ^ n11451;
  assign n11459 = n11458 ^ n11385;
  assign n11460 = ~n11445 & n11459;
  assign n11461 = n11460 ^ n11445;
  assign n11462 = ~n11433 & ~n11461;
  assign n11463 = ~n11425 & n11462;
  assign n11464 = ~n11417 & n11463;
  assign n11465 = ~n11413 & n11464;
  assign n11466 = n11465 ^ n9427;
  assign n11467 = n11466 ^ x482;
  assign n11304 = ~n11067 & n11303;
  assign n11297 = n11296 ^ n11069;
  assign n11305 = n11304 ^ n11297;
  assign n11306 = ~n11088 & ~n11305;
  assign n11307 = n11306 ^ n11297;
  assign n11308 = n11102 ^ n11056;
  assign n11309 = n11308 ^ n11095;
  assign n11310 = n11309 ^ n11050;
  assign n11311 = n11309 ^ n11051;
  assign n11312 = ~n11309 & n11311;
  assign n11313 = n11312 ^ n11309;
  assign n11314 = n11310 & ~n11313;
  assign n11315 = n11314 ^ n11312;
  assign n11316 = n11315 ^ n11309;
  assign n11317 = n11316 ^ n11051;
  assign n11318 = ~n11299 & n11317;
  assign n11319 = n11318 ^ n11051;
  assign n11320 = n11307 & n11319;
  assign n11329 = n11050 & n11076;
  assign n11321 = n11119 ^ n11091;
  assign n11322 = n11321 ^ n11300;
  assign n11323 = n11300 ^ n11050;
  assign n11324 = ~n11117 & n11323;
  assign n11325 = n11324 ^ n11050;
  assign n11326 = n11322 & ~n11325;
  assign n11327 = n11326 ^ n11321;
  assign n11328 = ~n11103 & ~n11327;
  assign n11330 = n11329 ^ n11328;
  assign n11331 = ~n11117 & ~n11330;
  assign n11332 = n11331 ^ n11328;
  assign n11333 = n11320 & n11332;
  assign n11334 = ~n11068 & n11333;
  assign n11335 = n11295 & n11334;
  assign n11336 = n11062 & n11335;
  assign n11337 = n11336 ^ n9812;
  assign n11338 = n11337 ^ x480;
  assign n11288 = n11287 ^ x479;
  assign n11589 = n11542 & ~n11588;
  assign n11593 = n11592 ^ n11578;
  assign n11605 = n11604 ^ n11593;
  assign n11606 = n11546 & n11605;
  assign n11607 = ~n11589 & ~n11606;
  assign n11608 = n11563 ^ n11561;
  assign n11609 = n11544 & n11608;
  assign n11617 = n11568 ^ n11540;
  assign n11618 = n11617 ^ n11591;
  assign n11619 = n11618 ^ n11592;
  assign n11620 = ~n11541 & ~n11619;
  assign n11621 = n11620 ^ n11592;
  assign n11611 = n11598 ^ n11592;
  assign n11612 = n11611 ^ n11577;
  assign n11613 = n11612 ^ n11551;
  assign n11610 = n11563 ^ n11553;
  assign n11614 = n11613 ^ n11610;
  assign n11615 = n11541 & n11614;
  assign n11616 = n11615 ^ n11610;
  assign n11622 = n11621 ^ n11616;
  assign n11623 = ~n11542 & n11622;
  assign n11624 = n11623 ^ n11616;
  assign n11625 = ~n11609 & ~n11624;
  assign n11626 = n11607 & n11625;
  assign n11627 = ~n11587 & n11626;
  assign n11628 = ~n11583 & n11627;
  assign n11629 = ~n11581 & n11628;
  assign n11630 = ~n11545 & n11629;
  assign n11631 = n11630 ^ n9850;
  assign n11632 = n11631 ^ x481;
  assign n11633 = ~n11288 & n11632;
  assign n11634 = n11633 ^ n11288;
  assign n11635 = n11634 ^ n11632;
  assign n11640 = n11338 & n11635;
  assign n11641 = ~n11467 & n11640;
  assign n11674 = n11641 ^ n11640;
  assign n11636 = n11338 & ~n11467;
  assign n11643 = n11633 ^ n11632;
  assign n11644 = n11636 & n11643;
  assign n12692 = n11674 ^ n11644;
  assign n11651 = n11636 ^ n11467;
  assign n11652 = n11633 & ~n11651;
  assign n11637 = n11636 ^ n11338;
  assign n11650 = n11633 & n11637;
  assign n11653 = n11652 ^ n11650;
  assign n11649 = n11633 & n11636;
  assign n11654 = n11653 ^ n11649;
  assign n11655 = n11654 ^ n11633;
  assign n13304 = n12692 ^ n11655;
  assign n13305 = n11248 & n13304;
  assign n13306 = n13305 ^ n11655;
  assign n13307 = n11207 & n13306;
  assign n11249 = n11207 & n11248;
  assign n11250 = n11249 ^ n11207;
  assign n11251 = n11250 ^ n11248;
  assign n11252 = n11251 ^ n11207;
  assign n11638 = n11637 ^ n11467;
  assign n11688 = ~n11634 & n11638;
  assign n13649 = n11688 ^ n11654;
  assign n13650 = n11252 & n13649;
  assign n11658 = n11640 ^ n11635;
  assign n11639 = n11635 & n11638;
  assign n11659 = n11658 ^ n11639;
  assign n11642 = n11641 ^ n11639;
  assign n11645 = n11644 ^ n11642;
  assign n11468 = n11467 ^ n11338;
  assign n11469 = n11288 & n11468;
  assign n11646 = n11645 ^ n11469;
  assign n13651 = n11659 ^ n11646;
  assign n13652 = n11249 & n13651;
  assign n11647 = n11252 & n11646;
  assign n13310 = n11659 ^ n11207;
  assign n11669 = n11646 ^ n11644;
  assign n11661 = ~n11634 & ~n11651;
  assign n11662 = n11661 ^ n11650;
  assign n11663 = n11662 ^ n11651;
  assign n11660 = n11659 ^ n11653;
  assign n11664 = n11663 ^ n11660;
  assign n11670 = n11669 ^ n11664;
  assign n11671 = n11670 ^ n11643;
  assign n13653 = n11671 ^ n11669;
  assign n13654 = n13653 ^ n11642;
  assign n13655 = ~n11248 & ~n13654;
  assign n13656 = n13655 ^ n11642;
  assign n13657 = n13656 ^ n11659;
  assign n13658 = n13310 & n13657;
  assign n13659 = n13658 ^ n13655;
  assign n13660 = n13659 ^ n11642;
  assign n13661 = n13660 ^ n11207;
  assign n13662 = ~n11659 & n13661;
  assign n13663 = n13662 ^ n11659;
  assign n13664 = n13663 ^ n11207;
  assign n11672 = n11671 ^ n11664;
  assign n13665 = n11672 ^ n11640;
  assign n11678 = n11645 ^ n11636;
  assign n11677 = n11649 ^ n11639;
  assign n11679 = n11678 ^ n11677;
  assign n11689 = n11688 ^ n11679;
  assign n11690 = n11689 ^ n11655;
  assign n11691 = n11690 ^ n11661;
  assign n13666 = n13665 ^ n11691;
  assign n13667 = n11248 & n13666;
  assign n13668 = n13667 ^ n13665;
  assign n13669 = n11207 & n13668;
  assign n13670 = ~n13664 & ~n13669;
  assign n13671 = ~n11647 & n13670;
  assign n13672 = ~n13652 & n13671;
  assign n13673 = ~n13650 & n13672;
  assign n13675 = n11689 ^ n11653;
  assign n11687 = n11654 ^ n11288;
  assign n11692 = n11691 ^ n11687;
  assign n12707 = n11692 ^ n11652;
  assign n13674 = n12707 ^ n11649;
  assign n13676 = n13675 ^ n13674;
  assign n13677 = ~n11207 & ~n13676;
  assign n13678 = n13677 ^ n13674;
  assign n13679 = ~n11248 & ~n13678;
  assign n13680 = n13673 & ~n13679;
  assign n13681 = ~n13307 & n13680;
  assign n13682 = n13681 ^ n11364;
  assign n13683 = n13682 ^ x511;
  assign n11746 = n10644 & ~n10683;
  assign n11747 = n10625 & ~n10692;
  assign n11754 = n11753 ^ n10635;
  assign n11755 = n11754 ^ n10642;
  assign n11756 = n11755 ^ n10633;
  assign n11757 = n10680 & ~n11756;
  assign n11758 = n11757 ^ n10633;
  assign n11749 = n10700 ^ n10694;
  assign n11748 = n10701 ^ n10622;
  assign n11750 = n11749 ^ n11748;
  assign n11751 = ~n10680 & n11750;
  assign n11752 = n11751 ^ n11748;
  assign n11759 = n11758 ^ n11752;
  assign n11760 = ~n10693 & n11759;
  assign n11761 = n11760 ^ n11758;
  assign n11762 = ~n11747 & ~n11761;
  assign n11764 = ~n10680 & n10696;
  assign n11763 = ~n10682 & ~n10719;
  assign n11765 = n11764 ^ n11763;
  assign n11766 = n11762 & ~n11765;
  assign n11768 = n10646 & n10681;
  assign n11767 = n10686 & ~n10693;
  assign n11769 = n11768 ^ n11767;
  assign n11770 = n11766 & ~n11769;
  assign n11771 = ~n11746 & n11770;
  assign n11772 = ~n10691 & n11771;
  assign n11773 = ~n10684 & n11772;
  assign n11774 = n11773 ^ n9220;
  assign n12452 = n11774 ^ x489;
  assign n12453 = n11466 ^ x484;
  assign n12487 = n11191 ^ n9729;
  assign n12488 = n12487 ^ n11195;
  assign n12489 = n12488 ^ n11192;
  assign n12484 = n9760 ^ n9729;
  assign n12485 = n12484 ^ n11202;
  assign n12486 = n12485 ^ n11199;
  assign n12490 = n12489 ^ n12486;
  assign n12491 = ~n9571 & ~n12490;
  assign n12492 = n12491 ^ n12489;
  assign n12493 = n12492 ^ n9486;
  assign n12494 = n12493 ^ x486;
  assign n11852 = n10165 ^ n10145;
  assign n11853 = n11852 ^ n11837;
  assign n11851 = n10154 ^ n10147;
  assign n11854 = n11853 ^ n11851;
  assign n11855 = n11854 ^ n11851;
  assign n11856 = ~n9968 & n11855;
  assign n11857 = n11856 ^ n11851;
  assign n11858 = n10164 & n11857;
  assign n11859 = n11858 ^ n11851;
  assign n11861 = ~n9934 & ~n10156;
  assign n11860 = n10167 & n10180;
  assign n11862 = n11861 ^ n11860;
  assign n11863 = ~n11859 & ~n11862;
  assign n11864 = ~n11850 & n11863;
  assign n11865 = ~n11846 & n11864;
  assign n11866 = n11843 & n11865;
  assign n11867 = ~n11833 & n11866;
  assign n11868 = ~n11828 & n11867;
  assign n11869 = ~n10175 & n11868;
  assign n11870 = ~n10183 & n11869;
  assign n11871 = n11870 ^ n9181;
  assign n12495 = n11871 ^ x488;
  assign n12496 = ~n12494 & ~n12495;
  assign n12506 = n12496 ^ n12494;
  assign n12458 = n10960 ^ n10934;
  assign n12459 = n10952 ^ n10805;
  assign n12460 = n10960 & n12459;
  assign n12461 = n12460 ^ n10805;
  assign n12462 = n12458 & n12461;
  assign n12463 = n12462 ^ n10960;
  assign n12469 = n10968 ^ n10966;
  assign n12470 = ~n10805 & n12469;
  assign n12471 = n12470 ^ n10966;
  assign n12465 = n11264 ^ n11253;
  assign n12464 = n11275 ^ n10985;
  assign n12466 = n12465 ^ n12464;
  assign n12467 = n10805 & n12466;
  assign n12468 = n12467 ^ n12464;
  assign n12472 = n12471 ^ n12468;
  assign n12473 = ~n10790 & ~n12472;
  assign n12474 = n12473 ^ n12471;
  assign n12475 = n12463 & ~n12474;
  assign n12476 = n10978 & n12475;
  assign n12477 = n11262 & n12476;
  assign n12478 = ~n11256 & n12477;
  assign n12479 = ~n10925 & n12478;
  assign n12480 = n12479 ^ n9459;
  assign n12481 = n12480 ^ x487;
  assign n12482 = n11247 ^ x485;
  assign n12483 = ~n12481 & ~n12482;
  assign n12507 = n12483 ^ n12482;
  assign n12508 = n12507 ^ n12481;
  assign n12509 = ~n12506 & ~n12508;
  assign n12545 = n12509 ^ n12508;
  assign n12531 = n12496 & ~n12508;
  assign n12497 = n12496 ^ n12495;
  assign n12498 = n12497 ^ n12494;
  assign n12526 = ~n12498 & ~n12508;
  assign n12535 = n12531 ^ n12526;
  assign n12546 = n12545 ^ n12535;
  assign n12520 = n12483 ^ n12481;
  assign n12523 = n12496 & ~n12520;
  assign n12524 = n12523 ^ n12520;
  assign n12521 = ~n12497 & ~n12520;
  assign n12514 = ~n12506 & ~n12507;
  assign n12502 = n12483 & ~n12497;
  assign n12515 = n12514 ^ n12502;
  assign n12516 = n12515 ^ n12506;
  assign n12503 = n12502 ^ n12483;
  assign n12500 = n12483 & n12496;
  assign n12499 = n12483 & ~n12498;
  assign n12501 = n12500 ^ n12499;
  assign n12504 = n12503 ^ n12501;
  assign n12505 = n12504 ^ n12502;
  assign n12510 = n12509 ^ n12505;
  assign n12517 = n12516 ^ n12510;
  assign n12522 = n12521 ^ n12517;
  assign n12525 = n12524 ^ n12522;
  assign n12773 = n12546 ^ n12525;
  assign n12774 = n12773 ^ n12522;
  assign n12775 = ~n12453 & n12774;
  assign n12776 = n12775 ^ n12773;
  assign n12777 = n12452 & ~n12776;
  assign n12538 = n12496 & ~n12507;
  assign n12778 = n12538 ^ n12514;
  assign n12528 = n12499 ^ n12498;
  assign n12527 = n12526 ^ n12525;
  assign n12529 = n12528 ^ n12527;
  assign n12779 = n12778 ^ n12529;
  assign n12780 = n12779 ^ n12507;
  assign n12781 = n12780 ^ n12504;
  assign n12782 = n12781 ^ n12531;
  assign n12783 = ~n12453 & n12782;
  assign n12784 = n12783 ^ n12531;
  assign n12785 = n12452 & n12784;
  assign n12547 = n12546 ^ n12529;
  assign n12544 = n12535 ^ n12525;
  assign n12548 = n12547 ^ n12544;
  assign n13446 = n12452 & n12548;
  assign n13447 = n13446 ^ n12544;
  assign n13448 = ~n12453 & n13447;
  assign n12454 = ~n12452 & ~n12453;
  assign n12456 = n12454 ^ n12453;
  assign n12518 = n12456 ^ n12452;
  assign n13450 = n12515 & ~n12518;
  assign n12455 = n12454 ^ n12452;
  assign n12457 = n12456 ^ n12455;
  assign n13449 = ~n12457 & n12781;
  assign n13451 = n13450 ^ n13449;
  assign n12557 = ~n12457 & n12523;
  assign n13452 = n13451 ^ n12557;
  assign n13453 = ~n13448 & ~n13452;
  assign n12796 = n12528 ^ n12520;
  assign n12797 = n12796 ^ n12521;
  assign n12794 = n12495 ^ n12494;
  assign n12795 = n12794 ^ n12482;
  assign n12798 = n12797 ^ n12795;
  assign n13455 = ~n12452 & ~n12798;
  assign n13454 = n12538 ^ n12499;
  assign n13456 = n13455 ^ n13454;
  assign n13457 = n12453 & n13456;
  assign n13458 = n13457 ^ n13454;
  assign n13459 = n13453 & ~n13458;
  assign n13460 = ~n12785 & n13459;
  assign n13461 = ~n12777 & n13460;
  assign n13462 = n13461 ^ n9570;
  assign n13684 = n13462 ^ x512;
  assign n13711 = n13683 & ~n13684;
  assign n13712 = n13711 ^ n13684;
  assign n13723 = n13712 ^ n13683;
  assign n13726 = ~n13708 & n13723;
  assign n13725 = ~n13708 & n13711;
  assign n13727 = n13726 ^ n13725;
  assign n13719 = ~n13708 & ~n13712;
  assign n13728 = n13727 ^ n13719;
  assign n13747 = n13728 ^ n13708;
  assign n13721 = n13648 & ~n13683;
  assign n13709 = n13708 ^ n13699;
  assign n13713 = n13709 & ~n13712;
  assign n13710 = ~n13684 & n13709;
  assign n13714 = n13713 ^ n13710;
  assign n13744 = n13721 ^ n13714;
  assign n13732 = n13723 ^ n13684;
  assign n13733 = n13706 & n13732;
  assign n13734 = n13733 ^ n13706;
  assign n13717 = n13706 & n13711;
  assign n13715 = n13714 ^ n13709;
  assign n13685 = n13684 ^ n13683;
  assign n13700 = n13699 ^ n13684;
  assign n13701 = n13700 ^ n13683;
  assign n13702 = n13701 ^ n13684;
  assign n13703 = ~n13685 & ~n13702;
  assign n13704 = n13703 ^ n13684;
  assign n13705 = n13648 & n13704;
  assign n13716 = n13715 ^ n13705;
  assign n13718 = n13717 ^ n13716;
  assign n13735 = n13734 ^ n13718;
  assign n13731 = n13716 ^ n13710;
  assign n13736 = n13735 ^ n13731;
  assign n13745 = n13744 ^ n13736;
  assign n13743 = n13710 ^ n13709;
  assign n13746 = n13745 ^ n13743;
  assign n13748 = n13747 ^ n13746;
  assign n13742 = n13733 ^ n13732;
  assign n13749 = n13748 ^ n13742;
  assign n13724 = n13707 & n13723;
  assign n13729 = n13728 ^ n13724;
  assign n13730 = n13729 ^ n13683;
  assign n13737 = n13736 ^ n13730;
  assign n13722 = n13721 ^ n13684;
  assign n13738 = n13737 ^ n13722;
  assign n13720 = n13719 ^ n13718;
  assign n13739 = n13738 ^ n13720;
  assign n13740 = n13739 ^ n13724;
  assign n13741 = n13740 ^ n13707;
  assign n13750 = n13749 ^ n13741;
  assign n13751 = n13647 & ~n13750;
  assign n13754 = n13646 & ~n13748;
  assign n13755 = n13754 ^ n13746;
  assign n13756 = n13645 & n13755;
  assign n13752 = n13645 & ~n13750;
  assign n13753 = n13646 & n13752;
  assign n13757 = n13756 ^ n13753;
  assign n13758 = n13749 ^ n13719;
  assign n13759 = n13758 ^ n13746;
  assign n13760 = n13645 & ~n13759;
  assign n13761 = n13760 ^ n13746;
  assign n13762 = n13646 & n13761;
  assign n13763 = n13646 ^ n13645;
  assign n13775 = n13740 ^ n13725;
  assign n13776 = n13775 ^ n13726;
  assign n13773 = n13749 ^ n13747;
  assign n13774 = n13773 ^ n13725;
  assign n13777 = n13776 ^ n13774;
  assign n13778 = n13776 ^ n13645;
  assign n13779 = ~n13763 & ~n13778;
  assign n13780 = n13779 ^ n13645;
  assign n13781 = n13777 & n13780;
  assign n13782 = n13781 ^ n13774;
  assign n13783 = ~n13713 & ~n13782;
  assign n13784 = ~n13718 & n13783;
  assign n13764 = n13745 ^ n13735;
  assign n13767 = n13764 ^ n13749;
  assign n13768 = n13767 ^ n13726;
  assign n13769 = n13768 ^ n13719;
  assign n13765 = n13764 ^ n13717;
  assign n13766 = n13765 ^ n13725;
  assign n13770 = n13769 ^ n13766;
  assign n13771 = ~n13646 & ~n13770;
  assign n13772 = n13771 ^ n13766;
  assign n13785 = n13784 ^ n13772;
  assign n13786 = ~n13763 & ~n13785;
  assign n13787 = n13786 ^ n13784;
  assign n13788 = ~n13762 & n13787;
  assign n13789 = n13733 ^ n13714;
  assign n13790 = n13789 ^ n13726;
  assign n13791 = ~n13646 & n13790;
  assign n13792 = n13791 ^ n13726;
  assign n13793 = ~n13645 & n13792;
  assign n13794 = n13788 & ~n13793;
  assign n13795 = ~n13757 & n13794;
  assign n13796 = ~n13751 & n13795;
  assign n13797 = n13796 ^ n11466;
  assign n15498 = n13797 ^ x578;
  assign n12533 = n12529 ^ n12502;
  assign n12534 = ~n12518 & ~n12533;
  assign n12786 = n12453 & n12501;
  assign n12787 = n12781 ^ n12525;
  assign n12788 = n12787 ^ n12521;
  assign n12789 = ~n12455 & n12788;
  assign n12790 = ~n12786 & ~n12789;
  assign n12791 = ~n12456 & n12515;
  assign n12519 = ~n12517 & ~n12518;
  assign n12792 = n12791 ^ n12519;
  assign n12793 = n12790 & ~n12792;
  assign n12799 = ~n12453 & ~n12798;
  assign n12800 = n12799 ^ n12535;
  assign n12801 = ~n12457 & n12800;
  assign n12802 = n12801 ^ n12535;
  assign n12803 = n12793 & ~n12802;
  assign n12804 = ~n12534 & n12803;
  assign n12805 = ~n12785 & n12804;
  assign n12806 = ~n12777 & n12805;
  assign n12807 = n12806 ^ n10834;
  assign n14488 = n12807 ^ x496;
  assign n13007 = n13005 ^ n12934;
  assign n13269 = n13007 ^ n12933;
  assign n13270 = n13268 & ~n13269;
  assign n13275 = n13274 ^ n13270;
  assign n14432 = ~n12933 & n12994;
  assign n14429 = n13022 & ~n13269;
  assign n14430 = n14429 ^ n13017;
  assign n14427 = n13005 & n13019;
  assign n14428 = n14427 ^ n13034;
  assign n14431 = n14430 ^ n14428;
  assign n14433 = n14432 ^ n14431;
  assign n14434 = n13013 & ~n14433;
  assign n14435 = n14434 ^ n14431;
  assign n14441 = n13008 ^ n12996;
  assign n14442 = n12933 & n14441;
  assign n14437 = n13004 & n13480;
  assign n13064 = n13004 & n13010;
  assign n14438 = n14437 ^ n13064;
  assign n13039 = n13038 ^ n13034;
  assign n13040 = n13039 ^ n13008;
  assign n14436 = n13007 & ~n13040;
  assign n14439 = n14438 ^ n14436;
  assign n14440 = n14439 ^ n13027;
  assign n14443 = n14442 ^ n14440;
  assign n14444 = ~n13013 & n14443;
  assign n14445 = n14444 ^ n14440;
  assign n14446 = n14435 & ~n14445;
  assign n14447 = n13035 ^ n13027;
  assign n14448 = n12933 & n14447;
  assign n14449 = n14448 ^ n13027;
  assign n14450 = n14449 ^ n13489;
  assign n14451 = ~n12934 & n14450;
  assign n14452 = n14451 ^ n13489;
  assign n14453 = n14446 & ~n14452;
  assign n14454 = ~n13275 & n14453;
  assign n14455 = n14454 ^ n11495;
  assign n14456 = n14455 ^ x498;
  assign n11656 = n11249 & n11655;
  assign n11648 = ~n11251 & n11641;
  assign n11657 = n11656 ^ n11648;
  assign n11665 = n11664 ^ n11639;
  assign n11666 = n11248 & ~n11665;
  assign n11667 = n11666 ^ n11639;
  assign n11668 = ~n11207 & n11667;
  assign n11673 = ~n11251 & n11672;
  assign n11675 = n11674 ^ n11670;
  assign n11676 = n11250 & ~n11675;
  assign n11681 = n11650 ^ n11639;
  assign n11680 = n11679 ^ n11660;
  assign n11682 = n11681 ^ n11680;
  assign n11683 = n11682 ^ n11632;
  assign n11684 = n11252 & ~n11683;
  assign n11702 = n11680 ^ n11645;
  assign n11703 = n11207 & n11702;
  assign n11693 = n11692 ^ n11649;
  assign n11694 = n11693 ^ n11688;
  assign n11685 = n11679 ^ n11655;
  assign n11686 = n11685 ^ n11650;
  assign n11695 = n11694 ^ n11686;
  assign n11696 = n11694 ^ n11207;
  assign n11697 = n11248 & n11696;
  assign n11698 = n11697 ^ n11207;
  assign n11699 = ~n11695 & n11698;
  assign n11700 = n11699 ^ n11686;
  assign n11701 = ~n11659 & ~n11700;
  assign n11704 = n11703 ^ n11701;
  assign n11705 = n11248 & ~n11704;
  assign n11706 = n11705 ^ n11701;
  assign n11707 = ~n11684 & n11706;
  assign n11708 = ~n11676 & n11707;
  assign n11709 = ~n11673 & n11708;
  assign n11710 = ~n11668 & n11709;
  assign n11711 = ~n11657 & n11710;
  assign n11712 = ~n11647 & n11711;
  assign n11713 = n11712 ^ n9933;
  assign n14457 = n11713 ^ x500;
  assign n12924 = n12923 ^ n12921;
  assign n12925 = ~n12916 & n12924;
  assign n12926 = n12925 ^ n12921;
  assign n12917 = n12903 & ~n12916;
  assign n12918 = n12917 ^ n12902;
  assign n12927 = n12926 ^ n12918;
  assign n12928 = ~n12915 & n12927;
  assign n12929 = n12928 ^ n12926;
  assign n12930 = n12914 & ~n12929;
  assign n12931 = n12930 ^ n10804;
  assign n14458 = n12931 ^ x497;
  assign n13497 = n12378 & ~n12425;
  assign n13509 = n12428 ^ n12387;
  assign n13510 = n13509 ^ n12397;
  assign n14461 = n12410 & ~n13510;
  assign n14462 = ~n12231 & n12399;
  assign n14467 = n12267 & n12382;
  assign n14463 = n12384 ^ n12366;
  assign n13503 = n12405 ^ n12367;
  assign n13504 = n13503 ^ n12368;
  assign n14464 = n14463 ^ n13504;
  assign n14465 = n12267 & n14464;
  assign n14466 = n14465 ^ n13504;
  assign n14468 = n14467 ^ n14466;
  assign n14469 = n12231 & n14468;
  assign n14470 = n14469 ^ n14466;
  assign n14471 = ~n12267 & ~n12395;
  assign n14472 = n14471 ^ n12388;
  assign n14473 = n12424 & ~n14472;
  assign n14474 = n14473 ^ n12388;
  assign n14475 = ~n14470 & n14474;
  assign n14476 = ~n14462 & n14475;
  assign n14477 = ~n14461 & n14476;
  assign n14478 = ~n13497 & n14477;
  assign n14479 = ~n12404 & n14478;
  assign n14480 = n14479 ^ n11536;
  assign n14481 = n14480 ^ x499;
  assign n14482 = n14458 & n14481;
  assign n14483 = n14457 & n14482;
  assign n14494 = ~n14456 & n14483;
  assign n14495 = n14494 ^ n14483;
  assign n14489 = n14456 & n14457;
  assign n14490 = ~n14458 & n14489;
  assign n14491 = n14490 ^ n14489;
  assign n11775 = n11774 ^ x491;
  assign n11785 = n11784 ^ n11436;
  assign n11786 = n11385 & n11785;
  assign n11787 = n11426 ^ n11407;
  assign n11788 = n11383 & ~n11787;
  assign n11789 = ~n11786 & ~n11788;
  assign n11790 = n11437 ^ n11391;
  assign n11791 = n11790 ^ n11400;
  assign n11792 = ~n11381 & n11791;
  assign n11793 = n11792 ^ n11400;
  assign n11794 = ~n11382 & n11793;
  assign n11795 = n11789 & ~n11794;
  assign n11796 = n11397 ^ n11386;
  assign n11797 = n11402 ^ n11384;
  assign n11798 = n11386 & n11797;
  assign n11799 = n11798 ^ n11384;
  assign n11800 = ~n11796 & n11799;
  assign n11801 = n11800 ^ n11397;
  assign n11802 = n11795 & n11801;
  assign n11803 = n11783 & n11802;
  assign n11804 = ~n11425 & n11803;
  assign n11805 = ~n11413 & n11804;
  assign n11806 = ~n11780 & n11805;
  assign n11807 = n11806 ^ n9249;
  assign n11808 = n11807 ^ x492;
  assign n11776 = n11127 ^ x494;
  assign n11809 = n11808 ^ n11776;
  assign n11716 = n11543 & n11600;
  assign n11722 = n11568 ^ n11551;
  assign n11723 = n11722 ^ n11560;
  assign n11724 = n11723 ^ n11612;
  assign n11725 = n11541 & ~n11724;
  assign n11726 = n11725 ^ n11612;
  assign n11717 = n11592 ^ n11576;
  assign n11718 = n11717 ^ n11578;
  assign n11719 = n11718 ^ n11599;
  assign n11720 = n11541 & ~n11719;
  assign n11721 = n11720 ^ n11599;
  assign n11727 = n11726 ^ n11721;
  assign n11728 = ~n11542 & n11727;
  assign n11729 = n11728 ^ n11721;
  assign n11730 = ~n11581 & ~n11729;
  assign n11731 = ~n11716 & n11730;
  assign n11732 = ~n11541 & n11558;
  assign n11733 = n11732 ^ n11560;
  assign n11734 = ~n11542 & n11733;
  assign n11735 = n11734 ^ n11560;
  assign n11736 = n11731 & ~n11735;
  assign n11738 = n11597 ^ n11594;
  assign n11739 = ~n11541 & ~n11738;
  assign n11740 = n11739 ^ n11594;
  assign n11741 = n11737 & ~n11740;
  assign n11742 = n11736 & ~n11741;
  assign n11743 = ~n11545 & n11742;
  assign n11744 = n11743 ^ n9280;
  assign n11745 = n11744 ^ x493;
  assign n11820 = n11808 ^ n11745;
  assign n11821 = n11809 & ~n11820;
  assign n11822 = ~n11775 & n11821;
  assign n11814 = ~n11775 & n11808;
  assign n11818 = n11814 ^ n11775;
  assign n11811 = ~n11776 & ~n11808;
  assign n11812 = ~n11775 & n11811;
  assign n11819 = n11818 ^ n11812;
  assign n11823 = n11822 ^ n11819;
  assign n11810 = ~n11775 & ~n11809;
  assign n11813 = n11812 ^ n11810;
  assign n11815 = n11814 ^ n11813;
  assign n11816 = n11745 & n11815;
  assign n11824 = n11823 ^ n11816;
  assign n11825 = n11824 ^ n11819;
  assign n11817 = n11816 ^ n11815;
  assign n11826 = n11825 ^ n11817;
  assign n11827 = n9778 ^ x495;
  assign n11872 = n11871 ^ x490;
  assign n11873 = n11827 & n11872;
  assign n11874 = n11873 ^ n11872;
  assign n11875 = n11874 ^ n11827;
  assign n11876 = n11826 & ~n11875;
  assign n11877 = ~n11745 & n11775;
  assign n11883 = n11808 & n11877;
  assign n11890 = n11883 ^ n11877;
  assign n11878 = n11811 ^ n11808;
  assign n11879 = n11877 & ~n11878;
  assign n11891 = n11890 ^ n11879;
  assign n11886 = n11810 ^ n11776;
  assign n11887 = n11886 ^ n11878;
  assign n11888 = n11887 ^ n11812;
  assign n11882 = n11814 ^ n11808;
  assign n11884 = n11883 ^ n11882;
  assign n11880 = n11879 ^ n11821;
  assign n11881 = n11880 ^ n11822;
  assign n11885 = n11884 ^ n11881;
  assign n11889 = n11888 ^ n11885;
  assign n11892 = n11891 ^ n11889;
  assign n11893 = ~n11872 & ~n11892;
  assign n11894 = n11893 ^ n11891;
  assign n11895 = ~n11827 & n11894;
  assign n11896 = n11873 ^ n11827;
  assign n11905 = ~n11745 & n11812;
  assign n11906 = n11905 ^ n11812;
  assign n11902 = n11877 ^ n11745;
  assign n11903 = n11902 ^ n11826;
  assign n11904 = n11903 ^ n11810;
  assign n11907 = n11906 ^ n11904;
  assign n11899 = n11891 ^ n11811;
  assign n11900 = n11899 ^ n11812;
  assign n11897 = n11889 ^ n11883;
  assign n11898 = n11897 ^ n11885;
  assign n11901 = n11900 ^ n11898;
  assign n11908 = n11907 ^ n11901;
  assign n11909 = n11896 & n11908;
  assign n11910 = ~n11895 & ~n11909;
  assign n11911 = n11907 ^ n11874;
  assign n11912 = n11875 ^ n11824;
  assign n11913 = n11907 & ~n11912;
  assign n11914 = n11913 ^ n11875;
  assign n11915 = ~n11911 & ~n11914;
  assign n11916 = n11915 ^ n11874;
  assign n11919 = n11882 ^ n11775;
  assign n11917 = n11900 ^ n11879;
  assign n11918 = n11917 ^ n11891;
  assign n11920 = n11919 ^ n11918;
  assign n11921 = n11920 ^ n11881;
  assign n11922 = n11921 ^ n11906;
  assign n11923 = n11827 & n11922;
  assign n11924 = n11923 ^ n11906;
  assign n11925 = n11872 & n11924;
  assign n11926 = n11872 ^ n11827;
  assign n11929 = n11889 ^ n11879;
  assign n11927 = n11907 ^ n11814;
  assign n11928 = n11927 ^ n11817;
  assign n11930 = n11929 ^ n11928;
  assign n11931 = n11872 & n11930;
  assign n11932 = n11931 ^ n11928;
  assign n11933 = n11926 & ~n11932;
  assign n11938 = ~n11872 & n11879;
  assign n11934 = n11883 ^ n11826;
  assign n11935 = n11934 ^ n11901;
  assign n11936 = n11872 & ~n11935;
  assign n11937 = n11936 ^ n11901;
  assign n11939 = n11938 ^ n11937;
  assign n11940 = n11939 ^ n11938;
  assign n11941 = n11824 & n11940;
  assign n11942 = n11941 ^ n11938;
  assign n11943 = ~n11926 & ~n11942;
  assign n11944 = n11943 ^ n11938;
  assign n11946 = n11874 & n11881;
  assign n11945 = n11875 & n11905;
  assign n11947 = n11946 ^ n11945;
  assign n11948 = ~n11944 & ~n11947;
  assign n11949 = ~n11933 & n11948;
  assign n11950 = ~n11925 & n11949;
  assign n11951 = ~n11916 & n11950;
  assign n11952 = n11910 & n11951;
  assign n11953 = ~n11876 & n11952;
  assign n11954 = n11953 ^ n10055;
  assign n14492 = n11954 ^ x501;
  assign n14493 = n14491 & ~n14492;
  assign n14496 = n14495 ^ n14493;
  assign n14497 = n14488 & n14496;
  assign n14498 = n14488 & n14492;
  assign n14484 = n14483 ^ n14482;
  assign n14499 = ~n14456 & n14484;
  assign n14500 = n14498 & n14499;
  assign n14485 = n14484 ^ n14457;
  assign n14459 = n14457 & ~n14458;
  assign n14460 = n14459 ^ n14458;
  assign n14486 = n14485 ^ n14460;
  assign n14487 = n14456 & n14486;
  assign n14507 = n14487 ^ n14486;
  assign n14541 = n14498 ^ n14488;
  assign n14776 = n14507 & n14541;
  assign n14505 = n14495 ^ n14491;
  assign n14758 = n14498 & n14505;
  assign n14520 = n14482 ^ n14481;
  assign n14517 = ~n14460 & ~n14481;
  assign n14518 = n14517 ^ n14460;
  assign n14521 = n14520 ^ n14518;
  assign n14523 = n14521 ^ n14490;
  assign n14522 = ~n14456 & ~n14521;
  assign n14524 = n14523 ^ n14522;
  assign n14542 = n14541 ^ n14492;
  assign n14544 = n14542 ^ n14488;
  assign n14545 = ~n14524 & n14544;
  assign n14759 = n14758 ^ n14545;
  assign n14509 = n14481 ^ n14456;
  assign n14510 = n14509 ^ n14457;
  assign n14501 = n14458 ^ n14457;
  assign n14502 = n14456 & ~n14501;
  assign n14511 = n14502 ^ n14458;
  assign n14512 = n14510 & n14511;
  assign n14513 = n14512 ^ n14458;
  assign n14514 = n14513 ^ n14483;
  assign n14504 = n14499 ^ n14484;
  assign n14506 = n14505 ^ n14504;
  assign n14508 = n14507 ^ n14506;
  assign n14515 = n14514 ^ n14508;
  assign n14503 = n14502 ^ n14491;
  assign n14516 = n14515 ^ n14503;
  assign n14760 = n14522 ^ n14516;
  assign n14761 = n14760 ^ n14495;
  assign n14762 = n14488 & n14761;
  assign n14763 = n14762 ^ n14495;
  assign n14764 = ~n14492 & n14763;
  assign n14525 = n14524 ^ n14490;
  assign n14755 = n14525 ^ n14515;
  assign n14756 = n14498 & ~n14755;
  assign n14531 = n14492 ^ n14488;
  assign n15506 = n14492 & n14513;
  assign n14519 = n14518 ^ n14516;
  assign n14773 = n14519 ^ n14494;
  assign n14552 = n14521 ^ n14459;
  assign n14553 = n14552 ^ n14524;
  assign n15505 = n14773 ^ n14553;
  assign n15507 = n15506 ^ n15505;
  assign n15222 = ~n14498 & n14524;
  assign n15502 = n14516 & ~n15222;
  assign n14532 = n14517 ^ n14515;
  assign n15503 = n15502 ^ n14532;
  assign n15499 = n15222 ^ n14553;
  assign n15500 = ~n14542 & ~n15499;
  assign n15501 = n15500 ^ n14522;
  assign n15504 = n15503 ^ n15501;
  assign n15508 = n15507 ^ n15504;
  assign n15509 = n14531 & ~n15508;
  assign n15510 = n15509 ^ n15504;
  assign n15512 = n14487 & ~n14492;
  assign n14533 = n14481 ^ n14457;
  assign n14534 = n14457 ^ n14456;
  assign n14535 = n14533 & n14534;
  assign n14536 = n14458 & n14535;
  assign n15511 = n14536 & ~n14542;
  assign n15513 = n15512 ^ n15511;
  assign n15514 = ~n15510 & ~n15513;
  assign n15515 = ~n14756 & n15514;
  assign n15516 = ~n14764 & n15515;
  assign n15517 = ~n14759 & n15516;
  assign n15518 = ~n14776 & n15517;
  assign n15519 = ~n14500 & n15518;
  assign n15520 = ~n14497 & n15519;
  assign n15521 = n15520 ^ n11631;
  assign n15522 = n15521 ^ x577;
  assign n15523 = ~n15498 & n15522;
  assign n12691 = ~n11251 & n11662;
  assign n12693 = n11248 & n12692;
  assign n12695 = n11671 ^ n11661;
  assign n12694 = n11649 ^ n11642;
  assign n12696 = n12695 ^ n12694;
  assign n12697 = n11249 & ~n12696;
  assign n12698 = ~n12693 & ~n12697;
  assign n12706 = n11672 ^ n11659;
  assign n12708 = n12707 ^ n12706;
  assign n12705 = n11689 ^ n11650;
  assign n12709 = n12708 ^ n12705;
  assign n12701 = n11689 ^ n11660;
  assign n12699 = n11679 ^ n11669;
  assign n12700 = n12699 ^ n11692;
  assign n12702 = n12701 ^ n12700;
  assign n12703 = n11248 & ~n12702;
  assign n12704 = n12703 ^ n12700;
  assign n12710 = n12709 ^ n12704;
  assign n12711 = n12710 ^ n12704;
  assign n12712 = ~n11248 & ~n12711;
  assign n12713 = n12712 ^ n12704;
  assign n12714 = n11207 & ~n12713;
  assign n12715 = n12714 ^ n12704;
  assign n12716 = n12698 & n12715;
  assign n12717 = ~n12691 & n12716;
  assign n12718 = ~n11668 & n12717;
  assign n12719 = ~n11657 & n12718;
  assign n12720 = n12719 ^ n10918;
  assign n14198 = n12720 ^ x537;
  assign n12033 = n12032 ^ x465;
  assign n11999 = n11998 ^ x460;
  assign n12079 = n10635 & n10648;
  assign n12080 = n12079 ^ n10615;
  assign n12081 = n10680 & n12080;
  assign n12082 = n12081 ^ n10615;
  assign n12084 = n10622 & ~n10680;
  assign n12083 = n10701 ^ n10627;
  assign n12085 = n12084 ^ n12083;
  assign n12086 = ~n10693 & n12085;
  assign n12087 = n12086 ^ n12083;
  assign n12088 = ~n12082 & ~n12087;
  assign n12098 = n11753 ^ n10621;
  assign n12099 = n12098 ^ n10716;
  assign n12100 = n10680 & ~n12099;
  assign n12101 = n12100 ^ n10716;
  assign n12090 = n12089 ^ n11746;
  assign n12091 = n12090 ^ n10681;
  assign n12092 = n10645 ^ n10585;
  assign n12093 = n12092 ^ n12089;
  assign n12094 = n12093 ^ n10585;
  assign n12095 = n12091 & ~n12094;
  assign n12096 = n12095 ^ n10681;
  assign n12097 = ~n10623 & ~n12096;
  assign n12102 = n12101 ^ n12097;
  assign n12103 = ~n10693 & ~n12102;
  assign n12104 = n12103 ^ n12101;
  assign n12105 = n12088 & ~n12104;
  assign n12106 = ~n12078 & n12105;
  assign n12107 = ~n10684 & n12106;
  assign n12108 = n12107 ^ n8852;
  assign n12109 = n12108 ^ x463;
  assign n12141 = n12140 ^ x461;
  assign n12142 = ~n12109 & n12141;
  assign n12152 = n12142 ^ n12109;
  assign n12039 = n9772 ^ n9400;
  assign n12040 = ~n9571 & n12039;
  assign n12041 = n12040 ^ n9772;
  assign n12035 = n9773 ^ n9734;
  assign n12036 = n12035 ^ n11200;
  assign n12037 = n9571 & n12036;
  assign n12038 = n12037 ^ n9768;
  assign n12042 = n12041 ^ n12038;
  assign n12043 = ~n9729 & ~n12042;
  assign n12044 = n12043 ^ n12038;
  assign n12045 = n12044 ^ n8662;
  assign n12046 = n12045 ^ x462;
  assign n12066 = n12065 ^ x464;
  assign n12067 = n12046 & ~n12066;
  assign n12068 = n12067 ^ n12046;
  assign n12069 = n12068 ^ n12066;
  assign n12154 = n12069 ^ n12046;
  assign n12155 = ~n12152 & ~n12154;
  assign n12190 = n12155 ^ n12154;
  assign n12171 = n12155 ^ n12152;
  assign n12166 = n12141 ^ n12109;
  assign n12167 = n12166 ^ n12046;
  assign n12168 = n12167 ^ n12066;
  assign n12165 = n12068 & ~n12141;
  assign n12169 = n12168 ^ n12165;
  assign n12160 = n12066 ^ n12046;
  assign n12162 = n12142 & n12160;
  assign n12163 = n12162 ^ n12142;
  assign n12143 = n12142 ^ n12141;
  assign n12161 = n12143 & n12160;
  assign n12164 = n12163 ^ n12161;
  assign n12170 = n12169 ^ n12164;
  assign n12172 = n12171 ^ n12170;
  assign n12148 = n12066 & n12142;
  assign n12149 = n12148 ^ n12141;
  assign n12146 = n12067 & n12142;
  assign n12147 = n12146 ^ n12143;
  assign n12150 = n12149 ^ n12147;
  assign n12189 = n12172 ^ n12150;
  assign n12191 = n12190 ^ n12189;
  assign n12188 = n12161 ^ n12146;
  assign n12192 = n12191 ^ n12188;
  assign n12193 = n12192 ^ n12147;
  assign n12653 = n12193 ^ n12191;
  assign n12175 = n12143 ^ n12109;
  assign n12205 = n12069 & n12175;
  assign n12206 = n12205 ^ n12155;
  assign n12654 = n12653 ^ n12206;
  assign n12655 = n11999 & n12654;
  assign n12656 = n12655 ^ n12653;
  assign n12657 = n12033 & n12656;
  assign n12034 = n12033 ^ n11999;
  assign n12157 = n12067 & ~n12152;
  assign n12158 = n12157 ^ n12152;
  assign n12153 = n12069 & ~n12152;
  assign n12156 = n12155 ^ n12153;
  assign n12159 = n12158 ^ n12156;
  assign n12174 = n12165 ^ n12159;
  assign n13192 = n12174 ^ n12157;
  assign n13193 = ~n12034 & ~n13192;
  assign n13894 = ~n11999 & n12170;
  assign n13895 = n13894 ^ n12164;
  assign n13896 = n13895 ^ n12164;
  assign n12665 = n12174 ^ n12162;
  assign n13898 = n12665 ^ n12190;
  assign n13899 = n13898 ^ n12193;
  assign n13900 = n11999 & n13899;
  assign n12176 = n12067 & n12175;
  assign n13897 = n12176 ^ n12150;
  assign n13901 = n13900 ^ n13897;
  assign n13902 = n13901 ^ n12164;
  assign n13903 = n13902 ^ n12164;
  assign n13904 = ~n13896 & ~n13903;
  assign n13905 = n13904 ^ n12164;
  assign n13906 = n12034 & ~n13905;
  assign n13907 = n13906 ^ n12164;
  assign n13909 = ~n12033 & n12153;
  assign n12658 = ~n11999 & ~n12033;
  assign n13908 = ~n12159 & n12658;
  assign n13910 = n13909 ^ n13908;
  assign n13911 = ~n13907 & ~n13910;
  assign n13912 = ~n13193 & n13911;
  assign n13913 = ~n12657 & n13912;
  assign n13914 = n13913 ^ n10557;
  assign n14199 = n13914 ^ x532;
  assign n13496 = n12268 & ~n12426;
  assign n13498 = n13497 ^ n13496;
  assign n13800 = n12267 & n12371;
  assign n13508 = n12377 ^ n12369;
  assign n13806 = n13508 ^ n12403;
  assign n13801 = ~n12403 & n12431;
  assign n13802 = n12398 ^ n12387;
  assign n13803 = n13802 ^ n12362;
  assign n13804 = ~n12410 & ~n13803;
  assign n13805 = ~n13801 & ~n13804;
  assign n13807 = n13806 ^ n13805;
  assign n13808 = n13807 ^ n13805;
  assign n13809 = ~n12267 & n13808;
  assign n13810 = n13809 ^ n13805;
  assign n13811 = n12231 & n13810;
  assign n13812 = n13811 ^ n13805;
  assign n13813 = ~n13800 & ~n13812;
  assign n13814 = n12365 ^ n12269;
  assign n13499 = n12398 ^ n12383;
  assign n13815 = n13499 ^ n12425;
  assign n13816 = ~n12365 & ~n13815;
  assign n13817 = n13816 ^ n12425;
  assign n13818 = n13814 & ~n13817;
  assign n13819 = n13818 ^ n12269;
  assign n13820 = n13813 & ~n13819;
  assign n13821 = ~n13498 & n13820;
  assign n13822 = ~n12409 & n13821;
  assign n13823 = ~n12404 & n13822;
  assign n13824 = n13823 ^ n10679;
  assign n14200 = n13824 ^ x533;
  assign n13006 = n13003 & n13005;
  assign n13011 = n13010 ^ n13008;
  assign n13012 = n13007 & n13011;
  assign n13028 = n13027 ^ n13019;
  assign n13029 = ~n13013 & n13028;
  assign n13041 = n13040 ^ n12997;
  assign n13030 = n13014 ^ n12994;
  assign n13031 = n13030 ^ n13022;
  assign n13042 = n13041 ^ n13031;
  assign n13043 = ~n12934 & ~n13042;
  assign n13044 = n13043 ^ n13031;
  assign n13045 = ~n12933 & n13044;
  assign n13046 = ~n13029 & ~n13045;
  assign n13047 = n13036 ^ n13032;
  assign n13048 = n13047 ^ n12933;
  assign n13049 = n13003 ^ n12996;
  assign n13050 = n13049 ^ n13039;
  assign n13051 = ~n12934 & ~n13050;
  assign n13052 = n13051 ^ n13039;
  assign n13053 = n13052 ^ n13047;
  assign n13054 = ~n13048 & ~n13053;
  assign n13055 = n13054 ^ n13051;
  assign n13056 = n13055 ^ n13039;
  assign n13057 = n13056 ^ n12933;
  assign n13058 = ~n13047 & n13057;
  assign n13059 = n13058 ^ n13047;
  assign n13060 = n13059 ^ n12933;
  assign n13061 = n13046 & n13060;
  assign n13062 = ~n13012 & n13061;
  assign n13063 = ~n13006 & n13062;
  assign n13067 = n12933 & n13015;
  assign n13069 = n13068 ^ n13067;
  assign n13066 = n13065 ^ n13064;
  assign n13070 = n13069 ^ n13066;
  assign n13071 = n13063 & ~n13070;
  assign n13072 = ~n13002 & n13071;
  assign n13073 = n13072 ^ n10789;
  assign n14201 = n13073 ^ x536;
  assign n14202 = ~n14200 & ~n14201;
  assign n14203 = n14202 ^ n14200;
  assign n14204 = n14203 ^ n14201;
  assign n13260 = ~n12904 & n12916;
  assign n13261 = n13260 ^ n12892;
  assign n13258 = ~n12913 & ~n12916;
  assign n13259 = n13258 ^ n12880;
  assign n13262 = n13261 ^ n13259;
  assign n13263 = n12915 & n13262;
  assign n14206 = n13263 ^ n13259;
  assign n14207 = n14206 ^ n11045;
  assign n14208 = n14207 ^ x534;
  assign n13159 = n11873 & ~n11903;
  assign n14209 = n11826 & n11874;
  assign n14210 = n11921 ^ n11898;
  assign n14211 = n11896 & ~n14210;
  assign n13160 = n11874 & n11900;
  assign n14216 = n11918 ^ n11888;
  assign n14217 = ~n11872 & ~n14216;
  assign n14218 = n14217 ^ n11888;
  assign n14213 = n11887 ^ n11820;
  assign n14214 = ~n11872 & ~n14213;
  assign n14212 = n11920 ^ n11901;
  assign n14215 = n14214 ^ n14212;
  assign n14219 = n14218 ^ n14215;
  assign n14220 = n11827 & n14219;
  assign n14221 = n14220 ^ n14218;
  assign n14222 = ~n11895 & n14221;
  assign n14223 = ~n13160 & n14222;
  assign n14224 = ~n14211 & n14223;
  assign n14225 = ~n14209 & n14224;
  assign n14227 = ~n11875 & n11906;
  assign n14226 = n11822 & ~n11926;
  assign n14228 = n14227 ^ n14226;
  assign n14229 = n14225 & ~n14228;
  assign n14230 = ~n11916 & n14229;
  assign n14231 = ~n13159 & n14230;
  assign n14232 = n14231 ^ n11036;
  assign n14233 = n14232 ^ x535;
  assign n14234 = n14208 & n14233;
  assign n14235 = n14234 ^ n14208;
  assign n14242 = ~n14204 & n14235;
  assign n14205 = n14204 ^ n14200;
  assign n14236 = n14235 ^ n14233;
  assign n14241 = ~n14205 & ~n14236;
  assign n14243 = n14242 ^ n14241;
  assign n14239 = ~n14204 & ~n14236;
  assign n14237 = n14236 ^ n14208;
  assign n14238 = ~n14205 & n14237;
  assign n14240 = n14239 ^ n14238;
  assign n14244 = n14243 ^ n14240;
  assign n14245 = ~n14199 & n14244;
  assign n14246 = n14245 ^ n14240;
  assign n14247 = n14198 & n14246;
  assign n14274 = ~n14203 & n14235;
  assign n14270 = n14202 & n14237;
  assign n14280 = n14274 ^ n14270;
  assign n14912 = n14198 & n14280;
  assign n14276 = ~n14205 & n14235;
  assign n14293 = n14276 ^ n14239;
  assign n14255 = ~n14203 & n14237;
  assign n14294 = n14293 ^ n14255;
  assign n14910 = ~n14198 & n14294;
  assign n14911 = n14910 ^ n14255;
  assign n14913 = n14912 ^ n14911;
  assign n14914 = n14199 & n14913;
  assign n14915 = n14914 ^ n14911;
  assign n14248 = n14198 & ~n14199;
  assign n14259 = ~n14203 & n14234;
  assign n14258 = n14202 & n14234;
  assign n14260 = n14259 ^ n14258;
  assign n15464 = n14276 ^ n14260;
  assign n15465 = n14248 & n15464;
  assign n14253 = n14199 ^ n14198;
  assign n14249 = n14248 ^ n14198;
  assign n14250 = n14249 ^ n14199;
  assign n15466 = n14204 & ~n14250;
  assign n14254 = n14202 & ~n14236;
  assign n14256 = n14255 ^ n14254;
  assign n14275 = n14274 ^ n14256;
  assign n14277 = n14276 ^ n14275;
  assign n14271 = n14270 ^ n14239;
  assign n14272 = n14271 ^ n14242;
  assign n14262 = ~n14204 & n14234;
  assign n14261 = n14260 ^ n14234;
  assign n14263 = n14262 ^ n14261;
  assign n14273 = n14272 ^ n14263;
  assign n14278 = n14277 ^ n14273;
  assign n14267 = n14208 ^ n14201;
  assign n14268 = n14267 ^ n14200;
  assign n14265 = n14259 ^ n14254;
  assign n14257 = n14256 ^ n14242;
  assign n14264 = n14263 ^ n14257;
  assign n14266 = n14265 ^ n14264;
  assign n14269 = n14268 ^ n14266;
  assign n14279 = n14278 ^ n14269;
  assign n15469 = n14279 ^ n14242;
  assign n15467 = n14239 & n14248;
  assign n15468 = n15467 ^ n14276;
  assign n15470 = n15469 ^ n15468;
  assign n15471 = ~n15466 & ~n15470;
  assign n15472 = n14253 & n15471;
  assign n15473 = ~n15465 & ~n15472;
  assign n14593 = n14262 ^ n14241;
  assign n14288 = n14202 & n14235;
  assign n15475 = n14593 ^ n14288;
  assign n14289 = n14254 ^ n14236;
  assign n14251 = n14241 ^ n14239;
  assign n14290 = n14289 ^ n14251;
  assign n14917 = n14290 ^ n14258;
  assign n15474 = n14917 ^ n14270;
  assign n15476 = n15475 ^ n15474;
  assign n15477 = n14198 & ~n15476;
  assign n15478 = n15477 ^ n15474;
  assign n15479 = n14199 & ~n15478;
  assign n15480 = n15473 & ~n15479;
  assign n15481 = n14270 ^ n14258;
  assign n15482 = n15481 ^ n14243;
  assign n15483 = n15482 ^ n14267;
  assign n15484 = n15483 ^ n14255;
  assign n15485 = n15484 ^ n14255;
  assign n15486 = ~n14198 & ~n15485;
  assign n15487 = n15486 ^ n14255;
  assign n15488 = ~n14199 & n15487;
  assign n15489 = n15488 ^ n14255;
  assign n15490 = n15480 & ~n15489;
  assign n15491 = ~n14915 & n15490;
  assign n15492 = ~n14247 & n15491;
  assign n15493 = n15492 ^ n11337;
  assign n15494 = n15493 ^ x576;
  assign n12725 = n10753 & n11128;
  assign n12726 = n11157 ^ n10754;
  assign n12727 = ~n11152 & n12726;
  assign n12728 = n10762 ^ n10756;
  assign n12729 = n12728 ^ n11151;
  assign n12730 = n11009 & ~n12729;
  assign n12731 = n12730 ^ n11151;
  assign n12732 = n11152 & n12731;
  assign n12733 = ~n11128 & n11134;
  assign n12734 = n12733 ^ n11133;
  assign n12735 = n11009 & n12734;
  assign n12742 = n11166 ^ n11145;
  assign n12741 = n11151 ^ n11143;
  assign n12743 = n12742 ^ n12741;
  assign n12744 = n12742 ^ n11009;
  assign n12745 = n11152 & ~n12744;
  assign n12746 = n12745 ^ n11009;
  assign n12747 = ~n12743 & ~n12746;
  assign n12748 = n12747 ^ n12741;
  assign n12749 = ~n11181 & ~n12748;
  assign n12736 = n12728 ^ n11164;
  assign n12737 = n12736 ^ n11162;
  assign n12738 = n12737 ^ n10759;
  assign n12739 = ~n11009 & n12738;
  assign n12740 = n12739 ^ n10759;
  assign n12750 = n12749 ^ n12740;
  assign n12751 = n11152 & n12750;
  assign n12752 = n12751 ^ n12749;
  assign n12753 = ~n12735 & n12752;
  assign n12754 = ~n12732 & n12753;
  assign n12755 = ~n12727 & n12754;
  assign n12756 = ~n12725 & n12755;
  assign n12757 = n11181 ^ n11141;
  assign n12758 = n12757 ^ n11137;
  assign n12759 = ~n11128 & n12758;
  assign n12760 = n12759 ^ n11137;
  assign n12761 = n11009 & n12760;
  assign n12762 = n12756 & ~n12761;
  assign n12763 = n11153 ^ n11009;
  assign n12764 = ~n10760 & ~n12763;
  assign n12765 = n12764 ^ n11155;
  assign n12766 = n12762 & ~n12765;
  assign n12767 = n12766 ^ n10881;
  assign n12768 = n12767 ^ x541;
  assign n12659 = n12658 ^ n12033;
  assign n12660 = n12206 ^ n12157;
  assign n12661 = ~n12659 & n12660;
  assign n12662 = n12153 ^ n12150;
  assign n12663 = n12662 ^ n12174;
  assign n12664 = n12658 & ~n12663;
  assign n12672 = n12193 ^ n12163;
  assign n12673 = n12672 ^ n12176;
  assign n12671 = n12653 ^ n12148;
  assign n12674 = n12673 ^ n12671;
  assign n12675 = n11999 & n12674;
  assign n12676 = n12675 ^ n12671;
  assign n12173 = n12172 ^ n12159;
  assign n12667 = n12206 ^ n12173;
  assign n12144 = n12069 & n12143;
  assign n12666 = n12665 ^ n12144;
  assign n12668 = n12667 ^ n12666;
  assign n12669 = ~n11999 & ~n12668;
  assign n12670 = n12669 ^ n12666;
  assign n12677 = n12676 ^ n12670;
  assign n12678 = n12034 & ~n12677;
  assign n12679 = n12678 ^ n12676;
  assign n12680 = ~n12664 & ~n12679;
  assign n12681 = ~n12661 & n12680;
  assign n12682 = n12173 ^ n12162;
  assign n12683 = ~n11999 & n12682;
  assign n12684 = n12683 ^ n12173;
  assign n12685 = n12033 & n12684;
  assign n12686 = n12681 & ~n12685;
  assign n12687 = ~n12657 & n12686;
  assign n12688 = n12172 & n12687;
  assign n12689 = n12688 ^ n10860;
  assign n12690 = n12689 ^ x540;
  assign n12721 = n12720 ^ x539;
  assign n12722 = ~n12690 & n12721;
  assign n12723 = n12722 ^ n12690;
  assign n12808 = n12807 ^ x542;
  assign n12812 = ~n12723 & ~n12808;
  assign n12813 = ~n12768 & n12812;
  assign n12814 = n12813 ^ n12812;
  assign n12809 = n12768 & ~n12808;
  assign n12810 = n12721 & n12809;
  assign n12811 = n12810 ^ n12809;
  assign n12815 = n12814 ^ n12811;
  assign n12769 = n12690 & ~n12768;
  assign n12770 = n12721 & n12769;
  assign n12771 = n12770 ^ n12769;
  assign n12724 = n12723 ^ n12721;
  assign n12772 = n12771 ^ n12724;
  assign n12816 = n12815 ^ n12772;
  assign n12817 = n12816 ^ n12814;
  assign n12932 = n12931 ^ x543;
  assign n13074 = n13073 ^ x538;
  assign n13075 = n13074 ^ n12932;
  assign n13076 = ~n12932 & ~n13075;
  assign n13077 = n13076 ^ n12932;
  assign n13078 = n13077 ^ n13074;
  assign n13079 = n12817 & ~n13078;
  assign n13086 = n12690 & n12810;
  assign n13080 = n12721 & n12808;
  assign n13081 = n12769 & n13080;
  assign n13096 = n13086 ^ n13081;
  assign n13087 = n13086 ^ n12810;
  assign n13097 = n13096 ^ n13087;
  assign n13098 = ~n13074 & n13097;
  assign n13099 = n13098 ^ n13087;
  assign n13100 = n13075 & n13099;
  assign n13105 = n12771 & n12808;
  assign n13083 = n12722 & ~n12808;
  assign n13101 = n13087 ^ n13083;
  assign n14307 = n13105 ^ n13101;
  assign n13090 = n12812 ^ n12723;
  assign n13091 = ~n12768 & ~n13090;
  assign n13131 = n13091 ^ n13090;
  assign n14305 = n13131 ^ n12815;
  assign n14306 = n14305 ^ n13091;
  assign n14308 = n14307 ^ n14306;
  assign n14309 = n12932 & ~n14308;
  assign n14310 = n14309 ^ n14306;
  assign n14311 = ~n13074 & ~n14310;
  assign n14312 = ~n13100 & ~n14311;
  assign n13084 = n13083 ^ n12722;
  assign n13082 = n13081 ^ n13080;
  assign n13085 = n13084 ^ n13082;
  assign n13088 = n13087 ^ n13085;
  assign n13089 = n13088 ^ n12813;
  assign n13092 = n13091 ^ n13089;
  assign n13093 = ~n12932 & n13092;
  assign n13094 = n13093 ^ n13091;
  assign n13095 = ~n13074 & n13094;
  assign n13106 = n13105 ^ n12771;
  assign n13107 = n12932 & n13106;
  assign n13102 = n13101 ^ n12815;
  assign n13103 = ~n12932 & n13102;
  assign n13104 = n13103 ^ n12815;
  assign n13108 = n13107 ^ n13104;
  assign n13109 = ~n13075 & n13108;
  assign n13110 = n13109 ^ n13104;
  assign n15130 = ~n13074 & n13088;
  assign n13127 = n13081 ^ n12770;
  assign n13111 = ~n12768 & n13084;
  assign n13128 = n13127 ^ n13111;
  assign n15131 = n15130 ^ n13128;
  assign n15132 = n13075 & n15131;
  assign n15133 = n15132 ^ n13128;
  assign n15134 = n13081 ^ n12932;
  assign n15135 = ~n13077 & ~n15134;
  assign n15136 = n15135 ^ n13076;
  assign n15137 = n15136 ^ n12932;
  assign n15138 = n15137 ^ n13074;
  assign n13133 = n13111 ^ n13084;
  assign n15141 = n13133 ^ n12813;
  assign n15139 = n12724 & ~n13077;
  assign n13143 = n12815 & n13074;
  assign n15140 = n15139 ^ n13143;
  assign n15142 = n15141 ^ n15140;
  assign n15143 = ~n15138 & ~n15142;
  assign n15144 = n15143 ^ n13074;
  assign n15145 = ~n15133 & ~n15144;
  assign n15146 = ~n13110 & n15145;
  assign n15147 = ~n13095 & n15146;
  assign n15148 = n14312 & n15147;
  assign n15149 = ~n13079 & n15148;
  assign n15150 = n15149 ^ n11287;
  assign n15495 = n15150 ^ x575;
  assign n15496 = ~n15494 & ~n15495;
  assign n15526 = n15496 ^ n15495;
  assign n15527 = n15526 ^ n15494;
  assign n15528 = n15523 & ~n15527;
  assign n15497 = n15496 ^ n15494;
  assign n15524 = n15523 ^ n15522;
  assign n15525 = ~n15497 & n15524;
  assign n15529 = n15528 ^ n15525;
  assign n13219 = n11161 ^ n11136;
  assign n13220 = n11009 & n13219;
  assign n13221 = n13220 ^ n11161;
  assign n13222 = ~n11152 & n13221;
  assign n13223 = n11138 ^ n10762;
  assign n13224 = n13223 ^ n11159;
  assign n13225 = ~n11154 & ~n11157;
  assign n13226 = n13225 ^ n12763;
  assign n13227 = n11159 & ~n13226;
  assign n13228 = n13227 ^ n12763;
  assign n13229 = n13224 & n13228;
  assign n13230 = n13229 ^ n13223;
  assign n13231 = ~n11128 & n13230;
  assign n13237 = n10743 & n11128;
  assign n13235 = n10759 ^ n10755;
  assign n13236 = n11153 & ~n13235;
  assign n13238 = n13237 ^ n13236;
  assign n13232 = n11153 ^ n11128;
  assign n13233 = n11138 ^ n10753;
  assign n13234 = n13232 & ~n13233;
  assign n13239 = n13238 ^ n13234;
  assign n13240 = ~n13231 & ~n13239;
  assign n13241 = n11181 ^ n11151;
  assign n13242 = n11154 & n13241;
  assign n13243 = n13242 ^ n11181;
  assign n13244 = n13240 & ~n13243;
  assign n13245 = ~n13222 & n13244;
  assign n13246 = n10754 & n11009;
  assign n13247 = n13246 ^ n11145;
  assign n13248 = ~n11128 & ~n13247;
  assign n13249 = n13248 ^ n11145;
  assign n13250 = n13245 & n13249;
  assign n13251 = n11151 & ~n12763;
  assign n13252 = n13251 ^ n12735;
  assign n13253 = n13250 & ~n13252;
  assign n13254 = ~n12732 & n13253;
  assign n13255 = ~n11149 & n13254;
  assign n13256 = n13255 ^ n9728;
  assign n13613 = n13256 ^ x519;
  assign n13463 = n13462 ^ x514;
  assign n13533 = n11826 & n11896;
  assign n13534 = n11920 ^ n11900;
  assign n13535 = ~n11875 & n13534;
  assign n13163 = n11874 & ~n11907;
  assign n13536 = n11891 ^ n11885;
  assign n13537 = ~n11926 & n13536;
  assign n13538 = n11906 ^ n11824;
  assign n13539 = n11873 & ~n13538;
  assign n13540 = ~n13537 & ~n13539;
  assign n13546 = ~n11872 & ~n11928;
  assign n13542 = n13534 ^ n11888;
  assign n13541 = n11905 ^ n11822;
  assign n13543 = n13542 ^ n13541;
  assign n13544 = ~n11872 & ~n13543;
  assign n13545 = n13544 ^ n13541;
  assign n13547 = n13546 ^ n13545;
  assign n13548 = ~n11926 & n13547;
  assign n13549 = n13548 ^ n13545;
  assign n13550 = n13540 & ~n13549;
  assign n13551 = ~n13159 & n13550;
  assign n13552 = ~n11876 & n13551;
  assign n13553 = ~n13163 & n13552;
  assign n13554 = ~n13535 & n13553;
  assign n13555 = ~n13533 & n13554;
  assign n13557 = n11872 & ~n11897;
  assign n13556 = n11873 & n11881;
  assign n13558 = n13557 ^ n13556;
  assign n13559 = n13555 & ~n13558;
  assign n13560 = ~n11933 & n13559;
  assign n13561 = ~n13160 & n13560;
  assign n13562 = n13561 ^ n9397;
  assign n13563 = n13562 ^ x517;
  assign n13495 = n13494 ^ x515;
  assign n13596 = n13563 ^ n13495;
  assign n13191 = n12176 & n12658;
  assign n12186 = n12173 ^ n12156;
  assign n13194 = n12186 & ~n12659;
  assign n13195 = n12205 & n12658;
  assign n13200 = n12191 ^ n12144;
  assign n13201 = n13200 ^ n12148;
  assign n13202 = n13201 ^ n12671;
  assign n13203 = ~n11999 & n13202;
  assign n13204 = n13203 ^ n12671;
  assign n12204 = n12176 ^ n12159;
  assign n13196 = n12204 ^ n12156;
  assign n12194 = n12193 ^ n12188;
  assign n13197 = n13196 ^ n12194;
  assign n13198 = ~n11999 & ~n13197;
  assign n13199 = n13198 ^ n12194;
  assign n13205 = n13204 ^ n13199;
  assign n13206 = n12034 & n13205;
  assign n13207 = n13206 ^ n13204;
  assign n13208 = ~n13195 & ~n13207;
  assign n13209 = ~n13194 & n13208;
  assign n13210 = n12192 ^ n12189;
  assign n13211 = ~n11999 & ~n13210;
  assign n13212 = n13211 ^ n12189;
  assign n13213 = n12033 & ~n13212;
  assign n13214 = n13209 & ~n13213;
  assign n13215 = ~n13193 & n13214;
  assign n13216 = ~n13191 & n13215;
  assign n13217 = n13216 ^ n8934;
  assign n13464 = n13217 ^ x518;
  assign n13576 = n13563 ^ n13464;
  assign n13599 = n13596 ^ n13576;
  assign n13500 = n13499 ^ n12403;
  assign n13501 = ~n12425 & ~n13500;
  assign n13511 = n13510 ^ n13508;
  assign n13502 = n12376 ^ n12370;
  assign n13505 = n13504 ^ n13502;
  assign n13506 = ~n12267 & n13505;
  assign n13507 = n13506 ^ n13504;
  assign n13512 = n13511 ^ n13507;
  assign n13513 = n13512 ^ n13507;
  assign n13514 = n12267 & ~n13513;
  assign n13515 = n13514 ^ n13507;
  assign n13516 = n12231 & n13515;
  assign n13517 = n13516 ^ n13507;
  assign n13518 = ~n13501 & ~n13517;
  assign n13521 = n12429 ^ n12412;
  assign n13519 = n12429 ^ n12399;
  assign n13520 = n13519 ^ n12362;
  assign n13522 = n13521 ^ n13520;
  assign n13523 = ~n12267 & n13522;
  assign n13524 = n13523 ^ n13520;
  assign n13525 = n12424 & ~n13524;
  assign n13526 = n13518 & ~n13525;
  assign n13527 = ~n13498 & n13526;
  assign n13528 = ~n12404 & n13527;
  assign n13529 = n13528 ^ n8449;
  assign n13530 = n13529 ^ x516;
  assign n13600 = n13576 ^ n13530;
  assign n13601 = ~n13464 & ~n13600;
  assign n13602 = n13601 ^ n13563;
  assign n13603 = ~n13599 & ~n13602;
  assign n13604 = n13603 ^ n13600;
  assign n13585 = n13530 ^ n13464;
  assign n13586 = n13585 ^ n13495;
  assign n13587 = n13530 & n13586;
  assign n13588 = n13587 ^ n13495;
  assign n13589 = ~n13563 & n13588;
  assign n13590 = n13589 ^ n13586;
  assign n13605 = n13604 ^ n13590;
  assign n13531 = ~n13495 & ~n13530;
  assign n13532 = n13531 ^ n13495;
  assign n13572 = n13464 & ~n13532;
  assign n13573 = n13572 ^ n13531;
  assign n13574 = ~n13563 & n13573;
  assign n13575 = n13574 ^ n13531;
  assign n13598 = n13575 ^ n13572;
  assign n13606 = n13605 ^ n13598;
  assign n13578 = n13531 ^ n13530;
  assign n13577 = ~n13532 & ~n13563;
  assign n13579 = n13578 ^ n13577;
  assign n13580 = ~n13576 & n13579;
  assign n13581 = ~n13575 & ~n13580;
  assign n13623 = n13606 ^ n13581;
  assign n13582 = n13572 ^ n13464;
  assign n13565 = n13495 & n13563;
  assign n13566 = n13565 ^ n13495;
  assign n13564 = n13563 ^ n13532;
  assign n13567 = n13566 ^ n13564;
  assign n13568 = n13567 ^ n13563;
  assign n13583 = n13582 ^ n13568;
  assign n13584 = ~n13575 & ~n13583;
  assign n13591 = n13590 ^ n13584;
  assign n13592 = n13581 & ~n13591;
  assign n13593 = n13592 ^ n13577;
  assign n13594 = n13593 ^ n13563;
  assign n13595 = n13594 ^ n13464;
  assign n13597 = n13596 ^ n13595;
  assign n13617 = n13597 ^ n13584;
  assign n13618 = n13617 ^ n13572;
  assign n13607 = n13606 ^ n13597;
  assign n13608 = n13607 ^ n13568;
  assign n13609 = n13608 ^ n13596;
  assign n13569 = n13568 ^ n13564;
  assign n13570 = ~n13464 & n13569;
  assign n13571 = n13570 ^ n13568;
  assign n13610 = n13609 ^ n13571;
  assign n13619 = n13618 ^ n13610;
  assign n13615 = n13565 & n13576;
  assign n13616 = n13615 ^ n13576;
  assign n13620 = n13619 ^ n13616;
  assign n13621 = n13606 ^ n13578;
  assign n13622 = n13620 & n13621;
  assign n13624 = n13623 ^ n13622;
  assign n13625 = n13463 & n13624;
  assign n13626 = n13625 ^ n13622;
  assign n13611 = ~n13463 & ~n13610;
  assign n13612 = n13611 ^ n13571;
  assign n13627 = n13626 ^ n13612;
  assign n13628 = ~n13613 & n13627;
  assign n15155 = n13628 ^ n13626;
  assign n15156 = n15155 ^ n11206;
  assign n15530 = n15156 ^ x574;
  assign n13161 = n11906 & ~n11926;
  assign n13162 = n11817 & n11827;
  assign n13164 = n11885 ^ n11879;
  assign n13165 = n13164 ^ n11928;
  assign n13166 = n11874 & ~n13165;
  assign n13168 = n11879 ^ n11816;
  assign n13167 = n11891 ^ n11824;
  assign n13169 = n13168 ^ n13167;
  assign n13170 = n13169 ^ n13167;
  assign n13171 = n11827 & n13170;
  assign n13172 = n13171 ^ n13167;
  assign n13173 = n11872 & ~n13172;
  assign n13174 = n13173 ^ n13167;
  assign n13175 = ~n13166 & n13174;
  assign n13176 = ~n11925 & n13175;
  assign n13177 = ~n13163 & n13176;
  assign n13178 = ~n13162 & n13177;
  assign n13179 = ~n13161 & n13178;
  assign n13180 = n11921 ^ n11889;
  assign n13181 = ~n11827 & ~n13180;
  assign n13182 = n13181 ^ n11889;
  assign n13183 = ~n11872 & ~n13182;
  assign n13184 = n13179 & ~n13183;
  assign n13185 = n11910 & n13184;
  assign n13186 = ~n13160 & n13185;
  assign n13187 = ~n13159 & n13186;
  assign n13188 = ~n11876 & n13187;
  assign n13189 = n13188 ^ n10250;
  assign n13190 = n13189 ^ x525;
  assign n13218 = n13217 ^ x520;
  assign n13257 = n13256 ^ x521;
  assign n13308 = n11252 ^ n11250;
  assign n13309 = n11689 & n13308;
  assign n13313 = n11672 & n13308;
  assign n13311 = ~n11207 & n13310;
  assign n13312 = n13311 ^ n12692;
  assign n13314 = n13313 ^ n13312;
  assign n13315 = n13314 ^ n11251;
  assign n13317 = ~n11250 & ~n12706;
  assign n13318 = n13308 & ~n13317;
  assign n13316 = n11655 ^ n11652;
  assign n13319 = n13318 ^ n13316;
  assign n13320 = n13314 & ~n13319;
  assign n13321 = n13320 ^ n13316;
  assign n13322 = ~n13315 & ~n13321;
  assign n13323 = n13322 ^ n11251;
  assign n13324 = ~n13309 & n13323;
  assign n13326 = n12705 ^ n11664;
  assign n13327 = n13326 ^ n11639;
  assign n13328 = n13327 ^ n11692;
  assign n13329 = n11207 & n13328;
  assign n13330 = n13329 ^ n11692;
  assign n13325 = n11207 & n11639;
  assign n13331 = n13330 ^ n13325;
  assign n13332 = n13331 ^ n13325;
  assign n13333 = ~n11649 & n13332;
  assign n13334 = n13333 ^ n13325;
  assign n13335 = n11248 & ~n13334;
  assign n13336 = n13335 ^ n13325;
  assign n13337 = n13324 & ~n13336;
  assign n13338 = ~n12691 & n13337;
  assign n13339 = ~n11648 & n13338;
  assign n13340 = ~n13307 & n13339;
  assign n13341 = ~n11647 & n13340;
  assign n13342 = n13341 ^ n10447;
  assign n13343 = n13342 ^ x523;
  assign n13349 = ~n13257 & ~n13343;
  assign n13350 = n13349 ^ n13257;
  assign n13264 = n13263 ^ n12915;
  assign n13265 = n13264 ^ n13261;
  assign n13266 = n13265 ^ n10372;
  assign n13267 = n13266 ^ x524;
  assign n13276 = n13047 & ~n13269;
  assign n13277 = n13039 ^ n13035;
  assign n13278 = n13005 & ~n13277;
  assign n13284 = n13283 ^ n13010;
  assign n13285 = n13284 ^ n12997;
  assign n13286 = n13285 ^ n12955;
  assign n13287 = n12934 & n13286;
  assign n13281 = n13023 ^ n13014;
  assign n13282 = n13281 ^ n12993;
  assign n13288 = n13287 ^ n13282;
  assign n13279 = ~n12933 & n13025;
  assign n13280 = n13279 ^ n13024;
  assign n13289 = n13288 ^ n13280;
  assign n13290 = n13013 & n13289;
  assign n13291 = n13290 ^ n13280;
  assign n13292 = ~n13278 & ~n13291;
  assign n13293 = ~n13276 & n13292;
  assign n13295 = n13027 ^ n13016;
  assign n13294 = n13034 ^ n13032;
  assign n13296 = n13295 ^ n13294;
  assign n13297 = ~n12933 & ~n13296;
  assign n13298 = n13297 ^ n13294;
  assign n13299 = n13013 & ~n13298;
  assign n13300 = n13293 & ~n13299;
  assign n13301 = ~n13275 & n13300;
  assign n13302 = n13301 ^ n10401;
  assign n13303 = n13302 ^ x522;
  assign n13351 = ~n13267 & n13303;
  assign n13367 = ~n13350 & n13351;
  assign n13344 = n13343 ^ n13303;
  assign n13345 = n13267 & n13344;
  assign n13374 = n13367 ^ n13345;
  assign n13352 = n13351 ^ n13267;
  assign n13363 = n13352 ^ n13303;
  assign n13372 = ~n13350 & n13363;
  assign n13365 = n13363 ^ n13267;
  assign n13366 = n13349 & n13365;
  assign n13368 = n13367 ^ n13366;
  assign n13360 = n13349 ^ n13343;
  assign n13364 = ~n13360 & n13363;
  assign n13369 = n13368 ^ n13364;
  assign n13357 = n13303 ^ n13257;
  assign n13358 = n13303 ^ n13267;
  assign n13359 = n13358 ^ n13343;
  assign n13361 = n13360 ^ n13359;
  assign n13362 = n13357 & n13361;
  assign n13370 = n13369 ^ n13362;
  assign n13371 = n13370 ^ n13368;
  assign n13373 = n13372 ^ n13371;
  assign n13375 = n13374 ^ n13373;
  assign n13353 = ~n13350 & ~n13352;
  assign n13354 = n13353 ^ n13350;
  assign n13346 = n13345 ^ n13303;
  assign n13355 = n13354 ^ n13346;
  assign n13347 = n13257 & ~n13346;
  assign n13348 = n13347 ^ n13257;
  assign n13356 = n13355 ^ n13348;
  assign n13376 = n13375 ^ n13356;
  assign n13377 = n13218 & ~n13376;
  assign n13378 = n13377 ^ n13375;
  assign n13379 = n13190 & n13378;
  assign n13380 = n13356 ^ n13353;
  assign n13381 = n13190 & ~n13380;
  assign n13382 = n13381 ^ n13356;
  assign n13383 = ~n13218 & ~n13382;
  assign n13384 = n13218 ^ n13190;
  assign n13387 = n13190 & n13366;
  assign n13385 = n13382 ^ n13353;
  assign n13386 = n13385 ^ n13356;
  assign n13388 = n13387 ^ n13386;
  assign n13389 = ~n13384 & n13388;
  assign n13390 = n13389 ^ n13386;
  assign n13391 = ~n13190 & ~n13218;
  assign n13392 = n13372 ^ n13367;
  assign n13393 = n13391 & n13392;
  assign n13394 = n13391 ^ n13384;
  assign n13403 = n13365 ^ n13343;
  assign n13404 = n13257 & n13403;
  assign n13400 = n13366 ^ n13349;
  assign n13397 = n13372 ^ n13370;
  assign n13396 = n13364 ^ n13363;
  assign n13398 = n13397 ^ n13396;
  assign n13399 = n13398 ^ n13356;
  assign n13401 = n13400 ^ n13399;
  assign n13395 = n13392 ^ n13354;
  assign n13402 = n13401 ^ n13395;
  assign n13405 = n13404 ^ n13402;
  assign n13406 = ~n13394 & n13405;
  assign n13407 = n13398 ^ n13218;
  assign n13416 = n13401 ^ n13352;
  assign n13408 = n13360 ^ n13257;
  assign n13410 = n13408 ^ n13375;
  assign n13411 = n13410 ^ n13404;
  assign n13409 = n13351 & ~n13408;
  assign n13412 = n13411 ^ n13409;
  assign n13413 = n13412 ^ n13370;
  assign n13414 = n13413 ^ n13408;
  assign n13415 = n13414 ^ n13353;
  assign n13417 = n13416 ^ n13415;
  assign n13418 = n13417 ^ n13409;
  assign n13419 = n13418 ^ n13364;
  assign n13420 = n13419 ^ n13347;
  assign n13421 = ~n13190 & n13420;
  assign n13422 = n13421 ^ n13419;
  assign n13423 = n13422 ^ n13398;
  assign n13424 = n13407 & n13423;
  assign n13425 = n13424 ^ n13421;
  assign n13426 = n13425 ^ n13419;
  assign n13427 = n13426 ^ n13218;
  assign n13428 = ~n13398 & n13427;
  assign n13429 = n13428 ^ n13398;
  assign n13430 = n13429 ^ n13218;
  assign n13431 = ~n13406 & ~n13430;
  assign n13432 = ~n13393 & n13431;
  assign n13433 = n13401 ^ n13398;
  assign n13434 = n13433 ^ n13414;
  assign n13435 = n13434 ^ n13348;
  assign n13436 = n13435 ^ n13395;
  assign n13437 = ~n13190 & n13436;
  assign n13438 = n13437 ^ n13395;
  assign n13439 = n13384 & ~n13438;
  assign n13440 = n13432 & ~n13439;
  assign n13441 = ~n13390 & n13440;
  assign n13442 = ~n13383 & n13441;
  assign n13443 = ~n13379 & n13442;
  assign n13444 = n13443 ^ n11247;
  assign n15531 = n13444 ^ x579;
  assign n15532 = n15530 & ~n15531;
  assign n15533 = n15529 & n15532;
  assign n15562 = n15495 ^ n15494;
  assign n15563 = n15522 ^ n15498;
  assign n15564 = n15563 ^ n15495;
  assign n15565 = n15562 & ~n15564;
  assign n15534 = n15523 ^ n15498;
  assign n15561 = ~n15526 & ~n15534;
  assign n15566 = n15565 ^ n15561;
  assign n15576 = n15531 & n15566;
  assign n15548 = ~n15497 & n15523;
  assign n15546 = n15524 ^ n15498;
  assign n15547 = ~n15497 & n15546;
  assign n15549 = n15548 ^ n15547;
  assign n15567 = n15566 ^ n15549;
  assign n15577 = n15576 ^ n15567;
  assign n15578 = n15530 & n15577;
  assign n15542 = n15532 ^ n15531;
  assign n15543 = n15542 ^ n15530;
  assign n15544 = n15543 ^ n15532;
  assign n15584 = n15563 ^ n15496;
  assign n15570 = n15527 ^ n15524;
  assign n15538 = n15528 ^ n15527;
  assign n15536 = n15524 & ~n15527;
  assign n15535 = ~n15527 & ~n15534;
  assign n15537 = n15536 ^ n15535;
  assign n15539 = n15538 ^ n15537;
  assign n15568 = n15567 ^ n15539;
  assign n15560 = n15535 ^ n15529;
  assign n15569 = n15568 ^ n15560;
  assign n15571 = n15570 ^ n15569;
  assign n15559 = n15496 & n15546;
  assign n15572 = n15571 ^ n15559;
  assign n15557 = n15496 & n15523;
  assign n15558 = n15557 ^ n15496;
  assign n15573 = n15572 ^ n15558;
  assign n15580 = n15573 ^ n15571;
  assign n15552 = ~n15526 & n15546;
  assign n15581 = n15580 ^ n15552;
  assign n15582 = n15581 ^ n15528;
  assign n15579 = n15549 ^ n15539;
  assign n15583 = n15582 ^ n15579;
  assign n15585 = n15584 ^ n15583;
  assign n15825 = n15531 & n15572;
  assign n15826 = n15825 ^ n15559;
  assign n15827 = n15585 & ~n15826;
  assign n15828 = n15544 & n15827;
  assign n15829 = n15828 ^ n15544;
  assign n15586 = n15585 ^ n15535;
  assign n15587 = ~n15542 & ~n15586;
  assign n15830 = n15567 ^ n15547;
  assign n15831 = n15531 & n15830;
  assign n15832 = n15831 ^ n15547;
  assign n15833 = n15530 & n15832;
  assign n15540 = n15532 ^ n15530;
  assign n15834 = n15573 ^ n15537;
  assign n15835 = n15834 ^ n15561;
  assign n15836 = n15540 & n15835;
  assign n15837 = n15548 ^ n15536;
  assign n15838 = ~n15543 & ~n15837;
  assign n15839 = ~n15525 & n15838;
  assign n15545 = n15525 ^ n15497;
  assign n15550 = n15549 ^ n15545;
  assign n15840 = n15550 ^ n15538;
  assign n15841 = n15543 & n15840;
  assign n15842 = n15542 & ~n15841;
  assign n15843 = ~n15839 & ~n15842;
  assign n15844 = ~n15836 & ~n15843;
  assign n15845 = n15557 ^ n15532;
  assign n15846 = n15550 ^ n15543;
  assign n15847 = n15557 & n15846;
  assign n15848 = n15847 ^ n15550;
  assign n15849 = n15845 & n15848;
  assign n15850 = n15849 ^ n15532;
  assign n15851 = n15844 & ~n15850;
  assign n15852 = n15552 ^ n15542;
  assign n15853 = n15580 ^ n15531;
  assign n15854 = ~n15552 & ~n15853;
  assign n15855 = n15854 ^ n15531;
  assign n15856 = ~n15852 & n15855;
  assign n15857 = n15856 ^ n15542;
  assign n15858 = n15851 & n15857;
  assign n15859 = ~n15833 & n15858;
  assign n15860 = ~n15587 & n15859;
  assign n15861 = ~n15829 & n15860;
  assign n15862 = ~n15578 & n15861;
  assign n15863 = ~n15533 & n15862;
  assign n15864 = n15863 ^ n13682;
  assign n15865 = n15864 ^ x607;
  assign n13445 = n13444 ^ x581;
  assign n13115 = n12814 & n12932;
  assign n13112 = n13111 ^ n13091;
  assign n13113 = n12932 & n13112;
  assign n13114 = n13113 ^ n13091;
  assign n13116 = n13115 ^ n13114;
  assign n13117 = ~n13074 & n13116;
  assign n13118 = n13117 ^ n13114;
  assign n13119 = n13085 ^ n12816;
  assign n13120 = n12932 & n13119;
  assign n13121 = n13120 ^ n13085;
  assign n13122 = n13075 & n13121;
  assign n13123 = n13074 & n13086;
  assign n13124 = n13123 ^ n13105;
  assign n13125 = n12932 & n13124;
  assign n13126 = n13125 ^ n13105;
  assign n13129 = n13078 ^ n12932;
  assign n13130 = n13128 & ~n13129;
  assign n13134 = n13133 ^ n13131;
  assign n13135 = n13134 ^ n13106;
  assign n13132 = n13131 ^ n13081;
  assign n13136 = n13135 ^ n13132;
  assign n13137 = n13136 ^ n13132;
  assign n13138 = ~n12932 & ~n13137;
  assign n13139 = n13138 ^ n13132;
  assign n13140 = ~n13074 & ~n13139;
  assign n13141 = n13140 ^ n13132;
  assign n13142 = ~n13130 & n13141;
  assign n13144 = n13143 ^ n13101;
  assign n13145 = n13075 & n13144;
  assign n13146 = n13145 ^ n13101;
  assign n13147 = n13142 & ~n13146;
  assign n13148 = ~n13126 & n13147;
  assign n13149 = ~n13122 & n13148;
  assign n13150 = ~n13118 & n13149;
  assign n13151 = ~n13110 & n13150;
  assign n13152 = ~n13100 & n13151;
  assign n13153 = ~n13095 & n13152;
  assign n13154 = ~n13079 & n13153;
  assign n13155 = n13154 ^ n12480;
  assign n13156 = n13155 ^ x583;
  assign n11189 = n11188 ^ x507;
  assign n11714 = n11713 ^ x502;
  assign n11715 = n11189 & n11714;
  assign n12451 = n12450 ^ x506;
  assign n12511 = ~n12453 & n12510;
  assign n12512 = n12511 ^ n12509;
  assign n12513 = ~n12457 & n12512;
  assign n12530 = n12454 & ~n12529;
  assign n12532 = ~n12456 & n12531;
  assign n12543 = n12520 ^ n12516;
  assign n12549 = n12548 ^ n12543;
  assign n12539 = n12538 ^ n12504;
  assign n12536 = n12535 ^ n12521;
  assign n12537 = n12536 ^ n12509;
  assign n12540 = n12539 ^ n12537;
  assign n12541 = n12453 & n12540;
  assign n12542 = n12541 ^ n12537;
  assign n12550 = n12549 ^ n12542;
  assign n12551 = ~n12457 & ~n12550;
  assign n12552 = n12551 ^ n12549;
  assign n12553 = ~n12534 & n12552;
  assign n12554 = ~n12532 & n12553;
  assign n12555 = ~n12530 & n12554;
  assign n12556 = n12453 & ~n12546;
  assign n12558 = n12557 ^ n12556;
  assign n12559 = n12555 & ~n12558;
  assign n12560 = ~n12519 & n12559;
  assign n12561 = ~n12513 & n12560;
  assign n12562 = n12561 ^ n10009;
  assign n12563 = n12562 ^ x505;
  assign n12564 = n12451 & ~n12563;
  assign n11955 = n11954 ^ x503;
  assign n12145 = ~n12034 & n12144;
  assign n12151 = ~n12033 & n12150;
  assign n12187 = n12186 ^ n12166;
  assign n12195 = n12194 ^ n12187;
  assign n12185 = n12141 ^ n12046;
  assign n12196 = n12195 ^ n12185;
  assign n12177 = n12176 ^ n12155;
  assign n12178 = n12176 ^ n12033;
  assign n12179 = ~n12034 & n12178;
  assign n12180 = n12179 ^ n12176;
  assign n12181 = n12177 & ~n12180;
  assign n12182 = n12181 ^ n12155;
  assign n12183 = n12174 & ~n12182;
  assign n12184 = ~n12173 & n12183;
  assign n12197 = n12196 ^ n12184;
  assign n12198 = n12197 ^ n12184;
  assign n12199 = ~n11999 & n12198;
  assign n12200 = n12199 ^ n12184;
  assign n12201 = n12034 & ~n12200;
  assign n12202 = n12201 ^ n12184;
  assign n12203 = n12162 ^ n11999;
  assign n12207 = n12206 ^ n12204;
  assign n12208 = n12207 ^ n12162;
  assign n12209 = n12162 ^ n12034;
  assign n12210 = ~n12162 & ~n12209;
  assign n12211 = n12210 ^ n12162;
  assign n12212 = ~n12208 & ~n12211;
  assign n12213 = n12212 ^ n12210;
  assign n12214 = n12213 ^ n12162;
  assign n12215 = n12214 ^ n12034;
  assign n12216 = n12203 & ~n12215;
  assign n12217 = n12216 ^ n12162;
  assign n12218 = n12202 & ~n12217;
  assign n12219 = ~n12151 & n12218;
  assign n12220 = ~n12145 & n12219;
  assign n12221 = n12163 ^ n12150;
  assign n12222 = n12221 ^ n12193;
  assign n12223 = n12033 & n12222;
  assign n12224 = n12223 ^ n12193;
  assign n12225 = n11999 & n12224;
  assign n12226 = n12220 & ~n12225;
  assign n12227 = n12226 ^ n10094;
  assign n12228 = n12227 ^ x504;
  assign n12229 = n11955 & n12228;
  assign n12574 = n12229 ^ n12228;
  assign n12575 = n12574 ^ n11955;
  assign n12581 = n12564 & ~n12575;
  assign n12577 = n12564 ^ n12563;
  assign n12578 = n12577 ^ n12451;
  assign n12579 = n12574 & n12578;
  assign n12565 = n12564 ^ n12451;
  assign n12576 = n12565 & ~n12575;
  assign n12580 = n12579 ^ n12576;
  assign n12582 = n12581 ^ n12580;
  assign n12572 = n12451 ^ n12228;
  assign n12573 = ~n11955 & n12572;
  assign n12583 = n12582 ^ n12573;
  assign n12598 = n12583 ^ n12577;
  assign n12567 = n12229 & n12565;
  assign n12595 = n12567 ^ n12229;
  assign n12593 = n12229 & n12564;
  assign n12230 = n12229 ^ n11955;
  assign n12590 = n12230 & n12578;
  assign n12591 = n12590 ^ n12578;
  assign n12587 = n12579 ^ n12575;
  assign n12570 = n12563 ^ n12451;
  assign n12571 = ~n11955 & ~n12570;
  assign n12584 = n12583 ^ n12571;
  assign n12566 = n12230 & n12565;
  assign n12568 = n12567 ^ n12566;
  assign n12569 = n12568 ^ n12565;
  assign n12585 = n12584 ^ n12569;
  assign n12586 = n12585 ^ n12582;
  assign n12588 = n12587 ^ n12586;
  assign n12589 = n12588 ^ n12579;
  assign n12592 = n12591 ^ n12589;
  assign n12594 = n12593 ^ n12592;
  assign n12596 = n12595 ^ n12594;
  assign n12597 = n12596 ^ n12585;
  assign n12599 = n12598 ^ n12597;
  assign n12600 = n11715 & n12599;
  assign n12601 = n11715 ^ n11189;
  assign n12602 = n12601 ^ n11714;
  assign n12603 = n12593 ^ n12590;
  assign n12604 = n12603 ^ n12599;
  assign n12605 = ~n12602 & n12604;
  assign n12606 = n12576 ^ n12569;
  assign n12607 = n12606 ^ n12588;
  assign n12608 = n12607 ^ n12585;
  assign n12609 = ~n11714 & ~n12608;
  assign n12610 = n12609 ^ n12585;
  assign n12611 = n11189 & n12610;
  assign n12612 = n12567 & ~n12602;
  assign n12613 = n12602 ^ n11189;
  assign n12617 = n12587 ^ n11955;
  assign n12616 = n12606 ^ n12583;
  assign n12618 = n12617 ^ n12616;
  assign n12619 = n12618 ^ n12581;
  assign n12615 = n12593 ^ n12564;
  assign n12620 = n12619 ^ n12615;
  assign n12621 = n12620 ^ n12592;
  assign n12614 = n12590 ^ n12566;
  assign n12622 = n12621 ^ n12614;
  assign n12623 = n12613 & ~n12622;
  assign n12625 = n11715 & n12579;
  assign n12624 = n12601 & n12603;
  assign n12626 = n12625 ^ n12624;
  assign n12627 = n11715 & n12568;
  assign n12628 = n11714 ^ n11189;
  assign n12638 = n12589 ^ n12581;
  assign n12639 = ~n12602 & ~n12638;
  assign n12635 = n12583 ^ n12576;
  assign n12636 = n11715 & n12635;
  assign n12637 = n12636 ^ n12618;
  assign n12640 = n12639 ^ n12637;
  assign n12629 = n12620 ^ n12596;
  assign n12630 = n12629 ^ n12592;
  assign n12631 = n12630 ^ n12581;
  assign n12632 = n12631 ^ n12571;
  assign n12633 = n11714 & n12632;
  assign n12634 = n12633 ^ n12631;
  assign n12641 = n12640 ^ n12634;
  assign n12642 = n12628 & n12641;
  assign n12643 = n12642 ^ n12640;
  assign n12644 = ~n12627 & ~n12643;
  assign n12645 = ~n12626 & n12644;
  assign n12646 = ~n12623 & n12645;
  assign n12647 = ~n12612 & n12646;
  assign n12648 = ~n12611 & n12647;
  assign n12649 = ~n12605 & n12648;
  assign n12650 = ~n12600 & n12649;
  assign n12651 = n12650 ^ n11871;
  assign n12652 = n12651 ^ x584;
  assign n13641 = n13156 ^ n12652;
  assign n13642 = n13445 & n13641;
  assign n13614 = n13613 ^ n13612;
  assign n13629 = n13628 ^ n13614;
  assign n13630 = n13629 ^ n12493;
  assign n13631 = n13630 ^ x582;
  assign n13632 = ~n13445 & n13631;
  assign n13633 = n13632 ^ n13631;
  assign n13643 = n13642 ^ n13633;
  assign n13157 = n12652 & n13156;
  assign n13639 = n13157 & n13633;
  assign n13634 = n13633 ^ n13445;
  assign n13636 = n12652 & n13634;
  assign n13637 = ~n13156 & n13636;
  assign n13158 = n13157 ^ n13156;
  assign n13635 = n13158 & n13634;
  assign n13638 = n13637 ^ n13635;
  assign n13640 = n13639 ^ n13638;
  assign n13644 = n13643 ^ n13640;
  assign n13799 = n13266 ^ x526;
  assign n13825 = n13824 ^ x531;
  assign n13826 = n13799 & ~n13825;
  assign n13827 = n13826 ^ n13825;
  assign n13828 = n13827 ^ n13799;
  assign n13829 = ~n12456 & n12527;
  assign n13830 = n12523 ^ n12453;
  assign n13831 = n12773 ^ n12509;
  assign n13832 = n13831 ^ n12779;
  assign n13833 = n12452 & n13832;
  assign n13834 = n13833 ^ n13831;
  assign n13835 = n13834 ^ n12523;
  assign n13836 = n13830 & ~n13835;
  assign n13837 = n13836 ^ n13833;
  assign n13838 = n13837 ^ n13831;
  assign n13839 = n13838 ^ n12453;
  assign n13840 = ~n12523 & ~n13839;
  assign n13841 = n13840 ^ n12523;
  assign n13842 = n13841 ^ n12453;
  assign n13843 = ~n13829 & ~n13842;
  assign n13844 = n12535 ^ n12517;
  assign n13845 = n13844 ^ n12523;
  assign n13846 = n13845 ^ n12521;
  assign n13847 = ~n12452 & ~n13846;
  assign n13848 = n13847 ^ n12521;
  assign n13849 = n12453 & n13848;
  assign n13850 = n13843 & ~n13849;
  assign n13857 = ~n12452 & n12778;
  assign n13851 = n12781 ^ n12500;
  assign n13852 = ~n12518 & n13851;
  assign n13853 = ~n12455 & n13454;
  assign n13854 = n13853 ^ n12780;
  assign n13855 = ~n13852 & ~n13854;
  assign n13856 = n12529 & n13855;
  assign n13858 = n13857 ^ n13856;
  assign n13859 = ~n12453 & ~n13858;
  assign n13860 = n13859 ^ n13856;
  assign n13861 = n13850 & n13860;
  assign n13862 = ~n12513 & n13861;
  assign n13863 = ~n12777 & n13862;
  assign n13864 = n13863 ^ n10584;
  assign n13865 = n13864 ^ x528;
  assign n13866 = n11141 & ~n11152;
  assign n13867 = n10747 ^ n10211;
  assign n13868 = n13867 ^ n10760;
  assign n13869 = n13868 ^ n10745;
  assign n13870 = n11153 & n13869;
  assign n13871 = n11154 & ~n13235;
  assign n13875 = ~n10759 & n13232;
  assign n13876 = n13875 ^ n11181;
  assign n13873 = n11128 & n12727;
  assign n13872 = ~n11167 & ~n13225;
  assign n13874 = n13873 ^ n13872;
  assign n13877 = n13876 ^ n13874;
  assign n13878 = n11009 & n13877;
  assign n13879 = ~n13871 & ~n13878;
  assign n13880 = ~n13870 & n13879;
  assign n13881 = ~n13866 & n13880;
  assign n13882 = ~n11009 & ~n12728;
  assign n13883 = n13882 ^ n11161;
  assign n13884 = ~n11128 & n13883;
  assign n13885 = n13884 ^ n11161;
  assign n13886 = n13881 & ~n13885;
  assign n13887 = ~n12765 & n13886;
  assign n13888 = ~n13252 & n13887;
  assign n13889 = ~n11149 & n13888;
  assign n13890 = n13889 ^ n10611;
  assign n13891 = n13890 ^ x529;
  assign n13892 = ~n13865 & n13891;
  assign n13915 = n13914 ^ x530;
  assign n13916 = n13189 ^ x527;
  assign n13917 = n13915 & ~n13916;
  assign n13925 = n13892 & n13917;
  assign n13926 = n13925 ^ n13917;
  assign n13893 = n13892 ^ n13891;
  assign n13923 = n13893 & n13917;
  assign n13920 = n13893 ^ n13865;
  assign n13921 = n13920 ^ n13891;
  assign n13922 = n13917 & ~n13921;
  assign n13924 = n13923 ^ n13922;
  assign n13927 = n13926 ^ n13924;
  assign n13918 = n13917 ^ n13916;
  assign n13919 = n13893 & ~n13918;
  assign n13928 = n13927 ^ n13919;
  assign n13929 = n13828 & n13928;
  assign n13930 = n13828 ^ n13826;
  assign n13933 = ~n13918 & n13920;
  assign n13931 = n13917 ^ n13915;
  assign n13932 = n13920 & n13931;
  assign n13934 = n13933 ^ n13932;
  assign n13935 = ~n13825 & n13934;
  assign n13936 = n13935 ^ n13932;
  assign n13937 = ~n13930 & n13936;
  assign n13938 = n13918 ^ n13915;
  assign n13941 = n13893 & n13938;
  assign n13942 = n13941 ^ n13893;
  assign n13940 = n13923 ^ n13919;
  assign n13943 = n13942 ^ n13940;
  assign n13939 = n13892 & n13938;
  assign n13944 = n13943 ^ n13939;
  assign n13945 = ~n13827 & n13944;
  assign n13953 = n13927 ^ n13920;
  assign n13954 = n13953 ^ n13934;
  assign n13950 = n13915 ^ n13865;
  assign n13951 = n13950 ^ n13891;
  assign n13952 = n13916 & n13951;
  assign n13955 = n13954 ^ n13952;
  assign n13956 = n13955 ^ n13944;
  assign n13967 = n13956 ^ n13943;
  assign n13947 = n13932 ^ n13931;
  assign n13968 = n13967 ^ n13947;
  assign n13969 = n13968 ^ n13941;
  assign n13946 = ~n13865 & n13916;
  assign n13948 = n13947 ^ n13946;
  assign n13949 = n13948 ^ n13944;
  assign n13961 = n13949 ^ n13932;
  assign n13965 = n13961 ^ n13865;
  assign n13962 = n13961 ^ n13922;
  assign n13958 = n13922 ^ n13921;
  assign n13957 = n13956 ^ n13949;
  assign n13959 = n13958 ^ n13957;
  assign n13960 = n13959 ^ n13925;
  assign n13963 = n13962 ^ n13960;
  assign n13964 = n13963 ^ n13946;
  assign n13966 = n13965 ^ n13964;
  assign n13970 = n13969 ^ n13966;
  assign n13971 = ~n13825 & n13970;
  assign n13972 = n13971 ^ n13966;
  assign n13973 = n13799 & n13972;
  assign n13974 = n13826 ^ n13799;
  assign n13975 = n13933 ^ n13923;
  assign n13976 = n13974 & n13975;
  assign n13977 = n13954 ^ n13826;
  assign n13978 = n13925 ^ n13828;
  assign n13979 = n13826 & ~n13978;
  assign n13980 = n13979 ^ n13828;
  assign n13981 = n13977 & ~n13980;
  assign n13982 = n13981 ^ n13954;
  assign n13983 = n13956 ^ n13939;
  assign n13984 = n13983 ^ n13941;
  assign n13985 = n13828 & n13984;
  assign n13992 = n13825 & ~n13964;
  assign n13993 = n13992 ^ n13963;
  assign n13986 = n13959 ^ n13927;
  assign n13987 = n13986 ^ n13919;
  assign n13988 = n13987 ^ n13922;
  assign n13989 = n13988 ^ n13960;
  assign n13990 = ~n13825 & n13989;
  assign n13991 = n13990 ^ n13960;
  assign n13994 = n13993 ^ n13991;
  assign n13995 = ~n13930 & n13994;
  assign n13996 = n13995 ^ n13991;
  assign n13997 = ~n13985 & n13996;
  assign n13998 = ~n13982 & n13997;
  assign n13999 = ~n13976 & n13998;
  assign n14000 = ~n13973 & n13999;
  assign n14001 = ~n13945 & n14000;
  assign n14002 = ~n13937 & n14001;
  assign n14003 = ~n13929 & n14002;
  assign n14004 = n14003 ^ n11774;
  assign n14005 = n14004 ^ x585;
  assign n13798 = n13797 ^ x580;
  assign n14006 = n14005 ^ n13798;
  assign n14007 = n13644 & ~n14006;
  assign n14008 = n13798 & n14005;
  assign n14009 = n13158 ^ n12652;
  assign n14010 = n14009 ^ n13156;
  assign n14011 = n13633 & n14010;
  assign n14017 = n14011 ^ n13635;
  assign n14013 = n13639 ^ n13633;
  assign n14012 = n14011 ^ n13644;
  assign n14014 = n14013 ^ n14012;
  assign n14015 = n14014 ^ n13637;
  assign n14016 = n14015 ^ n14011;
  assign n14018 = n14017 ^ n14016;
  assign n14019 = n14008 & n14018;
  assign n14020 = n14008 ^ n14005;
  assign n14021 = n14020 ^ n13798;
  assign n14022 = n13637 ^ n13636;
  assign n14023 = n14022 ^ n14014;
  assign n14024 = n14023 ^ n13637;
  assign n14025 = ~n14021 & n14024;
  assign n14046 = n13642 ^ n13641;
  assign n14036 = n13634 ^ n13631;
  assign n14037 = n13158 & ~n14036;
  assign n14038 = n14037 ^ n13158;
  assign n14035 = n14014 ^ n13635;
  assign n14039 = n14038 ^ n14035;
  assign n14033 = n13157 & n13632;
  assign n14040 = n14039 ^ n14033;
  assign n14027 = n13632 & ~n14009;
  assign n14041 = n14040 ^ n14027;
  assign n14042 = n14041 ^ n13632;
  assign n14029 = n13635 ^ n13634;
  assign n14030 = n14029 ^ n13636;
  assign n14028 = n14027 ^ n13640;
  assign n14031 = n14030 ^ n14028;
  assign n14026 = n14009 ^ n13643;
  assign n14032 = n14031 ^ n14026;
  assign n14034 = n14033 ^ n14032;
  assign n14043 = n14042 ^ n14034;
  assign n14044 = n14043 ^ n14037;
  assign n14045 = n14005 & ~n14044;
  assign n14047 = n14046 ^ n14045;
  assign n14048 = n13798 & n14047;
  assign n14049 = n14048 ^ n14046;
  assign n14050 = ~n14025 & ~n14049;
  assign n14057 = n14030 ^ n14017;
  assign n14052 = n14037 ^ n14036;
  assign n14051 = n14046 ^ n14044;
  assign n14053 = n14052 ^ n14051;
  assign n14054 = n14053 ^ n14040;
  assign n14058 = n14057 ^ n14054;
  assign n14055 = n14054 ^ n14044;
  assign n14056 = n14055 ^ n14016;
  assign n14059 = n14058 ^ n14056;
  assign n14060 = ~n14005 & n14059;
  assign n14061 = n14060 ^ n14058;
  assign n14062 = n14006 & n14061;
  assign n14063 = n14050 & ~n14062;
  assign n14064 = ~n14019 & n14063;
  assign n14065 = ~n14007 & n14064;
  assign n14066 = n14065 ^ n13462;
  assign n15901 = n14066 ^ x608;
  assign n15923 = ~n15865 & ~n15901;
  assign n14071 = n13190 & n13353;
  assign n14068 = n13190 & n13397;
  assign n14069 = n14068 ^ n13408;
  assign n14070 = n14069 ^ n13412;
  assign n14072 = n14071 ^ n14070;
  assign n14073 = ~n13218 & n14072;
  assign n14074 = n14073 ^ n14071;
  assign n14075 = n13394 ^ n13218;
  assign n14076 = n13417 ^ n13411;
  assign n14077 = n14076 ^ n13414;
  assign n14078 = ~n14075 & ~n14077;
  assign n14079 = ~n13218 & n13417;
  assign n14090 = n13433 ^ n13409;
  assign n14091 = n14090 ^ n13368;
  assign n14088 = n13413 ^ n13364;
  assign n14089 = n14088 ^ n13368;
  assign n14092 = n14091 ^ n14089;
  assign n14093 = ~n13190 & n14092;
  assign n14094 = n14093 ^ n14089;
  assign n14080 = n13413 ^ n13348;
  assign n14081 = n14080 ^ n13402;
  assign n14083 = n14081 ^ n13364;
  assign n14084 = n14083 ^ n13366;
  assign n14082 = n14081 ^ n13356;
  assign n14085 = n14084 ^ n14082;
  assign n14086 = ~n13190 & ~n14085;
  assign n14087 = n14086 ^ n14082;
  assign n14095 = n14094 ^ n14087;
  assign n14096 = ~n13384 & ~n14095;
  assign n14097 = n14096 ^ n14087;
  assign n14098 = ~n14079 & ~n14097;
  assign n14099 = ~n14078 & n14098;
  assign n14100 = ~n14074 & n14099;
  assign n14101 = ~n13379 & n14100;
  assign n14102 = n14101 ^ n10524;
  assign n14103 = n14102 ^ x547;
  assign n14105 = n12592 ^ n12581;
  assign n14106 = n11714 & ~n14105;
  assign n14107 = n14106 ^ n12592;
  assign n14108 = n11189 & ~n14107;
  assign n14104 = n12599 & n12601;
  assign n14109 = n14108 ^ n14104;
  assign n14110 = n12601 & n12619;
  assign n14111 = ~n12608 & n12613;
  assign n14112 = ~n12594 & n12613;
  assign n14113 = n12618 ^ n12585;
  assign n14114 = ~n12602 & n14113;
  assign n14119 = n12581 ^ n12568;
  assign n14120 = n11714 & n14119;
  assign n14117 = n12614 ^ n12600;
  assign n14115 = ~n12602 & n12620;
  assign n14116 = n14115 ^ n12596;
  assign n14118 = n14117 ^ n14116;
  assign n14121 = n14120 ^ n14118;
  assign n14122 = n12628 & ~n14121;
  assign n14123 = n14122 ^ n14118;
  assign n14124 = ~n14114 & n14123;
  assign n14126 = n11189 & n12616;
  assign n14125 = n12579 ^ n12567;
  assign n14127 = n14126 ^ n14125;
  assign n14128 = n11714 & n14127;
  assign n14129 = n14128 ^ n14125;
  assign n14130 = n14124 & ~n14129;
  assign n14131 = ~n14112 & n14130;
  assign n14132 = ~n14111 & n14131;
  assign n14133 = ~n14110 & n14132;
  assign n14134 = ~n14109 & n14133;
  assign n14135 = ~n12626 & n14134;
  assign n14136 = n14135 ^ n10210;
  assign n14137 = n14136 ^ x546;
  assign n14138 = n14103 & n14137;
  assign n14139 = n14138 ^ n14103;
  assign n14140 = n14139 ^ n14137;
  assign n14141 = n14140 ^ n14103;
  assign n14144 = n13463 & ~n13617;
  assign n14145 = n14144 ^ n13584;
  assign n14142 = ~n13463 & ~n13605;
  assign n14143 = n14142 ^ n13604;
  assign n14146 = n14145 ^ n14143;
  assign n14147 = n13613 & n14146;
  assign n14148 = n14147 ^ n14145;
  assign n14149 = ~n13606 & n14148;
  assign n14150 = n14149 ^ n9778;
  assign n14151 = n14150 ^ x545;
  assign n14152 = n13960 ^ n13954;
  assign n14153 = ~n13827 & ~n14152;
  assign n14154 = n13828 & n13933;
  assign n14155 = n13966 ^ n13927;
  assign n14156 = n14155 ^ n13954;
  assign n14157 = n13826 & n14156;
  assign n14158 = ~n13825 & n13967;
  assign n14159 = n14158 ^ n13943;
  assign n14160 = n13930 & n14159;
  assign n14168 = n13954 ^ n13940;
  assign n14169 = n14168 ^ n13939;
  assign n14170 = n14169 ^ n13960;
  assign n14161 = n13957 ^ n13944;
  assign n14162 = n13957 ^ n13799;
  assign n14163 = ~n13930 & n14162;
  assign n14164 = n14163 ^ n13799;
  assign n14165 = n14161 & ~n14164;
  assign n14166 = n14165 ^ n13944;
  assign n14167 = ~n13941 & ~n14166;
  assign n14171 = n14170 ^ n14167;
  assign n14172 = n14171 ^ n14167;
  assign n14173 = n13825 & ~n14172;
  assign n14174 = n14173 ^ n14167;
  assign n14175 = ~n13930 & ~n14174;
  assign n14176 = n14175 ^ n14167;
  assign n14178 = ~n13827 & n13969;
  assign n14177 = ~n13930 & n13961;
  assign n14179 = n14178 ^ n14177;
  assign n14180 = n14176 & ~n14179;
  assign n14181 = ~n14160 & n14180;
  assign n14182 = ~n14157 & n14181;
  assign n14183 = ~n14154 & n14182;
  assign n14184 = ~n13799 & n13923;
  assign n14185 = n14184 ^ n13922;
  assign n14186 = ~n13930 & n14185;
  assign n14187 = n14186 ^ n13922;
  assign n14188 = n14183 & ~n14187;
  assign n14189 = ~n14153 & n14188;
  assign n14190 = ~n13929 & n14189;
  assign n14191 = n14190 ^ n10740;
  assign n14192 = n14191 ^ x548;
  assign n14193 = n14151 & ~n14192;
  assign n14357 = n14141 & n14193;
  assign n14194 = n14193 ^ n14151;
  assign n14195 = n14194 ^ n14192;
  assign n14196 = n14195 ^ n14151;
  assign n14197 = n14141 & ~n14196;
  assign n14252 = n14250 & n14251;
  assign n14281 = n14280 ^ n14279;
  assign n14282 = n14253 & ~n14281;
  assign n14283 = ~n14252 & ~n14282;
  assign n14284 = n14199 & n14266;
  assign n14285 = n14284 ^ n14265;
  assign n14286 = n14198 & n14285;
  assign n14287 = n14283 & ~n14286;
  assign n14292 = n14262 ^ n14204;
  assign n14295 = n14294 ^ n14292;
  assign n14296 = n14295 ^ n14268;
  assign n14297 = ~n14198 & ~n14296;
  assign n14291 = n14290 ^ n14288;
  assign n14298 = n14297 ^ n14291;
  assign n14299 = ~n14199 & ~n14298;
  assign n14300 = n14299 ^ n14291;
  assign n14301 = n14287 & n14300;
  assign n14302 = ~n14247 & n14301;
  assign n14303 = n14302 ^ n11127;
  assign n14304 = n14303 ^ x544;
  assign n14313 = n13133 ^ n13106;
  assign n14314 = n12932 & n14313;
  assign n14315 = n14314 ^ n13133;
  assign n14316 = n13075 & n14315;
  assign n14317 = ~n13122 & ~n14316;
  assign n14318 = ~n13074 & n13133;
  assign n14319 = n14318 ^ n13085;
  assign n14320 = n13075 & n14319;
  assign n14321 = n14320 ^ n13085;
  assign n14323 = n13101 ^ n13081;
  assign n14324 = n14323 ^ n13086;
  assign n14322 = n13127 ^ n12814;
  assign n14325 = n14324 ^ n14322;
  assign n14326 = n14325 ^ n14322;
  assign n14327 = ~n12932 & n14326;
  assign n14328 = n14327 ^ n14322;
  assign n14329 = ~n13074 & n14328;
  assign n14330 = n14329 ^ n14322;
  assign n14331 = ~n14321 & ~n14330;
  assign n14332 = n14306 ^ n12813;
  assign n14333 = n12932 & ~n14332;
  assign n14334 = n14333 ^ n12813;
  assign n14335 = n13074 & n14334;
  assign n14336 = n14331 & ~n14335;
  assign n14337 = ~n13126 & n14336;
  assign n14338 = ~n13118 & n14337;
  assign n14339 = n14317 & n14338;
  assign n14340 = n14312 & n14339;
  assign n14341 = n14340 ^ n11008;
  assign n14342 = n14341 ^ x549;
  assign n14343 = n14304 & ~n14342;
  assign n14344 = n14343 ^ n14304;
  assign n14345 = n14197 & n14344;
  assign n14374 = n14139 & n14193;
  assign n14375 = n14374 ^ n14357;
  assign n14368 = ~n14140 & n14193;
  assign n14373 = n14368 ^ n14193;
  assign n14376 = n14375 ^ n14373;
  assign n14371 = n14357 ^ n14141;
  assign n14361 = n14141 & n14195;
  assign n14370 = n14361 ^ n14197;
  assign n14372 = n14371 ^ n14370;
  assign n14377 = n14376 ^ n14372;
  assign n15866 = n14377 ^ n14374;
  assign n14367 = n14138 & n14194;
  assign n15867 = n15866 ^ n14367;
  assign n15868 = ~n14342 & n15867;
  assign n15869 = n15868 ^ n14367;
  assign n15870 = ~n14304 & n15869;
  assign n15871 = ~n14345 & ~n15870;
  assign n14366 = n14343 ^ n14342;
  assign n15872 = n14366 ^ n14304;
  assign n14379 = n14139 & n14194;
  assign n14380 = n14379 ^ n14375;
  assign n14381 = n14380 ^ n14151;
  assign n14369 = n14368 ^ n14367;
  assign n14378 = n14377 ^ n14369;
  assign n14382 = n14381 ^ n14378;
  assign n14352 = n14151 ^ n14137;
  assign n14353 = n14192 ^ n14137;
  assign n14354 = ~n14352 & n14353;
  assign n14386 = n14382 ^ n14354;
  assign n14383 = n14382 ^ n14357;
  assign n14384 = n14383 ^ n14376;
  assign n14358 = n14357 ^ n14139;
  assign n14347 = n14151 ^ n14103;
  assign n14348 = n14347 ^ n14192;
  assign n14349 = n14348 ^ n14137;
  assign n14350 = n14349 ^ n14151;
  assign n14351 = n14350 ^ n14192;
  assign n14355 = n14354 ^ n14137;
  assign n14356 = n14351 & ~n14355;
  assign n14359 = n14358 ^ n14356;
  assign n14385 = n14384 ^ n14359;
  assign n14387 = n14386 ^ n14385;
  assign n15873 = n15872 ^ n14387;
  assign n14402 = n14380 ^ n14356;
  assign n15874 = n14402 ^ n14366;
  assign n15875 = ~n14387 & n15874;
  assign n15876 = n15875 ^ n14366;
  assign n15877 = n15873 & ~n15876;
  assign n15878 = n15877 ^ n15872;
  assign n14346 = n14342 ^ n14304;
  assign n14360 = n14359 ^ n14197;
  assign n14362 = n14361 ^ n14360;
  assign n14363 = ~n14342 & n14362;
  assign n14364 = n14363 ^ n14361;
  assign n14365 = n14346 & n14364;
  assign n15885 = n14356 ^ n14348;
  assign n14388 = n14387 ^ n14197;
  assign n14400 = n14388 ^ n14195;
  assign n14401 = n14400 ^ n14362;
  assign n14403 = n14402 ^ n14401;
  assign n14404 = n14403 ^ n14382;
  assign n14405 = n14404 ^ n14377;
  assign n15886 = n15885 ^ n14405;
  assign n15887 = n14342 & n15886;
  assign n15888 = n15887 ^ n14405;
  assign n14415 = ~n14140 & ~n14196;
  assign n14416 = n14415 ^ n14401;
  assign n15881 = n14416 ^ n14379;
  assign n14412 = n14138 & ~n14196;
  assign n15879 = n14412 ^ n14359;
  assign n15880 = n15879 ^ n14368;
  assign n15882 = n15881 ^ n15880;
  assign n15883 = n14342 & n15882;
  assign n15884 = n15883 ^ n15880;
  assign n15889 = n15888 ^ n15884;
  assign n15890 = ~n14304 & n15889;
  assign n15891 = n15890 ^ n15888;
  assign n15892 = ~n14365 & ~n15891;
  assign n15893 = ~n15878 & n15892;
  assign n15894 = n15871 & n15893;
  assign n15895 = ~n14357 & n15894;
  assign n15896 = n15895 ^ n11188;
  assign n15897 = n15896 ^ x605;
  assign n15924 = n15923 ^ n15897;
  assign n14526 = n14525 ^ n14519;
  assign n14527 = n14526 ^ n14507;
  assign n14528 = ~n14488 & n14527;
  assign n14529 = n14528 ^ n14507;
  assign n14530 = n14492 & n14529;
  assign n14753 = n14553 ^ n14515;
  assign n14754 = ~n14542 & n14753;
  assign n14757 = n14756 ^ n14754;
  assign n14765 = n14536 ^ n14487;
  assign n14766 = n14544 & n14765;
  assign n14543 = n14499 & ~n14542;
  assign n14546 = n14545 ^ n14543;
  assign n15215 = ~n14492 & n14495;
  assign n15216 = n14516 ^ n14487;
  assign n15217 = n15216 ^ n14524;
  assign n15218 = ~n14542 & ~n15217;
  assign n15219 = ~n15215 & ~n15218;
  assign n15227 = n14505 ^ n14499;
  assign n15228 = n14492 & n15227;
  assign n15220 = n14553 ^ n14532;
  assign n15221 = ~n14541 & ~n15220;
  assign n15223 = ~n14753 & n15222;
  assign n15224 = ~n14522 & n15223;
  assign n15225 = ~n15221 & ~n15224;
  assign n15226 = ~n14504 & ~n15225;
  assign n15229 = n15228 ^ n15226;
  assign n15230 = ~n14488 & ~n15229;
  assign n15231 = n15230 ^ n15226;
  assign n15232 = n14494 & ~n14531;
  assign n15233 = n15231 & ~n15232;
  assign n15234 = n15219 & n15233;
  assign n15235 = ~n14546 & n15234;
  assign n15236 = ~n14766 & n15235;
  assign n15237 = ~n14757 & n15236;
  assign n15238 = ~n14530 & n15237;
  assign n15239 = ~n14776 & n15238;
  assign n15240 = ~n14497 & n15239;
  assign n15241 = n15240 ^ n12329;
  assign n15607 = n15241 ^ x567;
  assign n14916 = n14250 & ~n14296;
  assign n14919 = n14276 ^ n14265;
  assign n14920 = n14919 ^ n14263;
  assign n14918 = n14917 ^ n14280;
  assign n14921 = n14920 ^ n14918;
  assign n14922 = n14921 ^ n14918;
  assign n14923 = n14198 & n14922;
  assign n14924 = n14923 ^ n14918;
  assign n14925 = n14199 & ~n14924;
  assign n14926 = n14925 ^ n14918;
  assign n14927 = ~n14916 & n14926;
  assign n14928 = n14279 ^ n14238;
  assign n14929 = ~n14198 & ~n14928;
  assign n14930 = n14929 ^ n14238;
  assign n14931 = ~n14199 & n14930;
  assign n14932 = n14927 & ~n14931;
  assign n14933 = ~n14915 & n14932;
  assign n14934 = ~n14247 & n14933;
  assign n14935 = n14934 ^ n12065;
  assign n15608 = n14935 ^ x562;
  assign n15609 = ~n13129 & ~n14305;
  assign n15610 = ~n13078 & n13127;
  assign n15613 = n12772 ^ n12721;
  assign n15612 = n13091 ^ n12813;
  assign n15614 = n15613 ^ n15612;
  assign n15615 = n13074 & ~n15614;
  assign n15611 = n13087 ^ n13081;
  assign n15616 = n15615 ^ n15611;
  assign n15617 = n13075 & n15616;
  assign n15618 = n15617 ^ n15611;
  assign n15624 = n13106 ^ n12816;
  assign n15625 = n15624 ^ n14305;
  assign n15619 = n14323 ^ n13085;
  assign n15620 = n15619 ^ n13111;
  assign n15621 = n15620 ^ n15612;
  assign n15622 = ~n13074 & n15621;
  assign n15623 = n15622 ^ n15612;
  assign n15626 = n15625 ^ n15623;
  assign n15627 = n15626 ^ n15623;
  assign n15628 = ~n13074 & ~n15627;
  assign n15629 = n15628 ^ n15623;
  assign n15630 = n15629 ^ n15623;
  assign n15631 = ~n13101 & ~n15630;
  assign n15632 = n15631 ^ n15623;
  assign n15633 = ~n12932 & ~n15632;
  assign n15634 = n15633 ^ n15623;
  assign n15635 = ~n15618 & ~n15634;
  assign n15636 = ~n13079 & n15635;
  assign n15637 = ~n15610 & n15636;
  assign n15638 = ~n15609 & n15637;
  assign n15639 = ~n12932 & n13111;
  assign n15640 = n15639 ^ n13086;
  assign n15641 = ~n13074 & n15640;
  assign n15642 = n15641 ^ n13086;
  assign n15643 = n15638 & ~n15642;
  assign n15644 = n14317 & n15643;
  assign n15645 = n15644 ^ n12847;
  assign n15646 = n15645 ^ x565;
  assign n14638 = n13375 & ~n14075;
  assign n14639 = n14638 ^ n13390;
  assign n15647 = n13392 ^ n13370;
  assign n15648 = n15647 ^ n14083;
  assign n15649 = ~n13394 & ~n15648;
  assign n14648 = n14080 ^ n14076;
  assign n15650 = n14648 ^ n13364;
  assign n15651 = n15650 ^ n13373;
  assign n15652 = n15650 ^ n13391;
  assign n15653 = ~n15650 & ~n15652;
  assign n15654 = n15653 ^ n15650;
  assign n15655 = n15651 & ~n15654;
  assign n15656 = n15655 ^ n15653;
  assign n15657 = n15656 ^ n15650;
  assign n15658 = n15657 ^ n13391;
  assign n15659 = ~n15649 & ~n15658;
  assign n15660 = n15659 ^ n15649;
  assign n15662 = n13433 ^ n13367;
  assign n15663 = n15662 ^ n13404;
  assign n15661 = n13399 ^ n13395;
  assign n15664 = n15663 ^ n15661;
  assign n15665 = n13190 & ~n15664;
  assign n15666 = n15665 ^ n15661;
  assign n15667 = n13384 & n15666;
  assign n15668 = ~n15660 & ~n15667;
  assign n15669 = ~n14078 & n15668;
  assign n15670 = ~n14639 & n15669;
  assign n15671 = n15670 ^ n12869;
  assign n15672 = n15671 ^ x564;
  assign n14608 = n13647 ^ n13646;
  assign n15100 = n13764 & ~n14608;
  assign n15101 = n13735 ^ n13716;
  assign n15102 = n13647 ^ n13645;
  assign n15103 = n15101 & ~n15102;
  assign n15105 = n13773 ^ n13745;
  assign n15104 = n13739 ^ n13731;
  assign n15106 = n15105 ^ n15104;
  assign n15107 = n13647 & n15106;
  assign n15113 = n13646 & n13729;
  assign n15108 = n13750 ^ n13727;
  assign n15109 = n15108 ^ n13717;
  assign n15110 = n15109 ^ n13736;
  assign n15111 = ~n13646 & ~n15110;
  assign n15112 = n15111 ^ n13736;
  assign n15114 = n15113 ^ n15112;
  assign n15115 = ~n13645 & n15114;
  assign n15116 = n15115 ^ n15112;
  assign n15117 = ~n15107 & ~n15116;
  assign n15118 = ~n13751 & n15117;
  assign n15119 = ~n15103 & n15118;
  assign n15120 = ~n15100 & n15119;
  assign n15121 = n13646 & n13739;
  assign n15122 = n15121 ^ n13733;
  assign n15123 = ~n13763 & n15122;
  assign n15124 = n15123 ^ n13733;
  assign n15125 = n15120 & ~n15124;
  assign n15126 = ~n13762 & n15125;
  assign n15127 = ~n13756 & n15126;
  assign n15128 = n15127 ^ n12266;
  assign n15674 = n15128 ^ x566;
  assign n15021 = n12592 ^ n12566;
  assign n15022 = n15021 ^ n12629;
  assign n15023 = n11189 & n15022;
  assign n15024 = n15023 ^ n12629;
  assign n15025 = n11714 & ~n15024;
  assign n15026 = ~n12602 & ~n12621;
  assign n15027 = n12563 ^ n12228;
  assign n15028 = n12573 ^ n12451;
  assign n15029 = n15027 & n15028;
  assign n15030 = n12601 & n15029;
  assign n15031 = n12603 & ~n12628;
  assign n15032 = n12590 ^ n12567;
  assign n15033 = n15032 ^ n12618;
  assign n15034 = n15033 ^ n12586;
  assign n15035 = ~n11714 & n15034;
  assign n15036 = n15035 ^ n15033;
  assign n15037 = ~n11189 & n15036;
  assign n15038 = ~n15031 & ~n15037;
  assign n15039 = ~n12636 & n15038;
  assign n15040 = ~n15030 & n15039;
  assign n15041 = ~n15026 & n15040;
  assign n15042 = ~n14111 & n15041;
  assign n15043 = ~n15025 & n15042;
  assign n15044 = ~n12611 & n15043;
  assign n15045 = ~n14109 & n15044;
  assign n15046 = n15045 ^ n12032;
  assign n15673 = n15046 ^ x563;
  assign n15675 = n15674 ^ n15673;
  assign n15676 = n15675 ^ n15672;
  assign n15677 = n15672 & n15676;
  assign n15905 = n15677 ^ n15673;
  assign n15906 = ~n15646 & n15905;
  assign n15907 = n15906 ^ n15676;
  assign n15702 = n15674 ^ n15672;
  assign n15703 = n15702 ^ n15646;
  assign n15684 = n15672 ^ n15646;
  assign n15685 = n15673 & ~n15684;
  assign n15686 = n15685 ^ n15672;
  assign n15687 = ~n15675 & n15686;
  assign n15704 = n15703 ^ n15687;
  assign n15908 = n15907 ^ n15704;
  assign n15909 = n15608 & ~n15908;
  assign n15910 = n15909 ^ n15907;
  assign n15697 = n15674 ^ n15646;
  assign n15688 = n15687 ^ n15686;
  assign n15678 = n15677 ^ n15672;
  assign n15695 = n15688 ^ n15678;
  assign n15718 = n15695 ^ n15673;
  assign n15719 = ~n15697 & n15718;
  assign n15682 = n15673 ^ n15672;
  assign n15693 = n15674 & ~n15682;
  assign n15711 = n15693 ^ n15673;
  assign n15698 = n15646 & n15697;
  assign n15699 = n15698 ^ n15672;
  assign n15712 = n15711 ^ n15699;
  assign n15720 = n15719 ^ n15712;
  assign n15721 = n15720 ^ n15673;
  assign n15722 = n15721 ^ n15674;
  assign n15708 = n15673 ^ n15646;
  assign n15723 = n15722 ^ n15708;
  assign n15710 = n15693 ^ n15674;
  assign n15713 = n15712 ^ n15675;
  assign n15700 = ~n15673 & ~n15699;
  assign n15701 = n15700 ^ n15697;
  assign n15705 = n15704 ^ n15701;
  assign n15714 = n15713 ^ n15705;
  assign n15715 = n15714 ^ n15673;
  assign n15716 = n15715 ^ n15672;
  assign n15717 = n15710 & n15716;
  assign n15724 = n15723 ^ n15717;
  assign n15902 = n15724 ^ n15701;
  assign n15903 = ~n15608 & n15902;
  assign n15904 = n15903 ^ n15724;
  assign n15911 = n15910 ^ n15904;
  assign n15912 = n15607 & ~n15911;
  assign n15913 = n15912 ^ n15910;
  assign n15914 = n15913 ^ n13698;
  assign n15915 = n15914 ^ x606;
  assign n15931 = n15915 ^ n15897;
  assign n15932 = ~n15924 & n15931;
  assign n15898 = n15865 & n15897;
  assign n15899 = n15898 ^ n15865;
  assign n15916 = n15901 & ~n15915;
  assign n15917 = n15916 ^ n15915;
  assign n15918 = n15917 ^ n15901;
  assign n15930 = n15899 & n15918;
  assign n15933 = n15932 ^ n15930;
  assign n15925 = n15915 ^ n15901;
  assign n15926 = n15925 ^ n15897;
  assign n15927 = n15926 ^ n15865;
  assign n15928 = ~n15924 & n15927;
  assign n15900 = n15899 ^ n15897;
  assign n15921 = ~n15900 & n15916;
  assign n15919 = n15918 ^ n15915;
  assign n15920 = ~n15900 & n15919;
  assign n15922 = n15921 ^ n15920;
  assign n15929 = n15928 ^ n15922;
  assign n15934 = n15933 ^ n15929;
  assign n14426 = n14191 ^ x550;
  assign n14537 = n14536 ^ n14532;
  assign n14538 = n14492 & n14537;
  assign n14539 = n14538 ^ n14536;
  assign n14540 = n14531 & n14539;
  assign n14547 = n14524 ^ n14495;
  assign n14548 = n14488 & ~n14547;
  assign n14549 = n14548 ^ n14495;
  assign n14550 = n14492 & n14549;
  assign n14551 = n14508 & ~n14542;
  assign n14554 = n14553 ^ n14522;
  assign n14555 = ~n14522 & ~n14542;
  assign n14556 = n14555 ^ n14492;
  assign n14557 = n14554 & ~n14556;
  assign n14558 = n14557 ^ n14553;
  assign n14559 = ~n14551 & ~n14558;
  assign n14560 = n14492 & n14494;
  assign n14561 = n14560 ^ n14516;
  assign n14562 = n14531 & n14561;
  assign n14563 = n14562 ^ n14516;
  assign n14565 = n14488 & n14515;
  assign n14564 = n14526 & n14541;
  assign n14566 = n14565 ^ n14564;
  assign n14567 = ~n14563 & ~n14566;
  assign n14568 = n14559 & n14567;
  assign n14569 = ~n14550 & n14568;
  assign n14570 = ~n14546 & n14569;
  assign n14571 = ~n14540 & n14570;
  assign n14572 = ~n14530 & n14571;
  assign n14573 = ~n14500 & n14572;
  assign n14574 = ~n14497 & n14573;
  assign n14575 = ~n14487 & n14574;
  assign n14576 = n14575 ^ n12140;
  assign n14577 = n14576 ^ x555;
  assign n14578 = n14275 ^ n14258;
  assign n14579 = n14249 & n14578;
  assign n14586 = ~n14198 & n14278;
  assign n14587 = n14586 ^ n14273;
  assign n14581 = n14251 ^ n14200;
  assign n14582 = n14581 ^ n14279;
  assign n14580 = n14272 ^ n14238;
  assign n14583 = n14582 ^ n14580;
  assign n14584 = n14198 & ~n14583;
  assign n14585 = n14584 ^ n14580;
  assign n14588 = n14587 ^ n14585;
  assign n14589 = ~n14199 & n14588;
  assign n14590 = n14589 ^ n14585;
  assign n14591 = ~n14579 & ~n14590;
  assign n14594 = n14593 ^ n14279;
  assign n14592 = n14291 ^ n14260;
  assign n14595 = n14594 ^ n14592;
  assign n14596 = n14595 ^ n14592;
  assign n14597 = ~n14198 & ~n14596;
  assign n14598 = n14597 ^ n14592;
  assign n14599 = ~n14253 & ~n14598;
  assign n14600 = n14599 ^ n14592;
  assign n14601 = n14591 & n14600;
  assign n14602 = n14601 ^ n12954;
  assign n14603 = n14602 ^ x553;
  assign n14604 = n13646 & n13764;
  assign n14605 = n14604 ^ n13750;
  assign n14606 = ~n13763 & ~n14605;
  assign n14607 = n14606 ^ n13750;
  assign n14609 = n13789 ^ n13716;
  assign n14610 = n14609 ^ n13726;
  assign n14611 = n14610 ^ n13746;
  assign n14612 = n14611 ^ n13739;
  assign n14613 = ~n14608 & n14612;
  assign n14614 = n13699 ^ n13648;
  assign n14615 = n14614 ^ n13737;
  assign n14616 = n14615 ^ n13747;
  assign n14617 = n14616 ^ n13747;
  assign n14618 = n13646 & ~n14617;
  assign n14619 = n14618 ^ n13747;
  assign n14620 = ~n13763 & ~n14619;
  assign n14621 = n14620 ^ n13747;
  assign n14622 = ~n14613 & n14621;
  assign n14624 = n13705 ^ n13701;
  assign n14623 = n13789 ^ n13720;
  assign n14625 = n14624 ^ n14623;
  assign n14626 = ~n13646 & ~n14625;
  assign n14627 = n14626 ^ n14623;
  assign n14628 = ~n13645 & n14627;
  assign n14629 = n14622 & ~n14628;
  assign n14630 = ~n13793 & n14629;
  assign n14631 = n14607 & n14630;
  assign n14632 = n14631 ^ n12986;
  assign n14633 = n14632 ^ x552;
  assign n14634 = ~n14603 & n14633;
  assign n14635 = n14634 ^ n14603;
  assign n14637 = n14341 ^ x551;
  assign n14640 = ~n13218 & n13367;
  assign n14641 = n13391 & ~n14083;
  assign n14642 = ~n14640 & ~n14641;
  assign n14649 = n14648 ^ n13371;
  assign n14644 = n13362 ^ n13359;
  assign n14643 = n14076 ^ n13398;
  assign n14645 = n14644 ^ n14643;
  assign n14646 = n13218 & n14645;
  assign n14647 = n14646 ^ n14643;
  assign n14650 = n14649 ^ n14647;
  assign n14651 = n14650 ^ n14647;
  assign n14652 = n13218 & n14651;
  assign n14653 = n14652 ^ n14647;
  assign n14654 = ~n13190 & ~n14653;
  assign n14655 = n14654 ^ n14647;
  assign n14656 = n14642 & n14655;
  assign n14657 = ~n14074 & n14656;
  assign n14658 = ~n13383 & n14657;
  assign n14659 = ~n14639 & n14658;
  assign n14660 = n14659 ^ n11998;
  assign n14661 = n14660 ^ x554;
  assign n14662 = n14637 & ~n14661;
  assign n14669 = n14662 ^ n14637;
  assign n14676 = ~n14635 & n14669;
  assign n14636 = n14635 ^ n14633;
  assign n14665 = n14636 ^ n14603;
  assign n14667 = n14662 & n14665;
  assign n14678 = n14676 ^ n14667;
  assign n14675 = n14634 & n14662;
  assign n14683 = n14678 ^ n14675;
  assign n14684 = n14683 ^ n14637;
  assign n14672 = n14636 & n14662;
  assign n14679 = n14678 ^ n14672;
  assign n14680 = n14679 ^ n14662;
  assign n14677 = n14676 ^ n14675;
  assign n14681 = n14680 ^ n14677;
  assign n14671 = n14634 & n14669;
  assign n14673 = n14672 ^ n14671;
  assign n14670 = n14636 & n14669;
  assign n14674 = n14673 ^ n14670;
  assign n14682 = n14681 ^ n14674;
  assign n14685 = n14684 ^ n14682;
  assign n14686 = n14685 ^ n14665;
  assign n14663 = n14662 ^ n14661;
  assign n14666 = ~n14663 & n14665;
  assign n14668 = n14667 ^ n14666;
  assign n14687 = n14686 ^ n14668;
  assign n14664 = n14636 & ~n14663;
  assign n14688 = n14687 ^ n14664;
  assign n14689 = n14688 ^ n14673;
  assign n14690 = n14577 & n14689;
  assign n14691 = n14690 ^ n14673;
  assign n14692 = ~n14426 & n14691;
  assign n14693 = n14577 & n14668;
  assign n14694 = n14693 ^ n14666;
  assign n14695 = ~n14426 & n14694;
  assign n14696 = n14426 & n14577;
  assign n14697 = n14696 ^ n14426;
  assign n14699 = n14634 & ~n14663;
  assign n14700 = n14699 ^ n14663;
  assign n14698 = n14666 ^ n14664;
  assign n14701 = n14700 ^ n14698;
  assign n14702 = n14701 ^ n14687;
  assign n14703 = n14697 & ~n14702;
  assign n14704 = n14577 ^ n14426;
  assign n14706 = n14675 ^ n14634;
  assign n14705 = n14699 ^ n14671;
  assign n14707 = n14706 ^ n14705;
  assign n14708 = n14707 ^ n14664;
  assign n14709 = ~n14426 & n14708;
  assign n14710 = n14709 ^ n14664;
  assign n14711 = n14704 & n14710;
  assign n14712 = ~n14703 & ~n14711;
  assign n14713 = n14699 ^ n14681;
  assign n14714 = ~n14426 & n14713;
  assign n14715 = n14714 ^ n14699;
  assign n14716 = n14577 & n14715;
  assign n14717 = n14697 & n14707;
  assign n14718 = n14663 ^ n14637;
  assign n14719 = ~n14635 & n14718;
  assign n14720 = n14719 ^ n14707;
  assign n14721 = n14720 ^ n14718;
  assign n14722 = n14721 ^ n14687;
  assign n14723 = n14722 ^ n14701;
  assign n14724 = n14723 ^ n14719;
  assign n14725 = ~n14704 & ~n14724;
  assign n14732 = n14674 ^ n14667;
  assign n14727 = n14685 ^ n14670;
  assign n14728 = n14727 ^ n14667;
  assign n14729 = n14728 ^ n14671;
  assign n14730 = n14729 ^ n14637;
  assign n14726 = n14685 ^ n14681;
  assign n14731 = n14730 ^ n14726;
  assign n14733 = n14732 ^ n14731;
  assign n14734 = n14577 & n14733;
  assign n14735 = n14734 ^ n14731;
  assign n14736 = n14426 & n14735;
  assign n14737 = ~n14725 & ~n14736;
  assign n14738 = ~n14717 & n14737;
  assign n14739 = n14705 ^ n14670;
  assign n14740 = n14739 ^ n14678;
  assign n14741 = n14577 & n14740;
  assign n14742 = n14741 ^ n14678;
  assign n14743 = ~n14426 & n14742;
  assign n14744 = n14738 & ~n14743;
  assign n14745 = ~n14716 & n14744;
  assign n14746 = n14712 & n14745;
  assign n14747 = ~n14695 & n14746;
  assign n14748 = ~n14692 & n14747;
  assign n14749 = n14748 ^ n13494;
  assign n15935 = n14749 ^ x609;
  assign n15129 = n15128 ^ x568;
  assign n15151 = n15150 ^ x573;
  assign n15152 = ~n15129 & ~n15151;
  assign n15315 = n15152 ^ n15129;
  assign n15157 = n15156 ^ x572;
  assign n14937 = n13986 ^ n13954;
  assign n14938 = n13799 & ~n14937;
  assign n14939 = n14938 ^ n13954;
  assign n14940 = n13825 & n14939;
  assign n15158 = n13941 & n13974;
  assign n15159 = n13983 ^ n13925;
  assign n15160 = ~n13930 & n15159;
  assign n15161 = ~n15158 & ~n15160;
  assign n15165 = n13932 ^ n13923;
  assign n15164 = n13966 ^ n13922;
  assign n15166 = n15165 ^ n15164;
  assign n15167 = n15165 ^ n13799;
  assign n15168 = ~n13930 & ~n15167;
  assign n15169 = n15168 ^ n13799;
  assign n15170 = n15166 & n15169;
  assign n15171 = n15170 ^ n15164;
  assign n15172 = n13986 & ~n15171;
  assign n15162 = n14168 ^ n13949;
  assign n15163 = ~n13799 & n15162;
  assign n15173 = n15172 ^ n15163;
  assign n15174 = ~n13930 & ~n15173;
  assign n15175 = n15174 ^ n15172;
  assign n15176 = n15161 & n15175;
  assign n15177 = n13969 ^ n13939;
  assign n15178 = n13825 & n15177;
  assign n15179 = n15178 ^ n13939;
  assign n15180 = n13930 & n15179;
  assign n15181 = n15176 & ~n15180;
  assign n15182 = ~n13973 & n15181;
  assign n15183 = ~n13937 & n15182;
  assign n15184 = ~n14940 & n15183;
  assign n15185 = ~n14160 & n15184;
  assign n15186 = n15185 ^ n12299;
  assign n15187 = n15186 ^ x571;
  assign n15188 = ~n15157 & n15187;
  assign n15192 = ~n12628 & n14113;
  assign n15198 = n12588 ^ n12568;
  assign n15199 = n15198 ^ n12597;
  assign n15200 = n15199 ^ n12629;
  assign n15201 = ~n11714 & ~n15200;
  assign n15202 = n15201 ^ n12629;
  assign n15194 = n12607 ^ n12580;
  assign n15193 = n12635 ^ n12566;
  assign n15195 = n15194 ^ n15193;
  assign n15196 = n11714 & ~n15195;
  assign n15197 = n15196 ^ n15193;
  assign n15203 = n15202 ^ n15197;
  assign n15204 = n11189 & ~n15203;
  assign n15205 = n15204 ^ n15197;
  assign n15206 = ~n15192 & ~n15205;
  assign n15207 = ~n12625 & n15206;
  assign n15208 = ~n14112 & n15207;
  assign n15209 = ~n14108 & n15208;
  assign n15210 = ~n15025 & n15209;
  assign n15211 = ~n14110 & n15210;
  assign n15212 = ~n12605 & n15211;
  assign n15213 = n15212 ^ n12356;
  assign n15214 = n15213 ^ x570;
  assign n15242 = n15241 ^ x569;
  assign n15243 = ~n15214 & ~n15242;
  assign n15257 = n15188 & n15243;
  assign n15189 = n15188 ^ n15157;
  assign n15256 = ~n15189 & n15243;
  assign n15258 = n15257 ^ n15256;
  assign n15190 = n15189 ^ n15187;
  assign n15191 = n15190 ^ n15157;
  assign n15255 = n15191 & n15243;
  assign n15259 = n15258 ^ n15255;
  assign n15260 = n15259 ^ n15243;
  assign n15936 = n15260 ^ n15257;
  assign n15937 = ~n15315 & n15936;
  assign n15244 = n15243 ^ n15214;
  assign n15245 = n15244 ^ n15242;
  assign n15246 = n15245 ^ n15214;
  assign n15250 = n15188 & ~n15246;
  assign n15938 = n15256 ^ n15250;
  assign n15939 = n15152 & n15938;
  assign n15284 = n15151 ^ n15129;
  assign n15265 = n15191 & ~n15245;
  assign n15248 = ~n15189 & ~n15246;
  assign n15266 = n15265 ^ n15248;
  assign n15263 = n15188 & ~n15244;
  assign n15269 = n15266 ^ n15263;
  assign n15270 = n15269 ^ n15188;
  assign n15267 = n15266 ^ n15257;
  assign n15268 = n15267 ^ n15250;
  assign n15271 = n15270 ^ n15268;
  assign n15943 = n15151 & n15271;
  assign n15247 = n15191 & ~n15246;
  assign n15249 = n15248 ^ n15247;
  assign n15251 = n15250 ^ n15249;
  assign n15252 = n15251 ^ n15246;
  assign n15940 = n15255 ^ n15252;
  assign n15941 = n15151 & ~n15940;
  assign n15942 = n15941 ^ n15252;
  assign n15944 = n15943 ^ n15942;
  assign n15945 = ~n15284 & ~n15944;
  assign n15946 = n15945 ^ n15942;
  assign n15153 = n15152 ^ n15151;
  assign n15154 = n15153 ^ n15129;
  assign n15275 = ~n15189 & ~n15244;
  assign n15261 = n15260 ^ n15190;
  assign n15253 = n15190 & ~n15244;
  assign n15254 = n15253 ^ n15252;
  assign n15262 = n15261 ^ n15254;
  assign n15291 = n15275 ^ n15262;
  assign n15947 = n15291 ^ n15253;
  assign n15948 = ~n15154 & ~n15947;
  assign n15276 = n15275 ^ n15253;
  assign n15273 = ~n15189 & ~n15245;
  assign n15274 = n15273 ^ n15265;
  assign n15277 = n15276 ^ n15274;
  assign n15278 = n15277 ^ n15242;
  assign n15264 = n15263 ^ n15262;
  assign n15272 = n15271 ^ n15264;
  assign n15279 = n15278 ^ n15272;
  assign n15949 = ~n15153 & ~n15279;
  assign n15954 = n15263 ^ n15249;
  assign n15955 = n15151 & n15954;
  assign n15956 = n15955 ^ n15954;
  assign n15953 = ~n15151 & n15249;
  assign n15957 = n15956 ^ n15953;
  assign n15950 = n15274 ^ n15252;
  assign n15951 = ~n15151 & ~n15950;
  assign n15952 = n15951 ^ n15252;
  assign n15958 = n15957 ^ n15952;
  assign n15959 = ~n15129 & ~n15958;
  assign n15960 = n15959 ^ n15952;
  assign n15961 = ~n15949 & n15960;
  assign n15282 = ~n15153 & n15257;
  assign n15281 = n15152 & ~n15279;
  assign n15283 = n15282 ^ n15281;
  assign n15966 = n15273 ^ n15253;
  assign n15967 = n15966 ^ n15259;
  assign n15968 = n15151 & n15967;
  assign n15969 = n15968 ^ n15966;
  assign n15962 = n15275 ^ n15269;
  assign n15963 = n15962 ^ n15291;
  assign n15964 = n15151 & ~n15963;
  assign n15965 = n15964 ^ n15291;
  assign n15970 = n15969 ^ n15965;
  assign n15971 = ~n15284 & ~n15970;
  assign n15972 = n15971 ^ n15965;
  assign n15973 = ~n15283 & n15972;
  assign n15974 = n15961 & n15973;
  assign n15975 = ~n15948 & n15974;
  assign n15976 = n15953 ^ n15250;
  assign n15977 = ~n15284 & n15976;
  assign n15978 = n15977 ^ n15250;
  assign n15979 = n15975 & ~n15978;
  assign n15980 = n15946 & n15979;
  assign n15981 = ~n15939 & n15980;
  assign n15982 = ~n15937 & n15981;
  assign n15983 = n15982 ^ n12450;
  assign n15984 = n15983 ^ x604;
  assign n15985 = ~n15935 & ~n15984;
  assign n15986 = n15985 ^ n15935;
  assign n15987 = n15934 & ~n15986;
  assign n15996 = n15925 ^ n15865;
  assign n15997 = n15985 ^ n15984;
  assign n15998 = n15897 ^ n15865;
  assign n15999 = ~n15997 & ~n15998;
  assign n16000 = n15996 & n15999;
  assign n15993 = n15898 & n15919;
  assign n15991 = n15922 ^ n15900;
  assign n15988 = n15898 ^ n15897;
  assign n15989 = ~n15917 & n15988;
  assign n15990 = n15989 ^ n15923;
  assign n15992 = n15991 ^ n15990;
  assign n15994 = n15993 ^ n15992;
  assign n15995 = ~n15986 & ~n15994;
  assign n16001 = n16000 ^ n15995;
  assign n16002 = n15984 ^ n15935;
  assign n16003 = n15934 ^ n15920;
  assign n16004 = n16003 ^ n15989;
  assign n16005 = n16004 ^ n15929;
  assign n16011 = n16005 ^ n15921;
  assign n16010 = n15898 & ~n15917;
  assign n16012 = n16011 ^ n16010;
  assign n16038 = n15984 & n16012;
  assign n16018 = n15897 & n15996;
  assign n16035 = n16018 ^ n15898;
  assign n16022 = n15992 ^ n15988;
  assign n16019 = n16018 ^ n16010;
  assign n16020 = n16019 ^ n15994;
  assign n16021 = n16020 ^ n15989;
  assign n16023 = n16022 ^ n16021;
  assign n16027 = n16023 ^ n16010;
  assign n16028 = n16027 ^ n16020;
  assign n16029 = n16028 ^ n15917;
  assign n16030 = n16029 ^ n16004;
  assign n16031 = n16030 ^ n15916;
  assign n16009 = n15928 ^ n15917;
  assign n16013 = n16012 ^ n16009;
  assign n16015 = n16013 ^ n15991;
  assign n16016 = n16015 ^ n16005;
  assign n16024 = n16023 ^ n16016;
  assign n16025 = n16024 ^ n15922;
  assign n16007 = n15934 ^ n15899;
  assign n16006 = n16005 ^ n15930;
  assign n16008 = n16007 ^ n16006;
  assign n16014 = n16013 ^ n16008;
  assign n16017 = n16016 ^ n16014;
  assign n16026 = n16025 ^ n16017;
  assign n16032 = n16031 ^ n16026;
  assign n16033 = n16032 ^ n15992;
  assign n16034 = n16033 ^ n16020;
  assign n16036 = n16035 ^ n16034;
  assign n16037 = n16036 ^ n16032;
  assign n16039 = n16038 ^ n16037;
  assign n16040 = n16002 & n16039;
  assign n16041 = n16040 ^ n16037;
  assign n16042 = ~n15997 & n16004;
  assign n16043 = ~n15984 & ~n16026;
  assign n16044 = n16043 ^ n16017;
  assign n16045 = n16044 ^ n15930;
  assign n16046 = ~n16002 & ~n16045;
  assign n16047 = n16046 ^ n15930;
  assign n16048 = ~n16042 & ~n16047;
  assign n16049 = ~n16041 & n16048;
  assign n16050 = n15984 & ~n16021;
  assign n16051 = n16050 ^ n15989;
  assign n16052 = ~n15935 & n16051;
  assign n16053 = n16049 & ~n16052;
  assign n16054 = ~n16001 & n16053;
  assign n16055 = n15997 ^ n15935;
  assign n16057 = n15989 & ~n16055;
  assign n16056 = n16023 & ~n16055;
  assign n16058 = n16057 ^ n16056;
  assign n16059 = n16054 & ~n16058;
  assign n16060 = ~n15987 & n16059;
  assign n16061 = n16060 ^ n13797;
  assign n17711 = n16061 ^ x676;
  assign n15280 = ~n15154 & ~n15279;
  assign n15321 = n15260 ^ n15248;
  assign n15302 = n15255 ^ n15250;
  assign n16139 = n15321 ^ n15302;
  assign n16140 = n16139 ^ n15271;
  assign n16141 = n16140 ^ n15271;
  assign n16142 = ~n15151 & n16141;
  assign n16143 = n16142 ^ n15271;
  assign n16144 = ~n15284 & n16143;
  assign n16145 = n16144 ^ n15271;
  assign n16147 = n15272 ^ n15256;
  assign n16148 = n16147 ^ n15249;
  assign n16146 = n15260 ^ n15258;
  assign n16149 = n16148 ^ n16146;
  assign n16150 = n15151 & ~n16149;
  assign n16151 = n16150 ^ n16146;
  assign n16152 = n16151 ^ n15947;
  assign n16153 = n15129 & ~n16152;
  assign n16154 = n16153 ^ n15947;
  assign n16155 = ~n16145 & n16154;
  assign n16156 = n15955 ^ n15263;
  assign n16157 = n15284 & n16156;
  assign n16158 = n16155 & ~n16157;
  assign n16159 = ~n15937 & n16158;
  assign n16160 = n15961 & n16159;
  assign n16161 = ~n15280 & n16160;
  assign n16162 = n16161 ^ n13824;
  assign n16802 = n16162 ^ x627;
  assign n15709 = n15708 ^ n15686;
  assign n15725 = n15724 ^ n15709;
  assign n15694 = n15693 ^ n15646;
  assign n15696 = n15695 ^ n15694;
  assign n15706 = n15705 ^ n15696;
  assign n15707 = n15706 ^ n15697;
  assign n15726 = n15725 ^ n15707;
  assign n15727 = n15608 & n15726;
  assign n15728 = n15727 ^ n15725;
  assign n15683 = n15682 ^ n15646;
  assign n15689 = n15688 ^ n15683;
  assign n15679 = n15678 ^ n15674;
  assign n15680 = n15646 & n15679;
  assign n15681 = n15680 ^ n15676;
  assign n15690 = n15689 ^ n15681;
  assign n15691 = ~n15608 & n15690;
  assign n15692 = n15691 ^ n15681;
  assign n15729 = n15728 ^ n15692;
  assign n15730 = n15607 & n15729;
  assign n15731 = n15730 ^ n15728;
  assign n15732 = n15731 ^ n13266;
  assign n16801 = n15732 ^ x622;
  assign n16803 = n16802 ^ n16801;
  assign n14751 = n12651 ^ x586;
  assign n14752 = n14150 ^ x591;
  assign n14767 = ~n14492 & n14499;
  assign n14768 = n14525 ^ n14506;
  assign n14769 = n14768 ^ n14532;
  assign n14770 = ~n14542 & ~n14769;
  assign n14771 = ~n14767 & ~n14770;
  assign n14772 = ~n14524 & n14541;
  assign n14774 = n14773 ^ n14507;
  assign n14775 = n14498 & ~n14774;
  assign n14777 = n14522 ^ n14515;
  assign n14778 = n14777 ^ n14487;
  assign n14779 = n14492 & n14778;
  assign n14780 = n14779 ^ n14487;
  assign n14781 = n14531 & n14780;
  assign n14782 = ~n14540 & ~n14781;
  assign n14783 = ~n14776 & n14782;
  assign n14784 = ~n14775 & n14783;
  assign n14785 = ~n14772 & n14784;
  assign n14786 = n14771 & n14785;
  assign n14787 = ~n14550 & n14786;
  assign n14788 = ~n14766 & n14787;
  assign n14789 = ~n14764 & n14788;
  assign n14790 = ~n14759 & n14789;
  assign n14791 = ~n14757 & n14790;
  assign n14792 = ~n14500 & n14791;
  assign n14793 = n14792 ^ n11744;
  assign n14794 = n14793 ^ x589;
  assign n14795 = n14303 ^ x590;
  assign n14799 = n14004 ^ x587;
  assign n14848 = ~n14795 & n14799;
  assign n14807 = n14610 ^ n13775;
  assign n14806 = n13789 ^ n13740;
  assign n14808 = n14807 ^ n14806;
  assign n14809 = ~n13645 & n14808;
  assign n14810 = n14809 ^ n14806;
  assign n14801 = n13746 ^ n13733;
  assign n14800 = n13768 ^ n13717;
  assign n14802 = n14801 ^ n14800;
  assign n14803 = n14802 ^ n14624;
  assign n14804 = n13646 & n14803;
  assign n14805 = n14804 ^ n14624;
  assign n14811 = n14810 ^ n14805;
  assign n14812 = n13763 & ~n14811;
  assign n14813 = n14812 ^ n14810;
  assign n14814 = n14607 & ~n14813;
  assign n14815 = ~n13757 & n14814;
  assign n14816 = ~n13751 & n14815;
  assign n14817 = n14816 ^ n11807;
  assign n14818 = n14817 ^ x588;
  assign n14847 = n14818 ^ n14799;
  assign n14849 = n14848 ^ n14847;
  assign n14850 = n14794 & ~n14849;
  assign n14859 = n14850 ^ n14847;
  assign n14819 = n14799 & n14818;
  assign n14860 = n14859 ^ n14819;
  assign n14796 = n14794 & n14795;
  assign n14797 = n14796 ^ n14795;
  assign n14820 = n14819 ^ n14799;
  assign n14828 = n14797 & n14820;
  assign n14844 = n14828 ^ n14820;
  assign n14833 = n14796 & n14819;
  assign n14840 = n14833 ^ n14819;
  assign n14798 = n14797 ^ n14794;
  assign n14837 = n14798 ^ n14795;
  assign n14838 = n14819 & n14837;
  assign n14836 = n14797 & n14819;
  assign n14839 = n14838 ^ n14836;
  assign n14841 = n14840 ^ n14839;
  assign n14824 = ~n14798 & n14799;
  assign n14842 = n14841 ^ n14824;
  assign n14835 = n14796 & n14820;
  assign n14843 = n14842 ^ n14835;
  assign n14845 = n14844 ^ n14843;
  assign n14857 = n14845 ^ n14833;
  assign n14821 = n14820 ^ n14818;
  assign n14822 = ~n14798 & ~n14821;
  assign n14858 = n14857 ^ n14822;
  assign n14861 = n14860 ^ n14858;
  assign n14855 = n14819 ^ n14818;
  assign n14868 = n14861 ^ n14855;
  assign n14864 = n14835 ^ n14796;
  assign n14826 = n14796 & ~n14821;
  assign n14834 = n14833 ^ n14826;
  assign n14865 = n14864 ^ n14834;
  assign n14823 = n14822 ^ n14798;
  assign n14825 = n14824 ^ n14823;
  assign n14827 = n14826 ^ n14825;
  assign n14866 = n14865 ^ n14827;
  assign n14856 = n14837 & n14855;
  assign n14862 = n14861 ^ n14856;
  assign n14863 = n14862 ^ n14826;
  assign n14867 = n14866 ^ n14863;
  assign n14869 = n14868 ^ n14867;
  assign n14846 = n14845 ^ n14834;
  assign n14851 = n14850 ^ n14846;
  assign n14870 = n14869 ^ n14851;
  assign n14871 = n14752 & ~n14870;
  assign n14872 = n14871 ^ n14869;
  assign n14873 = ~n14751 & ~n14872;
  assign n14874 = n14873 ^ n14872;
  assign n15382 = n14862 ^ n14858;
  assign n15383 = n14752 & ~n15382;
  assign n15384 = n15383 ^ n14858;
  assign n15385 = ~n14751 & n15384;
  assign n14852 = n14751 & n14752;
  assign n14853 = n14852 ^ n14751;
  assign n14880 = n14853 ^ n14752;
  assign n15386 = n14880 ^ n14751;
  assign n15387 = ~n14869 & n15386;
  assign n14899 = n14856 ^ n14842;
  assign n14900 = n14752 & n14899;
  assign n14901 = n14900 ^ n14856;
  assign n15388 = ~n14751 & n14901;
  assign n15389 = ~n15387 & ~n15388;
  assign n14876 = n14752 ^ n14751;
  assign n15390 = ~n14752 & ~n14862;
  assign n15391 = n15390 ^ n14856;
  assign n15392 = ~n14876 & n15391;
  assign n15393 = n14842 ^ n14825;
  assign n15394 = n14853 & ~n15393;
  assign n15395 = n14865 ^ n14822;
  assign n15396 = n14751 & n15395;
  assign n15397 = ~n15394 & ~n15396;
  assign n15405 = n14857 ^ n14839;
  assign n15400 = n14835 ^ n14825;
  assign n15401 = n15400 ^ n14841;
  assign n15398 = n14845 ^ n14835;
  assign n15399 = n15398 ^ n14836;
  assign n15402 = n15401 ^ n15399;
  assign n15403 = n14752 & ~n15402;
  assign n15404 = n15403 ^ n15399;
  assign n15406 = n15405 ^ n15404;
  assign n15407 = n15406 ^ n15404;
  assign n15408 = n14752 & n15407;
  assign n15409 = n15408 ^ n15404;
  assign n15410 = ~n14751 & n15409;
  assign n15411 = n15410 ^ n15404;
  assign n15412 = n15397 & ~n15411;
  assign n15413 = n14880 ^ n14828;
  assign n14885 = n14841 ^ n14826;
  assign n15414 = n14885 ^ n14852;
  assign n15415 = ~n14880 & ~n15414;
  assign n15416 = n15415 ^ n14852;
  assign n15417 = ~n15413 & ~n15416;
  assign n15418 = n15417 ^ n14828;
  assign n15419 = n15412 & ~n15418;
  assign n15420 = ~n15392 & n15419;
  assign n15421 = n15389 & n15420;
  assign n15422 = ~n15385 & n15421;
  assign n15423 = n14874 & n15422;
  assign n15424 = n15423 ^ n13189;
  assign n16804 = n15424 ^ x623;
  assign n16339 = n14008 ^ n13798;
  assign n16340 = n14054 ^ n14032;
  assign n16341 = n16340 ^ n14052;
  assign n16342 = n16339 & n16341;
  assign n16343 = n14030 ^ n14011;
  assign n16344 = n16343 ^ n14023;
  assign n16345 = n14005 & n16344;
  assign n16346 = n16345 ^ n14023;
  assign n16347 = n14006 & n16346;
  assign n16805 = n14043 ^ n14039;
  assign n16806 = n16805 ^ n14012;
  assign n16807 = ~n13798 & ~n16806;
  assign n16808 = n16807 ^ n14012;
  assign n16809 = ~n14005 & n16808;
  assign n16819 = ~n14042 & ~n16339;
  assign n16823 = n14039 & ~n16819;
  assign n16820 = n16819 ^ n13644;
  assign n16821 = n13798 & n16820;
  assign n16822 = n16821 ^ n13644;
  assign n16824 = n16823 ^ n16822;
  assign n16818 = n14008 & ~n14031;
  assign n16825 = n16824 ^ n16818;
  assign n16814 = n14040 ^ n13636;
  assign n16815 = n14020 & ~n16814;
  assign n16349 = ~n14020 & ~n14037;
  assign n16816 = n16815 ^ n16349;
  assign n16810 = n14037 ^ n13640;
  assign n16811 = n16810 ^ n14054;
  assign n16812 = ~n14021 & n16811;
  assign n16813 = n16812 ^ n14054;
  assign n16817 = n16816 ^ n16813;
  assign n16826 = n16825 ^ n16817;
  assign n16827 = ~n16809 & n16826;
  assign n16828 = ~n16347 & n16827;
  assign n16829 = ~n16342 & n16828;
  assign n16830 = n16829 ^ n13864;
  assign n16831 = n16830 ^ x624;
  assign n16832 = ~n16804 & ~n16831;
  assign n16869 = n16832 ^ n16831;
  assign n15020 = n14660 ^ x556;
  assign n15047 = n15046 ^ x561;
  assign n15048 = ~n15020 & ~n15047;
  assign n15051 = n15048 ^ n15047;
  assign n15068 = n15051 ^ n15020;
  assign n15078 = n15068 ^ n15048;
  assign n14936 = n14935 ^ x560;
  assign n14941 = n13966 ^ n13826;
  assign n14943 = n13959 ^ n13947;
  assign n14942 = n13891 ^ n13865;
  assign n14944 = n14943 ^ n14942;
  assign n14945 = n14944 ^ n13828;
  assign n14946 = ~n13966 & ~n14945;
  assign n14947 = n14946 ^ n13828;
  assign n14948 = n14941 & n14947;
  assign n14949 = n14948 ^ n13826;
  assign n14954 = n13961 ^ n13925;
  assign n14950 = n13968 ^ n13928;
  assign n14951 = n14950 ^ n13952;
  assign n14952 = n13825 & n14951;
  assign n14953 = n14952 ^ n14950;
  assign n14955 = n14954 ^ n14953;
  assign n14956 = n14955 ^ n14953;
  assign n14957 = n13825 & n14956;
  assign n14958 = n14957 ^ n14953;
  assign n14959 = n13930 & n14958;
  assign n14960 = n14959 ^ n14953;
  assign n14961 = ~n14949 & ~n14960;
  assign n14962 = ~n13976 & n14961;
  assign n14963 = ~n13945 & n14962;
  assign n14964 = ~n14153 & n14963;
  assign n14965 = ~n14940 & n14964;
  assign n14966 = ~n14160 & n14965;
  assign n14967 = ~n13929 & n14966;
  assign n14968 = n14967 ^ n12108;
  assign n14969 = n14968 ^ x559;
  assign n14970 = ~n14936 & ~n14969;
  assign n14971 = n14970 ^ n14936;
  assign n14972 = n14971 ^ n14969;
  assign n14976 = n13591 & n13613;
  assign n14977 = n14976 ^ n13590;
  assign n14973 = n13607 ^ n13604;
  assign n14974 = n13613 & n14973;
  assign n14975 = n14974 ^ n13604;
  assign n14978 = n14977 ^ n14975;
  assign n14979 = n13463 & ~n14978;
  assign n14980 = n14979 ^ n14977;
  assign n14981 = n14980 ^ n12045;
  assign n14982 = n14981 ^ x558;
  assign n14983 = n14576 ^ x557;
  assign n14984 = ~n14982 & n14983;
  assign n14985 = n14984 ^ n14982;
  assign n15007 = ~n14972 & ~n14985;
  assign n14986 = n14985 ^ n14983;
  assign n15012 = n15007 ^ n14986;
  assign n14996 = n14970 & n14986;
  assign n15010 = n15007 ^ n14996;
  assign n15003 = ~n14971 & ~n14985;
  assign n15004 = n15003 ^ n14971;
  assign n14989 = n14986 ^ n14982;
  assign n14999 = ~n14972 & n14989;
  assign n15000 = n14999 ^ n14989;
  assign n14993 = n14970 & n14984;
  assign n14992 = n14970 & ~n14985;
  assign n14994 = n14993 ^ n14992;
  assign n14995 = n14994 ^ n14970;
  assign n14997 = n14996 ^ n14995;
  assign n14990 = n14972 ^ n14936;
  assign n14991 = n14989 & ~n14990;
  assign n14998 = n14997 ^ n14991;
  assign n15001 = n15000 ^ n14998;
  assign n14988 = ~n14971 & n14984;
  assign n15002 = n15001 ^ n14988;
  assign n15005 = n15004 ^ n15002;
  assign n14987 = ~n14972 & n14986;
  assign n15006 = n15005 ^ n14987;
  assign n15011 = n15010 ^ n15006;
  assign n15013 = n15012 ^ n15011;
  assign n16094 = n15013 ^ n15005;
  assign n16095 = n16094 ^ n15001;
  assign n16096 = ~n15020 & n16095;
  assign n16097 = n16096 ^ n15001;
  assign n16098 = n15078 & n16097;
  assign n16099 = n14991 & n15078;
  assign n15014 = n15013 ^ n15003;
  assign n15015 = n15014 ^ n14996;
  assign n15016 = n15015 ^ n14983;
  assign n15008 = n15007 ^ n15006;
  assign n15009 = n15008 ^ n14992;
  assign n15017 = n15016 ^ n15009;
  assign n15018 = n15017 ^ n15003;
  assign n15019 = n15018 ^ n15001;
  assign n15049 = n15048 ^ n15020;
  assign n15050 = ~n15019 & ~n15049;
  assign n16100 = n14999 ^ n14988;
  assign n15058 = n15014 ^ n14990;
  assign n15057 = n15018 ^ n14991;
  assign n15059 = n15058 ^ n15057;
  assign n15080 = n15059 ^ n14997;
  assign n16101 = n16100 ^ n15080;
  assign n16102 = n15020 & ~n16101;
  assign n16103 = n16102 ^ n16100;
  assign n16104 = ~n15078 & n16103;
  assign n16105 = n15018 ^ n14987;
  assign n16106 = n16105 ^ n15007;
  assign n16107 = ~n15051 & ~n16106;
  assign n16108 = n14994 & n15078;
  assign n16109 = n16108 ^ n14992;
  assign n16110 = ~n16107 & ~n16109;
  assign n16112 = n15017 ^ n14996;
  assign n16111 = n15080 ^ n14987;
  assign n16113 = n16112 ^ n16111;
  assign n16114 = n16113 ^ n15001;
  assign n16115 = ~n15020 & n16114;
  assign n16116 = n16115 ^ n15001;
  assign n16117 = ~n15078 & n16116;
  assign n16118 = n16110 & ~n16117;
  assign n15055 = n14993 ^ n14991;
  assign n15056 = n15055 ^ n14988;
  assign n15060 = n15059 ^ n15056;
  assign n15061 = n15060 ^ n14984;
  assign n15062 = n15061 ^ n14991;
  assign n16119 = n15062 ^ n15010;
  assign n16120 = n15047 & ~n16119;
  assign n16121 = n16120 ^ n15062;
  assign n16122 = n15020 & ~n16121;
  assign n16123 = n16118 & ~n16122;
  assign n16124 = ~n16104 & n16123;
  assign n16125 = n15003 ^ n14987;
  assign n16126 = ~n15068 & n16125;
  assign n15063 = ~n15049 & ~n15062;
  assign n16127 = n16126 ^ n15063;
  assign n16128 = n16124 & ~n16127;
  assign n16129 = ~n15050 & n16128;
  assign n16130 = ~n16099 & n16129;
  assign n16131 = ~n16098 & n16130;
  assign n16132 = n16131 ^ n13914;
  assign n16834 = n16132 ^ x626;
  assign n16312 = n14374 ^ n14372;
  assign n16313 = n14344 & n16312;
  assign n16314 = n14370 ^ n14367;
  assign n16315 = n14342 & n16314;
  assign n16316 = n16315 ^ n14367;
  assign n16317 = ~n14304 & n16316;
  assign n16835 = n14379 ^ n14193;
  assign n16836 = n16835 ^ n15866;
  assign n16837 = n14343 & n16836;
  assign n16842 = n14343 & n14387;
  assign n14417 = n14344 & n14416;
  assign n16843 = n16842 ^ n14417;
  assign n16840 = n14343 & n14402;
  assign n16841 = n16840 ^ n15879;
  assign n16844 = n16843 ^ n16841;
  assign n16318 = n14415 ^ n14385;
  assign n16838 = n16318 ^ n14361;
  assign n16839 = ~n14342 & n16838;
  assign n16845 = n16844 ^ n16839;
  assign n16846 = ~n14304 & n16845;
  assign n16847 = n16846 ^ n16844;
  assign n16848 = ~n16837 & ~n16847;
  assign n16849 = n14378 ^ n14367;
  assign n16850 = ~n14304 & n16849;
  assign n16851 = n16850 ^ n14367;
  assign n16852 = n14342 & n16851;
  assign n16853 = n16848 & ~n16852;
  assign n16854 = ~n16317 & n16853;
  assign n16855 = ~n16313 & n16854;
  assign n16856 = ~n15878 & n16855;
  assign n16857 = ~n14345 & n16856;
  assign n16858 = n16857 ^ n13890;
  assign n16859 = n16858 ^ x625;
  assign n16860 = ~n16834 & n16859;
  assign n16881 = n16860 ^ n16834;
  assign n16893 = ~n16869 & ~n16881;
  assign n16861 = n16860 ^ n16859;
  assign n16873 = n16861 & ~n16869;
  assign n16894 = n16893 ^ n16873;
  assign n16870 = n16860 & ~n16869;
  assign n16833 = n16832 ^ n16804;
  assign n16867 = n16833 ^ n16831;
  assign n16868 = n16861 & ~n16867;
  assign n16871 = n16870 ^ n16868;
  assign n16895 = n16894 ^ n16871;
  assign n16896 = n16895 ^ n16804;
  assign n16888 = ~n16867 & ~n16881;
  assign n16889 = n16888 ^ n16867;
  assign n16886 = n16860 & ~n16867;
  assign n16887 = n16886 ^ n16868;
  assign n16890 = n16889 ^ n16887;
  assign n16891 = n16890 ^ n16886;
  assign n16892 = n16891 ^ n16888;
  assign n16897 = n16896 ^ n16892;
  assign n16882 = n16832 & ~n16881;
  assign n16898 = n16897 ^ n16882;
  assign n16899 = ~n16802 & ~n16898;
  assign n16900 = n16899 ^ n16897;
  assign n16866 = n16832 & n16861;
  assign n16883 = n16882 ^ n16866;
  assign n16879 = n16832 & n16860;
  assign n16880 = n16879 ^ n16832;
  assign n16884 = n16883 ^ n16880;
  assign n16874 = n16873 ^ n16870;
  assign n16875 = n16874 ^ n16861;
  assign n16872 = n16871 ^ n16866;
  assign n16876 = n16875 ^ n16872;
  assign n16877 = n16876 ^ n16833;
  assign n16864 = ~n16833 & n16860;
  assign n16862 = n16861 ^ n16834;
  assign n16863 = ~n16833 & n16862;
  assign n16865 = n16864 ^ n16863;
  assign n16878 = n16877 ^ n16865;
  assign n16885 = n16884 ^ n16878;
  assign n16901 = n16900 ^ n16885;
  assign n16902 = ~n16803 & n16901;
  assign n16903 = n16902 ^ n16885;
  assign n16904 = n16801 & n16802;
  assign n16905 = n16891 ^ n16864;
  assign n16906 = n16904 & ~n16905;
  assign n17433 = n16897 ^ n16888;
  assign n17434 = n17433 ^ n16890;
  assign n17435 = ~n16802 & n17434;
  assign n17436 = n17435 ^ n16890;
  assign n17437 = ~n16801 & ~n17436;
  assign n17712 = n16803 & n16879;
  assign n17713 = n16883 ^ n16876;
  assign n17714 = n16801 & n17713;
  assign n17715 = n17714 ^ n16876;
  assign n17716 = n16802 & n17715;
  assign n17717 = ~n17712 & ~n17716;
  assign n17719 = n16876 ^ n16871;
  assign n17718 = n16873 ^ n16863;
  assign n17720 = n17719 ^ n17718;
  assign n17721 = n16801 & n17720;
  assign n17722 = n17721 ^ n17718;
  assign n17723 = ~n16802 & n17722;
  assign n17724 = n16888 ^ n16868;
  assign n17725 = n17724 ^ n16893;
  assign n17726 = n17725 ^ n16893;
  assign n17727 = n16802 & n17726;
  assign n17728 = n17727 ^ n16893;
  assign n17729 = ~n16803 & n17728;
  assign n17730 = n17729 ^ n16893;
  assign n17731 = ~n17723 & ~n17730;
  assign n17733 = ~n16801 & n16886;
  assign n16914 = n16904 ^ n16801;
  assign n16915 = n16914 ^ n16802;
  assign n16916 = n16915 ^ n16801;
  assign n17732 = n16870 & n16916;
  assign n17734 = n17733 ^ n17732;
  assign n17735 = n17731 & ~n17734;
  assign n17736 = n17717 & n17735;
  assign n17737 = ~n17437 & n17736;
  assign n17738 = ~n16906 & n17737;
  assign n17739 = n16903 & n17738;
  assign n17740 = n16863 & n16914;
  assign n17439 = n16878 ^ n16876;
  assign n17440 = ~n16915 & ~n17439;
  assign n17741 = n17740 ^ n17440;
  assign n17742 = n17739 & ~n17741;
  assign n17743 = n17742 ^ n14004;
  assign n17744 = n17743 ^ x681;
  assign n17746 = n17711 & ~n17744;
  assign n17745 = n17744 ^ n17711;
  assign n17747 = n17746 ^ n17745;
  assign n14389 = ~n14366 & n14388;
  assign n14390 = n14378 ^ n14361;
  assign n14391 = n14343 & n14390;
  assign n14392 = n14376 ^ n14369;
  assign n14393 = n14392 ^ n14379;
  assign n14394 = n14344 & n14393;
  assign n14395 = n14366 & ~n14394;
  assign n14396 = ~n14344 & ~n14367;
  assign n14397 = ~n14380 & n14396;
  assign n14398 = ~n14395 & ~n14397;
  assign n14399 = ~n14391 & ~n14398;
  assign n14406 = n14405 ^ n14375;
  assign n14407 = n14342 & n14406;
  assign n14408 = n14407 ^ n14387;
  assign n14409 = ~n14304 & n14408;
  assign n14410 = n14409 ^ n14387;
  assign n14411 = n14399 & ~n14410;
  assign n14413 = n14412 ^ n14361;
  assign n14414 = ~n14366 & n14413;
  assign n14418 = n14417 ^ n14414;
  assign n14419 = n14411 & ~n14418;
  assign n14420 = ~n14389 & n14419;
  assign n14421 = ~n14365 & n14420;
  assign n14422 = ~n14345 & n14421;
  assign n14423 = n14422 ^ n13256;
  assign n14424 = n14423 ^ x615;
  assign n14067 = n14066 ^ x610;
  assign n14425 = n14424 ^ n14067;
  assign n15052 = n15017 ^ n14992;
  assign n15053 = ~n15051 & ~n15052;
  assign n15054 = ~n15011 & n15048;
  assign n15064 = n14999 & ~n15051;
  assign n15065 = n15048 & ~n15060;
  assign n15066 = n15056 ^ n14997;
  assign n15067 = n15066 ^ n15009;
  assign n15069 = n15068 ^ n15009;
  assign n15070 = n15009 & ~n15069;
  assign n15071 = n15070 ^ n15009;
  assign n15072 = ~n15067 & n15071;
  assign n15073 = n15072 ^ n15070;
  assign n15074 = n15073 ^ n15009;
  assign n15075 = n15074 ^ n15068;
  assign n15076 = ~n15065 & ~n15075;
  assign n15077 = n15076 ^ n15065;
  assign n15081 = n15080 ^ n14999;
  assign n15079 = n15062 ^ n14998;
  assign n15082 = n15081 ^ n15079;
  assign n15083 = ~n15020 & n15082;
  assign n15084 = n15083 ^ n15079;
  assign n15085 = n15078 & ~n15084;
  assign n15086 = ~n15077 & ~n15085;
  assign n15087 = ~n15064 & n15086;
  assign n15088 = ~n15063 & n15087;
  assign n15089 = ~n15054 & n15088;
  assign n15090 = ~n15015 & n15020;
  assign n15091 = n15090 ^ n14996;
  assign n15092 = n15078 & n15091;
  assign n15093 = n15089 & ~n15092;
  assign n15094 = ~n15053 & n15093;
  assign n15095 = ~n15050 & n15094;
  assign n15096 = n15095 ^ n13217;
  assign n15097 = n15096 ^ x614;
  assign n14829 = n14828 ^ n14827;
  assign n14830 = ~n14752 & ~n14829;
  assign n14831 = n14830 ^ n14828;
  assign n14832 = ~n14751 & n14831;
  assign n14854 = n14851 & n14853;
  assign n14875 = n14874 ^ n14854;
  assign n14877 = n14865 & ~n14876;
  assign n14886 = n14885 ^ n14838;
  assign n14887 = n14886 ^ n14869;
  assign n14888 = n14887 ^ n14818;
  assign n14881 = n14824 ^ n14799;
  assign n14882 = ~n14880 & ~n14881;
  assign n14878 = n14843 ^ n14838;
  assign n14879 = n14878 ^ n14833;
  assign n14883 = n14882 ^ n14879;
  assign n14884 = n14883 ^ n14751;
  assign n14889 = n14888 ^ n14884;
  assign n14890 = n14889 ^ n14884;
  assign n14891 = ~n14751 & ~n14890;
  assign n14892 = n14891 ^ n14884;
  assign n14893 = n14752 & ~n14892;
  assign n14894 = n14893 ^ n14884;
  assign n14895 = ~n14877 & n14894;
  assign n14896 = n14859 ^ n14827;
  assign n14897 = n14752 & n14896;
  assign n14898 = n14897 ^ n14827;
  assign n14902 = n14901 ^ n14898;
  assign n14903 = n14751 & ~n14902;
  assign n14904 = n14903 ^ n14901;
  assign n14905 = n14895 & ~n14904;
  assign n14906 = n14875 & n14905;
  assign n14907 = ~n14832 & n14906;
  assign n14908 = n14907 ^ n13562;
  assign n14909 = n14908 ^ x613;
  assign n15343 = n15097 ^ n14909;
  assign n15287 = ~n15151 & n15247;
  assign n15285 = n15151 & ~n15254;
  assign n15286 = n15285 ^ n15252;
  assign n15288 = n15287 ^ n15286;
  assign n15289 = n15284 & ~n15288;
  assign n15290 = n15289 ^ n15286;
  assign n15297 = ~n15151 & n15277;
  assign n15292 = n15291 ^ n15263;
  assign n15293 = n15292 ^ n15265;
  assign n15294 = n15293 ^ n15278;
  assign n15295 = n15151 & ~n15294;
  assign n15296 = n15295 ^ n15293;
  assign n15298 = n15297 ^ n15296;
  assign n15299 = ~n15284 & ~n15298;
  assign n15300 = n15299 ^ n15296;
  assign n15303 = n15302 ^ n15256;
  assign n15304 = n15303 ^ n15247;
  assign n15301 = n15273 ^ n15252;
  assign n15305 = n15304 ^ n15301;
  assign n15306 = n15301 ^ n15154;
  assign n15307 = n15301 & ~n15306;
  assign n15308 = n15307 ^ n15301;
  assign n15309 = ~n15305 & n15308;
  assign n15310 = n15309 ^ n15307;
  assign n15311 = n15310 ^ n15301;
  assign n15312 = n15311 ^ n15154;
  assign n15313 = n15300 & ~n15312;
  assign n15314 = n15313 ^ n15300;
  assign n15317 = ~n15129 & n15250;
  assign n15316 = n15256 & ~n15315;
  assign n15318 = n15317 ^ n15316;
  assign n15319 = n15314 & ~n15318;
  assign n15320 = ~n15151 & n15255;
  assign n15322 = n15321 ^ n15320;
  assign n15323 = ~n15284 & n15322;
  assign n15324 = n15323 ^ n15321;
  assign n15325 = n15319 & ~n15324;
  assign n15326 = n15290 & n15325;
  assign n15327 = ~n15283 & n15326;
  assign n15328 = ~n15280 & n15327;
  assign n15329 = n15328 ^ n13529;
  assign n15330 = n15329 ^ x612;
  assign n15344 = n15343 ^ n15330;
  assign n14750 = n14749 ^ x611;
  assign n15338 = n14909 ^ n14750;
  assign n15331 = n15330 ^ n14909;
  assign n15332 = n14750 & ~n15331;
  assign n15341 = n15338 ^ n15332;
  assign n15339 = n15338 ^ n15330;
  assign n15333 = n15332 ^ n15330;
  assign n15336 = n15097 ^ n14750;
  assign n15337 = n15333 & n15336;
  assign n15340 = n15339 ^ n15337;
  assign n15342 = n15341 ^ n15340;
  assign n15345 = n15344 ^ n15342;
  assign n15098 = n14909 & n15097;
  assign n15099 = ~n14750 & n15098;
  assign n15334 = n15333 ^ n15099;
  assign n15335 = n15334 ^ n15097;
  assign n15346 = n15345 ^ n15335;
  assign n17751 = n14067 & n15346;
  assign n17752 = n17751 ^ n15345;
  assign n15353 = n15330 & ~n15338;
  assign n15369 = ~n15097 & n15353;
  assign n15370 = n15369 ^ n15342;
  assign n15362 = n15336 ^ n15330;
  assign n15363 = ~n15330 & ~n15343;
  assign n15364 = n15363 ^ n15097;
  assign n15365 = ~n15362 & n15364;
  assign n15366 = n15365 ^ n15097;
  assign n15349 = n15330 ^ n15097;
  assign n15358 = n15349 ^ n15098;
  assign n15352 = n14909 & n15330;
  assign n15359 = n15358 ^ n15352;
  assign n15356 = ~n15349 & n15352;
  assign n15357 = n15356 ^ n15344;
  assign n15360 = n15359 ^ n15357;
  assign n15354 = n15353 ^ n15352;
  assign n15355 = n15354 ^ n15342;
  assign n15361 = n15360 ^ n15355;
  assign n15367 = n15366 ^ n15361;
  assign n15371 = n15370 ^ n15367;
  assign n15372 = n15371 ^ n15362;
  assign n17748 = n15372 ^ n14424;
  assign n15350 = ~n14750 & ~n15349;
  assign n15351 = n15350 ^ n15335;
  assign n15368 = n15367 ^ n15351;
  assign n15373 = n15372 ^ n15368;
  assign n15374 = n14424 & n15373;
  assign n15375 = n15374 ^ n15368;
  assign n17749 = n17748 ^ n15375;
  assign n17750 = n17749 ^ n15368;
  assign n17753 = n17752 ^ n17750;
  assign n17754 = ~n14425 & n17753;
  assign n17755 = n17754 ^ n17750;
  assign n17756 = n17755 ^ n13630;
  assign n17757 = n17756 ^ x678;
  assign n16451 = n15608 ^ n15607;
  assign n16455 = ~n15607 & ~n15705;
  assign n16456 = n16455 ^ n15704;
  assign n16452 = n15907 ^ n15723;
  assign n16453 = ~n15607 & n16452;
  assign n16454 = n16453 ^ n15907;
  assign n16457 = n16456 ^ n16454;
  assign n16458 = n16451 & ~n16457;
  assign n16459 = n16458 ^ n16456;
  assign n16460 = ~n15717 & n16459;
  assign n16461 = n16460 ^ n12931;
  assign n16462 = n16461 ^ x639;
  assign n16165 = n14426 & n14670;
  assign n16166 = n14679 & n14697;
  assign n15432 = n14697 ^ n14577;
  assign n16167 = n15432 ^ n14426;
  assign n16168 = n14673 & n16167;
  assign n15428 = n14707 ^ n14666;
  assign n15429 = ~n14426 & n15428;
  assign n15430 = n15429 ^ n14666;
  assign n15431 = ~n14704 & n15430;
  assign n16169 = n16168 ^ n15431;
  assign n16170 = ~n14704 & n14726;
  assign n16171 = n14719 ^ n14698;
  assign n16172 = ~n15432 & n16171;
  assign n16173 = ~n16170 & ~n16172;
  assign n16176 = n14577 & n14677;
  assign n16174 = n14696 & n14707;
  assign n15433 = n14722 ^ n14699;
  assign n16175 = n16174 ^ n15433;
  assign n16177 = n16176 ^ n16175;
  assign n16178 = ~n14426 & n16177;
  assign n16179 = n16178 ^ n16175;
  assign n16180 = n16173 & ~n16179;
  assign n16181 = ~n14703 & n16180;
  assign n16182 = ~n16169 & n16181;
  assign n16183 = ~n16166 & n16182;
  assign n16184 = ~n16165 & n16183;
  assign n16185 = n14719 ^ n14667;
  assign n16186 = n16185 ^ n14701;
  assign n16187 = ~n14426 & ~n16186;
  assign n16188 = n16187 ^ n14701;
  assign n16189 = n14577 & ~n16188;
  assign n16190 = n16184 & ~n16189;
  assign n16191 = ~n14692 & n16190;
  assign n16192 = n16191 ^ n13073;
  assign n16463 = n16192 ^ x634;
  assign n16464 = ~n16462 & n16463;
  assign n16465 = n16464 ^ n16463;
  assign n16319 = n15872 & n16318;
  assign n16320 = n14368 ^ n14361;
  assign n16321 = n14304 & n16320;
  assign n16322 = n14403 ^ n14379;
  assign n16323 = n14344 & n16322;
  assign n16324 = ~n16321 & ~n16323;
  assign n16325 = ~n16319 & n16324;
  assign n16326 = n14384 ^ n14374;
  assign n16327 = n16326 ^ n15879;
  assign n16328 = n16327 ^ n14416;
  assign n16329 = n14304 & n16328;
  assign n16330 = n16329 ^ n14416;
  assign n16331 = ~n14342 & n16330;
  assign n16332 = n16325 & ~n16331;
  assign n16333 = ~n16317 & n16332;
  assign n16334 = ~n16313 & n16333;
  assign n16335 = ~n14389 & n16334;
  assign n16336 = n15871 & n16335;
  assign n16337 = n16336 ^ n12767;
  assign n16338 = n16337 ^ x637;
  assign n16348 = n16339 ^ n14037;
  assign n16350 = n16349 ^ n13637;
  assign n16351 = n16350 ^ n14020;
  assign n16352 = n16348 & n16351;
  assign n16353 = n16352 ^ n16339;
  assign n16354 = n13798 & n14027;
  assign n16355 = n14052 ^ n14011;
  assign n16356 = n14008 & ~n16355;
  assign n16357 = ~n16354 & ~n16356;
  assign n16363 = ~n14005 & n14056;
  assign n16359 = n14043 ^ n14023;
  assign n16358 = n14042 ^ n14030;
  assign n16360 = n16359 ^ n16358;
  assign n16361 = n14005 & ~n16360;
  assign n16362 = n16361 ^ n16358;
  assign n16364 = n16363 ^ n16362;
  assign n16365 = ~n14006 & n16364;
  assign n16366 = n16365 ^ n16362;
  assign n16367 = n16357 & ~n16366;
  assign n16368 = ~n14019 & n16367;
  assign n16369 = ~n16353 & n16368;
  assign n16370 = ~n16347 & n16369;
  assign n16371 = ~n16342 & n16370;
  assign n16372 = n16371 ^ n12807;
  assign n16373 = n16372 ^ x638;
  assign n16374 = ~n16338 & ~n16373;
  assign n16375 = ~n15078 & n16094;
  assign n16376 = n16375 ^ n16104;
  assign n16384 = n16113 ^ n16100;
  assign n16385 = ~n15047 & n16384;
  assign n16386 = n16385 ^ n16100;
  assign n16387 = n16121 & ~n16386;
  assign n16380 = n15057 ^ n14996;
  assign n16377 = n15001 ^ n14992;
  assign n16378 = n16377 ^ n15059;
  assign n16379 = n16378 ^ n15010;
  assign n16381 = n16380 ^ n16379;
  assign n16382 = ~n15047 & n16381;
  assign n16383 = n16382 ^ n16379;
  assign n16388 = n16387 ^ n16383;
  assign n16389 = n15020 & n16388;
  assign n16390 = n16389 ^ n16383;
  assign n16391 = ~n16098 & n16390;
  assign n16392 = ~n16376 & n16391;
  assign n16393 = ~n15064 & n16392;
  assign n16394 = ~n15063 & n16393;
  assign n16395 = n16394 ^ n12689;
  assign n16396 = n16395 ^ x636;
  assign n15574 = n15544 & n15573;
  assign n15541 = ~n15539 & n15540;
  assign n15551 = ~n15531 & ~n15550;
  assign n15553 = n15552 ^ n15551;
  assign n15554 = ~n15544 & n15553;
  assign n15555 = n15554 ^ n15552;
  assign n15556 = ~n15541 & ~n15555;
  assign n15575 = n15574 ^ n15556;
  assign n16066 = ~n15531 & n15580;
  assign n16063 = n15550 ^ n15535;
  assign n16064 = n15531 & ~n16063;
  assign n16065 = n16064 ^ n15535;
  assign n16067 = n16066 ^ n16065;
  assign n16068 = ~n15530 & n16067;
  assign n16069 = n16068 ^ n16065;
  assign n16070 = n15539 & n15838;
  assign n16071 = n16070 ^ n15542;
  assign n16073 = n15549 ^ n15535;
  assign n16074 = n16073 ^ n15528;
  assign n16075 = n15543 & n16074;
  assign n16072 = n15561 ^ n15559;
  assign n16076 = n16075 ^ n16072;
  assign n16077 = ~n16070 & ~n16076;
  assign n16078 = n16077 ^ n16072;
  assign n16079 = n16071 & ~n16078;
  assign n16080 = n16079 ^ n15542;
  assign n16081 = n15565 ^ n15525;
  assign n16082 = n16081 ^ n15557;
  assign n16083 = n16082 ^ n15571;
  assign n16084 = n15531 & n16083;
  assign n16085 = n16084 ^ n15571;
  assign n16086 = n15530 & n16085;
  assign n16087 = n16080 & ~n16086;
  assign n16088 = ~n16069 & n16087;
  assign n16089 = ~n15829 & n16088;
  assign n16090 = n15575 & n16089;
  assign n16091 = ~n15533 & n16090;
  assign n16092 = n16091 ^ n12720;
  assign n16397 = n16092 ^ x635;
  assign n16398 = ~n16396 & ~n16397;
  assign n16415 = n16374 & n16398;
  assign n16399 = n16398 ^ n16397;
  assign n16401 = n16374 ^ n16338;
  assign n16409 = ~n16399 & ~n16401;
  assign n16468 = n16415 ^ n16409;
  assign n16469 = n16465 & n16468;
  assign n16477 = n16463 ^ n16462;
  assign n16404 = n16374 ^ n16373;
  assign n16408 = ~n16399 & ~n16404;
  assign n16402 = n16398 & ~n16401;
  assign n17758 = n16408 ^ n16402;
  assign n17759 = ~n16477 & n17758;
  assign n16418 = n16399 ^ n16396;
  assign n16419 = ~n16404 & ~n16418;
  assign n16448 = n16419 ^ n16397;
  assign n16423 = n16418 ^ n16397;
  assign n16441 = ~n16401 & ~n16423;
  assign n16424 = n16374 & ~n16423;
  assign n16422 = ~n16401 & ~n16418;
  assign n16425 = n16424 ^ n16422;
  assign n16446 = n16441 ^ n16425;
  assign n16400 = n16374 & ~n16399;
  assign n16411 = n16400 ^ n16399;
  assign n16442 = n16441 ^ n16411;
  assign n16416 = n16415 ^ n16398;
  assign n16405 = n16404 ^ n16338;
  assign n16406 = n16398 & ~n16405;
  assign n16414 = n16406 ^ n16402;
  assign n16417 = n16416 ^ n16414;
  assign n16420 = n16419 ^ n16417;
  assign n16437 = n16420 ^ n16409;
  assign n16428 = n16396 ^ n16373;
  assign n16429 = n16428 ^ n16397;
  assign n16430 = n16429 ^ n16338;
  assign n16410 = n16409 ^ n16408;
  assign n16412 = n16411 ^ n16410;
  assign n16413 = n16412 ^ n16406;
  assign n16421 = n16420 ^ n16413;
  assign n16426 = n16425 ^ n16421;
  assign n16403 = n16402 ^ n16400;
  assign n16407 = n16406 ^ n16403;
  assign n16427 = n16426 ^ n16407;
  assign n16431 = n16430 ^ n16427;
  assign n16436 = n16431 ^ n16410;
  assign n16438 = n16437 ^ n16436;
  assign n16439 = n16438 ^ n16429;
  assign n16440 = n16439 ^ n16415;
  assign n16443 = n16442 ^ n16440;
  assign n16434 = n16419 ^ n16405;
  assign n16432 = n16431 ^ n16419;
  assign n16433 = n16432 ^ n16413;
  assign n16435 = n16434 ^ n16433;
  assign n16444 = n16443 ^ n16435;
  assign n16445 = n16444 ^ n16431;
  assign n16447 = n16446 ^ n16445;
  assign n16449 = n16448 ^ n16447;
  assign n16476 = ~n16449 & n16464;
  assign n16478 = n16435 ^ n16400;
  assign n16479 = ~n16463 & ~n16478;
  assign n16480 = n16479 ^ n16435;
  assign n16481 = n16477 & ~n16480;
  assign n17760 = n16425 & n16464;
  assign n17366 = n16444 ^ n16406;
  assign n17767 = n17366 ^ n16432;
  assign n17768 = n17767 ^ n16468;
  assign n17769 = ~n16463 & ~n17768;
  assign n17761 = n16463 ^ n16446;
  assign n17762 = n16477 & n17761;
  assign n17763 = n17762 ^ n16463;
  assign n17764 = ~n16447 & ~n17763;
  assign n17765 = n17764 ^ n16445;
  assign n17766 = n16449 & n17765;
  assign n17770 = n17769 ^ n17766;
  assign n17771 = n16477 & ~n17770;
  assign n17772 = n17771 ^ n17766;
  assign n17773 = ~n17760 & n17772;
  assign n17774 = ~n16481 & n17773;
  assign n17775 = ~n16476 & n17774;
  assign n17776 = ~n17759 & n17775;
  assign n17503 = n16413 ^ n16403;
  assign n16473 = n16417 ^ n16412;
  assign n17777 = n17503 ^ n16473;
  assign n17778 = n16463 & n17777;
  assign n17779 = n17778 ^ n16473;
  assign n17780 = ~n16462 & ~n17779;
  assign n17781 = n17776 & ~n17780;
  assign n17782 = ~n16469 & n17781;
  assign n17783 = n17782 ^ n13155;
  assign n17784 = n17783 ^ x679;
  assign n17785 = n17757 & n17784;
  assign n17786 = n17785 ^ n17757;
  assign n17787 = n17786 ^ n17784;
  assign n17821 = n17787 ^ n17757;
  assign n15381 = n15096 ^ x616;
  assign n15425 = n15424 ^ x621;
  assign n15426 = n15381 & n15425;
  assign n15427 = n15426 ^ n15381;
  assign n15434 = ~n15432 & n15433;
  assign n15435 = n14698 ^ n14687;
  assign n15436 = n15435 ^ n14722;
  assign n15437 = n14697 & n15436;
  assign n15439 = n14683 ^ n14670;
  assign n15438 = n14728 ^ n14675;
  assign n15440 = n15439 ^ n15438;
  assign n15441 = n14426 & n15440;
  assign n15442 = n15441 ^ n15438;
  assign n15443 = n14577 & n15442;
  assign n15450 = ~n14577 & n14682;
  assign n15446 = n14683 ^ n14671;
  assign n15444 = n14720 ^ n14701;
  assign n15445 = n15444 ^ n14664;
  assign n15447 = n15446 ^ n15445;
  assign n15448 = n14426 & ~n15447;
  assign n15449 = n15448 ^ n15445;
  assign n15451 = n15450 ^ n15449;
  assign n15452 = ~n14704 & ~n15451;
  assign n15453 = n15452 ^ n15449;
  assign n15454 = ~n15443 & n15453;
  assign n15455 = ~n15437 & n15454;
  assign n15456 = ~n15434 & n15455;
  assign n15458 = ~n14701 & ~n14704;
  assign n15457 = n14696 & n14720;
  assign n15459 = n15458 ^ n15457;
  assign n15460 = n15456 & ~n15459;
  assign n15461 = ~n15431 & n15460;
  assign n15462 = n15461 ^ n13302;
  assign n15463 = n15462 ^ x618;
  assign n15588 = n15531 & n15557;
  assign n15593 = n15571 ^ n15565;
  assign n15591 = n15559 ^ n15537;
  assign n15592 = n15591 ^ n15529;
  assign n15594 = n15593 ^ n15592;
  assign n15595 = ~n15531 & n15594;
  assign n15596 = n15595 ^ n15592;
  assign n15589 = n15531 & ~n15583;
  assign n15590 = n15589 ^ n15579;
  assign n15597 = n15596 ^ n15590;
  assign n15598 = ~n15530 & ~n15597;
  assign n15599 = n15598 ^ n15590;
  assign n15600 = ~n15588 & n15599;
  assign n15601 = ~n15587 & n15600;
  assign n15602 = ~n15578 & n15601;
  assign n15603 = n15575 & n15602;
  assign n15604 = ~n15533 & n15603;
  assign n15605 = n15604 ^ n13342;
  assign n15606 = n15605 ^ x619;
  assign n15733 = n15732 ^ x620;
  assign n15734 = n14423 ^ x617;
  assign n15735 = n15733 & n15734;
  assign n15736 = n15735 ^ n15734;
  assign n15737 = n15736 ^ n15733;
  assign n15738 = ~n15606 & ~n15737;
  assign n15739 = ~n15463 & n15738;
  assign n15740 = n15739 ^ n15738;
  assign n15741 = n15427 & n15740;
  assign n15742 = n15463 & ~n15606;
  assign n15747 = n15742 ^ n15606;
  assign n15748 = n15747 ^ n15463;
  assign n15750 = n15735 & n15748;
  assign n15749 = n15736 & n15748;
  assign n15751 = n15750 ^ n15749;
  assign n15752 = n15751 ^ n15748;
  assign n15743 = n15742 ^ n15463;
  assign n15744 = ~n15737 & n15743;
  assign n15745 = n15744 ^ n15738;
  assign n15746 = n15745 ^ n15737;
  assign n15753 = n15752 ^ n15746;
  assign n15754 = n15753 ^ n15751;
  assign n15755 = ~n15425 & ~n15754;
  assign n15756 = n15755 ^ n15753;
  assign n15757 = n15381 & ~n15756;
  assign n15765 = n15753 ^ n15739;
  assign n15762 = n15606 & ~n15734;
  assign n15758 = n15735 ^ n15733;
  assign n15763 = n15762 ^ n15758;
  assign n15759 = n15742 & n15758;
  assign n15760 = n15759 ^ n15744;
  assign n15761 = n15760 ^ n15746;
  assign n15764 = n15763 ^ n15761;
  assign n15766 = n15765 ^ n15764;
  assign n15767 = ~n15381 & n15766;
  assign n15768 = n15767 ^ n15764;
  assign n15769 = ~n15425 & ~n15768;
  assign n15771 = n15759 ^ n15758;
  assign n15770 = n15764 ^ n15753;
  assign n15772 = n15771 ^ n15770;
  assign n15773 = n15426 ^ n15425;
  assign n15774 = n15772 & n15773;
  assign n15775 = n15425 ^ n15381;
  assign n15781 = n15735 & n15742;
  assign n15789 = n15781 ^ n15734;
  assign n15786 = n15735 & ~n15747;
  assign n15777 = n15736 & n15742;
  assign n15776 = n15736 & ~n15747;
  assign n15778 = n15777 ^ n15776;
  assign n15779 = n15778 ^ n15749;
  assign n15787 = n15786 ^ n15779;
  assign n15780 = n15779 ^ n15736;
  assign n15785 = n15780 ^ n15750;
  assign n15788 = n15787 ^ n15785;
  assign n15790 = n15789 ^ n15788;
  assign n15797 = n15790 ^ n15776;
  assign n15798 = n15797 ^ n15786;
  assign n15799 = n15798 ^ n15761;
  assign n15791 = n15790 ^ n15739;
  assign n15784 = n15777 ^ n15751;
  assign n15792 = n15791 ^ n15784;
  assign n15793 = n15792 ^ n15760;
  assign n15782 = n15781 ^ n15780;
  assign n15783 = n15782 ^ n15778;
  assign n15794 = n15793 ^ n15783;
  assign n15795 = n15425 & n15794;
  assign n15796 = n15795 ^ n15783;
  assign n15800 = n15799 ^ n15796;
  assign n15801 = n15800 ^ n15796;
  assign n15802 = n15425 & ~n15801;
  assign n15803 = n15802 ^ n15796;
  assign n15804 = n15775 & n15803;
  assign n15805 = n15804 ^ n15796;
  assign n15806 = n15797 ^ n15744;
  assign n15807 = n15806 ^ n15786;
  assign n15808 = n15381 & n15807;
  assign n15809 = n15808 ^ n15786;
  assign n15810 = ~n15425 & n15809;
  assign n15811 = ~n15805 & ~n15810;
  assign n15812 = ~n15774 & n15811;
  assign n15813 = ~n15769 & n15812;
  assign n15816 = ~n15381 & n15777;
  assign n15814 = n15381 & n15752;
  assign n15815 = n15814 ^ n15746;
  assign n15817 = n15816 ^ n15815;
  assign n15818 = n15425 & ~n15817;
  assign n15819 = n15818 ^ n15815;
  assign n15820 = n15813 & n15819;
  assign n15821 = ~n15757 & n15820;
  assign n15822 = ~n15741 & n15821;
  assign n15823 = n15822 ^ n13444;
  assign n17788 = n15823 ^ x677;
  assign n16942 = n15896 ^ x603;
  assign n16572 = n15543 & n15561;
  assign n16573 = ~n15542 & ~n15569;
  assign n16577 = n15580 ^ n15535;
  assign n16578 = n16577 ^ n15548;
  assign n16574 = ~n15532 & n15545;
  assign n16575 = n16574 ^ n15837;
  assign n16579 = n16578 ^ n16575;
  assign n16580 = n16579 ^ n16575;
  assign n16581 = n15531 & ~n16580;
  assign n16582 = n16581 ^ n16575;
  assign n16583 = ~n15544 & ~n16582;
  assign n16576 = n16575 ^ n15530;
  assign n16584 = n16583 ^ n16576;
  assign n16586 = n15531 & ~n15585;
  assign n16585 = n15528 & n15544;
  assign n16587 = n16586 ^ n16585;
  assign n16588 = n16584 & ~n16587;
  assign n16589 = ~n16573 & n16588;
  assign n16590 = ~n16572 & n16589;
  assign n16591 = n15559 ^ n15532;
  assign n16592 = n15557 ^ n15543;
  assign n16593 = ~n15559 & ~n16592;
  assign n16594 = n16593 ^ n15543;
  assign n16595 = n16591 & n16594;
  assign n16596 = n16595 ^ n15532;
  assign n16597 = n16590 & ~n16596;
  assign n16598 = ~n15833 & n16597;
  assign n16599 = ~n16069 & n16598;
  assign n16600 = n15556 & n16599;
  assign n16601 = n16600 ^ n11713;
  assign n16943 = n16601 ^ x598;
  assign n16944 = n16942 & n16943;
  assign n16945 = n16944 ^ n16942;
  assign n16194 = n14838 ^ n14828;
  assign n16195 = n14852 & n16194;
  assign n16196 = n14865 ^ n14839;
  assign n16197 = n15386 & n16196;
  assign n16517 = n15386 & ~n15400;
  assign n16518 = n14858 ^ n14835;
  assign n16519 = n16518 ^ n14834;
  assign n16520 = n16519 ^ n14834;
  assign n16521 = ~n14752 & n16520;
  assign n16522 = n16521 ^ n14834;
  assign n16523 = n14876 & n16522;
  assign n16524 = n16523 ^ n14834;
  assign n16525 = ~n16517 & ~n16524;
  assign n16207 = n14842 ^ n14836;
  assign n16527 = n16207 ^ n14838;
  assign n16526 = n14861 ^ n14841;
  assign n16528 = n16527 ^ n16526;
  assign n16529 = n16528 ^ n16526;
  assign n16530 = ~n14752 & n16529;
  assign n16531 = n16530 ^ n16526;
  assign n16532 = ~n14751 & ~n16531;
  assign n16533 = n16532 ^ n16526;
  assign n16534 = n16525 & n16533;
  assign n16535 = ~n16197 & n16534;
  assign n16536 = ~n14873 & n16535;
  assign n16537 = ~n16195 & n16536;
  assign n16538 = ~n15392 & n16537;
  assign n16539 = n14875 & n16538;
  assign n16540 = n15389 & n16539;
  assign n16541 = n16540 ^ n11954;
  assign n16946 = n16541 ^ x599;
  assign n16947 = n13639 & n14008;
  assign n16948 = n16340 ^ n14042;
  assign n16949 = ~n14021 & ~n16948;
  assign n16956 = n16340 & n16819;
  assign n16957 = ~n14039 & n16956;
  assign n16958 = ~n14008 & ~n14041;
  assign n16959 = ~n16957 & ~n16958;
  assign n16952 = n16341 ^ n14041;
  assign n16950 = n14030 ^ n14023;
  assign n16951 = n16950 ^ n13639;
  assign n16953 = n16952 ^ n16951;
  assign n16954 = n14005 & n16953;
  assign n16955 = n16954 ^ n16951;
  assign n16960 = n16959 ^ n16955;
  assign n16961 = ~n13798 & n16960;
  assign n16962 = n16961 ^ n16959;
  assign n16963 = ~n16342 & ~n16962;
  assign n16964 = ~n16949 & n16963;
  assign n16965 = ~n16947 & n16964;
  assign n16966 = n14005 & n14016;
  assign n16967 = n16966 ^ n14017;
  assign n16968 = ~n13798 & n16967;
  assign n16969 = n16968 ^ n14017;
  assign n16970 = n16965 & ~n16969;
  assign n16971 = ~n14007 & n16970;
  assign n16972 = ~n16353 & n16971;
  assign n16973 = n16972 ^ n12562;
  assign n16974 = n16973 ^ x601;
  assign n16975 = ~n16946 & n16974;
  assign n17001 = n16975 ^ n16974;
  assign n17002 = n17001 ^ n16946;
  assign n16983 = n16378 ^ n15007;
  assign n16982 = n15062 ^ n14993;
  assign n16984 = n16983 ^ n16982;
  assign n16985 = ~n15020 & n16984;
  assign n16986 = n16985 ^ n16982;
  assign n16976 = n16100 ^ n15005;
  assign n16977 = n16976 ^ n15017;
  assign n16978 = n16977 ^ n15002;
  assign n16979 = ~n15020 & n16978;
  assign n16980 = n16979 ^ n15002;
  assign n16981 = ~n15010 & ~n16980;
  assign n16987 = n16986 ^ n16981;
  assign n16988 = n15078 & n16987;
  assign n16989 = n16988 ^ n16986;
  assign n16990 = ~n15053 & n16989;
  assign n16991 = ~n16127 & n16990;
  assign n16992 = ~n16099 & n16991;
  assign n16993 = ~n16376 & n16992;
  assign n16994 = ~n15064 & n16993;
  assign n16995 = n16994 ^ n12227;
  assign n16996 = n16995 ^ x600;
  assign n16997 = n15983 ^ x602;
  assign n16998 = n16996 & ~n16997;
  assign n17006 = n16998 ^ n16997;
  assign n17018 = n17002 & ~n17006;
  assign n17010 = n16998 & n17001;
  assign n17007 = n17006 ^ n16996;
  assign n17008 = n17001 & n17007;
  assign n17017 = n17010 ^ n17008;
  assign n17019 = n17018 ^ n17017;
  assign n17020 = n17019 ^ n16946;
  assign n17014 = n16998 & n17002;
  assign n17011 = n17010 ^ n17001;
  assign n17003 = n16998 ^ n16996;
  assign n17005 = n17001 & n17003;
  assign n17009 = n17008 ^ n17005;
  assign n17012 = n17011 ^ n17009;
  assign n17004 = n17002 & n17003;
  assign n17013 = n17012 ^ n17004;
  assign n17015 = n17014 ^ n17013;
  assign n17016 = n17015 ^ n17005;
  assign n17021 = n17020 ^ n17016;
  assign n17037 = n16945 & n17021;
  assign n17022 = n17021 ^ n17014;
  assign n17023 = n16942 & n17022;
  assign n17024 = n17023 ^ n17021;
  assign n17025 = n16943 & n17024;
  assign n16999 = n16975 & n16998;
  assign n17000 = n16945 & n16999;
  assign n17026 = n17025 ^ n17000;
  assign n17032 = n16999 ^ n16975;
  assign n17030 = n16975 & ~n17006;
  assign n17029 = n16975 & n17007;
  assign n17031 = n17030 ^ n17029;
  assign n17033 = n17032 ^ n17031;
  assign n17034 = n17033 ^ n17030;
  assign n17027 = n16975 ^ n16946;
  assign n17028 = n17003 & ~n17027;
  assign n17035 = n17034 ^ n17028;
  assign n17269 = n17035 ^ n16946;
  assign n17046 = n16998 & ~n17027;
  assign n17047 = n17046 ^ n17029;
  assign n17044 = n17007 & ~n17027;
  assign n17045 = n17044 ^ n16999;
  assign n17048 = n17047 ^ n17045;
  assign n17270 = n17269 ^ n17048;
  assign n17271 = n17270 ^ n17028;
  assign n17272 = n16945 & ~n17271;
  assign n17273 = n16944 ^ n16943;
  assign n17274 = n17273 ^ n16942;
  assign n17275 = n17274 ^ n17004;
  assign n17276 = n17273 ^ n17012;
  assign n17277 = ~n17004 & ~n17276;
  assign n17278 = n17277 ^ n17273;
  assign n17279 = ~n17275 & n17278;
  assign n17280 = n17279 ^ n17274;
  assign n17281 = ~n17272 & n17280;
  assign n17789 = n16943 & n17033;
  assign n17790 = n17017 ^ n17013;
  assign n17791 = n16945 & n17790;
  assign n17792 = n17045 ^ n17030;
  assign n17793 = n17792 ^ n17028;
  assign n17794 = ~n16943 & ~n17793;
  assign n17038 = n16943 ^ n16942;
  assign n17795 = n17044 ^ n17030;
  assign n17796 = n17274 & ~n17795;
  assign n17797 = ~n17038 & ~n17796;
  assign n17798 = ~n17047 & ~n17797;
  assign n17799 = ~n17794 & ~n17798;
  assign n17800 = ~n17791 & ~n17799;
  assign n17801 = ~n17789 & n17800;
  assign n17803 = n17270 ^ n17010;
  assign n17804 = n17803 ^ n17014;
  assign n17802 = n17018 ^ n17005;
  assign n17805 = n17804 ^ n17802;
  assign n17806 = n17805 ^ n17802;
  assign n17807 = n16943 & ~n17806;
  assign n17808 = n17807 ^ n17802;
  assign n17809 = n17038 & n17808;
  assign n17810 = n17809 ^ n17802;
  assign n17811 = n17801 & ~n17810;
  assign n17812 = n17281 & n17811;
  assign n17813 = ~n17026 & n17812;
  assign n17814 = ~n17037 & n17813;
  assign n17815 = n17814 ^ n12651;
  assign n17816 = n17815 ^ x680;
  assign n17817 = ~n17788 & ~n17816;
  assign n17839 = n17817 ^ n17788;
  assign n17849 = n17821 & ~n17839;
  assign n17818 = n17817 ^ n17816;
  assign n17819 = n17818 ^ n17788;
  assign n17826 = n17786 & ~n17819;
  assign n17855 = n17849 ^ n17826;
  assign n17830 = ~n17787 & ~n17818;
  assign n17856 = n17855 ^ n17830;
  assign n17822 = ~n17818 & n17821;
  assign n17857 = n17856 ^ n17822;
  assign n17858 = n17857 ^ n17821;
  assign n17824 = n17785 & ~n17819;
  assign n17825 = n17824 ^ n17822;
  assign n17827 = n17826 ^ n17825;
  assign n17828 = n17827 ^ n17819;
  assign n17820 = ~n17787 & ~n17819;
  assign n17823 = n17822 ^ n17820;
  assign n17829 = n17828 ^ n17823;
  assign n17831 = n17830 ^ n17829;
  assign n17832 = n17831 ^ n17826;
  assign n17859 = n17858 ^ n17832;
  assign n17840 = n17786 & ~n17839;
  assign n17864 = n17859 ^ n17840;
  assign n17846 = n17786 & n17817;
  assign n17865 = n17864 ^ n17846;
  assign n17848 = ~n17787 & n17817;
  assign n17862 = n17848 ^ n17840;
  assign n17863 = n17862 ^ n17817;
  assign n17866 = n17865 ^ n17863;
  assign n17845 = ~n17787 & ~n17839;
  assign n18309 = n17866 ^ n17845;
  assign n18310 = n17747 & ~n18309;
  assign n17860 = n17747 & ~n17859;
  assign n18311 = n18310 ^ n17860;
  assign n17850 = n17849 ^ n17848;
  assign n17847 = n17846 ^ n17845;
  assign n17851 = n17850 ^ n17847;
  assign n17852 = n17744 & n17851;
  assign n17853 = n17852 ^ n17847;
  assign n17854 = n17711 & n17853;
  assign n18312 = n17786 & ~n17818;
  assign n18313 = ~n17745 & n18312;
  assign n17835 = n17785 & ~n17788;
  assign n17867 = n17866 ^ n17835;
  assign n17834 = n17824 ^ n17785;
  assign n17836 = n17835 ^ n17834;
  assign n17837 = n17836 ^ n17820;
  assign n18625 = n17867 ^ n17837;
  assign n18626 = n18625 ^ n17846;
  assign n18627 = n17747 & ~n18626;
  assign n18628 = n17746 & n17835;
  assign n18629 = n17849 ^ n17836;
  assign n18630 = n18629 ^ n17824;
  assign n18631 = n18630 ^ n17831;
  assign n18632 = n18631 ^ n17826;
  assign n18633 = n18632 ^ n17826;
  assign n18634 = ~n17711 & ~n18633;
  assign n18635 = n18634 ^ n17826;
  assign n18636 = ~n17744 & n18635;
  assign n18637 = n18636 ^ n17826;
  assign n18638 = n17866 ^ n17840;
  assign n18639 = n18638 ^ n17823;
  assign n18640 = ~n17744 & ~n18639;
  assign n18641 = n18640 ^ n18638;
  assign n18642 = n17711 & ~n18641;
  assign n18643 = ~n18637 & ~n18642;
  assign n18644 = ~n18628 & n18643;
  assign n18645 = ~n18627 & n18644;
  assign n18646 = n17862 ^ n17859;
  assign n18647 = ~n17711 & ~n18646;
  assign n18648 = n18647 ^ n17859;
  assign n18649 = ~n17744 & ~n18648;
  assign n18650 = n18645 & ~n18649;
  assign n18651 = ~n18313 & n18650;
  assign n18652 = ~n17854 & n18651;
  assign n18653 = n17744 & n17827;
  assign n18654 = n18653 ^ n17826;
  assign n18655 = n17711 & n18654;
  assign n18656 = n18652 & ~n18655;
  assign n18657 = ~n18311 & n18656;
  assign n18658 = n18657 ^ n16973;
  assign n18659 = n18658 ^ x697;
  assign n17326 = n15764 ^ n15746;
  assign n17327 = n15773 & n17326;
  assign n17321 = n15786 ^ n15772;
  assign n17568 = n17321 ^ n15770;
  assign n17569 = n15425 & n17568;
  assign n17570 = n17569 ^ n17321;
  assign n17571 = ~n15775 & n17570;
  assign n17572 = ~n15738 & ~n17571;
  assign n17573 = ~n15790 & n17572;
  assign n17574 = ~n15780 & n17573;
  assign n17575 = n17574 ^ n15776;
  assign n17576 = n17575 ^ n15776;
  assign n17577 = ~n15425 & ~n17576;
  assign n17578 = n17577 ^ n15776;
  assign n17579 = ~n15381 & n17578;
  assign n17580 = n17579 ^ n15776;
  assign n17586 = n15425 & n15792;
  assign n17582 = ~n15781 & n17572;
  assign n17581 = n15785 ^ n15761;
  assign n17583 = n17582 ^ n17581;
  assign n17584 = n15425 & n17583;
  assign n17585 = n17584 ^ n17581;
  assign n17587 = n17586 ^ n17585;
  assign n17588 = ~n15381 & ~n17587;
  assign n17589 = n17588 ^ n17585;
  assign n17590 = ~n17580 & n17589;
  assign n17328 = n15786 ^ n15744;
  assign n17329 = n15425 & n17328;
  assign n17330 = n17329 ^ n15786;
  assign n17591 = n15381 & n17330;
  assign n17592 = n17590 & ~n17591;
  assign n17593 = ~n17327 & n17592;
  assign n17594 = n15426 & n15749;
  assign n17316 = n15781 ^ n15749;
  assign n17317 = n17316 ^ n15772;
  assign n17318 = ~n15425 & n17317;
  assign n17319 = n17318 ^ n15772;
  assign n17320 = ~n15381 & n17319;
  assign n17595 = n17594 ^ n17320;
  assign n17596 = n17593 & ~n17595;
  assign n17597 = ~n15741 & n17596;
  assign n17598 = n17597 ^ n14660;
  assign n18402 = n17598 ^ x652;
  assign n17282 = n16945 & n17031;
  assign n17283 = n17271 ^ n17005;
  assign n17284 = ~n16943 & ~n17283;
  assign n17285 = n17284 ^ n17271;
  assign n17286 = n17038 & ~n17285;
  assign n17287 = ~n17037 & ~n17286;
  assign n17288 = n17033 & ~n17038;
  assign n17294 = n17047 ^ n16999;
  assign n17295 = n17294 ^ n17034;
  assign n17296 = n16942 & n17295;
  assign n17297 = n17296 ^ n17034;
  assign n17290 = n17046 ^ n17045;
  assign n17289 = n17014 ^ n17012;
  assign n17291 = n17290 ^ n17289;
  assign n17292 = ~n16942 & n17291;
  assign n17293 = n17292 ^ n17289;
  assign n17298 = n17297 ^ n17293;
  assign n17299 = n16943 & n17298;
  assign n17300 = n17299 ^ n17293;
  assign n17301 = ~n17288 & ~n17300;
  assign n17302 = n17287 & n17301;
  assign n17303 = ~n17282 & n17302;
  assign n17304 = n17019 ^ n17010;
  assign n17305 = n16943 & n17304;
  assign n17306 = n17305 ^ n17010;
  assign n17307 = ~n16942 & n17306;
  assign n17308 = n17303 & ~n17307;
  assign n17310 = n17021 & ~n17038;
  assign n17309 = n16944 & n17015;
  assign n17311 = n17310 ^ n17309;
  assign n17312 = n17308 & ~n17311;
  assign n17313 = n17281 & n17312;
  assign n17314 = n17313 ^ n15046;
  assign n18403 = n17314 ^ x657;
  assign n18404 = n18402 & n18403;
  assign n18405 = n18404 ^ n18402;
  assign n18406 = n18405 ^ n18403;
  assign n18502 = n18406 ^ n18402;
  assign n16133 = n16132 ^ x628;
  assign n16093 = n16092 ^ x633;
  assign n16134 = n16133 ^ n16093;
  assign n16135 = n15692 ^ n15607;
  assign n16136 = n16135 ^ n15730;
  assign n16137 = n16136 ^ n14207;
  assign n16138 = n16137 ^ x630;
  assign n16163 = n16162 ^ x629;
  assign n16164 = n16138 & n16163;
  assign n16223 = n16164 ^ n16138;
  assign n16224 = n16223 ^ n16163;
  assign n16193 = n16192 ^ x632;
  assign n16198 = n14853 & n14857;
  assign n16201 = ~n14752 & n14843;
  assign n16199 = n14752 & n14867;
  assign n16200 = n16199 ^ n14863;
  assign n16202 = n16201 ^ n16200;
  assign n16203 = ~n14751 & ~n16202;
  assign n16204 = n16203 ^ n16200;
  assign n16205 = ~n16198 & n16204;
  assign n16206 = n14752 & n14841;
  assign n16208 = n16207 ^ n16206;
  assign n16209 = ~n14751 & n16208;
  assign n16210 = n16209 ^ n16207;
  assign n16211 = n16205 & ~n16210;
  assign n16212 = ~n16197 & n16211;
  assign n16213 = ~n14873 & n16212;
  assign n16214 = ~n16195 & n16213;
  assign n16215 = ~n14832 & n16214;
  assign n16216 = ~n15385 & n16215;
  assign n16217 = n14874 & n16216;
  assign n16218 = n16217 ^ n14232;
  assign n16219 = n16218 ^ x631;
  assign n16220 = n16193 & n16219;
  assign n16221 = n16220 ^ n16193;
  assign n16225 = n16221 ^ n16219;
  assign n16239 = ~n16224 & ~n16225;
  assign n16238 = n16220 & ~n16224;
  assign n16240 = n16239 ^ n16238;
  assign n16243 = n16240 ^ n16224;
  assign n16226 = n16225 ^ n16193;
  assign n16227 = ~n16224 & n16226;
  assign n16244 = n16243 ^ n16227;
  assign n16232 = n16193 ^ n16163;
  assign n16233 = n16232 ^ n16219;
  assign n16234 = ~n16138 & n16219;
  assign n16235 = n16234 ^ n16193;
  assign n16236 = ~n16233 & ~n16235;
  assign n16231 = n16164 & n16226;
  assign n16237 = n16236 ^ n16231;
  assign n16241 = n16240 ^ n16237;
  assign n16229 = n16193 & n16223;
  assign n16230 = n16229 ^ n16223;
  assign n16242 = n16241 ^ n16230;
  assign n16245 = n16244 ^ n16242;
  assign n16222 = n16164 & n16221;
  assign n16228 = n16227 ^ n16222;
  assign n16246 = n16245 ^ n16228;
  assign n16247 = n16093 & ~n16246;
  assign n16248 = n16247 ^ n16228;
  assign n16249 = ~n16134 & n16248;
  assign n17253 = n16236 ^ n16163;
  assign n16261 = n16219 ^ n16193;
  assign n16262 = n16163 & n16261;
  assign n16254 = n16163 ^ n16138;
  assign n16255 = n16254 ^ n16193;
  assign n16256 = n16255 ^ n16219;
  assign n16257 = n16220 & ~n16256;
  assign n16258 = n16257 ^ n16238;
  assign n16259 = n16258 ^ n16164;
  assign n16279 = n16262 ^ n16259;
  assign n16263 = n16262 ^ n16193;
  assign n16264 = n16263 ^ n16225;
  assign n16265 = n16264 ^ n16244;
  assign n16266 = n16265 ^ n16246;
  assign n16253 = n16231 ^ n16222;
  assign n16260 = n16259 ^ n16253;
  assign n16267 = n16266 ^ n16260;
  assign n16280 = n16279 ^ n16267;
  assign n16281 = n16280 ^ n16238;
  assign n16272 = n16254 & ~n16263;
  assign n16273 = n16272 ^ n16230;
  assign n16274 = n16273 ^ n16266;
  assign n17252 = n16281 ^ n16274;
  assign n17254 = n17253 ^ n17252;
  assign n17255 = ~n16133 & ~n17254;
  assign n17256 = n17255 ^ n17252;
  assign n17245 = n16219 ^ n16138;
  assign n17246 = n17245 ^ n16227;
  assign n16282 = n16281 ^ n16234;
  assign n16283 = n16282 ^ n16227;
  assign n16293 = n16283 ^ n16260;
  assign n17244 = n16293 ^ n16280;
  assign n17247 = n17246 ^ n17244;
  assign n17248 = n17247 ^ n16255;
  assign n17240 = n16193 ^ n16138;
  assign n17239 = n16224 ^ n16221;
  assign n17241 = n17240 ^ n17239;
  assign n17242 = n17241 ^ n16281;
  assign n17243 = n17242 ^ n16255;
  assign n17249 = n17248 ^ n17243;
  assign n17250 = ~n16133 & ~n17249;
  assign n17251 = n17250 ^ n17243;
  assign n17257 = n17256 ^ n17251;
  assign n17258 = n16093 & ~n17257;
  assign n17259 = n17258 ^ n17251;
  assign n17260 = ~n16093 & n16133;
  assign n17261 = n17260 ^ n16133;
  assign n17262 = n16241 & n17261;
  assign n16268 = n16267 ^ n16253;
  assign n16269 = ~n16133 & n16268;
  assign n16270 = n16269 ^ n16253;
  assign n16271 = n16093 & n16270;
  assign n17263 = n17262 ^ n16271;
  assign n17264 = n17259 & ~n17263;
  assign n17265 = ~n16249 & n17264;
  assign n17266 = n17265 ^ n14935;
  assign n18407 = n17266 ^ x656;
  assign n16910 = n16801 & ~n16885;
  assign n16907 = n16879 ^ n16872;
  assign n16908 = n16801 & n16907;
  assign n16909 = n16908 ^ n16879;
  assign n16911 = n16910 ^ n16909;
  assign n16912 = n16802 & n16911;
  assign n16913 = n16912 ^ n16909;
  assign n18408 = n16802 & ~n16891;
  assign n18409 = n18408 ^ n16884;
  assign n18410 = n16801 & n18409;
  assign n18411 = n18410 ^ n16884;
  assign n18412 = n16916 ^ n16864;
  assign n17445 = n16864 & ~n16914;
  assign n18413 = n17445 ^ n17433;
  assign n18414 = n18412 & n18413;
  assign n18415 = n18414 ^ n16916;
  assign n18416 = ~n18411 & ~n18415;
  assign n18417 = n16887 & ~n16915;
  assign n18418 = n16890 ^ n16888;
  assign n18419 = n18418 ^ n16894;
  assign n18420 = ~n16914 & ~n18419;
  assign n18421 = n18420 ^ n18418;
  assign n18422 = ~n18417 & n18421;
  assign n18423 = n18416 & n18422;
  assign n18424 = n17717 & n18423;
  assign n18425 = ~n16913 & n18424;
  assign n18426 = ~n17741 & n18425;
  assign n18427 = n18426 ^ n14968;
  assign n18428 = n18427 ^ x655;
  assign n18429 = n18407 & ~n18428;
  assign n18430 = n18429 ^ n18428;
  assign n18431 = n18430 ^ n18407;
  assign n17893 = n15359 ^ n15098;
  assign n17894 = n14750 & n17893;
  assign n17895 = n17894 ^ n15098;
  assign n17892 = n15356 ^ n15350;
  assign n17896 = n17895 ^ n17892;
  assign n17897 = n17896 ^ n15340;
  assign n17898 = n14067 & ~n17897;
  assign n17899 = n17898 ^ n17896;
  assign n18432 = n17899 ^ n15369;
  assign n17890 = n14067 & n15367;
  assign n17891 = n17890 ^ n15361;
  assign n18433 = n18432 ^ n17891;
  assign n18434 = n14424 & n18433;
  assign n18435 = n18434 ^ n17899;
  assign n18436 = n18435 ^ n14981;
  assign n18437 = n18436 ^ x654;
  assign n16542 = n16541 ^ x597;
  assign n16543 = n16372 ^ x592;
  assign n16544 = n14670 & ~n14704;
  assign n16550 = n14665 ^ n14662;
  assign n16549 = n14685 ^ n14666;
  assign n16551 = n16550 ^ n16549;
  assign n16545 = n14731 ^ n14701;
  assign n16546 = n16545 ^ n14729;
  assign n16547 = ~n14426 & ~n16546;
  assign n16548 = n16547 ^ n14729;
  assign n16552 = n16551 ^ n16548;
  assign n16553 = n16552 ^ n16548;
  assign n16554 = n14426 & n16553;
  assign n16555 = n16554 ^ n16548;
  assign n16556 = n14577 & n16555;
  assign n16557 = n16556 ^ n16548;
  assign n16558 = ~n16544 & ~n16557;
  assign n16559 = n16167 ^ n14719;
  assign n16560 = n16549 ^ n14426;
  assign n16561 = n16167 & ~n16560;
  assign n16562 = n16561 ^ n14426;
  assign n16563 = n16559 & ~n16562;
  assign n16564 = n16563 ^ n14719;
  assign n16565 = n16558 & ~n16564;
  assign n16566 = ~n14716 & n16565;
  assign n16567 = n14712 & n16566;
  assign n16568 = ~n14695 & n16567;
  assign n16569 = ~n16169 & n16568;
  assign n16570 = n16569 ^ n14455;
  assign n16571 = n16570 ^ x594;
  assign n16602 = n16601 ^ x596;
  assign n16603 = ~n16571 & n16602;
  assign n16604 = n16461 ^ x593;
  assign n16605 = n15256 & n15284;
  assign n16606 = n15275 ^ n15260;
  assign n16607 = n16606 ^ n15271;
  assign n16608 = n15152 & n16607;
  assign n16613 = n15129 & n15276;
  assign n16609 = n15292 ^ n15273;
  assign n16610 = n16609 ^ n15268;
  assign n16611 = n15129 & ~n16610;
  assign n16612 = n16611 ^ n16609;
  assign n16614 = n16613 ^ n16612;
  assign n16615 = ~n15151 & ~n16614;
  assign n16616 = n16615 ^ n16612;
  assign n16617 = ~n16608 & n16616;
  assign n16618 = ~n16605 & n16617;
  assign n16619 = ~n15281 & n16618;
  assign n16620 = n15290 & n16619;
  assign n16621 = n15946 & n16620;
  assign n16622 = ~n15939 & n16621;
  assign n16623 = ~n16157 & n16622;
  assign n16624 = n15960 & n16623;
  assign n16625 = ~n15280 & n16624;
  assign n16626 = n16625 ^ n14480;
  assign n16627 = n16626 ^ x595;
  assign n16628 = ~n16604 & n16627;
  assign n16635 = n16628 ^ n16627;
  assign n16636 = n16635 ^ n16604;
  assign n16639 = n16603 & n16636;
  assign n16640 = n16639 ^ n16636;
  assign n16637 = ~n16602 & n16636;
  assign n16641 = n16640 ^ n16637;
  assign n16638 = ~n16571 & n16637;
  assign n16642 = n16641 ^ n16638;
  assign n16643 = n16543 & n16642;
  assign n16644 = n16643 ^ n16641;
  assign n16630 = n16628 ^ n16604;
  assign n16631 = n16603 & ~n16630;
  assign n16629 = n16603 & n16628;
  assign n16632 = n16631 ^ n16629;
  assign n16633 = n16543 & n16632;
  assign n16634 = n16633 ^ n16629;
  assign n16645 = n16644 ^ n16634;
  assign n16646 = n16542 & n16645;
  assign n16647 = n16646 ^ n16634;
  assign n16648 = ~n16602 & ~n16630;
  assign n16649 = n16571 & n16648;
  assign n16650 = n16649 ^ n16648;
  assign n16651 = n16650 ^ n16641;
  assign n16652 = ~n16543 & n16651;
  assign n16653 = n16652 ^ n16641;
  assign n16654 = n16542 & n16653;
  assign n16655 = ~n16602 & n16635;
  assign n16665 = ~n16571 & n16655;
  assign n16666 = n16665 ^ n16655;
  assign n16695 = n16543 ^ n16542;
  assign n16670 = n16631 ^ n16630;
  assign n16671 = n16670 ^ n16648;
  assign n17075 = ~n16543 & ~n16671;
  assign n17072 = n16665 ^ n16638;
  assign n17073 = n16543 & n17072;
  assign n17074 = n17073 ^ n16638;
  assign n17076 = n17075 ^ n17074;
  assign n17077 = n16695 & n17076;
  assign n17078 = n17077 ^ n17074;
  assign n16656 = ~n16542 & ~n16543;
  assign n16657 = n16656 ^ n16542;
  assign n16662 = n16632 ^ n16603;
  assign n16663 = n16662 ^ n16639;
  assign n17473 = ~n16657 & n16663;
  assign n16686 = n16655 ^ n16635;
  assign n16687 = n16686 ^ n16663;
  assign n16661 = n16638 ^ n16637;
  assign n16701 = n16687 ^ n16661;
  assign n16702 = n16701 ^ n16665;
  assign n17478 = n16702 ^ n16631;
  assign n17476 = n16701 ^ n16650;
  assign n16675 = ~n16602 & n16628;
  assign n16678 = ~n16571 & n16675;
  assign n16683 = n16678 ^ n16629;
  assign n16674 = n16629 ^ n16628;
  assign n16676 = n16675 ^ n16674;
  assign n16684 = n16683 ^ n16676;
  assign n16685 = n16684 ^ n16628;
  assign n17080 = n16685 ^ n16671;
  assign n17477 = n17476 ^ n17080;
  assign n17479 = n17478 ^ n17477;
  assign n17480 = ~n16543 & ~n17479;
  assign n17481 = n17480 ^ n17477;
  assign n17474 = n16684 ^ n16639;
  assign n17475 = ~n16543 & n17474;
  assign n17482 = n17481 ^ n17475;
  assign n17483 = n16542 & ~n17482;
  assign n17484 = n17483 ^ n17481;
  assign n17485 = ~n17473 & n17484;
  assign n16669 = n16657 ^ n16543;
  assign n17486 = n16669 ^ n16649;
  assign n16699 = n16685 ^ n16676;
  assign n16700 = n16699 ^ n16629;
  assign n17487 = n16700 ^ n16656;
  assign n17488 = ~n16649 & ~n17487;
  assign n17489 = n17488 ^ n16656;
  assign n17490 = ~n17486 & n17489;
  assign n17491 = n17490 ^ n16669;
  assign n17492 = n17485 & n17491;
  assign n17493 = ~n17078 & n17492;
  assign n17494 = ~n16666 & n17493;
  assign n17495 = ~n16654 & n17494;
  assign n17496 = ~n16647 & n17495;
  assign n17497 = n17496 ^ n14576;
  assign n18438 = n17497 ^ x653;
  assign n18439 = ~n18437 & ~n18438;
  assign n18442 = n18439 ^ n18437;
  assign n18443 = n18442 ^ n18438;
  assign n18444 = n18443 ^ n18437;
  assign n18475 = n18431 & ~n18444;
  assign n18469 = ~n18430 & n18439;
  assign n18445 = n18429 ^ n18407;
  assign n18468 = n18439 & n18445;
  assign n18470 = n18469 ^ n18468;
  assign n18473 = n18470 ^ n18439;
  assign n18440 = n18431 & n18439;
  assign n18474 = n18473 ^ n18440;
  assign n18476 = n18475 ^ n18474;
  assign n18477 = n18476 ^ n18440;
  assign n18466 = ~n18430 & ~n18444;
  assign n18446 = ~n18444 & n18445;
  assign n18467 = n18466 ^ n18446;
  assign n18471 = n18470 ^ n18467;
  assign n18472 = n18471 ^ n18438;
  assign n18478 = n18477 ^ n18472;
  assign n18695 = n18478 ^ n18469;
  assign n18696 = n18502 & ~n18695;
  assign n18460 = ~n18443 & n18445;
  assign n18455 = n18431 & ~n18443;
  assign n18461 = n18460 ^ n18455;
  assign n18448 = n18429 & ~n18443;
  assign n18459 = n18448 ^ n18443;
  assign n18462 = n18461 ^ n18459;
  assign n18463 = n18462 ^ n18438;
  assign n18454 = ~n18442 & n18445;
  assign n18456 = n18455 ^ n18454;
  assign n18450 = n18429 & ~n18442;
  assign n18457 = n18456 ^ n18450;
  assign n18458 = n18457 ^ n18448;
  assign n18464 = n18463 ^ n18458;
  assign n18494 = n18464 ^ n18455;
  assign n18700 = n18494 ^ n18443;
  assign n18698 = n18431 & ~n18442;
  assign n18699 = n18698 ^ n18462;
  assign n18701 = n18700 ^ n18699;
  assign n18697 = n18460 & ~n18502;
  assign n18702 = n18701 ^ n18697;
  assign n18703 = ~n18405 & ~n18702;
  assign n18704 = n18703 ^ n18701;
  assign n18705 = ~n18696 & n18704;
  assign n18453 = n18403 ^ n18402;
  assign n18706 = n18468 ^ n18450;
  assign n18707 = ~n18402 & n18706;
  assign n18708 = n18707 ^ n18450;
  assign n18709 = ~n18453 & n18708;
  assign n18710 = ~n18402 & ~n18462;
  assign n18711 = n18710 ^ n18467;
  assign n18712 = ~n18453 & n18711;
  assign n18713 = n18712 ^ n18467;
  assign n18714 = n18462 ^ n18440;
  assign n18715 = n18714 ^ n18474;
  assign n18716 = n18715 ^ n18454;
  assign n18717 = n18405 & ~n18716;
  assign n18719 = ~n18404 & ~n18477;
  assign n18500 = n18476 ^ n18466;
  assign n18720 = n18500 ^ n18468;
  assign n18441 = ~n18406 & n18440;
  assign n18721 = n18720 ^ n18441;
  assign n18722 = ~n18719 & n18721;
  assign n18723 = n18701 & ~n18722;
  assign n18718 = n18698 ^ n18457;
  assign n18724 = n18723 ^ n18718;
  assign n18725 = n18724 ^ n18718;
  assign n18726 = ~n18405 & ~n18725;
  assign n18727 = n18726 ^ n18718;
  assign n18728 = ~n18502 & n18727;
  assign n18729 = n18728 ^ n18718;
  assign n18730 = ~n18717 & ~n18729;
  assign n18731 = ~n18713 & n18730;
  assign n18732 = ~n18709 & n18731;
  assign n18733 = n18705 & n18732;
  assign n18734 = n18733 ^ n16995;
  assign n18735 = n18734 ^ x696;
  assign n17127 = n16013 ^ n16006;
  assign n17128 = ~n15984 & ~n17127;
  assign n17129 = n17128 ^ n16013;
  assign n17130 = ~n15935 & ~n17129;
  assign n17131 = n15985 & ~n16028;
  assign n17132 = n15930 ^ n15922;
  assign n17133 = ~n15997 & n17132;
  assign n17134 = n16002 & n16037;
  assign n17141 = n16008 ^ n15922;
  assign n17142 = ~n15984 & n17141;
  assign n17143 = n17142 ^ n15922;
  assign n17137 = n16030 ^ n15925;
  assign n17135 = n16010 ^ n15992;
  assign n17136 = n17135 ^ n16013;
  assign n17138 = n17137 ^ n17136;
  assign n17139 = n15984 & ~n17138;
  assign n17140 = n17139 ^ n17136;
  assign n17144 = n17143 ^ n17140;
  assign n17145 = ~n15935 & n17144;
  assign n17146 = n17145 ^ n17140;
  assign n17147 = ~n17134 & ~n17146;
  assign n17148 = ~n17133 & n17147;
  assign n17150 = n15985 & ~n16032;
  assign n17149 = ~n16002 & n16015;
  assign n17151 = n17150 ^ n17149;
  assign n17152 = n17148 & ~n17151;
  assign n17153 = ~n15995 & n17152;
  assign n17154 = ~n17131 & n17153;
  assign n17155 = ~n17130 & n17154;
  assign n17156 = ~n16056 & n17155;
  assign n17157 = ~n15987 & n17156;
  assign n17158 = n17157 ^ n15128;
  assign n17159 = n17158 ^ x664;
  assign n16450 = n16449 ^ n16435;
  assign n16466 = n16465 ^ n16462;
  assign n16467 = n16450 & n16466;
  assign n16470 = n16469 ^ n16467;
  assign n16471 = n16443 ^ n16422;
  assign n16472 = n16466 & ~n16471;
  assign n16474 = n16473 ^ n16410;
  assign n16475 = n16464 & ~n16474;
  assign n16482 = n16465 ^ n16441;
  assign n16483 = n16464 ^ n16408;
  assign n16484 = ~n16441 & ~n16483;
  assign n16485 = n16484 ^ n16464;
  assign n16486 = n16482 & n16485;
  assign n16487 = n16486 ^ n16465;
  assign n16488 = n16464 ^ n16462;
  assign n16489 = n16488 ^ n16424;
  assign n16491 = n16477 ^ n16422;
  assign n16490 = n16424 & ~n16477;
  assign n16492 = n16491 ^ n16490;
  assign n16493 = n16492 ^ n16477;
  assign n16494 = ~n16489 & ~n16493;
  assign n16495 = n16494 ^ n16488;
  assign n16496 = ~n16487 & n16495;
  assign n16497 = ~n16413 & ~n16463;
  assign n16498 = n16497 ^ n16432;
  assign n16499 = n16477 & ~n16498;
  assign n16500 = n16499 ^ n16432;
  assign n16501 = n16496 & n16500;
  assign n16502 = ~n16481 & n16501;
  assign n16503 = ~n16476 & n16502;
  assign n16504 = ~n16475 & n16503;
  assign n16505 = ~n16472 & n16504;
  assign n16506 = n16417 ^ n16400;
  assign n16507 = n16506 ^ n16488;
  assign n16508 = n16465 ^ n16414;
  assign n16509 = ~n16506 & ~n16508;
  assign n16510 = n16509 ^ n16465;
  assign n16511 = ~n16507 & n16510;
  assign n16512 = n16511 ^ n16488;
  assign n16513 = n16505 & n16512;
  assign n16514 = ~n16470 & n16513;
  assign n16515 = n16514 ^ n15150;
  assign n17160 = n16515 ^ x669;
  assign n16917 = n16876 & ~n16914;
  assign n16918 = n16917 ^ n16895;
  assign n16919 = ~n16916 & n16918;
  assign n16920 = n16919 ^ n16895;
  assign n16925 = n16897 ^ n16891;
  assign n16921 = n16893 ^ n16892;
  assign n16922 = n16921 ^ n16865;
  assign n16923 = ~n16802 & ~n16922;
  assign n16924 = n16923 ^ n16865;
  assign n16926 = n16925 ^ n16924;
  assign n16927 = n16926 ^ n16924;
  assign n16928 = ~n16802 & n16927;
  assign n16929 = n16928 ^ n16924;
  assign n16930 = n16801 & n16929;
  assign n16931 = n16930 ^ n16924;
  assign n16932 = ~n16920 & ~n16931;
  assign n16934 = n16870 & n16904;
  assign n16933 = n16866 & ~n16915;
  assign n16935 = n16934 ^ n16933;
  assign n16936 = n16932 & ~n16935;
  assign n16937 = ~n16913 & n16936;
  assign n16938 = ~n16906 & n16937;
  assign n16939 = n16903 & n16938;
  assign n16940 = n16939 ^ n15186;
  assign n16941 = n16940 ^ x667;
  assign n17036 = n16945 & n17035;
  assign n17050 = n17045 ^ n17034;
  assign n17049 = ~n16943 & n17048;
  assign n17051 = n17050 ^ n17049;
  assign n17039 = n17018 ^ n17014;
  assign n17040 = n17039 ^ n17008;
  assign n17041 = n17040 ^ n17027;
  assign n17042 = ~n16943 & ~n17041;
  assign n17043 = n17042 ^ n17027;
  assign n17052 = n17051 ^ n17043;
  assign n17053 = n17038 & ~n17052;
  assign n17054 = n17053 ^ n17051;
  assign n17055 = ~n17037 & ~n17054;
  assign n17056 = ~n17036 & n17055;
  assign n17057 = n17016 ^ n17012;
  assign n17058 = ~n16943 & n17057;
  assign n17059 = n17058 ^ n17012;
  assign n17060 = ~n16942 & n17059;
  assign n17061 = n17056 & ~n17060;
  assign n17063 = n16944 & n17021;
  assign n17062 = n16943 & n17017;
  assign n17064 = n17063 ^ n17062;
  assign n17065 = n17061 & ~n17064;
  assign n17066 = ~n17026 & n17065;
  assign n17067 = n17066 ^ n15213;
  assign n17068 = n17067 ^ x666;
  assign n17069 = n16941 & n17068;
  assign n17070 = n17069 ^ n16941;
  assign n15347 = n14424 & ~n15346;
  assign n15348 = n15347 ^ n15335;
  assign n15376 = n15375 ^ n15348;
  assign n15377 = n14425 & ~n15376;
  assign n15378 = n15377 ^ n15375;
  assign n15379 = n15378 ^ n15156;
  assign n17071 = n15379 ^ x668;
  assign n16659 = n16641 & n16656;
  assign n16703 = n16702 ^ n16700;
  assign n17085 = n16703 ^ n16641;
  assign n17081 = n17080 ^ n16683;
  assign n17079 = n16699 ^ n16649;
  assign n17082 = n17081 ^ n17079;
  assign n17083 = n16543 & ~n17082;
  assign n17084 = n17083 ^ n17079;
  assign n17086 = n17085 ^ n17084;
  assign n17087 = n17086 ^ n17084;
  assign n17088 = n16543 & n17087;
  assign n17089 = n17088 ^ n17084;
  assign n17090 = n16695 & n17089;
  assign n17091 = n17090 ^ n17084;
  assign n17092 = n16676 ^ n16638;
  assign n17093 = n17092 ^ n16687;
  assign n16664 = n16663 ^ n16661;
  assign n16667 = n16666 ^ n16664;
  assign n17094 = n17093 ^ n16667;
  assign n17095 = n17094 ^ n16639;
  assign n17096 = n17095 ^ n16639;
  assign n17097 = ~n16543 & n17096;
  assign n17098 = n17097 ^ n16639;
  assign n17099 = n16695 & n17098;
  assign n17100 = n17099 ^ n16639;
  assign n17101 = ~n17091 & ~n17100;
  assign n17102 = n16666 ^ n16661;
  assign n17103 = n16543 & n17102;
  assign n17104 = n17103 ^ n16666;
  assign n17105 = ~n16695 & n17104;
  assign n17106 = n17101 & ~n17105;
  assign n17107 = ~n16659 & n17106;
  assign n17108 = ~n17078 & n17107;
  assign n17109 = n16653 ^ n16634;
  assign n17110 = ~n16542 & n17109;
  assign n17111 = n17110 ^ n16653;
  assign n17112 = n17108 & ~n17111;
  assign n17113 = n17112 ^ n15241;
  assign n17114 = n17113 ^ x665;
  assign n17115 = n17071 & n17114;
  assign n17198 = n17115 ^ n17071;
  assign n17204 = n17070 & n17198;
  assign n17119 = n17115 ^ n17114;
  assign n17193 = n17119 ^ n17071;
  assign n17194 = ~n17068 & ~n17193;
  assign n17163 = n17071 ^ n17068;
  assign n17166 = ~n17114 & ~n17163;
  assign n17200 = n17194 ^ n17166;
  assign n17199 = n17069 & n17198;
  assign n17201 = n17200 ^ n17199;
  assign n17205 = n17204 ^ n17201;
  assign n17203 = n17199 ^ n17198;
  assign n17206 = n17205 ^ n17203;
  assign n17195 = n17194 ^ n17193;
  assign n17196 = ~n16941 & ~n17195;
  assign n17197 = n17196 ^ n17195;
  assign n18513 = n17206 ^ n17197;
  assign n18514 = n17160 & ~n18513;
  assign n18515 = n18514 ^ n17206;
  assign n18516 = ~n17159 & n18515;
  assign n17121 = n17071 ^ n16941;
  assign n17122 = ~n17068 & n17121;
  assign n17123 = n17122 ^ n16941;
  assign n17124 = n17114 & ~n17123;
  assign n17117 = n17069 ^ n17068;
  assign n17118 = n17115 & n17117;
  assign n17120 = n17119 ^ n17118;
  assign n17125 = n17124 ^ n17120;
  assign n17177 = n17125 ^ n17118;
  assign n17165 = n17117 & n17119;
  assign n17116 = n17070 & n17115;
  assign n17126 = n17125 ^ n17116;
  assign n17175 = n17165 ^ n17126;
  assign n17170 = n17070 & n17119;
  assign n17171 = n17170 ^ n17116;
  assign n17174 = n17171 ^ n17119;
  assign n17176 = n17175 ^ n17174;
  assign n17178 = n17177 ^ n17176;
  assign n17167 = n17166 ^ n17165;
  assign n17164 = n17163 ^ n17124;
  assign n17168 = n17167 ^ n17164;
  assign n17169 = n17168 ^ n17165;
  assign n17172 = n17171 ^ n17169;
  assign n17173 = n17172 ^ n17114;
  assign n17179 = n17178 ^ n17173;
  assign n17180 = n17179 ^ n17169;
  assign n17181 = n17159 & n17180;
  assign n17182 = n17181 ^ n17169;
  assign n17183 = ~n17160 & ~n17182;
  assign n17185 = n17179 ^ n17176;
  assign n17186 = n17160 & ~n17185;
  assign n17187 = n17186 ^ n17176;
  assign n17188 = n17159 & n17187;
  assign n17161 = n17159 & n17160;
  assign n17190 = n17161 ^ n17159;
  assign n17191 = n17190 ^ n17160;
  assign n17192 = n17191 ^ n17159;
  assign n18661 = ~n17068 & n17192;
  assign n18662 = n17114 ^ n16941;
  assign n18663 = n18662 ^ n17192;
  assign n18664 = n18661 ^ n17198;
  assign n18665 = n18663 & n18664;
  assign n18666 = n18665 ^ n17198;
  assign n18667 = n18661 & n18666;
  assign n17202 = n17201 ^ n17197;
  assign n18674 = n17202 ^ n17126;
  assign n18670 = n17167 ^ n17116;
  assign n17224 = n17199 ^ n17196;
  assign n18668 = n17224 ^ n17205;
  assign n18522 = n17170 ^ n17168;
  assign n18669 = n18668 ^ n18522;
  assign n18671 = n18670 ^ n18669;
  assign n18672 = n17160 & ~n18671;
  assign n18673 = n18672 ^ n18669;
  assign n18675 = n18674 ^ n18673;
  assign n18676 = n18675 ^ n18673;
  assign n18677 = ~n17160 & ~n18676;
  assign n18678 = n18677 ^ n18673;
  assign n18679 = ~n17159 & ~n18678;
  assign n18680 = n18679 ^ n18673;
  assign n18681 = ~n18667 & n18680;
  assign n18682 = ~n17188 & n18681;
  assign n18685 = n17160 & n17206;
  assign n18683 = n17160 & n17178;
  assign n18684 = n18683 ^ n17176;
  assign n18686 = n18685 ^ n18684;
  assign n18687 = n17159 & n18686;
  assign n18688 = n18687 ^ n18684;
  assign n18689 = n18682 & ~n18688;
  assign n18690 = ~n17183 & n18689;
  assign n18691 = ~n18516 & n18690;
  assign n18692 = n18691 ^ n15983;
  assign n18693 = n18692 ^ x698;
  assign n17900 = n17899 ^ n17891;
  assign n17901 = ~n14424 & ~n17900;
  assign n17902 = n17901 ^ n17899;
  assign n17903 = ~n15369 & n17902;
  assign n17904 = n17903 ^ n14150;
  assign n17905 = n17904 ^ x687;
  assign n17889 = n17815 ^ x682;
  assign n17906 = n17905 ^ n17889;
  assign n16250 = n16133 & n16240;
  assign n16251 = n16250 ^ n16238;
  assign n16252 = n16093 & n16251;
  assign n17541 = n16266 ^ n16242;
  assign n17542 = n16133 & n17541;
  assign n17543 = n17542 ^ n16242;
  assign n17544 = n16093 & n17543;
  assign n17545 = n17260 ^ n16093;
  assign n17907 = ~n17243 & ~n17545;
  assign n17908 = n16272 ^ n16219;
  assign n17909 = n17260 & ~n17908;
  assign n17910 = n16280 ^ n16134;
  assign n17911 = n17261 ^ n16258;
  assign n17912 = ~n16134 & ~n17911;
  assign n17913 = n17912 ^ n16258;
  assign n17914 = n17910 & n17913;
  assign n17915 = n17914 ^ n16280;
  assign n17916 = ~n17909 & ~n17915;
  assign n17917 = ~n17907 & n17916;
  assign n16286 = n16244 ^ n16241;
  assign n17918 = n16286 ^ n16229;
  assign n17919 = n16133 & ~n17918;
  assign n17920 = n17919 ^ n16286;
  assign n17921 = n16093 & ~n17920;
  assign n17922 = n17917 & ~n17921;
  assign n17923 = ~n17544 & n17922;
  assign n17924 = ~n16252 & n17923;
  assign n17925 = ~n17263 & n17924;
  assign n17926 = n17925 ^ n14303;
  assign n17927 = n17926 ^ x686;
  assign n17929 = n15928 & ~n15984;
  assign n17928 = n16014 ^ n16003;
  assign n17930 = n17929 ^ n17928;
  assign n17931 = ~n15935 & ~n17930;
  assign n17932 = n17931 ^ n17928;
  assign n17933 = n16034 ^ n16017;
  assign n17934 = n17933 ^ n16018;
  assign n17935 = n15984 & n17934;
  assign n17936 = n17935 ^ n16018;
  assign n17937 = n16002 & n17936;
  assign n17938 = n17932 & ~n17937;
  assign n17940 = n15993 & ~n16002;
  assign n17939 = n15930 & ~n16055;
  assign n17941 = n17940 ^ n17939;
  assign n17942 = n17938 & ~n17941;
  assign n17943 = ~n17131 & n17942;
  assign n17944 = ~n16058 & n17943;
  assign n17945 = ~n15987 & n17944;
  assign n17946 = n17945 ^ n14817;
  assign n17947 = n17946 ^ x684;
  assign n17948 = n17927 & ~n17947;
  assign n17988 = n17948 ^ n17947;
  assign n17949 = n17743 ^ x683;
  assign n17950 = ~n16695 & n17074;
  assign n16658 = n16655 & ~n16657;
  assign n16660 = n16659 ^ n16658;
  assign n17951 = n16676 ^ n16650;
  assign n17952 = ~n16669 & n17951;
  assign n16679 = n16678 ^ n16631;
  assign n17956 = n16699 ^ n16679;
  assign n16696 = n16687 ^ n16639;
  assign n17953 = n16701 ^ n16696;
  assign n17954 = ~n16543 & n17953;
  assign n17955 = n17954 ^ n16696;
  assign n17957 = n17956 ^ n17955;
  assign n17958 = n17957 ^ n17955;
  assign n17959 = ~n16543 & n17958;
  assign n17960 = n17959 ^ n17955;
  assign n17961 = n16695 & n17960;
  assign n17962 = n17961 ^ n17955;
  assign n17963 = ~n17952 & ~n17962;
  assign n17964 = n17092 ^ n16649;
  assign n17965 = n17964 ^ n16664;
  assign n17966 = n17965 ^ n17080;
  assign n17967 = n17966 ^ n17080;
  assign n17968 = n16543 & n17967;
  assign n17969 = n17968 ^ n17080;
  assign n17970 = n16695 & ~n17969;
  assign n17971 = n17970 ^ n17080;
  assign n17972 = n17963 & n17971;
  assign n17973 = n16678 ^ n16667;
  assign n17974 = n16542 & n17973;
  assign n17975 = n17974 ^ n16678;
  assign n17976 = ~n16543 & n17975;
  assign n17977 = n17972 & ~n17976;
  assign n17978 = ~n16660 & n17977;
  assign n17979 = ~n17950 & n17978;
  assign n17980 = ~n16647 & n17979;
  assign n17981 = n17980 ^ n14793;
  assign n17982 = n17981 ^ x685;
  assign n17983 = ~n17949 & ~n17982;
  assign n17984 = n17983 ^ n17982;
  assign n17993 = n17984 ^ n17949;
  assign n17994 = ~n17988 & ~n17993;
  assign n17989 = ~n17984 & ~n17988;
  assign n17986 = n17948 ^ n17927;
  assign n17987 = ~n17984 & n17986;
  assign n17990 = n17989 ^ n17987;
  assign n17985 = n17948 & ~n17984;
  assign n17991 = n17990 ^ n17985;
  assign n17992 = n17991 ^ n17984;
  assign n17995 = n17994 ^ n17992;
  assign n17996 = n17889 & ~n17995;
  assign n17997 = n17996 ^ n17994;
  assign n17998 = ~n17906 & n17997;
  assign n17999 = ~n17889 & n17905;
  assign n18000 = n17999 ^ n17905;
  assign n18001 = n18000 ^ n17889;
  assign n18002 = n17991 & n18001;
  assign n18017 = n17988 ^ n17927;
  assign n18014 = n17986 & ~n17993;
  assign n18015 = n18014 ^ n17994;
  assign n18012 = n17948 & ~n17993;
  assign n18013 = n18012 ^ n17993;
  assign n18016 = n18015 ^ n18013;
  assign n18018 = n18017 ^ n18016;
  assign n18008 = n17983 & ~n17988;
  assign n18007 = n17983 & n17986;
  assign n18009 = n18008 ^ n18007;
  assign n18005 = n17948 & n17983;
  assign n18006 = n18005 ^ n17983;
  assign n18010 = n18009 ^ n18006;
  assign n18011 = n18010 ^ n17992;
  assign n18019 = n18018 ^ n18011;
  assign n18003 = n17983 ^ n17949;
  assign n18004 = n17986 & ~n18003;
  assign n18020 = n18019 ^ n18004;
  assign n18021 = n17999 & n18020;
  assign n18023 = n17948 & ~n18003;
  assign n18026 = n18023 ^ n18004;
  assign n18030 = n18026 ^ n18008;
  assign n18022 = n18010 ^ n18005;
  assign n18024 = n18023 ^ n18022;
  assign n18025 = n18024 ^ n18008;
  assign n18027 = n18026 ^ n18025;
  assign n18028 = n17889 & n18027;
  assign n18029 = n18028 ^ n18026;
  assign n18031 = n18030 ^ n18029;
  assign n18032 = n18031 ^ n18029;
  assign n18033 = n17889 & n18032;
  assign n18034 = n18033 ^ n18029;
  assign n18035 = n17906 & n18034;
  assign n18036 = n18035 ^ n18029;
  assign n18038 = n17992 ^ n17985;
  assign n18039 = n18038 ^ n18015;
  assign n18037 = n18014 ^ n17992;
  assign n18040 = n18039 ^ n18037;
  assign n18041 = n17905 & n18040;
  assign n18042 = n18041 ^ n18037;
  assign n18043 = ~n17889 & ~n18042;
  assign n18044 = ~n18036 & ~n18043;
  assign n18047 = ~n17988 & ~n18003;
  assign n18048 = n18001 & n18047;
  assign n18045 = n17999 ^ n17889;
  assign n18046 = n18022 & ~n18045;
  assign n18049 = n18048 ^ n18046;
  assign n18050 = n18044 & ~n18049;
  assign n18051 = ~n18021 & n18050;
  assign n18052 = ~n18002 & n18051;
  assign n18054 = n17889 & ~n18016;
  assign n18053 = ~n17906 & n17987;
  assign n18055 = n18054 ^ n18053;
  assign n18056 = n18052 & ~n18055;
  assign n18057 = n18012 ^ n18009;
  assign n18058 = ~n17889 & n18057;
  assign n18059 = n18058 ^ n18012;
  assign n18060 = n17905 & n18059;
  assign n18061 = n18056 & ~n18060;
  assign n18062 = ~n17998 & n18061;
  assign n18063 = n18062 ^ n16541;
  assign n18660 = n18063 ^ x695;
  assign n18694 = n18693 ^ n18660;
  assign n18736 = n18735 ^ n18694;
  assign n18737 = ~n18659 & ~n18736;
  assign n15380 = n15379 ^ x670;
  assign n15824 = n15823 ^ x675;
  assign n16062 = n16061 ^ x674;
  assign n16275 = n16274 ^ n16242;
  assign n16276 = ~n16133 & n16275;
  assign n16277 = n16276 ^ n16242;
  assign n16278 = ~n16093 & n16277;
  assign n16295 = ~n16163 & n16219;
  assign n16296 = n16295 ^ n16138;
  assign n16297 = n16261 & n16296;
  assign n16298 = n16297 ^ n16163;
  assign n16299 = ~n16093 & n16298;
  assign n16291 = n16257 ^ n16220;
  assign n16292 = n16291 ^ n16283;
  assign n16294 = n16293 ^ n16292;
  assign n16300 = n16299 ^ n16294;
  assign n16288 = n16257 ^ n16256;
  assign n16289 = n16093 & n16288;
  assign n16284 = n16283 ^ n16231;
  assign n16285 = n16284 ^ n16238;
  assign n16287 = n16286 ^ n16285;
  assign n16290 = n16289 ^ n16287;
  assign n16301 = n16300 ^ n16290;
  assign n16302 = ~n16133 & ~n16301;
  assign n16303 = n16302 ^ n16300;
  assign n16304 = ~n16278 & ~n16303;
  assign n16305 = ~n16271 & n16304;
  assign n16306 = ~n16252 & n16305;
  assign n16307 = ~n16249 & n16306;
  assign n16308 = n16307 ^ n15493;
  assign n16309 = n16308 ^ x672;
  assign n16516 = n16515 ^ x671;
  assign n16724 = n16309 & n16516;
  assign n16725 = ~n16062 & n16724;
  assign n16310 = n16062 & ~n16309;
  assign n16311 = n16310 ^ n16309;
  assign n16722 = n16311 ^ n16062;
  assign n16747 = n16725 ^ n16722;
  assign n16668 = n16656 & n16667;
  assign n16677 = n16656 & n16676;
  assign n16680 = n16679 ^ n16677;
  assign n16672 = n16671 ^ n16649;
  assign n16673 = ~n16669 & ~n16672;
  assign n16681 = n16680 ^ n16673;
  assign n16682 = n16681 ^ n16669;
  assign n16688 = n16687 ^ n16685;
  assign n16689 = n16688 ^ n16656;
  assign n16690 = ~n16681 & ~n16689;
  assign n16691 = n16690 ^ n16656;
  assign n16692 = ~n16682 & n16691;
  assign n16693 = n16692 ^ n16669;
  assign n16694 = ~n16668 & n16693;
  assign n16697 = n16696 ^ n16648;
  assign n16698 = n16697 ^ n16629;
  assign n16704 = n16703 ^ n16698;
  assign n16705 = ~n16543 & n16704;
  assign n16706 = n16705 ^ n16698;
  assign n16707 = n16695 & n16706;
  assign n16708 = n16694 & ~n16707;
  assign n16709 = ~n16660 & n16708;
  assign n16710 = ~n16654 & n16709;
  assign n16711 = ~n16647 & n16710;
  assign n16712 = n16711 ^ n15521;
  assign n16713 = n16712 ^ x673;
  assign n16714 = ~n16516 & n16713;
  assign n16716 = n16714 ^ n16516;
  assign n16746 = ~n16716 & n16722;
  assign n16748 = n16747 ^ n16746;
  assign n16739 = n16713 ^ n16309;
  assign n16740 = n16739 ^ n16062;
  assign n16741 = n16740 ^ n16516;
  assign n16742 = n16741 ^ n16713;
  assign n16743 = n16716 ^ n16062;
  assign n16744 = ~n16742 & ~n16743;
  assign n16745 = n16744 ^ n16739;
  assign n16749 = n16748 ^ n16745;
  assign n16717 = n16716 ^ n16713;
  assign n16730 = n16310 & n16717;
  assign n16731 = n16730 ^ n16725;
  assign n16732 = n16731 ^ n16516;
  assign n16750 = n16749 ^ n16732;
  assign n16719 = n16717 ^ n16516;
  assign n16720 = n16310 & n16719;
  assign n16727 = n16720 ^ n16719;
  assign n16736 = n16727 ^ n16724;
  assign n16723 = n16717 & n16722;
  assign n16726 = n16725 ^ n16723;
  assign n16728 = n16727 ^ n16726;
  assign n16718 = ~n16311 & n16717;
  assign n16721 = n16720 ^ n16718;
  assign n16729 = n16728 ^ n16721;
  assign n16733 = n16732 ^ n16729;
  assign n16735 = n16733 ^ n16723;
  assign n16737 = n16736 ^ n16735;
  assign n16734 = n16733 ^ n16726;
  assign n16738 = n16737 ^ n16734;
  assign n16751 = n16750 ^ n16738;
  assign n16715 = ~n16311 & n16714;
  assign n16752 = n16751 ^ n16715;
  assign n16753 = n16752 ^ n16746;
  assign n16754 = n15824 & ~n16753;
  assign n16755 = n16754 ^ n16746;
  assign n16756 = n15380 & n16755;
  assign n16757 = n16751 ^ n16748;
  assign n16758 = n15380 & ~n15824;
  assign n16759 = n16758 ^ n15824;
  assign n16760 = ~n16757 & ~n16759;
  assign n16767 = n16748 ^ n16714;
  assign n16761 = n16310 ^ n16062;
  assign n16762 = n16714 & n16761;
  assign n16766 = n16762 ^ n16715;
  assign n16768 = n16767 ^ n16766;
  assign n16769 = n16768 ^ n16728;
  assign n16763 = n16762 ^ n16723;
  assign n16764 = n16763 ^ n16730;
  assign n16765 = n16764 ^ n16718;
  assign n16770 = n16769 ^ n16765;
  assign n16771 = n16758 & n16770;
  assign n16772 = n15824 ^ n15380;
  assign n16776 = n16747 ^ n16714;
  assign n16777 = ~n15380 & n16776;
  assign n16774 = n15380 & n16725;
  assign n16773 = n16738 ^ n16720;
  assign n16775 = n16774 ^ n16773;
  assign n16778 = n16777 ^ n16775;
  assign n16779 = n16772 & n16778;
  assign n16780 = n16779 ^ n16775;
  assign n16781 = ~n16771 & ~n16780;
  assign n16782 = ~n16760 & n16781;
  assign n16785 = n16761 ^ n16727;
  assign n16784 = n16762 ^ n16738;
  assign n16786 = n16785 ^ n16784;
  assign n16787 = ~n16772 & n16786;
  assign n16783 = ~n15380 & n16718;
  assign n16788 = n16787 ^ n16783;
  assign n16789 = n16782 & ~n16788;
  assign n16791 = n16786 ^ n16716;
  assign n16790 = n16751 ^ n16746;
  assign n16792 = n16791 ^ n16790;
  assign n16793 = n16792 ^ n16731;
  assign n16794 = ~n15380 & n16793;
  assign n16795 = n16794 ^ n16792;
  assign n16796 = n15824 & n16795;
  assign n16797 = n16789 & ~n16796;
  assign n16798 = ~n16756 & n16797;
  assign n16799 = n16798 ^ n16601;
  assign n18738 = n16799 ^ x694;
  assign n17438 = n16803 & n16874;
  assign n17449 = n17433 ^ n16886;
  assign n17450 = n16904 & ~n17449;
  assign n17451 = n17450 ^ n16893;
  assign n17452 = n17451 ^ n16933;
  assign n17444 = n16893 & n16914;
  assign n17446 = n17445 ^ n17444;
  assign n17443 = n16884 ^ n16865;
  assign n17447 = n17446 ^ n17443;
  assign n17441 = n16882 ^ n16879;
  assign n17442 = n16916 & n17441;
  assign n17448 = n17447 ^ n17442;
  assign n17453 = n17452 ^ n17448;
  assign n17454 = n16803 & n17453;
  assign n17455 = n17454 ^ n17452;
  assign n17456 = ~n17440 & ~n17455;
  assign n17457 = ~n17438 & n17456;
  assign n17463 = n16891 ^ n16871;
  assign n17464 = ~n16801 & ~n17463;
  assign n17465 = n17464 ^ n16891;
  assign n17458 = n17439 ^ n16879;
  assign n17459 = n17458 ^ n16866;
  assign n17460 = n17459 ^ n16888;
  assign n17461 = n16801 & ~n17460;
  assign n17462 = n17461 ^ n16888;
  assign n17466 = n17465 ^ n17462;
  assign n17467 = ~n16802 & ~n17466;
  assign n17468 = n17467 ^ n17462;
  assign n17469 = n17457 & ~n17468;
  assign n17470 = ~n17437 & n17469;
  assign n17471 = n17470 ^ n14191;
  assign n18135 = n17471 ^ x644;
  assign n18197 = n17904 ^ x641;
  assign n18204 = ~n18135 & ~n18197;
  assign n18205 = n18204 ^ n18135;
  assign n17322 = n15425 & n17321;
  assign n17323 = n17322 ^ n15772;
  assign n17324 = n15775 & n17323;
  assign n17325 = ~n15741 & ~n17324;
  assign n18136 = n15427 & ~n15746;
  assign n18137 = n15426 & n15763;
  assign n18142 = n15381 & n15788;
  assign n18143 = n18142 ^ n15785;
  assign n18138 = n15797 ^ n15780;
  assign n18139 = n18138 ^ n15745;
  assign n18140 = ~n15381 & n18139;
  assign n18141 = n18140 ^ n18138;
  assign n18144 = n18143 ^ n18141;
  assign n18145 = ~n15425 & n18144;
  assign n18146 = n18145 ^ n18141;
  assign n18147 = ~n17595 & ~n18146;
  assign n18148 = ~n18137 & n18147;
  assign n18149 = ~n18136 & n18148;
  assign n18151 = n15772 ^ n15759;
  assign n18152 = n18151 ^ n15776;
  assign n18150 = n15781 ^ n15750;
  assign n18153 = n18152 ^ n18150;
  assign n18154 = ~n15425 & n18153;
  assign n18155 = n18154 ^ n18150;
  assign n18156 = ~n15381 & n18155;
  assign n18157 = n18149 & ~n18156;
  assign n18158 = n15819 & n18157;
  assign n18159 = n17325 & n18158;
  assign n18160 = n18159 ^ n14102;
  assign n18161 = n18160 ^ x643;
  assign n18163 = n17270 ^ n17029;
  assign n18164 = n18163 ^ n17013;
  assign n18165 = ~n16943 & ~n18164;
  assign n18166 = n18165 ^ n18163;
  assign n18167 = n16942 & ~n18166;
  assign n18169 = n17033 & n17273;
  assign n18168 = n16943 & n16999;
  assign n18170 = n18169 ^ n18168;
  assign n18171 = ~n18167 & ~n18170;
  assign n18172 = ~n17038 & n17044;
  assign n18173 = n17034 ^ n17018;
  assign n18174 = ~n17274 & n18173;
  assign n18182 = n17792 ^ n17018;
  assign n18181 = n17039 ^ n17012;
  assign n18183 = n18182 ^ n18181;
  assign n18184 = ~n16943 & n18183;
  assign n18185 = n18184 ^ n18181;
  assign n18175 = n17017 ^ n17014;
  assign n18176 = n18175 ^ n17009;
  assign n18177 = ~n16943 & n18176;
  assign n18178 = n18177 ^ n17009;
  assign n18179 = n18178 ^ n17004;
  assign n18180 = ~n18178 & ~n18179;
  assign n18186 = n18185 ^ n18180;
  assign n18187 = n17038 & ~n18186;
  assign n18188 = n18187 ^ n18180;
  assign n18189 = ~n17025 & n18188;
  assign n18190 = ~n18174 & n18189;
  assign n18191 = ~n18172 & n18190;
  assign n18192 = n18171 & n18191;
  assign n18193 = n17287 & n18192;
  assign n18194 = n18193 ^ n14136;
  assign n18195 = n18194 ^ x642;
  assign n18202 = ~n18161 & ~n18195;
  assign n18203 = n18202 ^ n18195;
  assign n18214 = n18203 ^ n18161;
  assign n18217 = ~n18205 & ~n18214;
  assign n17358 = n16450 ^ n16441;
  assign n17359 = ~n16463 & n17358;
  assign n17360 = n17359 ^ n16441;
  assign n17361 = ~n16462 & n17360;
  assign n17511 = ~n16432 & n16465;
  assign n17507 = ~n16427 & ~n16462;
  assign n17508 = n17507 ^ n16471;
  assign n17509 = n16477 & ~n17508;
  assign n17510 = n17509 ^ n16471;
  assign n17512 = n17511 ^ n17510;
  assign n17502 = n16488 ^ n16439;
  assign n17504 = n17503 ^ n16488;
  assign n17505 = n17502 & n17504;
  assign n17499 = n16440 ^ n16407;
  assign n17500 = ~n16463 & n17499;
  assign n17501 = n17500 ^ n16415;
  assign n17506 = n17505 ^ n17501;
  assign n17513 = n17512 ^ n17506;
  assign n17514 = ~n16467 & n17513;
  assign n17515 = ~n17361 & n17514;
  assign n17516 = n17515 ^ n14341;
  assign n18252 = n17516 ^ x645;
  assign n18253 = n17926 ^ x640;
  assign n18206 = n18205 ^ n18197;
  assign n18216 = ~n18203 & ~n18206;
  assign n18232 = n18216 ^ n18203;
  assign n18162 = n18135 & n18161;
  assign n18196 = n18195 ^ n18162;
  assign n18221 = n18196 & n18197;
  assign n18226 = n18221 ^ n18197;
  assign n18225 = n18217 ^ n18205;
  assign n18227 = n18226 ^ n18225;
  assign n18219 = n18202 ^ n18161;
  assign n18220 = ~n18206 & ~n18219;
  assign n18222 = n18221 ^ n18220;
  assign n18218 = n18217 ^ n18216;
  assign n18223 = n18222 ^ n18218;
  assign n18215 = ~n18206 & ~n18214;
  assign n18224 = n18223 ^ n18215;
  assign n18228 = n18227 ^ n18224;
  assign n18229 = n18228 ^ n18202;
  assign n18198 = n18197 ^ n18161;
  assign n18209 = n18198 ^ n18135;
  assign n18210 = n18209 ^ n18197;
  assign n18211 = ~n18198 & ~n18210;
  assign n18212 = n18211 ^ n18209;
  assign n18213 = ~n18195 & n18212;
  assign n18230 = n18229 ^ n18213;
  assign n18207 = n18206 ^ n18135;
  assign n18208 = ~n18203 & ~n18207;
  assign n18231 = n18230 ^ n18208;
  assign n18233 = n18232 ^ n18231;
  assign n18234 = n18233 ^ n18223;
  assign n18235 = n18234 ^ n18225;
  assign n18199 = n18198 ^ n18195;
  assign n18200 = n18199 ^ n18135;
  assign n18201 = ~n18196 & ~n18200;
  assign n18236 = n18235 ^ n18201;
  assign n18237 = n18236 ^ n18226;
  assign n18262 = n18237 ^ n18204;
  assign n18246 = n18203 ^ n18201;
  assign n18247 = n18246 ^ n18211;
  assign n18242 = n18231 ^ n18228;
  assign n18248 = n18247 ^ n18242;
  assign n18261 = n18248 ^ n18230;
  assign n18263 = n18262 ^ n18261;
  assign n18249 = n18248 ^ n18208;
  assign n18244 = n18195 ^ n18135;
  assign n18245 = n18244 ^ n18161;
  assign n18250 = n18249 ^ n18245;
  assign n18240 = n18233 ^ n18224;
  assign n18238 = n18237 ^ n18229;
  assign n18239 = n18238 ^ n18235;
  assign n18241 = n18240 ^ n18239;
  assign n18243 = n18242 ^ n18241;
  assign n18251 = n18250 ^ n18243;
  assign n18265 = n18263 ^ n18251;
  assign n18266 = n18265 ^ n18239;
  assign n18267 = n18266 ^ n18208;
  assign n18264 = n18263 ^ n18207;
  assign n18268 = n18267 ^ n18264;
  assign n18269 = n18268 ^ n18237;
  assign n18270 = n18269 ^ n18233;
  assign n18271 = ~n18253 & ~n18270;
  assign n18272 = n18271 ^ n18233;
  assign n18273 = n18252 & n18272;
  assign n18254 = n18252 & n18253;
  assign n18743 = n18254 & ~n18265;
  assign n18281 = n18253 ^ n18252;
  assign n18739 = n18239 ^ n18220;
  assign n18740 = ~n18252 & ~n18739;
  assign n18741 = n18740 ^ n18220;
  assign n18742 = n18281 & n18741;
  assign n18744 = n18743 ^ n18742;
  assign n18255 = n18254 ^ n18253;
  assign n18256 = n18255 ^ n18252;
  assign n18259 = ~n18235 & ~n18256;
  assign n18257 = n18256 ^ n18253;
  assign n18258 = n18251 & n18257;
  assign n18260 = n18259 ^ n18258;
  assign n18747 = n18235 ^ n18220;
  assign n18748 = n18252 & ~n18747;
  assign n18745 = ~n18243 & ~n18252;
  assign n18746 = n18745 ^ n18242;
  assign n18749 = n18748 ^ n18746;
  assign n18750 = n18253 & n18749;
  assign n18751 = n18750 ^ n18746;
  assign n18752 = n18213 ^ n18209;
  assign n18753 = n18752 ^ n18249;
  assign n18754 = n18753 ^ n18249;
  assign n18755 = ~n18252 & n18754;
  assign n18756 = n18755 ^ n18249;
  assign n18757 = n18281 & ~n18756;
  assign n18758 = n18757 ^ n18249;
  assign n18759 = ~n18751 & n18758;
  assign n18760 = ~n18260 & n18759;
  assign n18761 = ~n18744 & n18760;
  assign n18762 = ~n18273 & n18761;
  assign n18763 = ~n18217 & n18762;
  assign n18764 = n18763 ^ n15896;
  assign n18765 = n18764 ^ x699;
  assign n18766 = n18738 & ~n18765;
  assign n18767 = n18766 ^ n18738;
  assign n18768 = n18737 & n18767;
  assign n18769 = ~n18659 & ~n18735;
  assign n18770 = n18769 ^ n18735;
  assign n18772 = n18660 & n18693;
  assign n18792 = ~n18770 & n18772;
  assign n18793 = n18792 ^ n18772;
  assign n18782 = n18769 ^ n18659;
  assign n18790 = n18772 & ~n18782;
  assign n18771 = n18770 ^ n18659;
  assign n18776 = ~n18771 & n18772;
  assign n18791 = n18790 ^ n18776;
  assign n18794 = n18793 ^ n18791;
  assign n18795 = n18794 ^ n18769;
  assign n18773 = n18772 ^ n18693;
  assign n18788 = n18769 & n18773;
  assign n18774 = n18773 ^ n18660;
  assign n18786 = n18769 & ~n18774;
  assign n18789 = n18788 ^ n18786;
  assign n18796 = n18795 ^ n18789;
  assign n18784 = ~n18770 & n18773;
  assign n18783 = ~n18774 & ~n18782;
  assign n18785 = n18784 ^ n18783;
  assign n18787 = n18786 ^ n18785;
  assign n18797 = n18796 ^ n18787;
  assign n18778 = ~n18771 & n18773;
  assign n18779 = n18778 ^ n18771;
  assign n18775 = ~n18771 & ~n18774;
  assign n18777 = n18776 ^ n18775;
  assign n18780 = n18779 ^ n18777;
  assign n18781 = n18780 ^ n18775;
  assign n18798 = n18797 ^ n18781;
  assign n18799 = n18798 ^ n18781;
  assign n18800 = ~n18765 & n18799;
  assign n18801 = n18800 ^ n18781;
  assign n18802 = ~n18738 & ~n18801;
  assign n18803 = n18802 ^ n18781;
  assign n18804 = ~n18768 & n18803;
  assign n18805 = n18765 ^ n18738;
  assign n18816 = ~n18693 & ~n18735;
  assign n18814 = n18772 ^ n18660;
  assign n18815 = ~n18770 & n18814;
  assign n18817 = n18816 ^ n18815;
  assign n18813 = n18796 ^ n18786;
  assign n18818 = n18817 ^ n18813;
  assign n18808 = n18773 & ~n18782;
  assign n18809 = n18808 ^ n18782;
  assign n18807 = n18790 ^ n18783;
  assign n18810 = n18809 ^ n18807;
  assign n18812 = n18810 ^ n18789;
  assign n18819 = n18818 ^ n18812;
  assign n18806 = n18794 ^ n18784;
  assign n18811 = n18810 ^ n18806;
  assign n18820 = n18819 ^ n18811;
  assign n18821 = n18765 & n18820;
  assign n18822 = n18821 ^ n18811;
  assign n18823 = n18805 & ~n18822;
  assign n18824 = n18804 & ~n18823;
  assign n18827 = ~n18765 & n18792;
  assign n18825 = n18765 & n18791;
  assign n18826 = n18825 ^ n18790;
  assign n18828 = n18827 ^ n18826;
  assign n18829 = ~n18805 & n18828;
  assign n18830 = n18829 ^ n18826;
  assign n18831 = n18824 & ~n18830;
  assign n18836 = n18765 & n18788;
  assign n18832 = n18815 ^ n18790;
  assign n18833 = n18832 ^ n18792;
  assign n18834 = ~n18765 & n18833;
  assign n18835 = n18834 ^ n18792;
  assign n18837 = n18836 ^ n18835;
  assign n18838 = n18738 & n18837;
  assign n18839 = n18838 ^ n18835;
  assign n18840 = n18831 & ~n18839;
  assign n18845 = n18767 ^ n18765;
  assign n18846 = n18845 ^ n18738;
  assign n18847 = n18808 & ~n18846;
  assign n18841 = n18792 ^ n18780;
  assign n18842 = ~n18738 & ~n18841;
  assign n18843 = n18842 ^ n18792;
  assign n18844 = n18765 & n18843;
  assign n18848 = n18847 ^ n18844;
  assign n18849 = n18840 & ~n18848;
  assign n18850 = n18818 ^ n18778;
  assign n18851 = n18850 ^ n18808;
  assign n18852 = ~n18765 & n18851;
  assign n18853 = n18852 ^ n18808;
  assign n18854 = n18805 & n18853;
  assign n18855 = n18849 & ~n18854;
  assign n18856 = n18855 ^ n17067;
  assign n18857 = n18856 ^ x762;
  assign n18889 = n18476 & n18502;
  assign n18890 = n18889 ^ n18709;
  assign n18891 = n18475 ^ n18456;
  assign n18892 = ~n18402 & n18891;
  assign n18893 = n18892 ^ n18475;
  assign n18894 = n18453 & n18893;
  assign n18451 = ~n18406 & n18450;
  assign n18895 = n18405 & n18456;
  assign n18900 = n18695 ^ n18474;
  assign n18901 = n18900 ^ n18471;
  assign n18902 = ~n18402 & ~n18901;
  assign n18903 = n18902 ^ n18471;
  assign n18479 = n18478 ^ n18440;
  assign n18896 = n18479 ^ n18468;
  assign n18897 = n18896 ^ n18714;
  assign n18898 = n18402 & n18897;
  assign n18899 = n18898 ^ n18714;
  assign n18904 = n18903 ^ n18899;
  assign n18905 = n18904 ^ n18899;
  assign n18906 = n18699 & ~n18905;
  assign n18907 = n18906 ^ n18899;
  assign n18908 = ~n18453 & n18907;
  assign n18909 = n18908 ^ n18899;
  assign n18910 = ~n18895 & n18909;
  assign n18911 = ~n18451 & n18910;
  assign n18912 = ~n18894 & n18911;
  assign n18913 = ~n18890 & n18912;
  assign n18914 = n18705 & n18913;
  assign n18915 = n18914 ^ n16132;
  assign n18916 = n18915 ^ x722;
  assign n17833 = n17747 & ~n17832;
  assign n18917 = n18312 ^ n17835;
  assign n18926 = n18917 ^ n17820;
  assign n18927 = n18926 ^ n17825;
  assign n18928 = ~n17711 & n18927;
  assign n18918 = n18917 ^ n17865;
  assign n18919 = n17865 ^ n17711;
  assign n18920 = ~n17744 & n18919;
  assign n18921 = n18920 ^ n17711;
  assign n18922 = ~n18918 & n18921;
  assign n18923 = n18922 ^ n18917;
  assign n18924 = ~n17820 & ~n18923;
  assign n18925 = ~n17849 & n18924;
  assign n18929 = n18928 ^ n18925;
  assign n18930 = ~n17744 & ~n18929;
  assign n18931 = n18930 ^ n18925;
  assign n18315 = n18309 ^ n17829;
  assign n18932 = n18315 ^ n18312;
  assign n18933 = n18932 ^ n18629;
  assign n18934 = n18933 ^ n17830;
  assign n18935 = ~n17744 & n18934;
  assign n18936 = n18935 ^ n17830;
  assign n18937 = n17711 & n18936;
  assign n18938 = n18931 & ~n18937;
  assign n18939 = ~n18649 & n18938;
  assign n18940 = ~n17833 & n18939;
  assign n18941 = ~n18655 & n18940;
  assign n18942 = n18941 ^ n16830;
  assign n18943 = n18942 ^ x720;
  assign n18360 = n18015 ^ n17987;
  assign n18361 = n18360 ^ n18020;
  assign n18362 = ~n17889 & n18361;
  assign n18363 = n18362 ^ n18020;
  assign n18364 = n17906 & n18363;
  assign n18858 = n18023 & ~n18045;
  assign n18859 = n18012 ^ n18010;
  assign n18860 = n18000 & n18859;
  assign n18863 = n18019 ^ n17985;
  assign n18864 = n18045 & ~n18863;
  assign n18379 = n18012 ^ n17989;
  assign n18380 = ~n18000 & ~n18379;
  assign n18865 = ~n17987 & n18380;
  assign n18866 = ~n18864 & ~n18865;
  assign n18867 = n18016 & ~n18866;
  assign n18861 = n18026 ^ n17989;
  assign n18862 = ~n17889 & n18861;
  assign n18868 = n18867 ^ n18862;
  assign n18869 = n17906 & ~n18868;
  assign n18870 = n18869 ^ n18867;
  assign n18871 = ~n18860 & n18870;
  assign n18872 = ~n18858 & n18871;
  assign n18873 = n18360 ^ n18007;
  assign n18874 = n18873 ^ n17991;
  assign n18875 = ~n17905 & n18874;
  assign n18876 = n18875 ^ n18047;
  assign n18877 = n17906 & n18876;
  assign n18878 = n18877 ^ n18047;
  assign n18879 = n18872 & ~n18878;
  assign n18880 = n18011 ^ n18009;
  assign n18881 = ~n17889 & ~n18880;
  assign n18882 = n18881 ^ n18009;
  assign n18883 = n17905 & n18882;
  assign n18884 = n18879 & ~n18883;
  assign n18885 = ~n18364 & n18884;
  assign n18886 = ~n18049 & n18885;
  assign n18887 = n18886 ^ n15424;
  assign n18888 = n18887 ^ x719;
  assign n18951 = ~n18231 & ~n18256;
  assign n18277 = n18254 & n18268;
  assign n18952 = n18951 ^ n18277;
  assign n18953 = n18240 & n18257;
  assign n18954 = n18747 ^ n18263;
  assign n18955 = n18954 ^ n18215;
  assign n18956 = n18955 ^ n18221;
  assign n18957 = n18252 & n18956;
  assign n18958 = n18957 ^ n18221;
  assign n18959 = ~n18281 & n18958;
  assign n18965 = n18249 ^ n18217;
  assign n18966 = n18965 ^ n18201;
  assign n18967 = n18966 ^ n18251;
  assign n18968 = n18253 & ~n18967;
  assign n18969 = n18968 ^ n18251;
  assign n18960 = n18263 ^ n18237;
  assign n18961 = n18960 ^ n18208;
  assign n18962 = n18961 ^ n18261;
  assign n18963 = ~n18253 & n18962;
  assign n18964 = n18963 ^ n18261;
  assign n18970 = n18969 ^ n18964;
  assign n18971 = ~n18252 & n18970;
  assign n18972 = n18971 ^ n18964;
  assign n18973 = ~n18959 & ~n18972;
  assign n18974 = ~n18258 & n18973;
  assign n18975 = ~n18953 & n18974;
  assign n18976 = ~n18239 & ~n18281;
  assign n18977 = n18975 & ~n18976;
  assign n18978 = ~n18952 & n18977;
  assign n18979 = ~n18742 & n18978;
  assign n18980 = n18979 ^ n16858;
  assign n18981 = n18980 ^ x721;
  assign n18985 = n18888 & ~n18981;
  assign n18986 = ~n18943 & n18985;
  assign n18987 = ~n18916 & n18986;
  assign n18988 = n18987 ^ n18986;
  assign n18998 = n18988 ^ n18985;
  assign n18944 = n18916 & ~n18943;
  assign n18945 = n18944 ^ n18916;
  assign n18996 = n18945 & n18985;
  assign n18997 = n18996 ^ n18987;
  assign n18999 = n18998 ^ n18997;
  assign n18994 = n18945 ^ n18943;
  assign n18948 = ~n18888 & ~n18916;
  assign n18993 = n18943 & n18948;
  assign n18995 = n18994 ^ n18993;
  assign n19000 = n18999 ^ n18995;
  assign n18989 = n18988 ^ n18944;
  assign n18982 = ~n18943 & n18981;
  assign n18983 = ~n18916 & n18982;
  assign n18984 = n18983 ^ n18982;
  assign n18990 = n18989 ^ n18984;
  assign n18949 = n18948 ^ n18888;
  assign n18946 = n18888 & n18945;
  assign n18947 = n18946 ^ n18945;
  assign n18950 = n18949 ^ n18947;
  assign n18991 = n18990 ^ n18950;
  assign n18992 = n18991 ^ n18984;
  assign n19001 = n19000 ^ n18992;
  assign n17267 = n17266 ^ x658;
  assign n17362 = n16422 & n16466;
  assign n17363 = n16436 ^ n16403;
  assign n17364 = ~n16463 & ~n17363;
  assign n17365 = ~n17362 & ~n17364;
  assign n17370 = n16412 ^ n16408;
  assign n17368 = n16471 ^ n16402;
  assign n17369 = n17368 ^ n16415;
  assign n17371 = n17370 ^ n17369;
  assign n17367 = n17366 ^ n16420;
  assign n17372 = n17371 ^ n17367;
  assign n17373 = ~n16462 & n17372;
  assign n17374 = n17373 ^ n17367;
  assign n17375 = n16463 & n17374;
  assign n17376 = ~n16490 & ~n17375;
  assign n17377 = n17365 & n17376;
  assign n17378 = ~n16470 & n17377;
  assign n17379 = ~n17361 & n17378;
  assign n17380 = ~n16476 & n17379;
  assign n17381 = n17380 ^ n15645;
  assign n17382 = n17381 ^ x661;
  assign n17337 = n15785 ^ n15740;
  assign n17338 = n17337 ^ n15759;
  assign n17336 = n15797 ^ n15760;
  assign n17339 = n17338 ^ n17336;
  assign n17340 = n15425 & n17339;
  assign n17341 = n17340 ^ n17336;
  assign n17331 = n15794 ^ n15771;
  assign n17332 = n17331 ^ n15797;
  assign n17333 = n17332 ^ n15782;
  assign n17334 = n15425 & ~n17333;
  assign n17335 = n17334 ^ n15782;
  assign n17342 = n17341 ^ n17335;
  assign n17343 = n17342 ^ n17341;
  assign n17344 = ~n17330 & ~n17343;
  assign n17345 = n17344 ^ n17341;
  assign n17346 = n15381 & ~n17345;
  assign n17347 = n17346 ^ n17341;
  assign n17348 = ~n17327 & ~n17347;
  assign n17349 = ~n15769 & n17348;
  assign n17350 = n17325 & n17349;
  assign n17351 = ~n15757 & n17350;
  assign n17352 = ~n17320 & n17351;
  assign n17353 = n17352 ^ n15671;
  assign n17354 = n17353 ^ x660;
  assign n17356 = n17158 ^ x662;
  assign n17315 = n17314 ^ x659;
  assign n17355 = n17354 ^ n17315;
  assign n17357 = n17356 ^ n17355;
  assign n17397 = ~n17354 & ~n17357;
  assign n17398 = n17397 ^ n17356;
  assign n17399 = ~n17382 & ~n17398;
  assign n17400 = n17399 ^ n17357;
  assign n17268 = n17113 ^ x663;
  assign n19014 = n17400 ^ n17268;
  assign n19007 = ~n17356 & n17382;
  assign n19008 = n19007 ^ n17354;
  assign n19009 = ~n17315 & ~n19008;
  assign n17383 = n17382 ^ n17356;
  assign n19010 = n19009 ^ n17383;
  assign n19011 = n19010 ^ n17400;
  assign n19012 = ~n17268 & n19011;
  assign n19013 = n19012 ^ n19010;
  assign n19015 = n19014 ^ n19013;
  assign n19016 = n19015 ^ n19010;
  assign n17388 = n17382 ^ n17354;
  assign n17393 = ~n17355 & ~n17382;
  assign n17394 = n17393 ^ n17356;
  assign n17395 = n17388 & n17394;
  assign n17426 = n17395 ^ n17355;
  assign n19004 = n17426 ^ n17268;
  assign n17421 = n17356 ^ n17315;
  assign n17422 = n17356 & ~n17388;
  assign n17423 = n17422 ^ n17354;
  assign n17424 = ~n17421 & ~n17423;
  assign n17420 = n17382 ^ n17355;
  assign n17425 = n17424 ^ n17420;
  assign n17427 = n17426 ^ n17425;
  assign n19002 = n17268 & n17427;
  assign n19003 = n19002 ^ n17425;
  assign n19005 = n19004 ^ n19003;
  assign n19006 = n19005 ^ n17425;
  assign n19017 = n19016 ^ n19006;
  assign n19018 = n17267 & n19017;
  assign n19019 = n19018 ^ n19006;
  assign n19020 = n19019 ^ n15732;
  assign n19021 = n19020 ^ x718;
  assign n17162 = n17126 & n17161;
  assign n17184 = n17183 ^ n17162;
  assign n18520 = n17176 & n17192;
  assign n18517 = n17160 ^ n17159;
  assign n18518 = n16941 & ~n18517;
  assign n18519 = n17194 & n18518;
  assign n18521 = n18520 ^ n18519;
  assign n19022 = n17118 & ~n18517;
  assign n19023 = n17166 ^ n17126;
  assign n19024 = ~n17160 & n19023;
  assign n17215 = n17204 ^ n17179;
  assign n19025 = n19024 ^ n17215;
  assign n19026 = n17159 & ~n19025;
  assign n19027 = n19026 ^ n17215;
  assign n19028 = ~n19022 & n19027;
  assign n19029 = n17159 & n17170;
  assign n17225 = n17160 & n17224;
  assign n19030 = n19029 ^ n17225;
  assign n19031 = n19028 & ~n19030;
  assign n19032 = ~n18688 & n19031;
  assign n19033 = ~n18521 & n19032;
  assign n19034 = ~n17184 & n19033;
  assign n19035 = ~n18516 & n19034;
  assign n19036 = n19035 ^ n16162;
  assign n19037 = n19036 ^ x723;
  assign n19038 = n19021 & ~n19037;
  assign n19039 = n19038 ^ n19021;
  assign n19040 = n19039 ^ n19037;
  assign n19041 = n19040 ^ n19021;
  assign n19042 = ~n19001 & ~n19041;
  assign n19043 = n18947 & n18981;
  assign n19044 = n19043 ^ n18947;
  assign n19045 = ~n19041 & n19044;
  assign n19050 = n18996 ^ n18946;
  assign n19051 = n19050 ^ n18999;
  assign n19046 = n18948 & n18982;
  assign n19047 = n19046 ^ n18948;
  assign n19048 = n19047 ^ n18993;
  assign n19049 = n19048 ^ n19044;
  assign n19052 = n19051 ^ n19049;
  assign n19053 = n19021 & n19052;
  assign n19054 = n19053 ^ n19049;
  assign n19055 = n19037 & n19054;
  assign n19056 = n19046 ^ n18983;
  assign n19057 = n19056 ^ n18988;
  assign n19058 = n19057 ^ n18991;
  assign n19059 = n19037 & ~n19058;
  assign n19060 = n19059 ^ n18991;
  assign n19061 = n19041 ^ n19039;
  assign n19062 = ~n19060 & n19061;
  assign n19063 = ~n19055 & ~n19062;
  assign n19064 = n19046 ^ n18996;
  assign n19065 = n19040 & n19064;
  assign n19076 = n19000 ^ n18991;
  assign n19077 = n19040 & ~n19076;
  assign n19067 = n19057 ^ n18999;
  assign n19068 = n19067 ^ n18987;
  assign n19066 = n19048 ^ n18996;
  assign n19069 = n19068 ^ n19066;
  assign n19070 = n19021 & n19069;
  assign n19071 = n19070 ^ n19066;
  assign n19072 = n19071 ^ n19043;
  assign n19073 = ~n19071 & ~n19072;
  assign n19074 = ~n19037 & n19073;
  assign n19075 = n19074 ^ n19037;
  assign n19078 = n19077 ^ n19075;
  assign n19082 = ~n18981 & n18993;
  assign n19083 = n19082 ^ n18993;
  assign n19079 = n19046 ^ n18990;
  assign n19080 = n19079 ^ n18992;
  assign n19081 = n19080 ^ n19044;
  assign n19084 = n19083 ^ n19081;
  assign n19085 = n19037 & ~n19084;
  assign n19086 = n19085 ^ n19083;
  assign n19087 = n19021 & n19086;
  assign n19088 = n19078 & ~n19087;
  assign n19089 = n19082 ^ n19048;
  assign n19090 = ~n19037 & n19089;
  assign n19091 = n19090 ^ n19048;
  assign n19092 = n19021 & n19091;
  assign n19093 = n19088 & ~n19092;
  assign n19094 = ~n19065 & n19093;
  assign n19095 = n19057 ^ n19000;
  assign n19096 = ~n19037 & n19095;
  assign n19097 = n19096 ^ n19000;
  assign n19098 = ~n19061 & n19097;
  assign n19099 = n19094 & ~n19098;
  assign n19100 = n19063 & n19099;
  assign n19101 = ~n19045 & n19100;
  assign n19102 = ~n19042 & n19101;
  assign n19103 = n19102 ^ n16940;
  assign n19104 = n19103 ^ x763;
  assign n19105 = n18857 & ~n19104;
  assign n19106 = n19105 ^ n18857;
  assign n17410 = n17398 ^ n17355;
  assign n17411 = n17410 ^ n17356;
  assign n17412 = n17382 & ~n17411;
  assign n17413 = n17412 ^ n17357;
  assign n17408 = n17356 ^ n17354;
  assign n17389 = n17382 ^ n17315;
  assign n17390 = ~n17356 & ~n17389;
  assign n17391 = n17390 ^ n17315;
  assign n17392 = ~n17388 & n17391;
  assign n17409 = n17408 ^ n17392;
  assign n17414 = n17413 ^ n17409;
  assign n17415 = n17268 & ~n17414;
  assign n17416 = n17415 ^ n17409;
  assign n17396 = n17395 ^ n17392;
  assign n17401 = n17400 ^ n17396;
  assign n17384 = n17354 & ~n17383;
  assign n17385 = n17384 ^ n17382;
  assign n17386 = ~n17357 & ~n17385;
  assign n17387 = n17386 ^ n17356;
  assign n17402 = n17401 ^ n17387;
  assign n17403 = ~n17268 & n17402;
  assign n17404 = n17403 ^ n17387;
  assign n17405 = n17404 ^ n17268;
  assign n17406 = n17405 ^ n17401;
  assign n17407 = n17406 ^ n17387;
  assign n17417 = n17416 ^ n17407;
  assign n17418 = n17267 & ~n17417;
  assign n17419 = n17418 ^ n17416;
  assign n17428 = n17427 ^ n17383;
  assign n17429 = n17428 ^ n17402;
  assign n17430 = n17419 & n17429;
  assign n17431 = n17430 ^ n16461;
  assign n17432 = n17431 ^ x689;
  assign n17472 = n17471 ^ x646;
  assign n17498 = n17497 ^ x651;
  assign n17517 = n17516 ^ x647;
  assign n17518 = n16036 ^ n16023;
  assign n17519 = ~n15997 & ~n17518;
  assign n17520 = n16034 ^ n16003;
  assign n17521 = n17520 ^ n16008;
  assign n17522 = ~n16002 & ~n17521;
  assign n17523 = n17522 ^ n16008;
  assign n17524 = ~n17519 & ~n17523;
  assign n17525 = n15932 & ~n15935;
  assign n17526 = n17525 ^ n16005;
  assign n17527 = n15984 & n17526;
  assign n17528 = n17524 & ~n17527;
  assign n17529 = n16051 ^ n16013;
  assign n17530 = ~n15935 & ~n17529;
  assign n17531 = n17530 ^ n16013;
  assign n17532 = n17528 & n17531;
  assign n17533 = ~n17130 & n17532;
  assign n17534 = ~n16001 & n17533;
  assign n17535 = ~n16056 & n17534;
  assign n17536 = n17535 ^ n14632;
  assign n17537 = n17536 ^ x648;
  assign n17538 = n17517 & ~n17537;
  assign n17539 = n17538 ^ n17517;
  assign n17546 = n16292 ^ n16286;
  assign n17547 = ~n17545 & ~n17546;
  assign n17550 = n17546 ^ n16274;
  assign n17549 = n16284 ^ n16227;
  assign n17551 = n17550 ^ n17549;
  assign n17548 = n17244 ^ n16258;
  assign n17552 = n17551 ^ n17548;
  assign n17553 = n16093 & ~n17552;
  assign n17554 = n17553 ^ n17548;
  assign n17555 = n17554 ^ n17239;
  assign n17556 = ~n16134 & ~n17555;
  assign n17557 = n17556 ^ n17239;
  assign n17558 = ~n17547 & n17557;
  assign n17559 = n16280 ^ n16231;
  assign n17560 = n16093 & n17559;
  assign n17561 = n17560 ^ n16231;
  assign n17562 = n16134 & n17561;
  assign n17563 = n17558 & ~n17562;
  assign n17564 = ~n17544 & n17563;
  assign n17565 = ~n16278 & n17564;
  assign n17566 = n17565 ^ n14602;
  assign n17567 = n17566 ^ x649;
  assign n17599 = n17598 ^ x650;
  assign n17600 = n17567 & ~n17599;
  assign n17601 = n17600 ^ n17567;
  assign n17626 = n17539 & n17601;
  assign n17602 = n17601 ^ n17599;
  assign n17540 = n17539 ^ n17537;
  assign n17605 = n17540 ^ n17517;
  assign n17609 = n17602 & ~n17605;
  assign n17627 = n17626 ^ n17609;
  assign n17628 = ~n17498 & n17627;
  assign n17629 = n17628 ^ n17626;
  assign n17616 = ~n17517 & ~n17567;
  assign n17617 = n17616 ^ n17540;
  assign n17613 = n17609 ^ n17605;
  assign n17611 = n17600 & ~n17605;
  assign n17606 = n17601 & ~n17605;
  assign n17612 = n17611 ^ n17606;
  assign n17614 = n17613 ^ n17612;
  assign n17608 = n17540 & n17600;
  assign n17610 = n17609 ^ n17608;
  assign n17615 = n17614 ^ n17610;
  assign n17618 = n17617 ^ n17615;
  assign n17619 = n17618 ^ n17611;
  assign n17603 = n17602 ^ n17567;
  assign n17604 = n17540 & ~n17603;
  assign n17607 = n17606 ^ n17604;
  assign n17620 = n17619 ^ n17607;
  assign n17621 = n17620 ^ n17517;
  assign n17622 = n17621 ^ n17615;
  assign n17623 = n17622 ^ n17606;
  assign n17624 = ~n17498 & ~n17623;
  assign n17625 = n17624 ^ n17606;
  assign n17630 = n17629 ^ n17625;
  assign n17631 = ~n17472 & n17630;
  assign n17632 = n17631 ^ n17625;
  assign n17637 = n17618 ^ n17614;
  assign n17633 = ~n17472 & ~n17498;
  assign n17638 = n17633 ^ n17498;
  assign n17639 = n17637 & ~n17638;
  assign n17634 = n17633 ^ n17472;
  assign n17635 = n17538 & n17602;
  assign n17636 = ~n17634 & n17635;
  assign n17640 = n17639 ^ n17636;
  assign n17642 = n17538 & n17600;
  assign n17641 = n17539 & n17602;
  assign n17643 = n17642 ^ n17641;
  assign n17644 = ~n17634 & n17643;
  assign n17646 = n17612 ^ n17601;
  assign n17645 = n17626 ^ n17619;
  assign n17647 = n17646 ^ n17645;
  assign n17648 = n17647 ^ n17642;
  assign n17649 = n17648 ^ n17538;
  assign n17650 = n17649 ^ n17635;
  assign n17651 = n17650 ^ n17619;
  assign n17652 = n17633 & n17651;
  assign n17653 = n17498 ^ n17472;
  assign n17659 = n17635 ^ n17517;
  assign n17655 = n17539 & n17600;
  assign n17656 = n17655 ^ n17647;
  assign n17657 = n17656 ^ n17643;
  assign n17654 = n17650 ^ n17626;
  assign n17658 = n17657 ^ n17654;
  assign n17660 = n17659 ^ n17658;
  assign n17661 = n17660 ^ n17647;
  assign n17662 = n17498 & ~n17661;
  assign n17663 = n17662 ^ n17660;
  assign n17664 = ~n17653 & n17663;
  assign n17675 = n17656 ^ n17641;
  assign n17672 = n17660 ^ n17635;
  assign n17673 = n17672 ^ n17642;
  assign n17674 = n17673 ^ n17650;
  assign n17676 = n17675 ^ n17674;
  assign n17677 = n17472 & n17676;
  assign n17678 = n17677 ^ n17675;
  assign n17667 = n17650 ^ n17611;
  assign n17668 = n17667 ^ n17610;
  assign n17665 = n17660 ^ n17641;
  assign n17666 = n17665 ^ n17626;
  assign n17669 = n17668 ^ n17666;
  assign n17670 = ~n17472 & ~n17669;
  assign n17671 = n17670 ^ n17666;
  assign n17679 = n17678 ^ n17671;
  assign n17680 = n17498 & ~n17679;
  assign n17681 = n17680 ^ n17678;
  assign n17682 = ~n17664 & n17681;
  assign n17683 = ~n17652 & n17682;
  assign n17684 = ~n17644 & n17683;
  assign n17685 = n17615 ^ n17608;
  assign n17686 = n17498 & ~n17685;
  assign n17687 = n17686 ^ n17608;
  assign n17688 = n17472 & n17687;
  assign n17689 = n17684 & ~n17688;
  assign n17690 = ~n17640 & n17689;
  assign n17691 = ~n17632 & n17690;
  assign n17692 = n17691 ^ n16570;
  assign n17693 = n17692 ^ x690;
  assign n17694 = n17432 & ~n17693;
  assign n17695 = n17694 ^ n17432;
  assign n16800 = n16799 ^ x692;
  assign n17189 = n17161 & ~n17168;
  assign n17207 = n17206 ^ n17202;
  assign n17208 = n17207 ^ n17199;
  assign n17209 = n17192 & ~n17208;
  assign n17210 = n17121 & ~n17163;
  assign n17211 = n17210 ^ n17197;
  assign n17212 = n17159 & ~n17211;
  assign n17213 = n17212 ^ n17171;
  assign n17214 = ~n17160 & n17213;
  assign n17220 = n17070 ^ n17068;
  assign n17221 = n17220 ^ n17206;
  assign n17222 = n17221 ^ n17185;
  assign n17223 = n17160 & n17222;
  assign n17226 = n17225 ^ n17223;
  assign n17227 = n17226 ^ n17204;
  assign n17216 = n17215 ^ n17195;
  assign n17217 = n17216 ^ n17124;
  assign n17218 = ~n17160 & n17217;
  assign n17219 = n17218 ^ n17124;
  assign n17228 = n17227 ^ n17219;
  assign n17229 = n17159 & n17228;
  assign n17230 = n17229 ^ n17219;
  assign n17231 = ~n17214 & ~n17230;
  assign n17232 = ~n17209 & n17231;
  assign n17233 = ~n17189 & n17232;
  assign n17234 = ~n17188 & n17233;
  assign n17235 = ~n17184 & n17234;
  assign n17236 = n17235 ^ n16626;
  assign n17237 = n17236 ^ x691;
  assign n17238 = n16800 & ~n17237;
  assign n17707 = n17238 ^ n17237;
  assign n17708 = n17695 & ~n17707;
  assign n17709 = n17708 ^ n17695;
  assign n17704 = n17238 ^ n16800;
  assign n17705 = n17695 & n17704;
  assign n17701 = n17238 & n17694;
  assign n17696 = n17695 ^ n17693;
  assign n17700 = n17238 & n17696;
  assign n17702 = n17701 ^ n17700;
  assign n17697 = n17696 ^ n17432;
  assign n17698 = n17238 & ~n17697;
  assign n17699 = n17698 ^ n17238;
  assign n17703 = n17702 ^ n17699;
  assign n17706 = n17705 ^ n17703;
  assign n17710 = n17709 ^ n17706;
  assign n17838 = n17837 ^ n17822;
  assign n17841 = n17840 ^ n17838;
  assign n17842 = n17711 & n17841;
  assign n17843 = n17842 ^ n17840;
  assign n17844 = n17744 & n17843;
  assign n17873 = n17864 ^ n17837;
  assign n17868 = n17867 ^ n17848;
  assign n17875 = n17873 ^ n17868;
  assign n17876 = n17875 ^ n17855;
  assign n17874 = n17873 ^ n17831;
  assign n17877 = n17876 ^ n17874;
  assign n17878 = n17711 & ~n17877;
  assign n17879 = n17878 ^ n17876;
  assign n17869 = n17868 ^ n17836;
  assign n17861 = n17847 ^ n17826;
  assign n17870 = n17869 ^ n17861;
  assign n17871 = ~n17711 & ~n17870;
  assign n17872 = n17871 ^ n17861;
  assign n17880 = n17879 ^ n17872;
  assign n17881 = ~n17744 & ~n17880;
  assign n17882 = n17881 ^ n17872;
  assign n17883 = ~n17860 & ~n17882;
  assign n17884 = ~n17854 & n17883;
  assign n17885 = ~n17844 & n17884;
  assign n17886 = ~n17833 & n17885;
  assign n17887 = n17886 ^ n16372;
  assign n17888 = n17887 ^ x688;
  assign n18064 = n18063 ^ x693;
  assign n18065 = ~n17888 & ~n18064;
  assign n18066 = n18065 ^ n17888;
  assign n18067 = n18066 ^ n18064;
  assign n18068 = n18067 ^ n17888;
  assign n18069 = n17710 & ~n18068;
  assign n18070 = n17708 ^ n17701;
  assign n18071 = ~n18066 & n18070;
  assign n18072 = n17707 ^ n16800;
  assign n18073 = n17694 & n18072;
  assign n18074 = n18065 & n18073;
  assign n18080 = n17696 & n18072;
  assign n18081 = n18080 ^ n17696;
  assign n18078 = n17696 & ~n17707;
  assign n18079 = n18078 ^ n17700;
  assign n18082 = n18081 ^ n18079;
  assign n18077 = ~n17697 & n18072;
  assign n18083 = n18082 ^ n18077;
  assign n18075 = n18073 ^ n17700;
  assign n18076 = n18075 ^ n17703;
  assign n18084 = n18083 ^ n18076;
  assign n18085 = ~n18066 & n18084;
  assign n18087 = n17694 & ~n17707;
  assign n18088 = n18087 ^ n17705;
  assign n18089 = n18088 ^ n17698;
  assign n18086 = ~n17697 & n17704;
  assign n18090 = n18089 ^ n18086;
  assign n18091 = ~n18068 & n18090;
  assign n18092 = n17694 & n17704;
  assign n18093 = n18092 ^ n17708;
  assign n18094 = n18093 ^ n17705;
  assign n18095 = n18065 & n18094;
  assign n18096 = n17710 ^ n17705;
  assign n18097 = n18096 ^ n18087;
  assign n18098 = n18097 ^ n18092;
  assign n18099 = n18098 ^ n18079;
  assign n18100 = n18099 ^ n18079;
  assign n18101 = n17888 & n18100;
  assign n18102 = n18101 ^ n18079;
  assign n18103 = n18064 & n18102;
  assign n18104 = n18103 ^ n18079;
  assign n18105 = ~n18095 & ~n18104;
  assign n18106 = ~n18091 & n18105;
  assign n18107 = ~n18085 & n18106;
  assign n18108 = ~n18074 & n18107;
  assign n18109 = n18064 ^ n17888;
  assign n18110 = n18080 ^ n17698;
  assign n18111 = n18064 & n18110;
  assign n18112 = n18111 ^ n18080;
  assign n18113 = ~n18109 & n18112;
  assign n18114 = n18108 & ~n18113;
  assign n18115 = n17703 ^ n17698;
  assign n18116 = ~n17888 & n18115;
  assign n18117 = n18116 ^ n17703;
  assign n18118 = ~n18064 & n18117;
  assign n18119 = n18114 & ~n18118;
  assign n18120 = ~n18071 & n18119;
  assign n18126 = n18078 ^ n17710;
  assign n18127 = n17888 & n18126;
  assign n18128 = n18127 ^ n17710;
  assign n18129 = n18064 & n18128;
  assign n18122 = n18086 ^ n17697;
  assign n18121 = n18077 ^ n17698;
  assign n18123 = n18122 ^ n18121;
  assign n18124 = n18123 ^ n18082;
  assign n18125 = ~n18067 & ~n18124;
  assign n18130 = n18129 ^ n18125;
  assign n18131 = n18120 & ~n18130;
  assign n18132 = ~n18069 & n18131;
  assign n18133 = n18132 ^ n17113;
  assign n18134 = n18133 ^ x761;
  assign n18320 = n17876 ^ n17857;
  assign n18321 = ~n17711 & ~n18320;
  assign n18322 = n18321 ^ n17876;
  assign n18316 = n18315 ^ n17873;
  assign n18314 = n17868 ^ n17864;
  assign n18317 = n18316 ^ n18314;
  assign n18318 = ~n17711 & ~n18317;
  assign n18319 = n18318 ^ n18314;
  assign n18323 = n18322 ^ n18319;
  assign n18324 = ~n17745 & ~n18323;
  assign n18325 = n18324 ^ n18322;
  assign n18326 = ~n18313 & n18325;
  assign n18327 = ~n17844 & n18326;
  assign n18328 = ~n18311 & n18327;
  assign n18329 = n18328 ^ n14066;
  assign n18330 = n18329 ^ x706;
  assign n18365 = ~n17889 & n18012;
  assign n18366 = n18365 ^ n18007;
  assign n18367 = n17906 & n18366;
  assign n18368 = n18367 ^ n18007;
  assign n18370 = n18001 & n18005;
  assign n18369 = n17889 & n18008;
  assign n18371 = n18370 ^ n18369;
  assign n18372 = ~n18368 & ~n18371;
  assign n18373 = n18019 & ~n18045;
  assign n18374 = n18047 ^ n18023;
  assign n18375 = n18000 & n18374;
  assign n18376 = n18022 ^ n18019;
  assign n18377 = n18376 ^ n18007;
  assign n18378 = n17999 & n18377;
  assign n18385 = n18038 ^ n17994;
  assign n18386 = n18385 ^ n17987;
  assign n18381 = n18016 ^ n17989;
  assign n18382 = n18045 & n18381;
  assign n18383 = ~n18380 & ~n18382;
  assign n18384 = ~n18014 & ~n18383;
  assign n18387 = n18386 ^ n18384;
  assign n18388 = n18387 ^ n18384;
  assign n18389 = n17889 & ~n18388;
  assign n18390 = n18389 ^ n18384;
  assign n18391 = n17906 & ~n18390;
  assign n18392 = n18391 ^ n18384;
  assign n18393 = ~n18378 & n18392;
  assign n18394 = ~n17998 & n18393;
  assign n18395 = ~n18375 & n18394;
  assign n18396 = ~n18373 & n18395;
  assign n18397 = n18372 & n18396;
  assign n18398 = ~n18046 & n18397;
  assign n18399 = ~n18364 & n18398;
  assign n18400 = n18399 ^ n14908;
  assign n18401 = n18400 ^ x709;
  assign n18523 = n17192 & ~n18522;
  assign n18524 = n17202 ^ n17176;
  assign n18525 = n18524 ^ n17222;
  assign n18526 = n17190 & ~n18525;
  assign n18527 = n17199 ^ n17191;
  assign n18528 = n17196 ^ n17161;
  assign n18529 = ~n17191 & ~n18528;
  assign n18530 = n18529 ^ n17161;
  assign n18531 = ~n18527 & ~n18530;
  assign n18532 = n18531 ^ n17199;
  assign n18534 = n17178 ^ n17175;
  assign n18535 = n17175 ^ n17160;
  assign n18536 = n18517 & n18535;
  assign n18537 = n18536 ^ n17160;
  assign n18538 = n18534 & ~n18537;
  assign n18539 = n18538 ^ n17178;
  assign n18540 = n17179 & ~n18539;
  assign n18533 = ~n17160 & ~n17172;
  assign n18541 = n18540 ^ n18533;
  assign n18542 = n18517 & ~n18541;
  assign n18543 = n18542 ^ n18540;
  assign n18544 = ~n18532 & n18543;
  assign n18547 = n17160 & n17205;
  assign n18545 = ~n16941 & n17192;
  assign n18546 = ~n17193 & n18545;
  assign n18548 = n18547 ^ n18546;
  assign n18549 = n18544 & ~n18548;
  assign n18550 = ~n18526 & n18549;
  assign n18551 = ~n18523 & n18550;
  assign n18552 = ~n18521 & n18551;
  assign n18553 = ~n18516 & n18552;
  assign n18554 = n18553 ^ n15329;
  assign n18555 = n18554 ^ x708;
  assign n18580 = ~n18401 & n18555;
  assign n18560 = n18401 ^ x708;
  assign n18561 = n18560 ^ n18554;
  assign n18588 = n18580 ^ n18561;
  assign n18447 = ~n18406 & n18446;
  assign n18449 = ~n18406 & n18448;
  assign n18452 = n18451 ^ n18449;
  assign n18485 = n18461 ^ n18458;
  assign n18486 = n18402 & n18485;
  assign n18487 = n18486 ^ n18461;
  assign n18480 = n18479 ^ n18474;
  assign n18481 = n18480 ^ n18466;
  assign n18465 = n18464 ^ n18454;
  assign n18482 = n18481 ^ n18465;
  assign n18483 = ~n18402 & n18482;
  assign n18484 = n18483 ^ n18465;
  assign n18488 = n18487 ^ n18484;
  assign n18489 = n18453 & ~n18488;
  assign n18490 = n18489 ^ n18487;
  assign n18491 = ~n18452 & ~n18490;
  assign n18492 = ~n18447 & n18491;
  assign n18493 = n18475 ^ n18462;
  assign n18495 = n18494 ^ n18493;
  assign n18496 = n18402 & n18495;
  assign n18497 = n18496 ^ n18494;
  assign n18498 = n18403 & ~n18497;
  assign n18499 = n18492 & ~n18498;
  assign n18503 = n18470 & ~n18502;
  assign n18501 = n18500 ^ n18478;
  assign n18504 = n18503 ^ n18501;
  assign n18505 = ~n18405 & ~n18504;
  assign n18506 = n18505 ^ n18501;
  assign n18507 = n18499 & n18506;
  assign n18508 = ~n18441 & n18507;
  assign n18509 = n18508 ^ n15096;
  assign n18510 = n18509 ^ x710;
  assign n18587 = ~n18510 & ~n18555;
  assign n18589 = n18588 ^ n18587;
  assign n18558 = n18510 ^ n18401;
  assign n18590 = n18589 ^ n18558;
  assign n18581 = ~n18510 & n18580;
  assign n18591 = n18590 ^ n18581;
  assign n18601 = n18591 ^ n18561;
  assign n18602 = n18601 ^ n18580;
  assign n18511 = n18401 & n18510;
  assign n18582 = n18581 ^ n18511;
  assign n18603 = n18602 ^ n18582;
  assign n18604 = n18603 ^ n18587;
  assign n18331 = ~n17614 & ~n17634;
  assign n18332 = n17660 ^ n17622;
  assign n18333 = ~n17472 & ~n18332;
  assign n18334 = n18333 ^ n17660;
  assign n18335 = n17498 & n18334;
  assign n18336 = ~n18331 & ~n18335;
  assign n18337 = n17655 ^ n17635;
  assign n18338 = n17633 & n18337;
  assign n18339 = n17675 ^ n17667;
  assign n18340 = ~n17638 & n18339;
  assign n18344 = ~n17472 & n17612;
  assign n18342 = n17618 ^ n17608;
  assign n18341 = n17643 ^ n17604;
  assign n18343 = n18342 ^ n18341;
  assign n18345 = n18344 ^ n18343;
  assign n18346 = n17653 & ~n18345;
  assign n18347 = n18346 ^ n18343;
  assign n18348 = ~n18340 & n18347;
  assign n18349 = ~n18338 & n18348;
  assign n18350 = n17673 ^ n17635;
  assign n18351 = ~n17472 & n18350;
  assign n18352 = n18351 ^ n17635;
  assign n18353 = n17498 & n18352;
  assign n18354 = n18349 & ~n18353;
  assign n18355 = ~n17639 & n18354;
  assign n18356 = n18336 & n18355;
  assign n18357 = ~n17632 & n18356;
  assign n18358 = n18357 ^ n14749;
  assign n18359 = n18358 ^ x707;
  assign n18610 = n18359 & n18602;
  assign n18564 = n18555 ^ n18510;
  assign n18565 = n18564 ^ n18359;
  assign n18572 = n18510 ^ n18359;
  assign n18573 = ~n18565 & ~n18572;
  assign n18605 = n18573 ^ n18565;
  assign n18606 = n18605 ^ n18510;
  assign n18611 = n18610 ^ n18606;
  assign n18607 = n18401 & ~n18606;
  assign n18608 = n18607 ^ n18565;
  assign n18562 = n18555 ^ n18359;
  assign n18563 = ~n18510 & n18562;
  assign n18566 = n18565 ^ n18563;
  assign n18567 = n18566 ^ n18401;
  assign n18568 = ~n18555 & ~n18567;
  assign n18569 = n18568 ^ n18555;
  assign n18592 = n18591 ^ n18569;
  assign n18583 = n18359 & n18582;
  assign n18584 = n18583 ^ n18511;
  assign n18570 = n18569 ^ n18359;
  assign n18577 = n18566 ^ n18510;
  assign n18578 = ~n18570 & n18577;
  assign n18579 = n18578 ^ n18563;
  assign n18585 = n18584 ^ n18579;
  assign n18574 = n18573 ^ n18510;
  assign n18575 = ~n18401 & ~n18574;
  assign n18576 = n18575 ^ n18565;
  assign n18586 = n18585 ^ n18576;
  assign n18593 = n18592 ^ n18586;
  assign n18512 = n18511 ^ n18510;
  assign n18556 = n18555 ^ n18512;
  assign n18571 = n18570 ^ n18556;
  assign n18594 = n18593 ^ n18571;
  assign n18595 = n18594 ^ n18510;
  assign n18596 = n18561 & n18595;
  assign n18597 = n18596 ^ n18562;
  assign n18609 = n18608 ^ n18597;
  assign n18612 = n18611 ^ n18609;
  assign n18613 = n18604 & ~n18612;
  assign n18614 = n18613 ^ n18580;
  assign n18615 = n18614 ^ n18608;
  assign n18616 = ~n18330 & n18615;
  assign n18617 = n18616 ^ n18608;
  assign n18274 = n18234 & n18255;
  assign n18275 = n18217 & ~n18256;
  assign n18276 = ~n18235 & n18257;
  assign n18278 = n18220 & ~n18257;
  assign n18279 = n18255 & n18267;
  assign n18280 = ~n18278 & ~n18279;
  assign n18291 = n18224 ^ n18218;
  assign n18292 = n18252 & n18291;
  assign n18283 = n18265 ^ n18249;
  assign n18282 = n18263 ^ n18231;
  assign n18284 = n18283 ^ n18282;
  assign n18285 = n18283 ^ n18252;
  assign n18286 = n18281 & n18285;
  assign n18287 = n18286 ^ n18252;
  assign n18288 = n18284 & ~n18287;
  assign n18289 = n18288 ^ n18282;
  assign n18290 = n18228 & ~n18289;
  assign n18293 = n18292 ^ n18290;
  assign n18294 = n18281 & ~n18293;
  assign n18295 = n18294 ^ n18290;
  assign n18296 = n18280 & n18295;
  assign n18297 = ~n18277 & n18296;
  assign n18298 = ~n18276 & n18297;
  assign n18299 = ~n18275 & n18298;
  assign n18300 = n18224 & ~n18252;
  assign n18301 = n18300 ^ n18223;
  assign n18302 = n18253 & n18301;
  assign n18303 = n18299 & ~n18302;
  assign n18304 = ~n18274 & n18303;
  assign n18305 = ~n18273 & n18304;
  assign n18306 = ~n18260 & n18305;
  assign n18307 = n18306 ^ n14423;
  assign n18308 = n18307 ^ x711;
  assign n18620 = n18617 ^ n18308;
  assign n18557 = ~n18359 & n18556;
  assign n18559 = n18558 ^ n18557;
  assign n18598 = n18597 ^ n18559;
  assign n18599 = n18330 & ~n18598;
  assign n18600 = n18599 ^ n18597;
  assign n18618 = n18617 ^ n18600;
  assign n18619 = ~n18308 & ~n18618;
  assign n18621 = n18620 ^ n18619;
  assign n18622 = n18621 ^ n15379;
  assign n18623 = n18622 ^ x764;
  assign n18624 = ~n18134 & n18623;
  assign n19113 = n18624 ^ n18623;
  assign n19114 = n19113 ^ n18134;
  assign n19118 = n19114 ^ n18623;
  assign n19119 = n19106 & ~n19118;
  assign n19120 = n19119 ^ n19106;
  assign n19116 = n19106 & n19113;
  assign n19115 = n19106 & n19114;
  assign n19117 = n19116 ^ n19115;
  assign n19121 = n19120 ^ n19117;
  assign n19148 = n19121 ^ n19118;
  assign n19107 = n19106 ^ n19104;
  assign n19131 = n19107 & n19113;
  assign n19138 = n19131 ^ n19115;
  assign n19136 = n19107 & n19114;
  assign n19133 = n19116 ^ n19113;
  assign n19108 = n19107 ^ n18857;
  assign n19111 = n18134 & ~n19108;
  assign n19130 = n18623 & n19111;
  assign n19132 = n19131 ^ n19130;
  assign n19134 = n19133 ^ n19132;
  assign n19137 = n19136 ^ n19134;
  assign n19139 = n19138 ^ n19137;
  assign n19109 = n18624 & ~n19108;
  assign n19110 = n19109 ^ n19108;
  assign n19112 = n19111 ^ n19110;
  assign n19140 = n19139 ^ n19112;
  assign n19141 = n19140 ^ n19119;
  assign n19142 = n19141 ^ n18857;
  assign n19129 = n19115 ^ n19111;
  assign n19135 = n19134 ^ n19129;
  assign n19143 = n19142 ^ n19135;
  assign n19144 = n19143 ^ n18134;
  assign n19125 = n19112 ^ n19109;
  assign n19126 = n19125 ^ n18624;
  assign n19123 = n18624 & n19107;
  assign n19122 = n19121 ^ n19112;
  assign n19124 = n19123 ^ n19122;
  assign n19127 = n19126 ^ n19124;
  assign n19128 = n19127 ^ n19122;
  assign n19145 = n19144 ^ n19128;
  assign n19146 = n19145 ^ n19122;
  assign n19147 = n19146 ^ n19119;
  assign n19149 = n19148 ^ n19147;
  assign n19150 = n19149 ^ n19112;
  assign n19299 = n17620 ^ n17609;
  assign n19300 = n17638 ^ n17472;
  assign n19301 = ~n19299 & ~n19300;
  assign n19302 = ~n17472 & ~n17657;
  assign n19303 = n19302 ^ n17654;
  assign n19304 = n17653 & ~n19303;
  assign n19305 = n19304 ^ n17654;
  assign n19306 = ~n19301 & n19305;
  assign n19308 = n17599 ^ n17567;
  assign n19309 = ~n17517 & n19308;
  assign n19307 = n17665 ^ n17607;
  assign n19310 = n19309 ^ n19307;
  assign n19311 = ~n17472 & n19310;
  assign n19312 = n19311 ^ n19307;
  assign n19313 = ~n17498 & n19312;
  assign n19314 = n19306 & ~n19313;
  assign n19315 = ~n17640 & n19314;
  assign n19316 = n18336 & n19315;
  assign n19320 = ~n17498 & n17643;
  assign n19317 = n18337 ^ n17608;
  assign n19318 = n17498 & n19317;
  assign n19319 = n19318 ^ n18337;
  assign n19321 = n19320 ^ n19319;
  assign n19322 = ~n17653 & n19321;
  assign n19323 = n19322 ^ n19319;
  assign n19324 = n19316 & ~n19323;
  assign n19325 = n19324 ^ n16192;
  assign n19326 = n19325 ^ x730;
  assign n19327 = n17431 ^ x735;
  assign n19151 = n16728 & ~n16759;
  assign n19328 = n16759 ^ n15380;
  assign n19329 = n19328 ^ n15824;
  assign n19330 = n16738 & n19329;
  assign n19158 = n16792 ^ n16768;
  assign n19331 = n19158 ^ n16748;
  assign n19332 = n19331 ^ n16730;
  assign n19333 = n19328 & n19332;
  assign n19334 = ~n16759 & ~n16790;
  assign n19152 = n16786 ^ n16715;
  assign n19153 = ~n16759 & n19152;
  assign n19335 = n16762 ^ n15380;
  assign n19336 = n16751 ^ n16716;
  assign n19337 = ~n15824 & n19336;
  assign n19338 = n19337 ^ n16746;
  assign n19339 = n19338 ^ n16762;
  assign n19340 = ~n19335 & n19339;
  assign n19341 = n19340 ^ n19337;
  assign n19342 = n19341 ^ n16746;
  assign n19343 = n19342 ^ n15380;
  assign n19344 = ~n16762 & ~n19343;
  assign n19345 = n19344 ^ n16762;
  assign n19346 = n19345 ^ n15380;
  assign n19347 = n16731 ^ n16720;
  assign n19348 = n19347 ^ n16724;
  assign n19349 = ~n15380 & n19348;
  assign n19350 = n19349 ^ n19347;
  assign n19351 = n16772 & n19350;
  assign n19352 = n19346 & ~n19351;
  assign n19353 = ~n19153 & n19352;
  assign n19354 = ~n19334 & n19353;
  assign n19355 = ~n16756 & n19354;
  assign n19356 = ~n19333 & n19355;
  assign n19357 = ~n19330 & n19356;
  assign n19359 = ~n16759 & n16762;
  assign n19358 = n16718 & ~n16772;
  assign n19360 = n19359 ^ n19358;
  assign n19361 = n19357 & ~n19360;
  assign n19362 = ~n19151 & n19361;
  assign n19363 = n19362 ^ n16092;
  assign n19364 = n19363 ^ x731;
  assign n19367 = n18251 ^ n18248;
  assign n19366 = n18235 ^ n18218;
  assign n19368 = n19367 ^ n19366;
  assign n19365 = n18747 ^ n18224;
  assign n19369 = n19368 ^ n19365;
  assign n19370 = n18253 & ~n19369;
  assign n19371 = n19370 ^ n19365;
  assign n19372 = ~n18252 & ~n19371;
  assign n19375 = n18247 ^ n18244;
  assign n19374 = n18268 ^ n18263;
  assign n19376 = n19375 ^ n19374;
  assign n19377 = n18252 & n19376;
  assign n19378 = n19377 ^ n19374;
  assign n19373 = ~n18236 & n18252;
  assign n19379 = n19378 ^ n19373;
  assign n19380 = n18253 & ~n19379;
  assign n19381 = n19380 ^ n19378;
  assign n19382 = ~n19372 & n19381;
  assign n19383 = ~n18274 & n19382;
  assign n19384 = ~n18952 & n19383;
  assign n19385 = ~n18744 & n19384;
  assign n19386 = ~n18258 & n19385;
  assign n19387 = n19386 ^ n16337;
  assign n19388 = n19387 ^ x733;
  assign n19389 = ~n19364 & ~n19388;
  assign n19390 = n19389 ^ n19364;
  assign n19391 = n17887 ^ x734;
  assign n19392 = n18701 ^ n18405;
  assign n19393 = n18470 ^ n18460;
  assign n19394 = n19393 ^ n18502;
  assign n19395 = n18701 & ~n19394;
  assign n19396 = n19395 ^ n18502;
  assign n19397 = ~n19392 & n19396;
  assign n19398 = n19397 ^ n18405;
  assign n19400 = n18716 ^ n18467;
  assign n19399 = n18478 ^ n18456;
  assign n19401 = n19400 ^ n19399;
  assign n19402 = n18402 & n19401;
  assign n19403 = n19402 ^ n19399;
  assign n19404 = ~n18453 & ~n19403;
  assign n19405 = ~n19398 & ~n19404;
  assign n19406 = ~n18713 & n19405;
  assign n19407 = ~n18894 & n19406;
  assign n19408 = ~n18890 & n19407;
  assign n19409 = ~n18452 & n19408;
  assign n19410 = ~n18475 & n19409;
  assign n19411 = n19410 ^ n16395;
  assign n19412 = n19411 ^ x732;
  assign n19413 = n19391 & ~n19412;
  assign n19415 = n19413 ^ n19391;
  assign n19435 = ~n19390 & n19415;
  assign n19436 = n19435 ^ n19390;
  assign n19418 = n19390 ^ n19388;
  assign n19420 = n19418 ^ n19364;
  assign n19416 = n19415 ^ n19412;
  assign n19432 = n19420 ^ n19416;
  assign n19425 = n19416 & ~n19420;
  assign n19422 = n19413 & ~n19420;
  assign n19426 = n19425 ^ n19422;
  assign n19421 = ~n19412 & ~n19420;
  assign n19423 = n19422 ^ n19421;
  assign n19424 = n19423 ^ n19420;
  assign n19427 = n19426 ^ n19424;
  assign n19419 = n19416 & ~n19418;
  assign n19428 = n19427 ^ n19419;
  assign n19429 = n19428 ^ n19423;
  assign n19417 = n19389 & n19416;
  assign n19430 = n19429 ^ n19417;
  assign n19431 = n19430 ^ n19422;
  assign n19433 = n19432 ^ n19431;
  assign n19414 = ~n19390 & n19413;
  assign n19434 = n19433 ^ n19414;
  assign n19437 = n19436 ^ n19434;
  assign n19438 = n19437 ^ n19435;
  assign n19439 = n19438 ^ n19423;
  assign n19440 = n19327 & ~n19439;
  assign n19441 = n19440 ^ n19423;
  assign n19442 = n19326 & n19441;
  assign n19443 = n19412 & ~n19418;
  assign n19444 = n19443 ^ n19419;
  assign n19445 = n19444 ^ n19433;
  assign n19446 = n19327 & n19445;
  assign n19447 = n19446 ^ n19444;
  assign n19448 = ~n19326 & n19447;
  assign n19456 = n19413 & ~n19418;
  assign n19457 = n19456 ^ n19418;
  assign n19458 = n19457 ^ n19443;
  assign n19451 = n19389 & n19415;
  assign n19452 = n19451 ^ n19417;
  assign n19449 = n19416 ^ n19391;
  assign n19450 = n19389 & ~n19449;
  assign n19453 = n19452 ^ n19450;
  assign n19454 = n19453 ^ n19389;
  assign n19455 = n19454 ^ n19451;
  assign n19459 = n19458 ^ n19455;
  assign n19460 = n19326 & ~n19327;
  assign n19461 = n19460 ^ n19326;
  assign n19462 = n19461 ^ n19327;
  assign n19463 = ~n19459 & n19462;
  assign n19464 = n19456 ^ n19433;
  assign n19465 = n19464 ^ n19417;
  assign n19466 = n19461 & n19465;
  assign n19467 = n19450 ^ n19327;
  assign n19470 = n19458 ^ n19426;
  assign n19468 = n19458 ^ n19456;
  assign n19469 = n19468 ^ n19427;
  assign n19471 = n19470 ^ n19469;
  assign n19472 = ~n19326 & ~n19471;
  assign n19473 = n19472 ^ n19469;
  assign n19474 = n19473 ^ n19450;
  assign n19475 = n19467 & n19474;
  assign n19476 = n19475 ^ n19472;
  assign n19477 = n19476 ^ n19469;
  assign n19478 = n19477 ^ n19327;
  assign n19479 = ~n19450 & n19478;
  assign n19480 = n19479 ^ n19450;
  assign n19481 = n19480 ^ n19327;
  assign n19482 = ~n19466 & ~n19481;
  assign n19483 = ~n19463 & n19482;
  assign n19487 = n19450 ^ n19444;
  assign n19488 = n19326 & n19487;
  assign n19489 = n19488 ^ n19444;
  assign n19484 = n19454 ^ n19435;
  assign n19485 = ~n19326 & n19484;
  assign n19486 = n19485 ^ n19435;
  assign n19490 = n19489 ^ n19486;
  assign n19491 = n19327 & n19490;
  assign n19492 = n19491 ^ n19486;
  assign n19493 = n19483 & ~n19492;
  assign n19494 = ~n19448 & n19493;
  assign n19498 = n19429 ^ n19426;
  assign n19499 = ~n19326 & ~n19498;
  assign n19500 = n19499 ^ n19426;
  assign n19495 = n19452 ^ n19434;
  assign n19496 = n19326 & n19495;
  assign n19497 = n19496 ^ n19434;
  assign n19501 = n19500 ^ n19497;
  assign n19502 = n19327 & n19501;
  assign n19503 = n19502 ^ n19497;
  assign n19504 = n19494 & ~n19503;
  assign n19505 = ~n19442 & n19504;
  assign n19506 = n19505 ^ n16515;
  assign n19507 = n19506 ^ x765;
  assign n19182 = n18764 ^ x701;
  assign n19154 = ~n15824 & ~n16749;
  assign n19155 = n19154 ^ n16748;
  assign n19156 = n16772 & n19155;
  assign n19157 = n19156 ^ n16748;
  assign n19168 = n16735 & ~n16759;
  assign n19159 = n16790 ^ n16734;
  assign n19160 = n19159 ^ n19158;
  assign n19161 = n19160 ^ n16764;
  assign n19162 = ~n15380 & ~n19161;
  assign n19163 = n19162 ^ n16764;
  assign n19164 = n19163 ^ n16721;
  assign n19165 = ~n19163 & ~n19164;
  assign n19166 = n15824 & n19165;
  assign n19167 = n19166 ^ n15824;
  assign n19169 = n19168 ^ n19167;
  assign n19170 = ~n19157 & ~n19169;
  assign n19171 = ~n19153 & n19170;
  assign n19172 = n15380 & n16767;
  assign n19173 = n19172 ^ n16768;
  assign n19174 = ~n15824 & n19173;
  assign n19175 = n19171 & ~n19174;
  assign n19176 = ~n19151 & n19175;
  assign n19177 = ~n16756 & n19176;
  assign n19178 = n19177 ^ n15864;
  assign n19179 = n19178 ^ x703;
  assign n19183 = ~n17268 & ~n17413;
  assign n19184 = n19183 ^ n17404;
  assign n19185 = ~n17267 & n19184;
  assign n19186 = n19185 ^ n17404;
  assign n19187 = ~n17267 & n17409;
  assign n19188 = n19187 ^ n17267;
  assign n19189 = n19188 ^ n17429;
  assign n19190 = n17268 & ~n19189;
  assign n19191 = n19190 ^ n17268;
  assign n19192 = ~n19186 & ~n19191;
  assign n19193 = n19192 ^ n15914;
  assign n19194 = n19193 ^ x702;
  assign n19180 = n18329 ^ x704;
  assign n19200 = n19194 ^ n19180;
  assign n19199 = n19180 & ~n19194;
  assign n19201 = n19200 ^ n19199;
  assign n19202 = n19179 & n19201;
  assign n19208 = n19182 & n19202;
  assign n19209 = n19208 ^ n19202;
  assign n19206 = ~n19180 & ~n19182;
  assign n19207 = n19194 & n19206;
  assign n19210 = n19209 ^ n19207;
  assign n19203 = n19202 ^ n19194;
  assign n19198 = ~n19179 & n19194;
  assign n19204 = n19203 ^ n19198;
  assign n19181 = n19179 & n19180;
  assign n19195 = n19182 & ~n19194;
  assign n19196 = n19181 & n19195;
  assign n19197 = n19196 ^ n19181;
  assign n19205 = n19204 ^ n19197;
  assign n19211 = n19210 ^ n19205;
  assign n19212 = n18358 ^ x705;
  assign n19213 = n18692 ^ x700;
  assign n19214 = n19212 & ~n19213;
  assign n19215 = n19214 ^ n19212;
  assign n19216 = n19215 ^ n19213;
  assign n19217 = n19216 ^ n19212;
  assign n19218 = n19211 & ~n19217;
  assign n19223 = n19207 ^ n19206;
  assign n19224 = ~n19179 & n19223;
  assign n19225 = n19224 ^ n19223;
  assign n19219 = n19202 ^ n19201;
  assign n19220 = n19219 ^ n19198;
  assign n19221 = n19182 & n19220;
  assign n19222 = n19221 ^ n19220;
  assign n19226 = n19225 ^ n19222;
  assign n19227 = n19226 ^ n19224;
  assign n19228 = n19216 & n19227;
  assign n19236 = n19200 ^ n19182;
  assign n19237 = n19182 ^ n19180;
  assign n19238 = n19179 & n19237;
  assign n19239 = n19238 ^ n19180;
  assign n19240 = n19236 & n19239;
  assign n19235 = n19211 ^ n19209;
  assign n19241 = n19240 ^ n19235;
  assign n19242 = n19241 ^ n19236;
  assign n19233 = n19201 ^ n19180;
  assign n19234 = n19233 ^ n19223;
  assign n19243 = n19242 ^ n19234;
  assign n19229 = n19181 ^ n19180;
  assign n19230 = n19229 ^ n19220;
  assign n19231 = ~n19182 & n19230;
  assign n19232 = n19231 ^ n19230;
  assign n19244 = n19243 ^ n19232;
  assign n19245 = ~n19217 & ~n19244;
  assign n19246 = n19196 & n19216;
  assign n19247 = n19240 ^ n19222;
  assign n19248 = n19247 ^ n19229;
  assign n19249 = n19248 ^ n19244;
  assign n19250 = n19249 ^ n19204;
  assign n19251 = n19250 ^ n19221;
  assign n19252 = ~n19212 & ~n19251;
  assign n19253 = n19252 ^ n19250;
  assign n19254 = n19213 & ~n19253;
  assign n19262 = n19242 ^ n19221;
  assign n19256 = n19219 ^ n19210;
  assign n19257 = n19256 ^ n19249;
  assign n19261 = n19257 ^ n19232;
  assign n19263 = n19262 ^ n19261;
  assign n19264 = ~n19212 & ~n19263;
  assign n19265 = n19264 ^ n19261;
  assign n19255 = n19224 ^ n19205;
  assign n19258 = n19257 ^ n19255;
  assign n19259 = n19212 & ~n19258;
  assign n19260 = n19259 ^ n19257;
  assign n19266 = n19265 ^ n19260;
  assign n19267 = n19213 & n19266;
  assign n19268 = n19267 ^ n19265;
  assign n19269 = ~n19254 & n19268;
  assign n19270 = ~n19246 & n19269;
  assign n19271 = ~n19245 & n19270;
  assign n19273 = n19196 & n19214;
  assign n19272 = n19209 & n19215;
  assign n19274 = n19273 ^ n19272;
  assign n19275 = n19271 & ~n19274;
  assign n19276 = ~n19228 & n19275;
  assign n19277 = ~n19218 & n19276;
  assign n19280 = n19210 ^ n19208;
  assign n19281 = n19280 ^ n19225;
  assign n19278 = n19262 ^ n19243;
  assign n19279 = n19278 ^ n19256;
  assign n19282 = n19281 ^ n19279;
  assign n19283 = ~n19213 & ~n19282;
  assign n19284 = n19283 ^ n19279;
  assign n19285 = n19212 & ~n19284;
  assign n19286 = n19277 & ~n19285;
  assign n19287 = n19250 ^ n19231;
  assign n19288 = ~n19212 & ~n19287;
  assign n19289 = n19288 ^ n19231;
  assign n19290 = ~n19213 & n19289;
  assign n19291 = n19286 & ~n19290;
  assign n19292 = n19231 ^ n19209;
  assign n19293 = ~n19213 & n19292;
  assign n19294 = n19293 ^ n19231;
  assign n19295 = ~n19212 & n19294;
  assign n19296 = n19291 & ~n19295;
  assign n19297 = n19296 ^ n17158;
  assign n19298 = n19297 ^ x760;
  assign n19509 = n19507 ^ n19298;
  assign n19508 = n19298 & ~n19507;
  assign n19510 = n19509 ^ n19508;
  assign n19511 = n19510 ^ n19507;
  assign n19512 = ~n19150 & n19511;
  assign n19516 = n19149 ^ n19127;
  assign n19517 = n19516 ^ n19119;
  assign n19518 = n19517 ^ n19131;
  assign n19519 = n19518 ^ n19143;
  assign n19520 = ~n19507 & n19519;
  assign n19521 = n19520 ^ n19143;
  assign n19513 = n19147 ^ n19135;
  assign n19514 = ~n19507 & ~n19513;
  assign n19515 = n19514 ^ n19135;
  assign n19522 = n19521 ^ n19515;
  assign n19523 = ~n19509 & n19522;
  assign n19524 = n19523 ^ n19521;
  assign n19525 = ~n19512 & ~n19524;
  assign n19527 = n19136 & ~n19298;
  assign n19526 = n19145 & n19510;
  assign n19528 = n19527 ^ n19526;
  assign n19529 = n19525 & ~n19528;
  assign n19531 = n19105 & n19114;
  assign n19532 = ~n19507 & n19531;
  assign n19530 = n19116 & n19509;
  assign n19533 = n19532 ^ n19530;
  assign n19534 = n19529 & ~n19533;
  assign n19535 = n19130 ^ n19111;
  assign n19536 = n19509 & n19535;
  assign n19537 = n19534 & ~n19536;
  assign n19541 = n19131 & ~n19507;
  assign n19538 = n19134 ^ n19123;
  assign n19539 = ~n19507 & n19538;
  assign n19540 = n19539 ^ n19123;
  assign n19542 = n19541 ^ n19540;
  assign n19543 = ~n19298 & n19542;
  assign n19544 = n19543 ^ n19540;
  assign n19545 = n19537 & ~n19544;
  assign n19546 = n19130 ^ n19127;
  assign n19547 = ~n19507 & n19546;
  assign n19548 = n19547 ^ n19127;
  assign n19549 = ~n19509 & n19548;
  assign n19550 = n19545 & ~n19549;
  assign n19551 = n19550 ^ n18692;
  assign n19552 = n18330 ^ n18308;
  assign n19557 = ~n18330 & n18593;
  assign n19558 = n19557 ^ n18330;
  assign n19555 = n18610 ^ n18580;
  assign n19556 = ~n18589 & ~n19555;
  assign n19559 = n19558 ^ n19556;
  assign n19553 = n18308 & ~n18586;
  assign n19554 = n19553 ^ n18576;
  assign n19560 = n19559 ^ n19554;
  assign n19561 = n19552 & n19560;
  assign n19562 = n19561 ^ n19554;
  assign n19563 = n19562 ^ n18436;
  assign n19564 = n19563 ^ x750;
  assign n19565 = n17702 & n18064;
  assign n19566 = n19565 ^ n17701;
  assign n19567 = n18109 & n19566;
  assign n19568 = ~n18074 & ~n19567;
  assign n19581 = n18087 ^ n17710;
  assign n19580 = n18083 ^ n18078;
  assign n19582 = n19581 ^ n19580;
  assign n19583 = ~n17888 & n19582;
  assign n19584 = n19583 ^ n19580;
  assign n19574 = n18090 ^ n16800;
  assign n19571 = n18087 ^ n17703;
  assign n19572 = n19571 ^ n17700;
  assign n19573 = n19572 ^ n17705;
  assign n19575 = n19574 ^ n19573;
  assign n19570 = n17693 ^ n17432;
  assign n19576 = n19575 ^ n19570;
  assign n19569 = n18124 ^ n18092;
  assign n19577 = n19576 ^ n19569;
  assign n19578 = n17888 & ~n19577;
  assign n19579 = n19578 ^ n19569;
  assign n19585 = n19584 ^ n19579;
  assign n19586 = n19585 ^ n19579;
  assign n19587 = ~n18086 & ~n19586;
  assign n19588 = n19587 ^ n19579;
  assign n19589 = ~n18064 & n19588;
  assign n19590 = n19589 ^ n19579;
  assign n19591 = ~n18113 & n19590;
  assign n19592 = n17706 & n18064;
  assign n19593 = n19592 ^ n17703;
  assign n19594 = ~n17888 & n19593;
  assign n19595 = n19591 & ~n19594;
  assign n19596 = ~n18066 & n18121;
  assign n19597 = n19596 ^ n18118;
  assign n19598 = n19595 & ~n19597;
  assign n19599 = n19568 & n19598;
  assign n19600 = ~n18069 & n19599;
  assign n19601 = ~n17708 & n19600;
  assign n19602 = n19601 ^ n17497;
  assign n19603 = n19602 ^ x749;
  assign n19604 = ~n19564 & n19603;
  assign n19605 = n19604 ^ n19564;
  assign n19606 = n19605 ^ n19603;
  assign n19607 = n19606 ^ n19564;
  assign n19642 = n19036 ^ x725;
  assign n19643 = n19325 ^ x728;
  assign n19644 = ~n19642 & n19643;
  assign n19647 = n19644 ^ n19642;
  assign n19608 = n19013 ^ n19003;
  assign n19609 = ~n17267 & n19608;
  assign n19610 = n19609 ^ n19013;
  assign n19611 = n19610 ^ n16137;
  assign n19612 = n19611 ^ x726;
  assign n19613 = n18023 ^ n17993;
  assign n19614 = n19613 ^ n17994;
  assign n19615 = n17999 & ~n19614;
  assign n19616 = n18047 ^ n18004;
  assign n19617 = ~n18045 & n19616;
  assign n19620 = ~n17905 & n17991;
  assign n19618 = n17990 & n18001;
  assign n19619 = n19618 ^ n18015;
  assign n19621 = n19620 ^ n19619;
  assign n19622 = ~n17889 & n19621;
  assign n19623 = n19622 ^ n19619;
  assign n19625 = n18026 ^ n18022;
  assign n19624 = n18019 ^ n18005;
  assign n19626 = n19625 ^ n19624;
  assign n19627 = n19626 ^ n19624;
  assign n19628 = ~n17905 & n19627;
  assign n19629 = n19628 ^ n19624;
  assign n19630 = n17906 & n19629;
  assign n19631 = n19630 ^ n19624;
  assign n19632 = ~n19623 & ~n19631;
  assign n19633 = ~n19617 & n19632;
  assign n19634 = ~n19615 & n19633;
  assign n19635 = ~n18060 & n19634;
  assign n19636 = ~n18883 & n19635;
  assign n19637 = ~n17998 & n19636;
  assign n19638 = n19637 ^ n16218;
  assign n19639 = n19638 ^ x727;
  assign n19640 = n19612 & n19639;
  assign n19665 = n19640 ^ n19612;
  assign n19666 = ~n19647 & n19665;
  assign n19653 = n19612 & ~n19642;
  assign n19667 = n19666 ^ n19653;
  assign n19684 = n19667 ^ n19644;
  assign n19641 = n19640 ^ n19639;
  assign n19669 = n19641 ^ n19612;
  assign n19663 = n19640 & n19644;
  assign n19681 = n19669 ^ n19663;
  assign n19670 = ~n19647 & ~n19669;
  assign n19671 = n19670 ^ n19663;
  assign n19677 = n19671 ^ n19642;
  assign n19648 = n19647 ^ n19643;
  assign n19650 = n19639 & n19648;
  assign n19645 = n19644 ^ n19643;
  assign n19658 = n19650 ^ n19645;
  assign n19678 = n19677 ^ n19658;
  assign n19656 = n19643 ^ n19612;
  assign n19676 = n19656 ^ n19642;
  assign n19679 = n19678 ^ n19676;
  assign n19654 = n19653 ^ n19647;
  assign n19649 = n19641 & n19648;
  assign n19651 = n19650 ^ n19649;
  assign n19646 = n19641 & n19645;
  assign n19652 = n19651 ^ n19646;
  assign n19655 = n19654 ^ n19652;
  assign n19680 = n19679 ^ n19655;
  assign n19682 = n19681 ^ n19680;
  assign n19662 = n19640 & ~n19647;
  assign n19683 = n19682 ^ n19662;
  assign n19685 = n19684 ^ n19683;
  assign n19686 = n19685 ^ n19656;
  assign n19664 = n19663 ^ n19662;
  assign n19668 = n19667 ^ n19664;
  assign n19672 = n19671 ^ n19668;
  assign n19673 = n19672 ^ n19654;
  assign n19674 = n19673 ^ n19668;
  assign n19675 = n19674 ^ n19666;
  assign n19687 = n19686 ^ n19675;
  assign n19661 = n19643 ^ n19639;
  assign n19688 = n19687 ^ n19661;
  assign n19659 = n19639 ^ n19612;
  assign n19660 = n19658 & n19659;
  assign n19689 = n19688 ^ n19660;
  assign n19690 = n19689 ^ n19642;
  assign n19699 = n19690 ^ n19658;
  assign n19696 = n19676 ^ n19639;
  assign n19697 = n19696 ^ n19643;
  assign n19657 = n19656 ^ n19655;
  assign n19691 = n19690 ^ n19657;
  assign n19692 = n19691 ^ n19651;
  assign n19693 = n19692 ^ n19649;
  assign n19694 = n19693 ^ n19654;
  assign n19695 = n19694 ^ n19687;
  assign n19698 = n19697 ^ n19695;
  assign n19700 = n19699 ^ n19698;
  assign n19701 = n18915 ^ x724;
  assign n19702 = n19363 ^ x729;
  assign n19703 = n19701 & n19702;
  assign n19704 = n19703 ^ n19701;
  assign n19705 = n19704 ^ n19702;
  assign n19706 = n19705 ^ n19701;
  assign n19707 = n19700 & n19706;
  assign n19708 = n19689 ^ n19673;
  assign n19709 = ~n19701 & ~n19708;
  assign n19710 = n19709 ^ n19673;
  assign n19711 = n19710 ^ n19689;
  assign n19712 = n19711 ^ n19673;
  assign n19713 = n19702 & n19712;
  assign n19714 = n19702 ^ n19701;
  assign n19720 = n19698 ^ n19692;
  assign n19721 = n19720 ^ n19685;
  assign n19722 = n19721 ^ n19654;
  assign n19717 = n19685 ^ n19649;
  assign n19718 = n19717 ^ n19668;
  assign n19719 = n19718 ^ n19683;
  assign n19723 = n19722 ^ n19719;
  assign n19724 = ~n19702 & ~n19723;
  assign n19725 = n19724 ^ n19719;
  assign n19715 = ~n19695 & ~n19702;
  assign n19716 = n19715 ^ n19694;
  assign n19726 = n19725 ^ n19716;
  assign n19727 = ~n19714 & ~n19726;
  assign n19728 = n19727 ^ n19725;
  assign n19729 = ~n19713 & ~n19728;
  assign n19730 = ~n19707 & n19729;
  assign n19731 = n19730 ^ n17266;
  assign n19732 = n19731 ^ x752;
  assign n19733 = n19083 ^ n19044;
  assign n19734 = n19039 & n19733;
  assign n19735 = n19082 ^ n19043;
  assign n19736 = n19040 & n19735;
  assign n19737 = ~n19734 & ~n19736;
  assign n19738 = n19051 & n19061;
  assign n19741 = n19043 ^ n18986;
  assign n19742 = n19741 ^ n19079;
  assign n19739 = n19049 ^ n18992;
  assign n19740 = n19739 ^ n19056;
  assign n19743 = n19742 ^ n19740;
  assign n19744 = ~n19021 & ~n19743;
  assign n19745 = n19744 ^ n19740;
  assign n19746 = ~n19037 & ~n19745;
  assign n19747 = ~n19738 & ~n19746;
  assign n19748 = n18997 ^ n18991;
  assign n19749 = n19748 ^ n19046;
  assign n19750 = n19749 ^ n19083;
  assign n19751 = n19750 ^ n19083;
  assign n19752 = n19021 & ~n19751;
  assign n19753 = n19752 ^ n19083;
  assign n19754 = n19037 & n19753;
  assign n19755 = n19754 ^ n19083;
  assign n19756 = n19747 & ~n19755;
  assign n19757 = n19063 & n19756;
  assign n19758 = n19737 & n19757;
  assign n19759 = ~n19042 & n19758;
  assign n19760 = n19759 ^ n18427;
  assign n19761 = n19760 ^ x751;
  assign n19762 = n19732 & n19761;
  assign n19763 = n19762 ^ n19732;
  assign n19765 = n19763 ^ n19761;
  assign n19766 = n19765 ^ n19732;
  assign n19767 = n19607 & n19766;
  assign n19764 = n19607 & n19763;
  assign n19768 = n19767 ^ n19764;
  assign n19773 = n18737 & n18738;
  assign n19769 = n18832 ^ n18787;
  assign n19770 = n19769 ^ n18807;
  assign n19771 = n18738 & n19770;
  assign n19772 = n19771 ^ n18807;
  assign n19774 = n19773 ^ n19772;
  assign n19775 = ~n18765 & n19774;
  assign n19776 = n19775 ^ n19772;
  assign n19778 = n18784 & ~n18846;
  assign n19777 = ~n18780 & ~n18805;
  assign n19779 = n19778 ^ n19777;
  assign n19780 = ~n19776 & ~n19779;
  assign n19781 = ~n18844 & n19780;
  assign n19782 = ~n18765 & n18813;
  assign n19783 = n19782 ^ n18796;
  assign n19784 = ~n18738 & n19783;
  assign n19785 = n19781 & ~n19784;
  assign n19786 = n18794 ^ n18776;
  assign n19787 = n18738 & n19786;
  assign n19788 = n19787 ^ n18794;
  assign n19789 = ~n18765 & n19788;
  assign n19790 = n19785 & ~n19789;
  assign n19791 = ~n18839 & n19790;
  assign n19796 = ~n18738 & n18850;
  assign n19792 = n18788 ^ n18775;
  assign n19793 = n19792 ^ n18815;
  assign n19794 = ~n18738 & n19793;
  assign n19795 = n19794 ^ n18815;
  assign n19797 = n19796 ^ n19795;
  assign n19798 = n18765 & n19797;
  assign n19799 = n19798 ^ n19795;
  assign n19800 = n19791 & ~n19799;
  assign n19801 = ~n18854 & n19800;
  assign n19802 = n19801 ^ n17314;
  assign n19803 = n19802 ^ x753;
  assign n19804 = n18509 ^ x712;
  assign n19805 = n19020 ^ x716;
  assign n19806 = n18307 ^ x713;
  assign n19807 = ~n19805 & ~n19806;
  assign n19808 = n19807 ^ n19806;
  assign n19809 = n19808 ^ n19805;
  assign n19810 = n16734 ^ n16718;
  assign n19811 = n19810 ^ n16723;
  assign n19812 = n16758 & n19811;
  assign n19813 = n16790 ^ n16748;
  assign n19814 = n15824 & ~n19813;
  assign n19815 = n16784 & n19328;
  assign n19816 = ~n19814 & ~n19815;
  assign n19817 = n16786 ^ n16729;
  assign n19818 = n19817 ^ n19158;
  assign n19819 = n15824 & n19818;
  assign n19820 = n19819 ^ n19158;
  assign n19821 = n15380 & n19820;
  assign n19822 = n19816 & ~n19821;
  assign n19823 = ~n19812 & n19822;
  assign n19825 = ~n15380 & n16730;
  assign n19824 = n16734 & ~n16759;
  assign n19826 = n19825 ^ n19824;
  assign n19827 = n19823 & ~n19826;
  assign n19828 = ~n19174 & n19827;
  assign n19829 = ~n19334 & n19828;
  assign n19830 = ~n19151 & n19829;
  assign n19831 = n19830 ^ n15605;
  assign n19832 = n19831 ^ x715;
  assign n19834 = n18337 & ~n19300;
  assign n19835 = ~n17638 & ~n17648;
  assign n19840 = n17672 ^ n17647;
  assign n19841 = n19840 ^ n17650;
  assign n19839 = n17619 ^ n17610;
  assign n19842 = n19841 ^ n19839;
  assign n19843 = ~n17472 & ~n19842;
  assign n19844 = n19843 ^ n19839;
  assign n19836 = n17620 ^ n17616;
  assign n19837 = n17472 & ~n19836;
  assign n19838 = n19837 ^ n17620;
  assign n19845 = n19844 ^ n19838;
  assign n19846 = n17498 & n19845;
  assign n19847 = n19846 ^ n19838;
  assign n19848 = ~n19835 & n19847;
  assign n19849 = ~n19834 & n19848;
  assign n19850 = ~n17498 & ~n17645;
  assign n19851 = n19850 ^ n17619;
  assign n19852 = ~n17472 & ~n19851;
  assign n19853 = n19849 & ~n19852;
  assign n19854 = ~n18335 & n19853;
  assign n19855 = ~n17664 & n19854;
  assign n19856 = ~n19323 & n19855;
  assign n19857 = n19856 ^ n15462;
  assign n19858 = n19857 ^ x714;
  assign n19859 = ~n19832 & n19858;
  assign n19860 = n19859 ^ n19858;
  assign n19861 = ~n19809 & n19860;
  assign n19862 = n19861 ^ n19809;
  assign n19833 = ~n19809 & ~n19832;
  assign n19863 = n19862 ^ n19833;
  assign n19864 = ~n19804 & ~n19863;
  assign n19865 = n18887 ^ x717;
  assign n19866 = n19865 ^ n19804;
  assign n19867 = n19859 ^ n19832;
  assign n19882 = n19806 & ~n19867;
  assign n19893 = n19882 ^ n19833;
  assign n19892 = ~n19809 & n19859;
  assign n19894 = n19893 ^ n19892;
  assign n19895 = n19894 ^ n19882;
  assign n19886 = n19807 & n19859;
  assign n19887 = n19886 ^ n19807;
  assign n19883 = n19882 ^ n19867;
  assign n19874 = ~n19808 & n19859;
  assign n19873 = ~n19808 & n19860;
  assign n19875 = n19874 ^ n19873;
  assign n19868 = n19867 ^ n19858;
  assign n19872 = ~n19808 & n19868;
  assign n19876 = n19875 ^ n19872;
  assign n19877 = n19876 ^ n19808;
  assign n19884 = n19883 ^ n19877;
  assign n19881 = n19807 & n19868;
  assign n19885 = n19884 ^ n19881;
  assign n19888 = n19887 ^ n19885;
  assign n19889 = n19888 ^ n19877;
  assign n19890 = n19889 ^ n19860;
  assign n19869 = n19807 ^ n19805;
  assign n19870 = n19868 & ~n19869;
  assign n19871 = n19870 ^ n19861;
  assign n19878 = n19877 ^ n19871;
  assign n19879 = n19878 ^ n19873;
  assign n19880 = n19879 ^ n19870;
  assign n19891 = n19890 ^ n19880;
  assign n19896 = n19895 ^ n19891;
  assign n19897 = n19896 ^ n19873;
  assign n19898 = n19897 ^ n19877;
  assign n19899 = n19866 & ~n19898;
  assign n19900 = n19899 ^ n19877;
  assign n19901 = ~n19864 & n19900;
  assign n19902 = n19804 & n19865;
  assign n19903 = n19902 ^ n19865;
  assign n19904 = n19903 ^ n19804;
  assign n19905 = n19888 & ~n19904;
  assign n19907 = n19859 & ~n19869;
  assign n19906 = n19882 ^ n19861;
  assign n19908 = n19907 ^ n19906;
  assign n19909 = n19908 ^ n19884;
  assign n19910 = n19804 & n19909;
  assign n19911 = n19910 ^ n19884;
  assign n19912 = n19911 ^ n19870;
  assign n19913 = n19865 & n19912;
  assign n19914 = n19913 ^ n19870;
  assign n19915 = ~n19905 & ~n19914;
  assign n19916 = n19901 & n19915;
  assign n19917 = n19881 ^ n19874;
  assign n19918 = ~n19804 & n19917;
  assign n19919 = n19918 ^ n19881;
  assign n19920 = n19865 & n19919;
  assign n19921 = n19916 & ~n19920;
  assign n19927 = n19865 & n19881;
  assign n19922 = n19886 ^ n19872;
  assign n19923 = n19865 & n19922;
  assign n19924 = n19923 ^ n19872;
  assign n19925 = n19924 ^ n19886;
  assign n19926 = n19925 ^ n19872;
  assign n19928 = n19927 ^ n19926;
  assign n19929 = ~n19804 & n19928;
  assign n19930 = n19929 ^ n19926;
  assign n19931 = n19921 & ~n19930;
  assign n19932 = ~n19865 & n19876;
  assign n19933 = n19932 ^ n19872;
  assign n19934 = ~n19804 & n19933;
  assign n19935 = n19931 & ~n19934;
  assign n19936 = n19907 ^ n19893;
  assign n19937 = ~n19804 & n19936;
  assign n19938 = n19937 ^ n19907;
  assign n19939 = ~n19865 & n19938;
  assign n19940 = n19935 & ~n19939;
  assign n19942 = n19902 ^ n19804;
  assign n19943 = n19892 & n19942;
  assign n19941 = n19804 & n19924;
  assign n19944 = n19943 ^ n19941;
  assign n19945 = n19940 & ~n19944;
  assign n19946 = n19945 ^ n17598;
  assign n19947 = n19946 ^ x748;
  assign n19948 = n19803 & ~n19947;
  assign n19949 = n19948 ^ n19947;
  assign n19950 = n19768 & ~n19949;
  assign n19954 = ~n19605 & n19762;
  assign n19955 = n19954 ^ n19605;
  assign n19952 = ~n19605 & n19763;
  assign n19951 = ~n19605 & n19766;
  assign n19953 = n19952 ^ n19951;
  assign n19956 = n19955 ^ n19953;
  assign n19957 = n19956 ^ n19951;
  assign n19958 = ~n19949 & ~n19957;
  assign n19962 = n19606 & n19762;
  assign n19963 = n19962 ^ n19606;
  assign n19960 = n19606 & n19763;
  assign n19959 = n19606 & n19766;
  assign n19961 = n19960 ^ n19959;
  assign n19964 = n19963 ^ n19961;
  assign n19965 = n19947 & n19964;
  assign n19966 = n19947 ^ n19803;
  assign n19977 = n19962 ^ n19954;
  assign n19972 = n19768 ^ n19607;
  assign n19968 = n19604 & n19762;
  assign n19969 = n19968 ^ n19954;
  assign n19970 = n19969 ^ n19762;
  assign n19971 = n19970 ^ n19962;
  assign n19973 = n19972 ^ n19971;
  assign n19978 = n19977 ^ n19973;
  assign n19974 = n19973 ^ n19765;
  assign n19967 = n19964 ^ n19956;
  assign n19975 = n19974 ^ n19967;
  assign n19976 = n19975 ^ n19971;
  assign n19979 = n19978 ^ n19976;
  assign n19980 = n19979 ^ n19976;
  assign n19981 = ~n19947 & n19980;
  assign n19982 = n19981 ^ n19976;
  assign n19983 = ~n19966 & n19982;
  assign n19984 = n19983 ^ n19976;
  assign n19985 = ~n19965 & ~n19984;
  assign n19988 = n19732 ^ n19564;
  assign n19989 = n19988 ^ n19761;
  assign n19990 = n19603 & n19989;
  assign n19987 = n19604 & n19766;
  assign n19991 = n19990 ^ n19987;
  assign n19992 = n19991 ^ n19972;
  assign n19986 = ~n19947 & n19959;
  assign n19993 = n19992 ^ n19986;
  assign n19994 = n19803 & n19993;
  assign n19995 = n19994 ^ n19992;
  assign n19997 = n19992 ^ n19767;
  assign n19998 = n19997 ^ n19975;
  assign n19996 = n19959 ^ n19952;
  assign n19999 = n19998 ^ n19996;
  assign n20000 = n19803 & n19999;
  assign n20001 = n20000 ^ n19996;
  assign n20002 = n19947 & n20001;
  assign n20003 = ~n19995 & ~n20002;
  assign n20004 = n19985 & n20003;
  assign n20005 = n19947 & n19954;
  assign n20006 = n20005 ^ n19968;
  assign n20007 = ~n19966 & n20006;
  assign n20008 = n20007 ^ n19968;
  assign n20009 = n20004 & ~n20008;
  assign n20010 = n19987 ^ n19764;
  assign n20011 = n20010 ^ n19962;
  assign n20012 = ~n19947 & n20011;
  assign n20013 = n20012 ^ n19962;
  assign n20014 = n19803 & n20013;
  assign n20015 = n20009 & ~n20014;
  assign n20016 = ~n19958 & n20015;
  assign n20017 = n19960 ^ n19956;
  assign n20018 = n20017 ^ n19973;
  assign n20019 = ~n19947 & ~n20018;
  assign n20020 = n20019 ^ n19973;
  assign n20021 = n19803 & n20020;
  assign n20022 = n20016 & ~n20021;
  assign n20023 = ~n19950 & n20022;
  assign n20024 = n19960 ^ n19951;
  assign n20025 = ~n19803 & n20024;
  assign n20026 = n20025 ^ n19951;
  assign n20027 = n19947 & n20026;
  assign n20028 = n20023 & ~n20027;
  assign n20029 = n20028 ^ n18509;
  assign n20030 = n20029 ^ x808;
  assign n20031 = n19682 ^ n19666;
  assign n20032 = n19701 & ~n20031;
  assign n20035 = n19720 ^ n19670;
  assign n20036 = n20035 ^ n19717;
  assign n20037 = n20036 ^ n19722;
  assign n20038 = ~n19702 & n20037;
  assign n20039 = n20038 ^ n20036;
  assign n20033 = n19680 & ~n19702;
  assign n20034 = n20033 ^ n19655;
  assign n20040 = n20039 ^ n20034;
  assign n20041 = ~n19714 & n20040;
  assign n20042 = n20041 ^ n20034;
  assign n20043 = ~n20032 & n20042;
  assign n20044 = ~n19707 & n20043;
  assign n20045 = n20044 ^ n17926;
  assign n20046 = n20045 ^ x782;
  assign n20056 = n19572 ^ n18092;
  assign n20057 = n20056 ^ n18083;
  assign n20054 = n18124 ^ n18078;
  assign n20055 = n20054 ^ n17698;
  assign n20058 = n20057 ^ n20055;
  assign n20059 = n18064 & ~n20058;
  assign n20060 = n20059 ^ n20055;
  assign n20048 = n18086 ^ n18080;
  assign n20049 = n20048 ^ n17708;
  assign n20050 = n20049 ^ n18075;
  assign n20047 = n18123 ^ n18086;
  assign n20051 = n20050 ^ n20047;
  assign n20052 = ~n18064 & ~n20051;
  assign n20053 = n20052 ^ n20047;
  assign n20061 = n20060 ^ n20053;
  assign n20062 = ~n18109 & n20061;
  assign n20063 = n20062 ^ n20053;
  assign n20064 = ~n18129 & n20063;
  assign n20065 = ~n18071 & n20064;
  assign n20066 = n18078 ^ n18073;
  assign n20067 = n17888 & n20066;
  assign n20068 = n20067 ^ n18078;
  assign n20069 = n18064 & n20068;
  assign n20070 = n20065 & ~n20069;
  assign n20071 = ~n17888 & n18097;
  assign n20072 = n20071 ^ n18087;
  assign n20073 = ~n18064 & n20072;
  assign n20074 = n20070 & ~n20073;
  assign n20075 = ~n19594 & n20074;
  assign n20076 = n19568 & n20075;
  assign n20077 = ~n18069 & n20076;
  assign n20078 = n20077 ^ n17981;
  assign n20079 = n20078 ^ x781;
  assign n20080 = ~n20046 & ~n20079;
  assign n20081 = n20080 ^ n20079;
  assign n20082 = n20081 ^ n20046;
  assign n20083 = n19250 ^ n19208;
  assign n20084 = n19217 & n20083;
  assign n20085 = n20084 ^ n19216;
  assign n20086 = n19261 ^ n19226;
  assign n20087 = ~n20084 & n20086;
  assign n20088 = n20087 ^ n19261;
  assign n20089 = ~n20085 & n20088;
  assign n20090 = n20089 ^ n19216;
  assign n20091 = n19261 ^ n19243;
  assign n20092 = n19215 & n20091;
  assign n20094 = n19235 ^ n19222;
  assign n20093 = n19232 ^ n19224;
  assign n20095 = n20094 ^ n20093;
  assign n20096 = n20093 ^ n19214;
  assign n20097 = ~n20093 & ~n20096;
  assign n20098 = n20097 ^ n20093;
  assign n20099 = n20095 & ~n20098;
  assign n20100 = n20099 ^ n20097;
  assign n20101 = n20100 ^ n20093;
  assign n20102 = n20101 ^ n19214;
  assign n20103 = ~n20092 & ~n20102;
  assign n20104 = n20103 ^ n20092;
  assign n20105 = ~n20090 & ~n20104;
  assign n20106 = n19213 ^ n19212;
  assign n20107 = ~n19213 & n19247;
  assign n20108 = n20107 ^ n19222;
  assign n20109 = ~n20106 & n20108;
  assign n20110 = n20105 & ~n20109;
  assign n20111 = n19211 ^ n19208;
  assign n20112 = n19213 & n20111;
  assign n20113 = n20112 ^ n19208;
  assign n20114 = n19212 & n20113;
  assign n20115 = n20110 & ~n20114;
  assign n20116 = ~n19246 & n20115;
  assign n20117 = ~n19295 & n20116;
  assign n20118 = ~n19274 & n20117;
  assign n20119 = ~n19210 & n20118;
  assign n20120 = n20119 ^ n17946;
  assign n20121 = n20120 ^ x780;
  assign n20122 = ~n19041 & n19083;
  assign n20123 = n19048 ^ n18990;
  assign n20124 = ~n19037 & n20123;
  assign n20125 = ~n20122 & ~n20124;
  assign n20126 = n18999 ^ n18991;
  assign n20127 = ~n19061 & ~n20126;
  assign n20133 = n18992 ^ n18987;
  assign n20128 = n19056 ^ n18997;
  assign n20129 = n20128 ^ n19050;
  assign n20130 = n20129 ^ n19095;
  assign n20131 = ~n19037 & n20130;
  assign n20132 = n20131 ^ n19095;
  assign n20134 = n20133 ^ n20132;
  assign n20135 = n20134 ^ n20132;
  assign n20136 = n19037 & ~n20135;
  assign n20137 = n20136 ^ n20132;
  assign n20138 = ~n19021 & n20137;
  assign n20139 = n20138 ^ n20132;
  assign n20140 = ~n20127 & ~n20139;
  assign n20141 = n20125 & n20140;
  assign n20142 = ~n19092 & n20141;
  assign n20143 = ~n19065 & n20142;
  assign n20144 = ~n19062 & n20143;
  assign n20145 = n19737 & n20144;
  assign n20146 = ~n19045 & n20145;
  assign n20147 = ~n19042 & n20146;
  assign n20148 = n20147 ^ n17743;
  assign n20149 = n20148 ^ x779;
  assign n20150 = ~n20121 & n20149;
  assign n20152 = n20150 ^ n20149;
  assign n20153 = n20152 ^ n20121;
  assign n20173 = ~n20082 & n20153;
  assign n20157 = ~n20081 & n20149;
  assign n20158 = n20157 ^ n20081;
  assign n20155 = n20150 ^ n20121;
  assign n20156 = ~n20081 & ~n20155;
  assign n20159 = n20158 ^ n20156;
  assign n20154 = n20080 & n20153;
  assign n20160 = n20159 ^ n20154;
  assign n20174 = n20173 ^ n20160;
  assign n20183 = n20174 ^ n20082;
  assign n20178 = n20157 ^ n20149;
  assign n20175 = n20174 ^ n20153;
  assign n20164 = n20080 ^ n20046;
  assign n20170 = ~n20155 & ~n20164;
  assign n20165 = n20152 & ~n20164;
  assign n20171 = n20170 ^ n20165;
  assign n20172 = n20171 ^ n20164;
  assign n20176 = n20175 ^ n20172;
  assign n20167 = ~n20046 & ~n20121;
  assign n20168 = n20167 ^ n20079;
  assign n20169 = n20149 & n20168;
  assign n20177 = n20176 ^ n20169;
  assign n20179 = n20178 ^ n20177;
  assign n20162 = ~n20121 & n20157;
  assign n20163 = n20162 ^ n20157;
  assign n20166 = n20165 ^ n20163;
  assign n20180 = n20179 ^ n20166;
  assign n20181 = n20180 ^ n20152;
  assign n20151 = ~n20082 & n20150;
  assign n20161 = n20160 ^ n20151;
  assign n20182 = n20181 ^ n20161;
  assign n20184 = n20183 ^ n20182;
  assign n20185 = n20184 ^ n20175;
  assign n20190 = n19557 ^ n19556;
  assign n20186 = n18584 ^ n18563;
  assign n20187 = n20186 ^ n18576;
  assign n20188 = n18308 & n20187;
  assign n20189 = n20188 ^ n20186;
  assign n20191 = n20190 ^ n20189;
  assign n20192 = ~n19552 & ~n20191;
  assign n20193 = n20192 ^ n20189;
  assign n20194 = ~n18578 & ~n20193;
  assign n20195 = n20194 ^ n17904;
  assign n20196 = n20195 ^ x783;
  assign n20197 = n18767 & n18786;
  assign n20198 = n18796 ^ n18776;
  assign n20199 = ~n18805 & n20198;
  assign n20200 = ~n20197 & ~n20199;
  assign n20207 = n18832 ^ n18818;
  assign n20202 = n18808 ^ n18785;
  assign n20203 = n20202 ^ n18775;
  assign n20201 = n18787 ^ n18778;
  assign n20204 = n20203 ^ n20201;
  assign n20205 = n18765 & n20204;
  assign n20206 = n20205 ^ n20201;
  assign n20208 = n20207 ^ n20206;
  assign n20209 = n20208 ^ n20206;
  assign n20210 = ~n18765 & n20209;
  assign n20211 = n20210 ^ n20206;
  assign n20212 = ~n18738 & n20211;
  assign n20213 = n20212 ^ n20206;
  assign n20214 = n20200 & ~n20213;
  assign n20215 = n18845 ^ n18794;
  assign n20216 = n18810 ^ n18766;
  assign n20217 = ~n18845 & n20216;
  assign n20218 = n20217 ^ n18810;
  assign n20219 = n20215 & ~n20218;
  assign n20220 = n20219 ^ n18794;
  assign n20221 = n20214 & ~n20220;
  assign n20222 = n18832 ^ n18788;
  assign n20223 = n20222 ^ n18841;
  assign n20224 = n18765 & ~n20223;
  assign n20225 = n20224 ^ n18841;
  assign n20226 = n18805 & ~n20225;
  assign n20227 = n20221 & ~n20226;
  assign n20228 = ~n19799 & n20227;
  assign n20229 = ~n18848 & n20228;
  assign n20230 = n20229 ^ n17815;
  assign n20231 = n20230 ^ x778;
  assign n20232 = n20196 & n20231;
  assign n20233 = n20232 ^ n20231;
  assign n20234 = n20233 ^ n20196;
  assign n20235 = n20185 & ~n20234;
  assign n20236 = n20080 & n20150;
  assign n20237 = n20236 ^ n20166;
  assign n20238 = n20232 ^ n20196;
  assign n20239 = n20237 & n20238;
  assign n20240 = n20179 ^ n20162;
  assign n20241 = n20240 ^ n20176;
  assign n20242 = n20196 & n20241;
  assign n20243 = n20242 ^ n20176;
  assign n20244 = n20231 & n20243;
  assign n20245 = n20181 ^ n20176;
  assign n20246 = n20245 ^ n20159;
  assign n20247 = n20238 & ~n20246;
  assign n20248 = n20185 ^ n20156;
  assign n20249 = n20248 ^ n20170;
  assign n20250 = n20249 ^ n20149;
  assign n20251 = n20250 ^ n20174;
  assign n20258 = n20251 ^ n20156;
  assign n20259 = n20258 ^ n20240;
  assign n20252 = n20173 ^ n20170;
  assign n20253 = ~n20233 & ~n20252;
  assign n20254 = n20175 & n20253;
  assign n20255 = n20174 & ~n20232;
  assign n20256 = ~n20254 & ~n20255;
  assign n20257 = ~n20251 & ~n20256;
  assign n20260 = n20259 ^ n20257;
  assign n20261 = n20260 ^ n20257;
  assign n20262 = ~n20196 & n20261;
  assign n20263 = n20262 ^ n20257;
  assign n20264 = ~n20231 & ~n20263;
  assign n20265 = n20264 ^ n20257;
  assign n20266 = ~n20247 & n20265;
  assign n20267 = n20236 ^ n20163;
  assign n20268 = n20267 ^ n20154;
  assign n20269 = ~n20196 & n20268;
  assign n20270 = n20269 ^ n20154;
  assign n20271 = n20270 ^ n20151;
  assign n20272 = n20270 ^ n20231;
  assign n20273 = ~n20270 & ~n20272;
  assign n20274 = n20273 ^ n20270;
  assign n20275 = n20271 & ~n20274;
  assign n20276 = n20275 ^ n20273;
  assign n20277 = n20276 ^ n20270;
  assign n20278 = n20277 ^ n20231;
  assign n20279 = n20266 & ~n20278;
  assign n20280 = n20279 ^ n20266;
  assign n20281 = ~n20244 & n20280;
  assign n20282 = n20175 ^ n20156;
  assign n20283 = n20282 ^ n20245;
  assign n20284 = n20196 & ~n20283;
  assign n20285 = n20284 ^ n20245;
  assign n20286 = ~n20231 & n20285;
  assign n20287 = n20281 & ~n20286;
  assign n20288 = ~n20239 & n20287;
  assign n20289 = ~n20235 & n20288;
  assign n20290 = n20289 ^ n18887;
  assign n20291 = n20290 ^ x813;
  assign n20292 = n20030 & ~n20291;
  assign n20293 = n20292 ^ n20291;
  assign n20294 = n20293 ^ n20030;
  assign n20332 = ~n19702 & ~n19710;
  assign n20333 = ~n19675 & n19703;
  assign n20334 = n19691 & n19706;
  assign n20335 = n19698 ^ n19652;
  assign n20336 = n20335 ^ n19689;
  assign n20337 = n19641 & n19706;
  assign n20338 = n20337 ^ n19704;
  assign n20339 = n20336 & n20338;
  assign n20342 = n19672 ^ n19662;
  assign n20340 = n19660 ^ n19645;
  assign n20341 = n20340 ^ n19699;
  assign n20343 = n20342 ^ n20341;
  assign n20344 = ~n19702 & n20343;
  assign n20345 = n20344 ^ n20341;
  assign n20346 = ~n19714 & n20345;
  assign n20347 = ~n20339 & ~n20346;
  assign n20348 = ~n20334 & n20347;
  assign n20349 = ~n19707 & n20348;
  assign n20350 = ~n20333 & n20349;
  assign n20351 = n19706 ^ n19685;
  assign n20352 = n19689 ^ n19664;
  assign n20353 = n20352 ^ n19701;
  assign n20354 = n19706 & ~n20353;
  assign n20355 = n20354 ^ n19701;
  assign n20356 = ~n20351 & ~n20355;
  assign n20357 = n20356 ^ n19685;
  assign n20358 = n20350 & n20357;
  assign n20359 = n20340 ^ n19683;
  assign n20360 = ~n19701 & ~n20359;
  assign n20361 = n20360 ^ n19683;
  assign n20362 = ~n19702 & ~n20361;
  assign n20363 = n20358 & ~n20362;
  assign n20364 = ~n20332 & n20363;
  assign n20365 = n20364 ^ n16308;
  assign n20366 = n20365 ^ x768;
  assign n20367 = ~n18068 & n18092;
  assign n20368 = ~n18066 & n19573;
  assign n20369 = n18064 ^ n17708;
  assign n20371 = n20048 ^ n18121;
  assign n20370 = n20047 ^ n17700;
  assign n20372 = n20371 ^ n20370;
  assign n20373 = n17888 & ~n20372;
  assign n20374 = n20373 ^ n20370;
  assign n20375 = n20374 ^ n17708;
  assign n20376 = n20369 & ~n20375;
  assign n20377 = n20376 ^ n20373;
  assign n20378 = n20377 ^ n20370;
  assign n20379 = n20378 ^ n18064;
  assign n20380 = ~n17708 & ~n20379;
  assign n20381 = n20380 ^ n17708;
  assign n20382 = n20381 ^ n18064;
  assign n20383 = ~n20368 & ~n20382;
  assign n20384 = ~n20367 & n20383;
  assign n20385 = n20048 ^ n17703;
  assign n20386 = n20385 ^ n17705;
  assign n20387 = n20386 ^ n17701;
  assign n20388 = n18064 & n20387;
  assign n20389 = n20388 ^ n17701;
  assign n20390 = ~n18109 & n20389;
  assign n20391 = n20384 & ~n20390;
  assign n20392 = ~n20069 & n20391;
  assign n20393 = ~n20073 & n20392;
  assign n20394 = ~n18130 & n20393;
  assign n20395 = ~n19597 & n20394;
  assign n20396 = n20395 ^ n16712;
  assign n20397 = n20396 ^ x769;
  assign n20398 = n20366 & ~n20397;
  assign n20401 = n20398 ^ n20397;
  assign n20419 = n20401 ^ n20366;
  assign n20295 = n19256 ^ n19232;
  assign n20296 = n19215 & n20295;
  assign n20297 = ~n19254 & ~n20296;
  assign n20300 = ~n19216 & ~n19226;
  assign n20301 = ~n19262 & n20300;
  assign n20302 = ~n19209 & n20301;
  assign n20298 = n19250 ^ n19205;
  assign n20299 = n20298 ^ n19225;
  assign n20303 = n20302 ^ n20299;
  assign n20304 = ~n19213 & n20303;
  assign n20305 = n20304 ^ n20299;
  assign n20306 = n20106 & ~n20305;
  assign n20311 = n19257 ^ n19210;
  assign n20312 = n20311 ^ n19224;
  assign n20310 = n19242 ^ n19208;
  assign n20313 = n20312 ^ n20310;
  assign n20314 = ~n19213 & ~n20313;
  assign n20315 = n20314 ^ n20310;
  assign n20316 = n20315 ^ n19231;
  assign n20317 = ~n20315 & ~n20316;
  assign n20318 = ~n19212 & n20317;
  assign n20319 = n20318 ^ n19212;
  assign n20307 = n19224 ^ n19208;
  assign n20308 = n20307 ^ n19225;
  assign n20309 = n19215 & n20308;
  assign n20320 = n20319 ^ n20309;
  assign n20321 = ~n20306 & n20320;
  assign n20322 = ~n19273 & n20321;
  assign n20323 = ~n19290 & n20322;
  assign n20324 = ~n20114 & n20323;
  assign n20325 = n20297 & n20324;
  assign n20326 = ~n19246 & n20325;
  assign n20327 = ~n19245 & n20326;
  assign n20328 = n20327 ^ n16061;
  assign n20329 = n20328 ^ x770;
  assign n20407 = ~n20329 & n20397;
  assign n20408 = ~n20366 & n20407;
  assign n20421 = n20419 ^ n20408;
  assign n20330 = n19506 ^ x767;
  assign n20331 = ~n20329 & ~n20330;
  assign n20413 = n20331 ^ n20330;
  assign n20420 = ~n20413 & n20419;
  assign n20422 = n20421 ^ n20420;
  assign n20414 = n20413 ^ n20329;
  assign n20416 = n20398 & ~n20414;
  assign n20399 = n20398 ^ n20366;
  assign n20415 = n20399 & ~n20414;
  assign n20417 = n20416 ^ n20415;
  assign n20418 = n20417 ^ n20414;
  assign n20423 = n20422 ^ n20418;
  assign n20400 = n20331 & n20399;
  assign n20410 = n20407 ^ n20400;
  assign n20411 = n20410 ^ n20408;
  assign n20405 = n20401 ^ n20331;
  assign n20403 = n20331 & ~n20397;
  assign n20402 = n20401 ^ n20400;
  assign n20404 = n20403 ^ n20402;
  assign n20406 = n20405 ^ n20404;
  assign n20409 = n20408 ^ n20406;
  assign n20412 = n20411 ^ n20409;
  assign n20424 = n20423 ^ n20412;
  assign n20425 = n18622 ^ x766;
  assign n20426 = n19888 & n19903;
  assign n20427 = ~n19804 & n19884;
  assign n20428 = n20427 ^ n19874;
  assign n20429 = ~n19865 & n20428;
  assign n20430 = n20429 ^ n19874;
  assign n20431 = ~n20426 & ~n20430;
  assign n20432 = n19927 ^ n19881;
  assign n20433 = n20432 ^ n19884;
  assign n20434 = ~n19866 & n20433;
  assign n20435 = n20434 ^ n19884;
  assign n20436 = n19889 ^ n19863;
  assign n20437 = n19865 & n20436;
  assign n20438 = n20437 ^ n19863;
  assign n20439 = n19804 & ~n20438;
  assign n20440 = n19907 ^ n19863;
  assign n20441 = ~n19942 & ~n20440;
  assign n20442 = n20441 ^ n19908;
  assign n20443 = ~n19903 & n20442;
  assign n20444 = n20443 ^ n19908;
  assign n20450 = ~n19865 & n19882;
  assign n20445 = n19891 ^ n19871;
  assign n20446 = n20445 ^ n19877;
  assign n20447 = n20446 ^ n19871;
  assign n20448 = ~n19865 & ~n20447;
  assign n20449 = n20448 ^ n19871;
  assign n20451 = n20450 ^ n20449;
  assign n20452 = ~n19804 & n20451;
  assign n20453 = n20452 ^ n20449;
  assign n20454 = ~n20444 & ~n20453;
  assign n20455 = ~n20439 & n20454;
  assign n20456 = ~n20435 & n20455;
  assign n20457 = n20431 & n20456;
  assign n20458 = ~n19934 & n20457;
  assign n20459 = ~n19944 & n20458;
  assign n20460 = n20459 ^ n15823;
  assign n20461 = n20460 ^ x771;
  assign n20462 = ~n20425 & n20461;
  assign n20463 = n20462 ^ n20425;
  assign n20464 = n20463 ^ n20461;
  assign n20465 = n20464 ^ n20425;
  assign n20466 = ~n20424 & n20465;
  assign n20482 = n20397 ^ n20330;
  assign n20488 = n20482 ^ n20408;
  assign n20489 = n20488 ^ n20416;
  assign n20490 = n20489 ^ n20401;
  assign n20467 = n20397 ^ n20366;
  assign n20468 = n20467 ^ n20329;
  assign n20469 = ~n20329 & n20468;
  assign n20483 = n20482 ^ n20469;
  assign n20479 = n20422 ^ n20411;
  assign n20471 = n20331 ^ n20329;
  assign n20472 = ~n20401 & ~n20471;
  assign n20473 = n20472 ^ n20471;
  assign n20474 = n20473 ^ n20412;
  assign n20480 = n20479 ^ n20474;
  assign n20481 = n20480 ^ n20415;
  assign n20484 = n20483 ^ n20481;
  assign n20485 = n20484 ^ n20468;
  assign n20486 = n20329 & ~n20485;
  assign n20478 = n20467 ^ n20330;
  assign n20487 = n20486 ^ n20478;
  assign n20491 = n20490 ^ n20487;
  assign n20492 = n20491 ^ n20406;
  assign n20470 = n20469 ^ n20408;
  assign n20475 = n20474 ^ n20470;
  assign n20476 = n20475 ^ n20403;
  assign n20493 = n20492 ^ n20476;
  assign n20494 = n20493 ^ n20484;
  assign n20498 = n20494 ^ n20413;
  assign n20477 = n20476 ^ n20420;
  assign n20495 = n20494 ^ n20477;
  assign n20496 = n20495 ^ n20406;
  assign n20497 = n20496 ^ n20484;
  assign n20499 = n20498 ^ n20497;
  assign n20500 = n20464 & n20499;
  assign n20501 = n20424 ^ n20422;
  assign n20502 = n20501 ^ n20481;
  assign n20503 = n20461 & n20502;
  assign n20504 = n20503 ^ n20501;
  assign n20505 = n20464 ^ n20462;
  assign n20506 = ~n20504 & n20505;
  assign n20507 = ~n20425 & n20497;
  assign n20508 = n20507 ^ n20496;
  assign n20509 = n20461 & n20508;
  assign n20510 = ~n20506 & ~n20509;
  assign n20511 = ~n20461 & n20489;
  assign n20512 = n20511 ^ n20416;
  assign n20513 = ~n20425 & n20512;
  assign n20514 = n20513 ^ n20416;
  assign n20515 = n20510 & ~n20514;
  assign n20516 = ~n20500 & n20515;
  assign n20517 = ~n20466 & n20516;
  assign n20518 = n20494 ^ n20476;
  assign n20519 = n20518 ^ n20475;
  assign n20520 = n20425 & ~n20519;
  assign n20521 = n20520 ^ n20475;
  assign n20522 = ~n20461 & ~n20521;
  assign n20523 = n20517 & ~n20522;
  assign n20524 = n20523 ^ n19831;
  assign n20525 = n20524 ^ x811;
  assign n20526 = n20195 ^ x737;
  assign n20563 = n18766 & n18789;
  assign n20564 = n18806 ^ n18769;
  assign n20565 = n20564 ^ n20201;
  assign n20566 = n18767 & n20565;
  assign n20567 = n18815 ^ n18775;
  assign n20568 = n20567 ^ n18810;
  assign n20569 = ~n18805 & ~n20568;
  assign n20570 = ~n20566 & ~n20569;
  assign n20571 = ~n20563 & n20570;
  assign n20572 = ~n18765 & n18777;
  assign n20573 = n20572 ^ n18775;
  assign n20574 = ~n18738 & n20573;
  assign n20575 = n20571 & ~n20574;
  assign n20576 = ~n19784 & n20575;
  assign n20577 = ~n19789 & n20576;
  assign n20578 = ~n18830 & n20577;
  assign n20579 = ~n20226 & n20578;
  assign n20580 = ~n18848 & n20579;
  assign n20581 = ~n18854 & n20580;
  assign n20582 = n20581 ^ n18194;
  assign n20583 = n20582 ^ x738;
  assign n20629 = ~n20526 & ~n20583;
  assign n20527 = n18997 ^ n18992;
  assign n20528 = n19038 & ~n20527;
  assign n20534 = n19079 ^ n18999;
  assign n20533 = n19082 ^ n18990;
  assign n20535 = n20534 ^ n20533;
  assign n20536 = ~n19037 & n20535;
  assign n20537 = n20536 ^ n20533;
  assign n20530 = n19040 & n20128;
  assign n20531 = n20530 ^ n20126;
  assign n20529 = n19048 ^ n19043;
  assign n20532 = n20531 ^ n20529;
  assign n20538 = n20537 ^ n20532;
  assign n20539 = ~n19061 & ~n20538;
  assign n20540 = n20539 ^ n20532;
  assign n20541 = ~n19734 & n20540;
  assign n20542 = ~n19045 & n20541;
  assign n20543 = ~n20528 & n20542;
  assign n20544 = ~n19021 & n19083;
  assign n20545 = n20544 ^ n19000;
  assign n20546 = n19037 & n20545;
  assign n20547 = n20546 ^ n19000;
  assign n20548 = n20543 & ~n20547;
  assign n20549 = n19050 ^ n19039;
  assign n20550 = n19041 ^ n18986;
  assign n20551 = ~n19050 & n20550;
  assign n20552 = n20551 ^ n19041;
  assign n20553 = n20549 & ~n20552;
  assign n20554 = n20553 ^ n19039;
  assign n20555 = n20548 & ~n20554;
  assign n20556 = ~n19098 & n20555;
  assign n20557 = n20556 ^ n17471;
  assign n20558 = n20557 ^ x740;
  assign n20559 = n20526 & ~n20558;
  assign n20560 = n20559 ^ n20526;
  assign n20561 = n20560 ^ n20558;
  assign n20562 = n20561 ^ n20526;
  assign n20634 = n20629 ^ n20562;
  assign n20584 = n19873 & ~n19942;
  assign n20585 = n20584 ^ n20440;
  assign n20586 = ~n19903 & ~n20585;
  assign n20587 = n20586 ^ n20440;
  assign n20588 = n19888 ^ n19886;
  assign n20589 = n19804 & n20588;
  assign n20590 = n20589 ^ n19886;
  assign n20591 = ~n19865 & n20590;
  assign n20592 = n20587 & ~n20591;
  assign n20593 = n19903 ^ n19877;
  assign n20594 = n19942 ^ n19833;
  assign n20595 = n19877 & ~n20594;
  assign n20596 = n20595 ^ n19942;
  assign n20597 = ~n20593 & n20596;
  assign n20598 = n20597 ^ n19903;
  assign n20604 = n20445 ^ n19886;
  assign n20605 = n20604 ^ n19894;
  assign n20606 = n20605 ^ n19863;
  assign n20607 = n20606 ^ n19863;
  assign n20608 = n19804 & n20607;
  assign n20600 = n19895 ^ n19878;
  assign n20599 = n19896 ^ n19893;
  assign n20601 = n20600 ^ n20599;
  assign n20602 = ~n19804 & ~n20601;
  assign n20603 = n20602 ^ n20599;
  assign n20609 = n20608 ^ n20603;
  assign n20610 = n20609 ^ n20608;
  assign n20611 = n19863 & ~n20610;
  assign n20612 = n20611 ^ n20608;
  assign n20613 = ~n19865 & ~n20612;
  assign n20614 = n20613 ^ n20608;
  assign n20615 = ~n20598 & ~n20614;
  assign n20616 = n20431 & n20615;
  assign n20617 = ~n19930 & n20616;
  assign n20618 = n20592 & n20617;
  assign n20619 = n20618 ^ n18160;
  assign n20620 = n20619 ^ x739;
  assign n20621 = ~n20583 & n20620;
  assign n20624 = n20621 ^ n20583;
  assign n20628 = ~n20562 & ~n20624;
  assign n20630 = n20629 ^ n20628;
  assign n20626 = ~n20562 & n20621;
  assign n20625 = n20561 & ~n20624;
  assign n20627 = n20626 ^ n20625;
  assign n20631 = n20630 ^ n20627;
  assign n20622 = n20621 ^ n20620;
  assign n20623 = ~n20562 & n20622;
  assign n20632 = n20631 ^ n20623;
  assign n20633 = n20632 ^ n20625;
  assign n20635 = n20634 ^ n20633;
  assign n20636 = n20635 ^ n20625;
  assign n20637 = n20045 ^ x736;
  assign n20638 = n19327 & n19500;
  assign n20639 = n19468 ^ n19425;
  assign n20640 = n19460 & ~n20639;
  assign n20641 = n19437 ^ n19326;
  assign n20643 = n19455 ^ n19450;
  assign n20642 = n19454 ^ n19434;
  assign n20644 = n20643 ^ n20642;
  assign n20645 = ~n19327 & n20644;
  assign n20646 = n20645 ^ n20642;
  assign n20647 = n20646 ^ n19437;
  assign n20648 = n20641 & ~n20647;
  assign n20649 = n20648 ^ n20645;
  assign n20650 = n20649 ^ n20642;
  assign n20651 = n20650 ^ n19326;
  assign n20652 = n19437 & ~n20651;
  assign n20653 = n20652 ^ n19437;
  assign n20654 = n20653 ^ n19326;
  assign n20655 = ~n20640 & ~n20654;
  assign n20661 = n19444 ^ n19434;
  assign n20660 = n19455 ^ n19428;
  assign n20662 = n20661 ^ n20660;
  assign n20656 = n19456 ^ n19452;
  assign n20657 = n20656 ^ n19443;
  assign n20658 = ~n19326 & n20657;
  assign n20659 = n20658 ^ n19443;
  assign n20663 = n20662 ^ n20659;
  assign n20664 = n20663 ^ n20659;
  assign n20665 = ~n19326 & ~n20664;
  assign n20666 = n20665 ^ n20659;
  assign n20667 = ~n19327 & n20666;
  assign n20668 = n20667 ^ n20659;
  assign n20669 = n20655 & ~n20668;
  assign n20670 = n19327 ^ n19326;
  assign n20674 = ~n19327 & n19423;
  assign n20671 = n19444 ^ n19438;
  assign n20672 = ~n19326 & ~n20671;
  assign n20673 = n20672 ^ n19444;
  assign n20675 = n20674 ^ n20673;
  assign n20676 = ~n20670 & n20675;
  assign n20677 = n20676 ^ n20673;
  assign n20678 = n20669 & ~n20677;
  assign n20679 = ~n20638 & n20678;
  assign n20680 = n20679 ^ n17516;
  assign n20681 = n20680 ^ x741;
  assign n20682 = ~n20637 & n20681;
  assign n20683 = n20682 ^ n20637;
  assign n20684 = ~n20636 & ~n20683;
  assign n20685 = n20683 ^ n20681;
  assign n20686 = n20685 ^ n20637;
  assign n20687 = n20622 & n20686;
  assign n20688 = n20560 & n20687;
  assign n20689 = n20559 & n20687;
  assign n20692 = n20559 & n20583;
  assign n20693 = n20692 ^ n20559;
  assign n20694 = n20693 ^ n20627;
  assign n20690 = n20620 ^ n20526;
  assign n20691 = n20690 ^ n20558;
  assign n20695 = n20694 ^ n20691;
  assign n20696 = ~n20683 & n20695;
  assign n20697 = ~n20689 & ~n20696;
  assign n20703 = n20583 ^ n20558;
  assign n20704 = n20703 ^ n20634;
  assign n20723 = n20704 ^ n20560;
  assign n20707 = n20622 ^ n20583;
  assign n20722 = n20559 & n20707;
  assign n20724 = n20723 ^ n20722;
  assign n20698 = n20559 & ~n20624;
  assign n20725 = n20724 ^ n20698;
  assign n20714 = n20561 & n20707;
  assign n20715 = n20714 ^ n20625;
  assign n20726 = n20725 ^ n20715;
  assign n20713 = n20631 ^ n20561;
  assign n20716 = n20715 ^ n20713;
  assign n20717 = n20716 ^ n20626;
  assign n20708 = n20560 & n20707;
  assign n20709 = n20708 ^ n20627;
  assign n20701 = n20620 ^ n20558;
  assign n20702 = n20583 ^ n20526;
  assign n20705 = n20704 ^ n20702;
  assign n20706 = n20701 & n20705;
  assign n20710 = n20709 ^ n20706;
  assign n20699 = n20698 ^ n20693;
  assign n20700 = n20699 ^ n20692;
  assign n20711 = n20710 ^ n20700;
  assign n20712 = n20711 ^ n20708;
  assign n20718 = n20717 ^ n20712;
  assign n20719 = n20718 ^ n20625;
  assign n20720 = ~n20637 & n20719;
  assign n20721 = n20720 ^ n20625;
  assign n20727 = n20726 ^ n20721;
  assign n20728 = n20727 ^ n20721;
  assign n20729 = n20637 & ~n20728;
  assign n20730 = n20729 ^ n20721;
  assign n20731 = ~n20681 & n20730;
  assign n20732 = n20731 ^ n20721;
  assign n20733 = n20697 & ~n20732;
  assign n20734 = ~n20688 & n20733;
  assign n20736 = n20631 & n20685;
  assign n20735 = ~n20635 & n20637;
  assign n20737 = n20736 ^ n20735;
  assign n20738 = n20734 & ~n20737;
  assign n20739 = ~n20684 & n20738;
  assign n20742 = n20682 & n20714;
  assign n20740 = n20716 ^ n20628;
  assign n20741 = n20686 & n20740;
  assign n20743 = n20742 ^ n20741;
  assign n20744 = n20739 & ~n20743;
  assign n20746 = n20704 ^ n20692;
  assign n20747 = n20746 ^ n20710;
  assign n20748 = n20686 & ~n20747;
  assign n20745 = n20686 & n20698;
  assign n20749 = n20748 ^ n20745;
  assign n20750 = n20744 & ~n20749;
  assign n20751 = n20750 ^ n18307;
  assign n20752 = n20751 ^ x809;
  assign n20753 = ~n20525 & ~n20752;
  assign n20986 = n20753 ^ n20525;
  assign n20987 = n20986 ^ n20752;
  assign n20990 = n20987 ^ n20525;
  assign n20754 = n18133 ^ x759;
  assign n20755 = n19731 ^ x754;
  assign n20814 = n19297 ^ x758;
  assign n20791 = n19802 ^ x755;
  assign n20840 = n20814 ^ n20791;
  assign n20793 = n19893 & n19902;
  assign n20794 = n19870 & ~n19942;
  assign n20795 = n20794 ^ n19879;
  assign n20796 = ~n19903 & ~n20795;
  assign n20797 = n20796 ^ n19879;
  assign n20798 = ~n20793 & n20797;
  assign n20800 = n19874 & n19942;
  assign n20799 = ~n19865 & n19896;
  assign n20801 = n20800 ^ n20799;
  assign n20802 = n20798 & ~n20801;
  assign n20803 = ~n20439 & n20802;
  assign n20804 = ~n20435 & n20803;
  assign n20805 = ~n19941 & n20804;
  assign n20806 = ~n19920 & n20805;
  assign n20807 = ~n19939 & n20806;
  assign n20808 = n20592 & n20807;
  assign n20809 = n20808 ^ n17353;
  assign n20810 = n20809 ^ x756;
  assign n20841 = n20840 ^ n20810;
  assign n20761 = n19427 ^ n19421;
  assign n20762 = n20761 ^ n19434;
  assign n20756 = n19484 ^ n19458;
  assign n20757 = n20756 ^ n19433;
  assign n20758 = n20757 ^ n19388;
  assign n20759 = ~n19327 & ~n20758;
  assign n20760 = n20759 ^ n19454;
  assign n20763 = n20762 ^ n20760;
  assign n20764 = n20763 ^ n20760;
  assign n20765 = n19327 & ~n20764;
  assign n20766 = n20765 ^ n20760;
  assign n20767 = ~n19326 & n20766;
  assign n20768 = n20767 ^ n20760;
  assign n20770 = n19435 ^ n19417;
  assign n20771 = n20770 ^ n19327;
  assign n20774 = n20771 ^ n19326;
  assign n20775 = n20771 ^ n19458;
  assign n20776 = n20775 ^ n20761;
  assign n20777 = ~n20774 & ~n20776;
  assign n20773 = ~n19420 & n19461;
  assign n20778 = n20777 ^ n20773;
  assign n20769 = n19428 & n19461;
  assign n20772 = n20771 ^ n20769;
  assign n20779 = n20778 ^ n20772;
  assign n20780 = n20779 ^ n19327;
  assign n20781 = n20780 ^ n19326;
  assign n20782 = n20781 ^ n20771;
  assign n20783 = ~n20768 & n20782;
  assign n20784 = n19497 ^ n19489;
  assign n20785 = ~n19327 & n20784;
  assign n20786 = n20785 ^ n19489;
  assign n20787 = n20783 & ~n20786;
  assign n20788 = ~n19442 & n20787;
  assign n20789 = n20788 ^ n17381;
  assign n20790 = n20789 ^ x757;
  assign n20815 = n20814 ^ n20790;
  assign n20842 = n20810 & ~n20815;
  assign n20843 = n20842 ^ n20814;
  assign n20844 = ~n20841 & ~n20843;
  assign n20839 = n20791 & n20815;
  assign n20845 = n20844 ^ n20839;
  assign n20828 = n20814 ^ n20810;
  assign n20829 = ~n20791 & ~n20828;
  assign n20830 = n20829 ^ n20815;
  assign n20812 = n20790 & ~n20791;
  assign n20826 = n20812 & ~n20814;
  assign n20813 = n20812 ^ n20791;
  assign n20827 = n20826 ^ n20813;
  assign n20831 = n20830 ^ n20827;
  assign n20846 = n20845 ^ n20831;
  assign n20847 = ~n20755 & n20846;
  assign n20818 = ~n20810 & n20814;
  assign n20819 = n20818 ^ n20810;
  assign n20836 = n20828 ^ n20790;
  assign n20837 = n20819 & n20836;
  assign n20821 = ~n20810 & n20812;
  assign n20835 = n20821 ^ n20813;
  assign n20838 = n20837 ^ n20835;
  assign n20848 = n20847 ^ n20838;
  assign n20811 = n20810 ^ n20790;
  assign n20820 = n20819 ^ n20814;
  assign n20822 = n20821 ^ n20820;
  assign n20816 = n20815 ^ n20813;
  assign n20817 = ~n20810 & n20816;
  assign n20823 = n20822 ^ n20817;
  assign n20824 = n20811 & ~n20823;
  assign n20792 = n20791 ^ n20790;
  assign n20825 = n20824 ^ n20792;
  assign n20832 = n20831 ^ n20825;
  assign n20833 = n20755 & n20832;
  assign n20834 = n20833 ^ n20825;
  assign n20849 = n20848 ^ n20834;
  assign n20850 = n20754 & ~n20849;
  assign n20851 = n20850 ^ n20754;
  assign n20852 = n20851 ^ n20834;
  assign n20853 = n20852 ^ n19020;
  assign n20854 = n20853 ^ x812;
  assign n20855 = n20680 ^ x743;
  assign n20881 = n19691 & n19704;
  assign n20883 = n19643 ^ n19642;
  assign n20884 = ~n19639 & ~n20883;
  assign n20885 = n20884 ^ n19643;
  assign n20886 = ~n19696 & n20885;
  assign n20882 = n19699 ^ n19652;
  assign n20887 = n20886 ^ n20882;
  assign n20888 = ~n19705 & n20887;
  assign n20889 = n20031 ^ n19664;
  assign n20890 = n19714 & ~n20889;
  assign n20891 = n19706 & n19720;
  assign n20892 = ~n20890 & ~n20891;
  assign n20893 = n19698 ^ n19649;
  assign n20894 = n19701 & n20893;
  assign n20895 = n20886 ^ n19662;
  assign n20896 = n19703 & n20895;
  assign n20897 = ~n20894 & ~n20896;
  assign n20898 = n20892 & n20897;
  assign n20899 = ~n20888 & n20898;
  assign n20900 = ~n20881 & n20899;
  assign n20901 = ~n19713 & n20900;
  assign n20902 = ~n20332 & n20901;
  assign n20903 = n20902 ^ n17566;
  assign n20904 = n20903 ^ x745;
  assign n20911 = n20855 & n20904;
  assign n20912 = n20911 ^ n20904;
  assign n20856 = n19216 & ~n19243;
  assign n20866 = n19226 ^ n19196;
  assign n20867 = n20866 ^ n19242;
  assign n20868 = n20867 ^ n19241;
  assign n20869 = n19213 & n20868;
  assign n20870 = n20869 ^ n19241;
  assign n20857 = n19222 ^ n19205;
  assign n20858 = n20857 ^ n19211;
  assign n20859 = n20857 ^ n19213;
  assign n20860 = n19212 & n20859;
  assign n20861 = n20860 ^ n19213;
  assign n20862 = n20858 & ~n20861;
  assign n20863 = n20862 ^ n19211;
  assign n20864 = ~n20307 & ~n20863;
  assign n20865 = n19249 & n20864;
  assign n20871 = n20870 ^ n20865;
  assign n20872 = n19212 & ~n20871;
  assign n20873 = n20872 ^ n20865;
  assign n20874 = ~n20856 & n20873;
  assign n20875 = n20297 & n20874;
  assign n20876 = ~n19295 & n20875;
  assign n20877 = ~n19245 & n20876;
  assign n20878 = ~n19274 & n20877;
  assign n20879 = n20878 ^ n17536;
  assign n20880 = n20879 ^ x744;
  assign n20905 = n19946 ^ x746;
  assign n20906 = ~n20904 & n20905;
  assign n20907 = ~n20880 & n20906;
  assign n20908 = n20907 ^ n20906;
  assign n20909 = ~n20855 & n20908;
  assign n20910 = n20909 ^ n20908;
  assign n20913 = n20912 ^ n20910;
  assign n20914 = n19602 ^ x747;
  assign n20915 = n20557 ^ x742;
  assign n20916 = ~n20914 & ~n20915;
  assign n20917 = n20916 ^ n20914;
  assign n20918 = n20913 & ~n20917;
  assign n20926 = n20906 ^ n20905;
  assign n20925 = n20905 & n20912;
  assign n20927 = n20926 ^ n20925;
  assign n20928 = n20880 & n20927;
  assign n20929 = n20928 ^ n20927;
  assign n20921 = n20906 ^ n20904;
  assign n20919 = ~n20880 & ~n20905;
  assign n20920 = ~n20904 & n20919;
  assign n20922 = n20921 ^ n20920;
  assign n20923 = ~n20855 & ~n20922;
  assign n20924 = n20923 ^ n20922;
  assign n20930 = n20929 ^ n20924;
  assign n20931 = n20917 ^ n20915;
  assign n20932 = n20931 ^ n20914;
  assign n20933 = ~n20930 & ~n20932;
  assign n20949 = ~n20855 & n20920;
  assign n20950 = n20949 ^ n20920;
  assign n20945 = n20880 & n20925;
  assign n20946 = n20945 ^ n20925;
  assign n20947 = n20946 ^ n20923;
  assign n20948 = n20947 ^ n20929;
  assign n20951 = n20950 ^ n20948;
  assign n20942 = n20855 & n20907;
  assign n20943 = n20942 ^ n20907;
  assign n20937 = n20920 ^ n20919;
  assign n20934 = n20912 & n20919;
  assign n20938 = n20937 ^ n20934;
  assign n20939 = n20938 ^ n20911;
  assign n20940 = n20939 ^ n20927;
  assign n20935 = n20934 ^ n20912;
  assign n20936 = n20935 ^ n20925;
  assign n20941 = n20940 ^ n20936;
  assign n20944 = n20943 ^ n20941;
  assign n20952 = n20951 ^ n20944;
  assign n20953 = ~n20915 & n20952;
  assign n20954 = n20953 ^ n20944;
  assign n20955 = n20931 ^ n20916;
  assign n20956 = n20954 & ~n20955;
  assign n20959 = n20949 ^ n20909;
  assign n20960 = ~n20917 & n20959;
  assign n20961 = n20960 ^ n20959;
  assign n20957 = n20942 ^ n20924;
  assign n20958 = n20915 & ~n20957;
  assign n20962 = n20961 ^ n20958;
  assign n20963 = ~n20956 & ~n20962;
  assign n20964 = ~n20933 & n20963;
  assign n20965 = ~n20918 & n20964;
  assign n20967 = n20943 ^ n20934;
  assign n20966 = n20938 ^ n20910;
  assign n20968 = n20967 ^ n20966;
  assign n20969 = n20914 & n20968;
  assign n20970 = n20969 ^ n20966;
  assign n20971 = ~n20915 & n20970;
  assign n20972 = n20965 & ~n20971;
  assign n20974 = ~n20917 & n20940;
  assign n20973 = n20928 & ~n20932;
  assign n20975 = n20974 ^ n20973;
  assign n20976 = n20972 & ~n20975;
  assign n20978 = n20929 & ~n20931;
  assign n20977 = ~n20932 & n20940;
  assign n20979 = n20978 ^ n20977;
  assign n20980 = n20976 & ~n20979;
  assign n20981 = n20980 ^ n19857;
  assign n20982 = n20981 ^ x810;
  assign n20983 = n20854 & ~n20982;
  assign n20998 = n20983 ^ n20854;
  assign n21007 = ~n20990 & n20998;
  assign n21008 = n21007 ^ n20990;
  assign n20984 = n20983 ^ n20982;
  assign n21003 = ~n20984 & ~n20986;
  assign n21004 = n21003 ^ n20984;
  assign n20999 = ~n20987 & n20998;
  assign n21000 = n20999 ^ n20987;
  assign n20993 = n20753 & n20983;
  assign n20992 = n20983 & ~n20986;
  assign n20994 = n20993 ^ n20992;
  assign n20995 = n20994 ^ n20983;
  assign n20991 = n20983 & ~n20990;
  assign n20996 = n20995 ^ n20991;
  assign n20988 = n20984 ^ n20854;
  assign n20989 = ~n20987 & n20988;
  assign n20997 = n20996 ^ n20989;
  assign n21001 = n21000 ^ n20997;
  assign n20985 = n20753 & ~n20984;
  assign n21002 = n21001 ^ n20985;
  assign n21005 = n21004 ^ n21002;
  assign n21006 = n21005 ^ n20991;
  assign n21009 = n21008 ^ n21006;
  assign n21010 = n20294 & ~n21009;
  assign n21029 = n20291 & n20997;
  assign n21014 = n20992 ^ n20986;
  assign n21020 = n21014 ^ n20988;
  assign n21012 = ~n20986 & n20998;
  assign n21013 = n21012 ^ n21003;
  assign n21018 = n21013 ^ n20989;
  assign n21019 = n21018 ^ n21009;
  assign n21021 = n21020 ^ n21019;
  assign n21022 = n21021 ^ n20991;
  assign n21023 = n21022 ^ n21007;
  assign n21024 = n21023 ^ n20992;
  assign n21025 = n21024 ^ n21001;
  assign n21015 = n21014 ^ n21013;
  assign n21011 = n21007 ^ n21005;
  assign n21016 = n21015 ^ n21011;
  assign n21017 = n21016 ^ n20996;
  assign n21026 = n21025 ^ n21017;
  assign n21027 = ~n20291 & n21026;
  assign n21028 = n21027 ^ n21017;
  assign n21030 = n21029 ^ n21028;
  assign n21031 = ~n20030 & ~n21030;
  assign n21032 = n21031 ^ n21028;
  assign n21034 = n20291 ^ n20030;
  assign n21035 = n20753 & n20998;
  assign n21036 = ~n21034 & n21035;
  assign n21033 = ~n20293 & ~n21009;
  assign n21037 = n21036 ^ n21033;
  assign n21038 = n21032 & ~n21037;
  assign n21039 = n20030 & n20994;
  assign n21040 = n21039 ^ n20993;
  assign n21041 = n20291 & n21040;
  assign n21042 = n21038 & ~n21041;
  assign n21043 = n21012 ^ n20985;
  assign n21044 = ~n20030 & n21043;
  assign n21045 = n21044 ^ n20985;
  assign n21046 = n20291 & n21045;
  assign n21047 = n21042 & ~n21046;
  assign n21048 = n20999 ^ n20985;
  assign n21049 = n20291 & n21048;
  assign n21050 = n21049 ^ n20999;
  assign n21051 = n21034 & n21050;
  assign n21052 = n21047 & ~n21051;
  assign n21053 = n20997 ^ n20991;
  assign n21054 = ~n20291 & n21053;
  assign n21055 = n21054 ^ n20991;
  assign n21056 = ~n20030 & n21055;
  assign n21057 = n21052 & ~n21056;
  assign n21062 = n20993 & ~n21034;
  assign n21060 = ~n20293 & n21003;
  assign n21058 = n21015 ^ n20999;
  assign n21059 = ~n20293 & ~n21058;
  assign n21061 = n21060 ^ n21059;
  assign n21063 = n21062 ^ n21061;
  assign n21064 = n21057 & ~n21063;
  assign n21065 = ~n21010 & n21064;
  assign n21066 = n21035 ^ n21003;
  assign n21067 = n21066 ^ n21001;
  assign n21068 = ~n20291 & ~n21067;
  assign n21069 = n21068 ^ n21001;
  assign n21070 = n21034 & ~n21069;
  assign n21071 = n21065 & ~n21070;
  assign n21072 = n21071 ^ n19946;
  assign n21073 = n19551 ^ x796;
  assign n21228 = ~n20754 & ~n20755;
  assign n21229 = ~n20790 & n20814;
  assign n21230 = n21229 ^ n20819;
  assign n21231 = n21230 ^ n20837;
  assign n21232 = n21231 ^ n20821;
  assign n21233 = n21232 ^ n20823;
  assign n21234 = n21233 ^ n20841;
  assign n21235 = n21228 & ~n21234;
  assign n21236 = ~n20827 & ~n20828;
  assign n21237 = n21236 ^ n20839;
  assign n21238 = n21237 ^ n20755;
  assign n21239 = n21237 ^ n20754;
  assign n21240 = n21237 & n21239;
  assign n21241 = n21240 ^ n21237;
  assign n21242 = ~n21238 & n21241;
  assign n21243 = n21242 ^ n21240;
  assign n21244 = n21243 ^ n21237;
  assign n21245 = n21244 ^ n20754;
  assign n21246 = n20845 ^ n20829;
  assign n21247 = n21246 ^ n20824;
  assign n21248 = n21245 & ~n21247;
  assign n21249 = n21248 ^ n20754;
  assign n21250 = ~n21235 & ~n21249;
  assign n21252 = n20791 & n21231;
  assign n21253 = n20817 ^ n20813;
  assign n21254 = ~n21252 & n21253;
  assign n21251 = n20844 ^ n20814;
  assign n21255 = n21254 ^ n21251;
  assign n21256 = ~n20754 & ~n21255;
  assign n21257 = n21256 ^ n21251;
  assign n21258 = n20755 & ~n21257;
  assign n21259 = n21250 & ~n21258;
  assign n21260 = n21259 ^ n19193;
  assign n21261 = n21260 ^ x798;
  assign n21262 = n20686 & n20699;
  assign n21265 = n20723 ^ n20558;
  assign n21263 = n20706 ^ n20702;
  assign n21264 = n21263 ^ n20715;
  assign n21266 = n21265 ^ n21264;
  assign n21267 = n20682 & n21266;
  assign n21268 = n20745 ^ n20722;
  assign n21269 = n20681 & ~n21268;
  assign n21274 = n20685 & n20710;
  assign n21273 = n20637 & n20698;
  assign n21275 = n21274 ^ n21273;
  assign n21271 = ~n20681 & n20698;
  assign n21270 = n20708 ^ n20692;
  assign n21272 = n21271 ^ n21270;
  assign n21276 = n21275 ^ n21272;
  assign n21277 = ~n21269 & n21276;
  assign n21278 = ~n21267 & ~n21277;
  assign n21280 = n20633 & ~n20683;
  assign n21279 = ~n20562 & n20687;
  assign n21281 = n21280 ^ n21279;
  assign n21282 = n21278 & ~n21281;
  assign n21283 = n20717 ^ n20715;
  assign n21284 = n20681 & n21283;
  assign n21285 = n21284 ^ n20717;
  assign n21286 = n20637 & n21285;
  assign n21287 = n21282 & ~n21286;
  assign n21288 = ~n20683 & n20699;
  assign n21289 = n21288 ^ n20742;
  assign n21290 = n21287 & ~n21289;
  assign n21291 = ~n20737 & n21290;
  assign n21292 = n20627 & n20682;
  assign n21293 = n21292 ^ n20688;
  assign n21294 = n21291 & ~n21293;
  assign n21295 = ~n21262 & n21294;
  assign n21296 = n21295 ^ n18764;
  assign n21297 = n21296 ^ x797;
  assign n21298 = ~n21261 & ~n21297;
  assign n21299 = n21298 ^ n21297;
  assign n21074 = n20148 ^ x777;
  assign n21075 = n20328 ^ x772;
  assign n21076 = n20460 ^ x773;
  assign n21077 = n19434 ^ n19427;
  assign n21078 = n21077 ^ n19459;
  assign n21079 = n19460 & n21078;
  assign n21085 = n19454 ^ n19428;
  assign n21086 = n21085 ^ n19426;
  assign n21080 = n19468 ^ n19453;
  assign n21081 = n21080 ^ n19431;
  assign n21082 = ~n19326 & n21081;
  assign n21083 = n21082 ^ n19431;
  assign n21084 = ~n19414 & n21083;
  assign n21087 = n21086 ^ n21084;
  assign n21088 = n21087 ^ n21084;
  assign n21089 = n19327 & ~n21088;
  assign n21090 = n21089 ^ n21084;
  assign n21091 = n20670 & ~n21090;
  assign n21092 = n21091 ^ n21084;
  assign n21093 = ~n21079 & n21092;
  assign n21094 = ~n19448 & n21093;
  assign n21095 = ~n20677 & n21094;
  assign n21096 = ~n19442 & n21095;
  assign n21097 = n21096 ^ n17783;
  assign n21098 = n21097 ^ x775;
  assign n21099 = n21076 & n21098;
  assign n21100 = n21099 ^ n21076;
  assign n21102 = n20230 ^ x776;
  assign n21103 = n18619 ^ n18600;
  assign n21104 = n21103 ^ n17756;
  assign n21105 = n21104 ^ x774;
  assign n21106 = ~n21102 & n21105;
  assign n21107 = n21106 ^ n21102;
  assign n21139 = n21100 & ~n21107;
  assign n21140 = n21139 ^ n21099;
  assign n21125 = n21107 ^ n21098;
  assign n21126 = n21076 & ~n21125;
  assign n21141 = n21140 ^ n21126;
  assign n21112 = n21106 ^ n21105;
  assign n21128 = n21099 & n21112;
  assign n21119 = n21105 ^ n21102;
  assign n21120 = n21119 ^ n21098;
  assign n21129 = n21128 ^ n21120;
  assign n21121 = ~n21076 & ~n21120;
  assign n21127 = n21126 ^ n21121;
  assign n21130 = n21129 ^ n21127;
  assign n21142 = n21141 ^ n21130;
  assign n21101 = n21100 ^ n21098;
  assign n21113 = ~n21101 & n21112;
  assign n21143 = n21142 ^ n21113;
  assign n21133 = n21102 ^ n21098;
  assign n21135 = n21105 ^ n21098;
  assign n21136 = n21135 ^ n21076;
  assign n21137 = n21133 & n21136;
  assign n21134 = n21076 & n21133;
  assign n21138 = n21137 ^ n21134;
  assign n21144 = n21143 ^ n21138;
  assign n21117 = n21099 ^ n21098;
  assign n21118 = n21106 & n21117;
  assign n21122 = n21121 ^ n21118;
  assign n21114 = n21113 ^ n21101;
  assign n21110 = ~n21101 & n21106;
  assign n21108 = n21107 ^ n21105;
  assign n21109 = ~n21101 & n21108;
  assign n21111 = n21110 ^ n21109;
  assign n21115 = n21114 ^ n21111;
  assign n21116 = n21115 ^ n21113;
  assign n21123 = n21122 ^ n21116;
  assign n21145 = n21144 ^ n21123;
  assign n21154 = ~n21075 & n21145;
  assign n21155 = n21154 ^ n21144;
  assign n21149 = n21099 & n21108;
  assign n21150 = n21149 ^ n21137;
  assign n21132 = n21118 ^ n21117;
  assign n21146 = n21145 ^ n21132;
  assign n21124 = n21123 ^ n21115;
  assign n21131 = n21130 ^ n21124;
  assign n21147 = n21146 ^ n21131;
  assign n21148 = n21147 ^ n21137;
  assign n21151 = n21150 ^ n21148;
  assign n21152 = ~n21075 & n21151;
  assign n21153 = n21152 ^ n21148;
  assign n21156 = n21155 ^ n21153;
  assign n21157 = n21074 & ~n21156;
  assign n21158 = n21157 ^ n21153;
  assign n21163 = n21146 ^ n21116;
  assign n21159 = ~n21074 & ~n21075;
  assign n21160 = n21159 ^ n21075;
  assign n21164 = n21160 ^ n21074;
  assign n21165 = ~n21163 & ~n21164;
  assign n21162 = ~n21075 & n21109;
  assign n21166 = n21165 ^ n21162;
  assign n21161 = ~n21143 & ~n21160;
  assign n21167 = n21166 ^ n21161;
  assign n21168 = ~n21158 & ~n21167;
  assign n21170 = n21100 & n21108;
  assign n21171 = n21170 ^ n21134;
  assign n21172 = n21171 ^ n21142;
  assign n21173 = ~n21164 & ~n21172;
  assign n21169 = n21139 & ~n21160;
  assign n21174 = n21173 ^ n21169;
  assign n21175 = n21168 & ~n21174;
  assign n21179 = ~n21144 & ~n21160;
  assign n21176 = n21075 ^ n21074;
  assign n21177 = n21100 & ~n21176;
  assign n21178 = n21106 & n21177;
  assign n21180 = n21179 ^ n21178;
  assign n21181 = n21175 & ~n21180;
  assign n21182 = n21170 ^ n21141;
  assign n21183 = n21074 & n21182;
  assign n21184 = n21183 ^ n21118;
  assign n21185 = n21075 & n21184;
  assign n21186 = n21185 ^ n21118;
  assign n21187 = n21181 & ~n21186;
  assign n21188 = n21187 ^ n18329;
  assign n21189 = n21188 ^ x800;
  assign n21190 = n20415 ^ n20409;
  assign n21191 = ~n20463 & n21190;
  assign n21192 = n20422 & n20464;
  assign n21193 = n20417 & n20462;
  assign n21194 = n20465 & n20485;
  assign n21201 = n20499 ^ n20492;
  assign n21202 = n21201 ^ n20400;
  assign n21197 = ~n20463 & ~n20477;
  assign n21198 = n21197 ^ n20494;
  assign n21199 = n21198 ^ n20400;
  assign n21195 = n20420 ^ n20406;
  assign n21196 = n20462 & n21195;
  assign n21200 = n21199 ^ n21196;
  assign n21203 = n21202 ^ n21200;
  assign n21204 = n21203 ^ n21200;
  assign n21205 = ~n20461 & n21204;
  assign n21206 = n21205 ^ n21200;
  assign n21207 = n20425 & ~n21206;
  assign n21208 = n21207 ^ n21200;
  assign n21209 = ~n21194 & n21208;
  assign n21210 = ~n21193 & n21209;
  assign n21211 = ~n21192 & n21210;
  assign n21213 = ~n20425 & ~n20474;
  assign n21212 = n20472 & n20505;
  assign n21214 = n21213 ^ n21212;
  assign n21215 = n21211 & ~n21214;
  assign n21216 = ~n21191 & n21215;
  assign n21217 = n20423 ^ n20411;
  assign n21218 = n21217 ^ n20422;
  assign n21219 = n20425 & ~n21218;
  assign n21220 = n21219 ^ n20422;
  assign n21221 = ~n20461 & n21220;
  assign n21222 = n21216 & ~n21221;
  assign n21223 = n21222 ^ n19178;
  assign n21224 = n21223 ^ x799;
  assign n21225 = n21189 & ~n21224;
  assign n21315 = n21225 ^ n21189;
  assign n21316 = ~n21299 & n21315;
  assign n21317 = n21316 ^ n21299;
  assign n21226 = n21225 ^ n21224;
  assign n21311 = ~n21226 & ~n21299;
  assign n21304 = n21224 ^ n21189;
  assign n21305 = n21298 & ~n21304;
  assign n21312 = n21311 ^ n21305;
  assign n21308 = n21305 ^ n21298;
  assign n21307 = n21225 & n21298;
  assign n21309 = n21308 ^ n21307;
  assign n21313 = n21312 ^ n21309;
  assign n21303 = n21225 & ~n21299;
  assign n21306 = n21305 ^ n21303;
  assign n21310 = n21309 ^ n21306;
  assign n21314 = n21313 ^ n21310;
  assign n21318 = n21317 ^ n21314;
  assign n21227 = n21226 ^ n21189;
  assign n21300 = n21299 ^ n21261;
  assign n21301 = n21300 ^ n21297;
  assign n21302 = n21227 & ~n21301;
  assign n21319 = n21318 ^ n21302;
  assign n21320 = ~n21073 & ~n21319;
  assign n21321 = ~n21261 & n21315;
  assign n21322 = n20916 & n20936;
  assign n21323 = n20949 ^ n20946;
  assign n21324 = n21323 ^ n20943;
  assign n21325 = ~n20955 & n21324;
  assign n21335 = n20938 ^ n20924;
  assign n21336 = n21335 ^ n20925;
  assign n21334 = n20904 ^ n20880;
  assign n21337 = n21336 ^ n21334;
  assign n21328 = n20966 ^ n20940;
  assign n21333 = n21328 ^ n20942;
  assign n21338 = n21337 ^ n21333;
  assign n21339 = n20914 & ~n21338;
  assign n21340 = n21339 ^ n21333;
  assign n21329 = n21328 ^ n20938;
  assign n21330 = ~n20931 & n21329;
  assign n21331 = n21330 ^ n20938;
  assign n21326 = n20957 ^ n20928;
  assign n21327 = ~n20917 & ~n21326;
  assign n21332 = n21331 ^ n21327;
  assign n21341 = n21340 ^ n21332;
  assign n21342 = ~n20915 & n21341;
  assign n21343 = n21342 ^ n21332;
  assign n21344 = ~n20960 & ~n21343;
  assign n21345 = ~n20979 & n21344;
  assign n21346 = ~n21325 & n21345;
  assign n21347 = ~n21322 & n21346;
  assign n21351 = n20945 ^ n20934;
  assign n21348 = n20950 ^ n20923;
  assign n21349 = n20915 & n21348;
  assign n21350 = n21349 ^ n20950;
  assign n21352 = n21351 ^ n21350;
  assign n21353 = n21352 ^ n21350;
  assign n21354 = n20915 & n21353;
  assign n21355 = n21354 ^ n21350;
  assign n21356 = ~n20914 & n21355;
  assign n21357 = n21356 ^ n21350;
  assign n21358 = n21347 & ~n21357;
  assign n21359 = n21358 ^ n18358;
  assign n21360 = n21359 ^ x801;
  assign n21361 = n21073 & n21360;
  assign n21362 = n21361 ^ n21360;
  assign n21363 = n21362 ^ n21073;
  assign n21364 = n21321 & ~n21363;
  assign n21365 = ~n21320 & ~n21364;
  assign n21370 = n21321 ^ n21305;
  assign n21369 = ~n21301 & n21315;
  assign n21371 = n21370 ^ n21369;
  assign n21372 = n21371 ^ n21303;
  assign n21366 = n21316 ^ n21315;
  assign n21367 = n21366 ^ n21321;
  assign n21368 = n21367 ^ n21302;
  assign n21373 = n21372 ^ n21368;
  assign n21374 = ~n21073 & n21373;
  assign n21375 = n21374 ^ n21368;
  assign n21376 = n21360 & n21375;
  assign n21377 = n21365 & ~n21376;
  assign n21384 = n21302 ^ n21300;
  assign n21380 = ~n21300 & n21304;
  assign n21383 = n21380 ^ n21368;
  assign n21385 = n21384 ^ n21383;
  assign n21379 = n21225 & ~n21300;
  assign n21381 = n21380 ^ n21379;
  assign n21382 = n21381 ^ n21369;
  assign n21386 = n21385 ^ n21382;
  assign n21378 = n21225 & ~n21301;
  assign n21387 = n21386 ^ n21378;
  assign n21388 = n21360 ^ n21073;
  assign n21389 = ~n21387 & n21388;
  assign n21390 = n21389 ^ n21378;
  assign n21400 = n21372 ^ n21307;
  assign n21401 = n21400 ^ n21309;
  assign n21396 = n21305 ^ n21297;
  assign n21393 = n21385 ^ n21378;
  assign n21394 = n21393 ^ n21369;
  assign n21392 = n21383 ^ n21305;
  assign n21395 = n21394 ^ n21392;
  assign n21397 = n21396 ^ n21395;
  assign n21391 = n21316 ^ n21309;
  assign n21398 = n21397 ^ n21391;
  assign n21399 = n21398 ^ n21311;
  assign n21402 = n21401 ^ n21399;
  assign n21403 = ~n21360 & ~n21402;
  assign n21404 = n21403 ^ n21399;
  assign n21405 = n21073 & ~n21404;
  assign n21406 = ~n21390 & ~n21405;
  assign n21407 = n21377 & n21406;
  assign n21414 = n21379 & ~n21388;
  assign n21410 = n21367 ^ n21307;
  assign n21411 = ~n21073 & n21410;
  assign n21412 = n21411 ^ n21367;
  assign n21413 = n21388 & n21412;
  assign n21415 = n21414 ^ n21413;
  assign n21408 = n21316 ^ n21311;
  assign n21409 = ~n21363 & n21408;
  assign n21416 = n21415 ^ n21409;
  assign n21417 = n21407 & ~n21416;
  assign n21418 = n21417 ^ n19297;
  assign n21419 = n19987 ^ n19964;
  assign n21420 = n19948 ^ n19803;
  assign n21421 = n21419 & n21420;
  assign n21422 = n19961 & n19966;
  assign n21423 = ~n19949 & n19968;
  assign n21424 = ~n19949 & n19975;
  assign n21425 = n19977 ^ n19956;
  assign n21426 = n21425 ^ n19959;
  assign n21427 = n21426 ^ n19990;
  assign n21428 = n21427 ^ n19990;
  assign n21429 = n19947 & ~n21428;
  assign n21430 = n21429 ^ n19990;
  assign n21431 = ~n19966 & n21430;
  assign n21432 = n21431 ^ n19990;
  assign n21433 = ~n21424 & ~n21432;
  assign n21434 = ~n21423 & n21433;
  assign n21435 = ~n19950 & n21434;
  assign n21436 = ~n21422 & n21435;
  assign n21437 = ~n21421 & n21436;
  assign n21439 = n19967 ^ n19962;
  assign n21440 = ~n19947 & ~n21439;
  assign n21441 = n21440 ^ n19962;
  assign n21438 = ~n19947 & n19951;
  assign n21442 = n21441 ^ n21438;
  assign n21443 = n21442 ^ n21438;
  assign n21444 = ~n19954 & ~n21443;
  assign n21445 = n21444 ^ n21438;
  assign n21446 = ~n19803 & ~n21445;
  assign n21447 = n21446 ^ n21438;
  assign n21448 = n21437 & ~n21447;
  assign n21453 = ~n19947 & n19960;
  assign n21449 = n19975 ^ n19764;
  assign n21450 = n21449 ^ n19952;
  assign n21451 = n19947 & n21450;
  assign n21452 = n21451 ^ n19952;
  assign n21454 = n21453 ^ n21452;
  assign n21455 = ~n19803 & n21454;
  assign n21456 = n21455 ^ n21452;
  assign n21457 = n21448 & ~n21456;
  assign n21458 = n21457 ^ n18915;
  assign n21459 = n21361 ^ n21073;
  assign n21460 = n21302 & n21459;
  assign n21468 = n21316 ^ n21312;
  assign n21469 = n21073 & n21468;
  assign n21463 = n21391 ^ n21307;
  assign n21464 = n21463 ^ n21318;
  assign n21461 = n21397 ^ n21318;
  assign n21462 = n21461 ^ n21368;
  assign n21465 = n21464 ^ n21462;
  assign n21466 = n21073 & ~n21465;
  assign n21467 = n21466 ^ n21462;
  assign n21470 = n21469 ^ n21467;
  assign n21471 = ~n21388 & n21470;
  assign n21472 = n21471 ^ n21467;
  assign n21473 = ~n21460 & ~n21472;
  assign n21479 = ~n21073 & n21303;
  assign n21478 = n21307 & ~n21363;
  assign n21480 = n21479 ^ n21478;
  assign n21476 = n21309 & n21362;
  assign n21474 = n21397 ^ n21382;
  assign n21475 = ~n21388 & ~n21474;
  assign n21477 = n21476 ^ n21475;
  assign n21481 = n21480 ^ n21477;
  assign n21482 = n21473 & ~n21481;
  assign n21483 = n21393 ^ n21311;
  assign n21484 = n21073 & ~n21483;
  assign n21485 = n21484 ^ n21311;
  assign n21486 = n21388 & n21485;
  assign n21487 = n21482 & ~n21486;
  assign n21488 = ~n21416 & n21487;
  assign n21489 = n21488 ^ n20328;
  assign n21490 = n21149 ^ n21130;
  assign n21491 = ~n21160 & ~n21490;
  assign n21492 = n21110 & ~n21164;
  assign n21500 = n21182 ^ n21109;
  assign n21501 = n21500 ^ n21131;
  assign n21502 = n21501 ^ n21148;
  assign n21503 = n21074 & ~n21502;
  assign n21504 = n21503 ^ n21148;
  assign n21495 = n21139 ^ n21111;
  assign n21496 = n21495 ^ n21150;
  assign n21493 = n21163 ^ n21144;
  assign n21494 = n21493 ^ n21172;
  assign n21497 = n21496 ^ n21494;
  assign n21498 = ~n21074 & ~n21497;
  assign n21499 = n21498 ^ n21494;
  assign n21505 = n21504 ^ n21499;
  assign n21506 = n21176 & ~n21505;
  assign n21507 = n21506 ^ n21504;
  assign n21508 = ~n21492 & ~n21507;
  assign n21509 = ~n21174 & n21508;
  assign n21510 = ~n21491 & n21509;
  assign n21511 = n21510 ^ n17887;
  assign n21544 = n21458 ^ x820;
  assign n21512 = ~n20425 & ~n20477;
  assign n21513 = n21512 ^ n20491;
  assign n21514 = n20461 & n21513;
  assign n21515 = n21514 ^ n20491;
  assign n21522 = n20473 ^ n20329;
  assign n21523 = n21522 ^ n20519;
  assign n21521 = n20366 ^ n20330;
  assign n21524 = n21523 ^ n21521;
  assign n21517 = n20474 ^ n20424;
  assign n21516 = n20480 ^ n20420;
  assign n21518 = n21517 ^ n21516;
  assign n21519 = n20461 & ~n21518;
  assign n21520 = n21519 ^ n21516;
  assign n21525 = n21524 ^ n21520;
  assign n21526 = n21525 ^ n21520;
  assign n21527 = n20461 & ~n21526;
  assign n21528 = n21527 ^ n21520;
  assign n21529 = ~n20505 & ~n21528;
  assign n21530 = n21529 ^ n21520;
  assign n21531 = ~n21191 & n21530;
  assign n21532 = n20472 ^ n20416;
  assign n21533 = n21532 ^ n20400;
  assign n21534 = n20505 & n21533;
  assign n21535 = n21534 ^ n21532;
  assign n21536 = n21531 & ~n21535;
  assign n21537 = ~n21515 & n21536;
  assign n21538 = n20462 & ~n20494;
  assign n21539 = n21538 ^ n21197;
  assign n21540 = n21537 & ~n21539;
  assign n21541 = ~n20522 & n21540;
  assign n21542 = n21541 ^ n19363;
  assign n21543 = n21542 ^ x825;
  assign n21545 = n21544 ^ n21543;
  assign n21616 = n20850 ^ n20848;
  assign n21617 = n21616 ^ n19611;
  assign n21618 = n21617 ^ x822;
  assign n21619 = n19149 ^ n19121;
  assign n21620 = n21619 ^ n19111;
  assign n21621 = n19510 & n21620;
  assign n21622 = n19115 & n19509;
  assign n21623 = n19145 ^ n19109;
  assign n21624 = n21623 ^ n19134;
  assign n21625 = ~n19298 & n21624;
  assign n21626 = ~n21622 & ~n21625;
  assign n21627 = n19531 ^ n19116;
  assign n21628 = n21627 ^ n19136;
  assign n21629 = n19298 & n21628;
  assign n21630 = n21629 ^ n19136;
  assign n21631 = ~n19507 & n21630;
  assign n21632 = n21626 & ~n21631;
  assign n21633 = ~n21621 & n21632;
  assign n21634 = n19150 ^ n19131;
  assign n21635 = n21634 ^ n19109;
  assign n21636 = n21635 ^ n19139;
  assign n21637 = ~n19507 & ~n21636;
  assign n21638 = n21637 ^ n19139;
  assign n21639 = n19298 & n21638;
  assign n21640 = n21633 & ~n21639;
  assign n21641 = ~n19124 & ~n19298;
  assign n21642 = n21641 ^ n19122;
  assign n21643 = ~n19509 & ~n21642;
  assign n21644 = n21640 & ~n21643;
  assign n21645 = n19535 ^ n19145;
  assign n21646 = ~n19298 & n21645;
  assign n21647 = n21646 ^ n19145;
  assign n21648 = ~n19509 & n21647;
  assign n21649 = n21644 & ~n21648;
  assign n21650 = n19136 ^ n19119;
  assign n21651 = ~n19298 & n21650;
  assign n21652 = n21651 ^ n19136;
  assign n21653 = ~n19507 & n21652;
  assign n21654 = n21649 & ~n21653;
  assign n21655 = ~n19549 & n21654;
  assign n21656 = n21655 ^ n19036;
  assign n21657 = n21656 ^ x821;
  assign n21658 = n21618 & ~n21657;
  assign n21546 = n20233 & n20245;
  assign n21549 = n20184 & n20253;
  assign n21550 = ~n20154 & n21549;
  assign n21551 = n20248 ^ n20159;
  assign n21552 = ~n20232 & n21551;
  assign n21553 = ~n21550 & ~n21552;
  assign n21554 = ~n20267 & ~n21553;
  assign n21547 = n20240 ^ n20166;
  assign n21548 = n20196 & n21547;
  assign n21555 = n21554 ^ n21548;
  assign n21556 = ~n20231 & ~n21555;
  assign n21557 = n21556 ^ n21554;
  assign n21558 = ~n21546 & n21557;
  assign n21559 = n20231 ^ n20196;
  assign n21560 = n20184 ^ n20161;
  assign n21561 = n21560 ^ n20251;
  assign n21562 = n21561 ^ n20162;
  assign n21563 = ~n20231 & n21562;
  assign n21564 = n21563 ^ n20162;
  assign n21565 = ~n21559 & n21564;
  assign n21566 = n21558 & ~n21565;
  assign n21567 = n20171 & ~n20231;
  assign n21568 = n21567 ^ n20165;
  assign n21569 = n20196 & n21568;
  assign n21570 = n21566 & ~n21569;
  assign n21571 = ~n20286 & n21570;
  assign n21572 = n20236 ^ n20173;
  assign n21573 = n20196 & n21572;
  assign n21574 = n21573 ^ n20236;
  assign n21575 = ~n20231 & n21574;
  assign n21576 = n21571 & ~n21575;
  assign n21577 = n21576 ^ n19638;
  assign n21578 = n21577 ^ x823;
  assign n21579 = n20938 ^ n20929;
  assign n21580 = n21579 ^ n20942;
  assign n21581 = ~n20917 & n21580;
  assign n21582 = n20950 ^ n20928;
  assign n21583 = ~n20955 & n21582;
  assign n21586 = n20966 ^ n20957;
  assign n21584 = n20936 ^ n20909;
  assign n21585 = n21584 ^ n20967;
  assign n21587 = n21586 ^ n21585;
  assign n21588 = n20914 & ~n21587;
  assign n21589 = n21588 ^ n21585;
  assign n21590 = ~n20915 & n21589;
  assign n21591 = ~n21583 & ~n21590;
  assign n21592 = n20947 ^ n20915;
  assign n21593 = n20949 ^ n20945;
  assign n21594 = n21593 ^ n21584;
  assign n21595 = ~n20914 & n21594;
  assign n21596 = n21595 ^ n21584;
  assign n21597 = n21596 ^ n20947;
  assign n21598 = ~n21592 & n21597;
  assign n21599 = n21598 ^ n21595;
  assign n21600 = n21599 ^ n21584;
  assign n21601 = n21600 ^ n20915;
  assign n21602 = ~n20947 & ~n21601;
  assign n21603 = n21602 ^ n20947;
  assign n21604 = n21603 ^ n20915;
  assign n21605 = n21591 & n21604;
  assign n21606 = ~n21581 & n21605;
  assign n21607 = ~n20915 & n21593;
  assign n21608 = n21607 ^ n20949;
  assign n21609 = n20914 & n21608;
  assign n21610 = n21606 & ~n21609;
  assign n21611 = ~n20974 & n21610;
  assign n21612 = ~n20971 & n21611;
  assign n21613 = ~n20979 & n21612;
  assign n21614 = n21613 ^ n19325;
  assign n21615 = n21614 ^ x824;
  assign n21673 = ~n21578 & ~n21615;
  assign n21686 = n21658 & n21673;
  assign n21687 = n21686 ^ n21673;
  assign n21659 = n21658 ^ n21618;
  assign n21660 = n21615 & n21659;
  assign n21683 = n21660 ^ n21659;
  assign n21674 = n21673 ^ n21615;
  assign n21675 = n21659 & ~n21674;
  assign n21684 = n21683 ^ n21675;
  assign n21663 = n21658 ^ n21657;
  assign n21664 = n21663 ^ n21618;
  assign n21665 = n21615 & n21664;
  assign n21678 = n21578 & n21665;
  assign n21679 = n21678 ^ n21665;
  assign n21680 = n21679 ^ n21674;
  assign n21661 = ~n21578 & n21660;
  assign n21676 = n21675 ^ n21661;
  assign n21669 = n21615 ^ n21578;
  assign n21670 = n21578 & n21618;
  assign n21671 = n21670 ^ n21657;
  assign n21672 = n21669 & n21671;
  assign n21677 = n21676 ^ n21672;
  assign n21681 = n21680 ^ n21677;
  assign n21667 = n21615 & ~n21663;
  assign n21668 = n21667 ^ n21663;
  assign n21682 = n21681 ^ n21668;
  assign n21685 = n21684 ^ n21682;
  assign n21688 = n21687 ^ n21685;
  assign n21666 = n21665 ^ n21664;
  assign n21689 = n21688 ^ n21666;
  assign n21662 = n21661 ^ n21660;
  assign n21690 = n21689 ^ n21662;
  assign n21691 = n21545 & n21690;
  assign n21692 = n21615 & n21658;
  assign n21697 = n21692 ^ n21658;
  assign n21698 = n21697 ^ n21686;
  assign n21695 = n21578 & n21667;
  assign n21696 = n21695 ^ n21667;
  assign n21699 = n21698 ^ n21696;
  assign n21694 = n21685 ^ n21661;
  assign n21700 = n21699 ^ n21694;
  assign n21693 = n21692 ^ n21682;
  assign n21701 = n21700 ^ n21693;
  assign n21702 = ~n21543 & n21701;
  assign n21703 = n21702 ^ n21693;
  assign n21704 = n21544 & n21703;
  assign n21705 = ~n21691 & ~n21704;
  assign n21706 = ~n21543 & n21544;
  assign n21707 = n21706 ^ n21543;
  assign n21714 = n21707 ^ n21544;
  assign n21708 = ~n21578 & n21692;
  assign n21709 = n21708 ^ n21692;
  assign n21710 = n21709 ^ n21696;
  assign n21711 = n21710 ^ n21695;
  assign n21712 = n21711 ^ n21672;
  assign n21713 = ~n21707 & ~n21712;
  assign n21715 = n21714 ^ n21713;
  assign n21716 = ~n21686 & n21715;
  assign n21717 = n21716 ^ n21714;
  assign n21718 = n21705 & ~n21717;
  assign n21719 = n21699 ^ n21686;
  assign n21720 = ~n21544 & n21719;
  assign n21721 = n21720 ^ n21686;
  assign n21722 = n21543 & n21721;
  assign n21723 = n21718 & ~n21722;
  assign n21729 = n21706 ^ n21544;
  assign n21730 = n21689 & n21729;
  assign n21724 = n21684 ^ n21679;
  assign n21725 = n21724 ^ n21676;
  assign n21726 = ~n21544 & n21725;
  assign n21727 = n21726 ^ n21676;
  assign n21728 = n21543 & n21727;
  assign n21731 = n21730 ^ n21728;
  assign n21732 = n21723 & ~n21731;
  assign n21737 = n21679 & n21729;
  assign n21733 = n21708 ^ n21695;
  assign n21734 = ~n21543 & n21733;
  assign n21735 = n21734 ^ n21695;
  assign n21736 = n21545 & n21735;
  assign n21738 = n21737 ^ n21736;
  assign n21739 = n21732 & ~n21738;
  assign n21740 = n21739 ^ n20045;
  assign n21741 = ~n21142 & ~n21164;
  assign n21742 = n21172 ^ n21130;
  assign n21743 = ~n21160 & n21742;
  assign n21744 = n21074 & n21127;
  assign n21745 = n21744 ^ n21126;
  assign n21746 = ~n21176 & n21745;
  assign n21747 = n21176 ^ n21118;
  assign n21748 = n21146 ^ n21111;
  assign n21749 = n21748 ^ n21074;
  assign n21750 = ~n21118 & ~n21749;
  assign n21751 = n21750 ^ n21074;
  assign n21752 = n21747 & ~n21751;
  assign n21753 = n21752 ^ n21118;
  assign n21754 = ~n21746 & ~n21753;
  assign n21755 = ~n21743 & n21754;
  assign n21756 = ~n21741 & n21755;
  assign n21757 = n21182 ^ n21144;
  assign n21758 = n21757 ^ n21123;
  assign n21759 = n21075 & n21758;
  assign n21760 = n21759 ^ n21123;
  assign n21761 = ~n21074 & ~n21760;
  assign n21762 = n21756 & ~n21761;
  assign n21763 = n21130 ^ n21128;
  assign n21764 = n21074 & ~n21763;
  assign n21765 = n21764 ^ n21130;
  assign n21766 = n21075 & ~n21765;
  assign n21767 = n21762 & ~n21766;
  assign n21768 = n21170 ^ n21116;
  assign n21769 = ~n21074 & ~n21768;
  assign n21770 = n21769 ^ n21170;
  assign n21771 = ~n21075 & n21770;
  assign n21772 = n21767 & ~n21771;
  assign n21773 = ~n21180 & n21772;
  assign n21774 = n21773 ^ n18658;
  assign n21775 = n21708 ^ n21681;
  assign n21776 = n21714 & ~n21775;
  assign n21777 = n21707 ^ n21688;
  assign n21778 = n21729 ^ n21690;
  assign n21779 = ~n21688 & ~n21778;
  assign n21780 = n21779 ^ n21729;
  assign n21781 = ~n21777 & n21780;
  assign n21782 = n21781 ^ n21707;
  assign n21783 = ~n21776 & n21782;
  assign n21784 = n21686 & ~n21707;
  assign n21785 = n21544 & n21578;
  assign n21786 = n21785 ^ n21706;
  assign n21787 = n21665 & n21786;
  assign n21788 = ~n21784 & ~n21787;
  assign n21791 = n21706 ^ n21615;
  assign n21792 = n21578 & ~n21791;
  assign n21793 = n21792 ^ n21615;
  assign n21794 = ~n21663 & ~n21793;
  assign n21789 = n21681 ^ n21675;
  assign n21790 = n21789 ^ n21686;
  assign n21795 = n21794 ^ n21790;
  assign n21796 = n21795 ^ n21790;
  assign n21797 = n21707 & n21796;
  assign n21798 = n21797 ^ n21790;
  assign n21799 = ~n21729 & ~n21798;
  assign n21800 = n21799 ^ n21790;
  assign n21801 = n21543 & n21677;
  assign n21802 = n21801 ^ n21676;
  assign n21803 = n21545 & n21802;
  assign n21804 = n21800 & ~n21803;
  assign n21805 = n21710 ^ n21707;
  assign n21806 = n21729 ^ n21684;
  assign n21807 = n21707 & ~n21806;
  assign n21808 = n21807 ^ n21684;
  assign n21809 = ~n21805 & n21808;
  assign n21810 = n21809 ^ n21710;
  assign n21811 = n21804 & ~n21810;
  assign n21812 = n21698 ^ n21678;
  assign n21813 = ~n21544 & n21812;
  assign n21814 = n21813 ^ n21698;
  assign n21815 = ~n21543 & n21814;
  assign n21816 = n21811 & ~n21815;
  assign n21817 = n21788 & n21816;
  assign n21818 = ~n21738 & n21817;
  assign n21819 = n21783 & n21818;
  assign n21820 = n21819 ^ n20903;
  assign n21821 = n20154 & ~n20196;
  assign n21822 = n21821 ^ n20170;
  assign n21823 = ~n20231 & n21822;
  assign n21824 = n21823 ^ n20170;
  assign n21825 = n20267 ^ n20162;
  assign n21826 = n21825 ^ n20181;
  assign n21827 = n21826 ^ n20258;
  assign n21828 = ~n20231 & n21827;
  assign n21829 = n21828 ^ n20258;
  assign n21830 = n20196 & n21829;
  assign n21831 = ~n21824 & ~n21830;
  assign n21832 = n20173 & ~n21559;
  assign n21833 = n20184 ^ n20160;
  assign n21834 = n20233 & n21833;
  assign n21835 = n20169 & n20231;
  assign n21836 = n21835 ^ n20176;
  assign n21837 = n21559 & n21836;
  assign n21838 = n21837 ^ n20176;
  assign n21843 = n20157 & ~n20231;
  assign n21839 = n20185 ^ n20154;
  assign n21840 = n21839 ^ n20180;
  assign n21841 = ~n20231 & n21840;
  assign n21842 = n21841 ^ n20180;
  assign n21844 = n21843 ^ n21842;
  assign n21845 = ~n20196 & n21844;
  assign n21846 = n21845 ^ n21842;
  assign n21847 = ~n21838 & ~n21846;
  assign n21848 = ~n21575 & n21847;
  assign n21849 = ~n21834 & n21848;
  assign n21850 = ~n21832 & n21849;
  assign n21851 = n21831 & n21850;
  assign n21852 = ~n20235 & n21851;
  assign n21853 = n21852 ^ n18400;
  assign n21854 = n20755 ^ n20754;
  assign n21858 = n21254 ^ n21237;
  assign n21859 = ~n20755 & ~n21858;
  assign n21860 = n21859 ^ n21254;
  assign n21855 = n21251 ^ n21234;
  assign n21856 = ~n20755 & ~n21855;
  assign n21857 = n21856 ^ n21251;
  assign n21861 = n21860 ^ n21857;
  assign n21862 = ~n21854 & n21861;
  assign n21863 = n21862 ^ n21857;
  assign n21864 = ~n21247 & n21863;
  assign n21865 = n21864 ^ n17431;
  assign n21866 = n21865 ^ x831;
  assign n21867 = n21614 ^ x826;
  assign n21868 = n21866 & ~n21867;
  assign n21869 = n21868 ^ n21866;
  assign n21870 = n21542 ^ x827;
  assign n21902 = ~n20635 & n20681;
  assign n21903 = n20708 ^ n20698;
  assign n21904 = n20681 & n21903;
  assign n21905 = n21904 ^ n20698;
  assign n21906 = n20637 & n21905;
  assign n21907 = ~n21902 & ~n21906;
  assign n21913 = ~n20637 & ~n21263;
  assign n21909 = n20711 ^ n20632;
  assign n21908 = n20740 ^ n20724;
  assign n21910 = n21909 ^ n21908;
  assign n21911 = n20637 & ~n21910;
  assign n21912 = n21911 ^ n21908;
  assign n21914 = n21913 ^ n21912;
  assign n21915 = n20681 & ~n21914;
  assign n21916 = n21915 ^ n21912;
  assign n21918 = n20637 & n20714;
  assign n21917 = n20686 & n20717;
  assign n21919 = n21918 ^ n21917;
  assign n21920 = n21916 & ~n21919;
  assign n21921 = ~n21289 & n21920;
  assign n21922 = n21907 & n21921;
  assign n21923 = ~n20684 & n21922;
  assign n21924 = ~n20749 & n21923;
  assign n21925 = ~n21262 & n21924;
  assign n21926 = n21925 ^ n19387;
  assign n21927 = n21926 ^ x829;
  assign n21941 = n21927 ^ n21870;
  assign n21928 = n21511 ^ x830;
  assign n21942 = n21941 ^ n21928;
  assign n21943 = ~n21870 & n21942;
  assign n21871 = n19962 ^ n19951;
  assign n21872 = n21871 ^ n19971;
  assign n21873 = n19948 & n21872;
  assign n21874 = n19947 & n19968;
  assign n21880 = n21449 ^ n19971;
  assign n21881 = n21880 ^ n19954;
  assign n21882 = n21881 ^ n19987;
  assign n21883 = n21882 ^ n19964;
  assign n21884 = n19947 & n21883;
  assign n21885 = n21884 ^ n19964;
  assign n21876 = n19997 ^ n19996;
  assign n21875 = n19952 ^ n19767;
  assign n21877 = n21876 ^ n21875;
  assign n21878 = ~n19947 & n21877;
  assign n21879 = n21878 ^ n21875;
  assign n21886 = n21885 ^ n21879;
  assign n21887 = n19966 & n21886;
  assign n21888 = n21887 ^ n21879;
  assign n21889 = ~n21874 & ~n21888;
  assign n21890 = ~n20014 & n21889;
  assign n21891 = ~n19958 & n21890;
  assign n21892 = ~n21873 & n21891;
  assign n21893 = ~n21456 & n21892;
  assign n21894 = ~n21423 & n21893;
  assign n21895 = ~n20027 & n21894;
  assign n21896 = n19956 & n21895;
  assign n21897 = n21896 ^ n19411;
  assign n21898 = n21897 ^ x828;
  assign n21899 = n21870 & n21898;
  assign n21900 = n21899 ^ n21870;
  assign n21901 = n21900 ^ n21898;
  assign n21929 = n21927 & ~n21928;
  assign n21936 = ~n21901 & n21929;
  assign n21944 = n21943 ^ n21936;
  assign n21932 = n21899 ^ n21898;
  assign n21938 = n21929 & n21932;
  assign n21930 = n21929 ^ n21927;
  assign n21933 = n21930 ^ n21928;
  assign n21934 = n21932 & n21933;
  assign n21939 = n21938 ^ n21934;
  assign n21945 = n21944 ^ n21939;
  assign n21946 = n21945 ^ n21938;
  assign n21947 = n21946 ^ n21901;
  assign n21931 = ~n21901 & n21930;
  assign n21935 = n21934 ^ n21931;
  assign n21937 = n21936 ^ n21935;
  assign n21940 = n21939 ^ n21937;
  assign n21948 = n21947 ^ n21940;
  assign n21949 = n21869 & ~n21948;
  assign n21958 = n21899 & ~n21927;
  assign n21950 = n21929 ^ n21928;
  assign n21959 = n21958 ^ n21950;
  assign n21952 = n21900 & n21933;
  assign n21953 = n21952 ^ n21938;
  assign n21954 = n21953 ^ n21933;
  assign n21955 = n21954 ^ n21944;
  assign n21951 = n21900 & ~n21950;
  assign n21956 = n21955 ^ n21951;
  assign n21957 = n21956 ^ n21948;
  assign n21960 = n21959 ^ n21957;
  assign n21961 = n21960 ^ n21945;
  assign n21962 = n21961 ^ n21952;
  assign n21963 = ~n21867 & n21962;
  assign n21964 = n21963 ^ n21952;
  assign n21965 = ~n21866 & n21964;
  assign n21966 = ~n21949 & ~n21965;
  assign n21968 = n21899 & n21928;
  assign n21969 = n21968 ^ n21955;
  assign n21967 = n21900 & n21929;
  assign n21970 = n21969 ^ n21967;
  assign n21971 = n21868 ^ n21867;
  assign n21972 = n21970 & ~n21971;
  assign n21973 = n21868 & n21934;
  assign n21977 = n21969 ^ n21930;
  assign n21974 = n21939 ^ n21932;
  assign n21975 = n21974 ^ n21960;
  assign n21976 = n21975 ^ n21931;
  assign n21978 = n21977 ^ n21976;
  assign n21979 = ~n21867 & n21978;
  assign n21982 = n21968 ^ n21946;
  assign n21980 = n21867 & n21940;
  assign n21981 = n21980 ^ n21939;
  assign n21983 = n21982 ^ n21981;
  assign n21984 = n21983 ^ n21981;
  assign n21985 = ~n21867 & n21984;
  assign n21986 = n21985 ^ n21981;
  assign n21987 = n21971 ^ n21869;
  assign n21988 = n21986 & n21987;
  assign n21989 = n21988 ^ n21981;
  assign n21990 = ~n21979 & ~n21989;
  assign n21991 = n21958 ^ n21946;
  assign n21992 = n21991 ^ n21951;
  assign n21993 = n21992 ^ n21951;
  assign n21994 = n21867 & n21993;
  assign n21995 = n21994 ^ n21951;
  assign n21996 = n21987 & n21995;
  assign n21997 = n21996 ^ n21951;
  assign n21998 = n21990 & ~n21997;
  assign n21999 = ~n21973 & n21998;
  assign n22000 = n21958 ^ n21899;
  assign n22001 = n22000 ^ n21969;
  assign n22002 = n22001 ^ n21975;
  assign n22003 = n21866 & n22002;
  assign n22004 = n22003 ^ n21975;
  assign n22005 = n21867 & n22004;
  assign n22006 = n21999 & ~n22005;
  assign n22007 = ~n21972 & n22006;
  assign n22008 = n21967 ^ n21948;
  assign n22009 = ~n21867 & ~n22008;
  assign n22010 = n22009 ^ n21948;
  assign n22011 = n21987 & ~n22010;
  assign n22012 = n22007 & ~n22011;
  assign n22017 = n21968 ^ n21958;
  assign n22018 = n21869 & n22017;
  assign n22013 = n21967 ^ n21960;
  assign n22014 = n21867 & n22013;
  assign n22015 = n22014 ^ n21960;
  assign n22016 = n21987 & n22015;
  assign n22019 = n22018 ^ n22016;
  assign n22020 = n22012 & ~n22019;
  assign n22021 = n21966 & n22020;
  assign n22022 = n22021 ^ n20789;
  assign n22023 = n20681 & ~n20725;
  assign n22024 = n22023 ^ n20632;
  assign n22025 = ~n20637 & n22024;
  assign n22026 = n22025 ^ n20632;
  assign n22027 = n20747 ^ n20722;
  assign n22028 = n22027 ^ n20709;
  assign n22029 = n22028 ^ n21264;
  assign n22030 = ~n20637 & n22029;
  assign n22031 = n22030 ^ n22028;
  assign n22032 = ~n20681 & ~n22031;
  assign n22033 = ~n22026 & ~n22032;
  assign n22034 = n21907 & n22033;
  assign n22035 = ~n20743 & n22034;
  assign n22036 = ~n21293 & n22035;
  assign n22037 = ~n21262 & n22036;
  assign n22038 = n22037 ^ n18980;
  assign n22039 = n21865 ^ x785;
  assign n22040 = n19145 ^ n19123;
  assign n22041 = n19510 & n22040;
  assign n22046 = n19138 ^ n19130;
  assign n22047 = ~n19298 & n22046;
  assign n22048 = n22047 ^ n19130;
  assign n22049 = ~n21630 & ~n22048;
  assign n22042 = n19531 ^ n19137;
  assign n22043 = n22042 ^ n19517;
  assign n22044 = ~n19298 & n22043;
  assign n22045 = n22044 ^ n19517;
  assign n22050 = n22049 ^ n22045;
  assign n22051 = ~n19507 & ~n22050;
  assign n22052 = n22051 ^ n22045;
  assign n22053 = ~n21648 & ~n22052;
  assign n22054 = ~n19536 & n22053;
  assign n22055 = ~n22041 & n22054;
  assign n22056 = n19125 ^ n19117;
  assign n22057 = ~n19298 & ~n22056;
  assign n22058 = n22057 ^ n19117;
  assign n22059 = ~n19509 & n22058;
  assign n22060 = n22055 & ~n22059;
  assign n22061 = n19508 ^ n19122;
  assign n22062 = n19510 ^ n19127;
  assign n22063 = ~n19122 & ~n22062;
  assign n22064 = n22063 ^ n19127;
  assign n22065 = ~n22061 & ~n22064;
  assign n22066 = n22065 ^ n19508;
  assign n22067 = n22060 & ~n22066;
  assign n22068 = n19132 ^ n19127;
  assign n22069 = n19298 & n22068;
  assign n22070 = n22069 ^ n19127;
  assign n22071 = ~n19509 & n22070;
  assign n22072 = n22067 & ~n22071;
  assign n22073 = ~n21653 & n22072;
  assign n22074 = n22073 ^ n17236;
  assign n22075 = n22074 ^ x787;
  assign n22076 = ~n22039 & ~n22075;
  assign n22079 = n20936 & ~n20955;
  assign n22080 = n20915 & n20943;
  assign n22081 = n21579 ^ n20957;
  assign n22082 = n20916 & ~n22081;
  assign n22083 = n20917 & ~n22082;
  assign n22084 = n22083 ^ n20916;
  assign n22086 = n20959 ^ n20928;
  assign n22085 = n20927 ^ n20910;
  assign n22087 = n22086 ^ n22085;
  assign n22088 = n22083 & ~n22087;
  assign n22089 = n22088 ^ n22085;
  assign n22090 = ~n22084 & n22089;
  assign n22091 = n22090 ^ n20916;
  assign n22093 = n21584 ^ n20943;
  assign n22094 = n22093 ^ n21328;
  assign n22092 = n21335 ^ n20950;
  assign n22095 = n22094 ^ n22092;
  assign n22096 = ~n20915 & ~n22095;
  assign n22097 = n22096 ^ n22092;
  assign n22098 = n20914 & ~n22097;
  assign n22099 = ~n22091 & ~n22098;
  assign n22100 = ~n20978 & n22099;
  assign n22101 = ~n20975 & n22100;
  assign n22102 = ~n22080 & n22101;
  assign n22103 = ~n22079 & n22102;
  assign n22104 = n20914 & n21593;
  assign n22105 = n22104 ^ n20949;
  assign n22106 = n20915 & n22105;
  assign n22107 = n22103 & ~n22106;
  assign n22108 = ~n21357 & n22107;
  assign n22109 = n22108 ^ n17692;
  assign n22110 = n22109 ^ x786;
  assign n22111 = ~n20505 & n21532;
  assign n22112 = n20409 & n20464;
  assign n22113 = n20465 & ~n20487;
  assign n22119 = n20499 ^ n20474;
  assign n22114 = n20492 ^ n20474;
  assign n22115 = n22114 ^ n20494;
  assign n22116 = n22115 ^ n20404;
  assign n22117 = n20461 & ~n22116;
  assign n22118 = n22117 ^ n22115;
  assign n22120 = n22119 ^ n22118;
  assign n22121 = n22120 ^ n22118;
  assign n22122 = ~n20461 & ~n22121;
  assign n22123 = n22122 ^ n22118;
  assign n22124 = ~n20505 & n22123;
  assign n22125 = n22124 ^ n22118;
  assign n22126 = ~n21539 & ~n22125;
  assign n22127 = ~n22113 & n22126;
  assign n22128 = ~n22112 & n22127;
  assign n22130 = n20411 & ~n20425;
  assign n22129 = n20415 & n20505;
  assign n22131 = n22130 ^ n22129;
  assign n22132 = n22128 & ~n22131;
  assign n22133 = ~n21221 & n22132;
  assign n22134 = ~n22111 & n22133;
  assign n22135 = n22134 ^ n16799;
  assign n22136 = n22135 ^ x788;
  assign n22139 = ~n22110 & n22136;
  assign n22140 = n22139 ^ n22136;
  assign n22145 = n22076 & n22140;
  assign n22146 = n22145 ^ n22140;
  assign n22077 = n22076 ^ n22075;
  assign n22143 = ~n22077 & n22140;
  assign n22141 = n22076 ^ n22039;
  assign n22142 = n22140 & ~n22141;
  assign n22144 = n22143 ^ n22142;
  assign n22147 = n22146 ^ n22144;
  assign n22078 = n22077 ^ n22039;
  assign n22137 = n22136 ^ n22110;
  assign n22138 = ~n22078 & n22137;
  assign n22148 = n22147 ^ n22138;
  assign n22149 = n22148 ^ n22078;
  assign n22150 = n22149 ^ n22147;
  assign n22151 = n22150 ^ n22143;
  assign n22152 = n21511 ^ x784;
  assign n22153 = ~n20161 & n20196;
  assign n22154 = n22153 ^ n20181;
  assign n22155 = ~n20231 & n22154;
  assign n22156 = n22155 ^ n20181;
  assign n22168 = n20231 & n20249;
  assign n22162 = n20282 ^ n20157;
  assign n22163 = n22162 ^ n21827;
  assign n22160 = n20079 ^ n20046;
  assign n22161 = n22160 ^ n20149;
  assign n22164 = n22163 ^ n22161;
  assign n22158 = n20166 ^ n20159;
  assign n22157 = n20181 ^ n20156;
  assign n22159 = n22158 ^ n22157;
  assign n22165 = n22164 ^ n22159;
  assign n22166 = n20231 & n22165;
  assign n22167 = n22166 ^ n22159;
  assign n22169 = n22168 ^ n22167;
  assign n22170 = n20196 & ~n22169;
  assign n22171 = n22170 ^ n22167;
  assign n22172 = ~n22156 & n22171;
  assign n22173 = ~n20244 & n22172;
  assign n22174 = ~n21569 & n22173;
  assign n22175 = ~n20239 & n22174;
  assign n22176 = ~n20235 & n22175;
  assign n22177 = ~n21575 & n22176;
  assign n22178 = n22177 ^ n18063;
  assign n22179 = n22178 ^ x789;
  assign n22180 = n22152 & ~n22179;
  assign n22181 = n22180 ^ n22179;
  assign n22182 = n22181 ^ n22152;
  assign n22183 = ~n22151 & n22182;
  assign n22206 = n22145 ^ n22076;
  assign n22184 = n22140 ^ n22110;
  assign n22204 = n22076 & n22184;
  assign n22203 = n22076 & n22139;
  assign n22205 = n22204 ^ n22203;
  assign n22207 = n22206 ^ n22205;
  assign n22199 = n22146 ^ n22136;
  assign n22195 = n22110 ^ n22075;
  assign n22196 = n22039 & n22195;
  assign n22197 = n22196 ^ n22075;
  assign n22198 = n22136 & ~n22197;
  assign n22200 = n22199 ^ n22198;
  assign n22189 = n22136 ^ n22039;
  assign n22190 = n22189 ^ n22110;
  assign n22191 = ~n22075 & ~n22136;
  assign n22192 = n22191 ^ n22110;
  assign n22193 = n22190 & n22192;
  assign n22185 = n22184 ^ n22136;
  assign n22186 = ~n22077 & ~n22185;
  assign n22187 = n22186 ^ n22142;
  assign n22188 = n22187 ^ n22146;
  assign n22194 = n22193 ^ n22188;
  assign n22201 = n22200 ^ n22194;
  assign n22202 = n22201 ^ n22142;
  assign n22208 = n22207 ^ n22202;
  assign n22209 = n22208 ^ n22193;
  assign n22210 = n22180 ^ n22152;
  assign n22211 = ~n22209 & ~n22210;
  assign n22212 = n22211 ^ n22193;
  assign n22213 = n22179 & n22212;
  assign n22214 = n22213 ^ n22182;
  assign n22215 = ~n22183 & ~n22214;
  assign n22227 = n22075 ^ n22039;
  assign n22228 = n22227 ^ n22198;
  assign n22225 = n22202 ^ n22141;
  assign n22218 = ~n22077 & n22139;
  assign n22219 = n22218 ^ n22143;
  assign n22220 = n22219 ^ n22149;
  assign n22221 = n22220 ^ n22039;
  assign n22217 = n22186 ^ n22148;
  assign n22222 = n22221 ^ n22217;
  assign n22216 = n22143 ^ n22138;
  assign n22223 = n22222 ^ n22216;
  assign n22224 = n22223 ^ n22142;
  assign n22226 = n22225 ^ n22224;
  assign n22229 = n22228 ^ n22226;
  assign n22230 = n22152 & ~n22229;
  assign n22231 = n22230 ^ n22226;
  assign n22232 = ~n22179 & n22231;
  assign n22233 = n22215 & ~n22232;
  assign n22234 = n22152 & n22203;
  assign n22235 = n22234 ^ n22200;
  assign n22236 = n22179 & n22235;
  assign n22237 = n22236 ^ n22200;
  assign n22238 = n22233 & ~n22237;
  assign n22239 = n22152 & n22204;
  assign n22240 = n22239 ^ n22203;
  assign n22241 = n22179 & n22240;
  assign n22242 = n22241 ^ n22203;
  assign n22243 = n22238 & ~n22242;
  assign n22244 = n22225 ^ n22145;
  assign n22245 = n22244 ^ n22222;
  assign n22246 = n22152 & n22245;
  assign n22247 = n22246 ^ n22222;
  assign n22248 = n22179 & ~n22247;
  assign n22249 = n22243 & ~n22248;
  assign n22250 = n22249 ^ n20396;
  assign n22251 = ~n22179 & ~n22222;
  assign n22252 = n22141 ^ n22140;
  assign n22253 = ~n22181 & ~n22252;
  assign n22254 = ~n22251 & ~n22253;
  assign n22255 = n22179 ^ n22152;
  assign n22257 = n22223 ^ n22194;
  assign n22258 = n22257 ^ n22203;
  assign n22256 = n22149 ^ n22138;
  assign n22259 = n22258 ^ n22256;
  assign n22260 = n22179 & n22259;
  assign n22261 = n22260 ^ n22256;
  assign n22262 = n22255 & ~n22261;
  assign n22263 = n22254 & ~n22262;
  assign n22264 = n22218 ^ n22150;
  assign n22265 = n22210 & ~n22264;
  assign n22266 = n22152 ^ n22142;
  assign n22269 = n22205 ^ n22186;
  assign n22267 = n22207 ^ n22145;
  assign n22268 = n22267 ^ n22194;
  assign n22270 = n22269 ^ n22268;
  assign n22271 = ~n22179 & n22270;
  assign n22272 = n22271 ^ n22268;
  assign n22273 = n22272 ^ n22142;
  assign n22274 = ~n22266 & n22273;
  assign n22275 = n22274 ^ n22271;
  assign n22276 = n22275 ^ n22268;
  assign n22277 = n22276 ^ n22152;
  assign n22278 = ~n22142 & ~n22277;
  assign n22279 = n22278 ^ n22142;
  assign n22280 = n22279 ^ n22152;
  assign n22281 = ~n22265 & n22280;
  assign n22282 = n22263 & n22281;
  assign n22283 = ~n22179 & n22187;
  assign n22284 = n22283 ^ n22142;
  assign n22285 = ~n22152 & n22284;
  assign n22286 = n22282 & ~n22285;
  assign n22287 = n22225 ^ n22186;
  assign n22288 = n22152 & ~n22287;
  assign n22289 = n22288 ^ n22225;
  assign n22290 = n22179 & ~n22289;
  assign n22291 = n22286 & ~n22290;
  assign n22292 = n22291 ^ n20078;
  assign n22293 = n19966 & n19997;
  assign n22294 = ~n19949 & n19953;
  assign n22295 = n21419 ^ n19962;
  assign n22296 = ~n19803 & n22295;
  assign n22297 = ~n22294 & ~n22296;
  assign n22298 = ~n22293 & n22297;
  assign n22299 = n21880 ^ n19996;
  assign n22300 = n22299 ^ n19956;
  assign n22301 = n19803 & ~n22300;
  assign n22302 = n22301 ^ n19956;
  assign n22303 = n19947 & ~n22302;
  assign n22304 = n22298 & ~n22303;
  assign n22305 = ~n20021 & n22304;
  assign n22306 = ~n20008 & n22305;
  assign n22307 = ~n21873 & n22306;
  assign n22308 = ~n21423 & n22307;
  assign n22309 = ~n19950 & n22308;
  assign n22310 = ~n20027 & n22309;
  assign n22311 = n22310 ^ n18734;
  assign n22312 = n21391 ^ n21379;
  assign n22313 = n22312 ^ n21372;
  assign n22314 = n21361 & n22313;
  assign n22315 = ~n21394 & ~n21459;
  assign n22316 = n22315 ^ n21392;
  assign n22317 = ~n21362 & n22316;
  assign n22318 = n22317 ^ n21392;
  assign n22319 = ~n22314 & ~n22318;
  assign n22320 = n21391 ^ n21305;
  assign n22321 = n21391 ^ n21073;
  assign n22322 = n21360 & n22321;
  assign n22323 = n22322 ^ n21073;
  assign n22324 = n22320 & ~n22323;
  assign n22325 = n22324 ^ n21305;
  assign n22326 = ~n21461 & ~n22325;
  assign n22327 = ~n21303 & n22326;
  assign n22328 = ~n21360 & ~n22327;
  assign n22329 = n22319 & ~n22328;
  assign n22330 = ~n21486 & n22329;
  assign n22331 = ~n21413 & n22330;
  assign n22332 = n22331 ^ n20879;
  assign n22333 = n19509 & n21623;
  assign n22339 = n21627 ^ n19141;
  assign n22340 = n19507 & ~n22339;
  assign n22341 = n22340 ^ n21627;
  assign n22335 = n19531 ^ n19119;
  assign n22334 = n21619 ^ n19116;
  assign n22336 = n22335 ^ n22334;
  assign n22337 = n19507 & n22336;
  assign n22338 = n22337 ^ n22334;
  assign n22342 = n22341 ^ n22338;
  assign n22343 = ~n19298 & n22342;
  assign n22344 = n22343 ^ n22338;
  assign n22345 = ~n22333 & ~n22344;
  assign n22346 = n19535 & n22345;
  assign n22347 = ~n19507 & n22346;
  assign n22348 = n22347 ^ n22345;
  assign n22349 = ~n21643 & n22348;
  assign n22350 = ~n22071 & n22349;
  assign n22351 = ~n19544 & n22350;
  assign n22352 = ~n21653 & n22351;
  assign n22353 = ~n19549 & n22352;
  assign n22354 = n22353 ^ n18554;
  assign n22355 = n20292 & ~n21002;
  assign n22363 = n21021 ^ n20999;
  assign n22358 = n21021 ^ n21011;
  assign n22359 = n22358 ^ n20993;
  assign n22356 = n21035 ^ n21006;
  assign n22357 = n22356 ^ n21007;
  assign n22360 = n22359 ^ n22357;
  assign n22361 = ~n20291 & n22360;
  assign n22362 = n22361 ^ n22357;
  assign n22364 = n22363 ^ n22362;
  assign n22365 = n22364 ^ n22362;
  assign n22366 = n20291 & n22365;
  assign n22367 = n22366 ^ n22362;
  assign n22368 = n21034 & n22367;
  assign n22369 = n22368 ^ n22362;
  assign n22371 = n20992 & ~n21034;
  assign n22370 = ~n20291 & ~n21015;
  assign n22372 = n22371 ^ n22370;
  assign n22373 = ~n22369 & ~n22372;
  assign n22374 = n20291 & ~n21019;
  assign n22375 = n22374 ^ n21009;
  assign n22376 = n20030 & ~n22375;
  assign n22377 = n22373 & ~n22376;
  assign n22378 = ~n22355 & n22377;
  assign n22379 = ~n21051 & n22378;
  assign n22380 = ~n21056 & n22379;
  assign n22381 = n21066 ^ n20996;
  assign n22382 = n20291 & n22381;
  assign n22383 = n22382 ^ n20996;
  assign n22384 = n21034 & n22383;
  assign n22385 = n22380 & ~n22384;
  assign n22386 = ~n21010 & n22385;
  assign n22387 = ~n21070 & n22386;
  assign n22388 = n22387 ^ n20809;
  assign n22389 = n21074 & ~n21155;
  assign n22390 = n21182 ^ n21128;
  assign n22391 = n21159 & n22390;
  assign n22392 = n21757 ^ n21129;
  assign n22393 = n22392 ^ n21748;
  assign n22394 = n22393 ^ n21074;
  assign n22395 = n21112 ^ n21109;
  assign n22396 = n22395 ^ n21143;
  assign n22397 = n22396 ^ n21098;
  assign n22398 = n22397 ^ n22393;
  assign n22399 = n22397 ^ n21075;
  assign n22400 = n22397 & n22399;
  assign n22401 = n22400 ^ n22397;
  assign n22402 = n22398 & n22401;
  assign n22403 = n22402 ^ n22400;
  assign n22404 = n22403 ^ n22397;
  assign n22405 = n22404 ^ n21075;
  assign n22406 = n22394 & n22405;
  assign n22407 = n22406 ^ n22393;
  assign n22408 = ~n22391 & n22407;
  assign n22409 = n21139 ^ n21123;
  assign n22410 = n22409 ^ n21113;
  assign n22411 = n22410 ^ n21146;
  assign n22412 = n22411 ^ n21146;
  assign n22413 = n21074 & ~n22412;
  assign n22414 = n22413 ^ n21146;
  assign n22415 = n21075 & n22414;
  assign n22416 = n22415 ^ n21146;
  assign n22417 = n22408 & ~n22416;
  assign n22418 = ~n21169 & n22417;
  assign n22419 = ~n22389 & n22418;
  assign n22420 = ~n21492 & n22419;
  assign n22421 = ~n21766 & n22420;
  assign n22422 = ~n21771 & n22421;
  assign n22423 = ~n21491 & n22422;
  assign n22424 = ~n21186 & n22423;
  assign n22425 = n22424 ^ n18942;
  assign n22426 = n21660 & n21714;
  assign n22427 = n21688 ^ n21681;
  assign n22428 = n22427 ^ n21667;
  assign n22429 = n22428 ^ n21676;
  assign n22430 = ~n21707 & ~n22429;
  assign n22431 = n21690 & n21706;
  assign n22433 = n21710 ^ n21698;
  assign n22434 = n22433 ^ n21685;
  assign n22432 = n22427 ^ n21709;
  assign n22435 = n22434 ^ n22432;
  assign n22436 = n22435 ^ n22432;
  assign n22437 = n21543 & n22436;
  assign n22438 = n22437 ^ n22432;
  assign n22439 = ~n21545 & ~n22438;
  assign n22440 = n22439 ^ n22432;
  assign n22441 = ~n22431 & n22440;
  assign n22442 = ~n22430 & n22441;
  assign n22443 = ~n22426 & n22442;
  assign n22444 = ~n21736 & n22443;
  assign n22445 = ~n21815 & n22444;
  assign n22446 = n21788 & n22445;
  assign n22447 = ~n21728 & n22446;
  assign n22448 = n22447 ^ n20365;
  assign n22449 = n21310 & n21362;
  assign n22450 = n21461 ^ n21367;
  assign n22451 = n21361 & n22450;
  assign n22455 = n21398 ^ n21307;
  assign n22454 = n21393 ^ n21368;
  assign n22456 = n22455 ^ n22454;
  assign n22457 = ~n21360 & n22456;
  assign n22458 = n22457 ^ n22454;
  assign n22452 = n21314 & ~n21360;
  assign n22453 = n22452 ^ n21310;
  assign n22459 = n22458 ^ n22453;
  assign n22460 = n21073 & ~n22459;
  assign n22461 = n22460 ^ n22458;
  assign n22462 = ~n22451 & n22461;
  assign n22463 = ~n22449 & n22462;
  assign n22465 = n21394 ^ n21316;
  assign n22464 = n21378 ^ n21368;
  assign n22466 = n22465 ^ n22464;
  assign n22467 = n21073 & ~n22466;
  assign n22468 = n22467 ^ n22464;
  assign n22469 = ~n21360 & n22468;
  assign n22470 = n22463 & ~n22469;
  assign n22471 = ~n21414 & n22470;
  assign n22472 = n22471 ^ n20120;
  assign n22473 = n21868 & n22017;
  assign n22474 = n22001 ^ n21978;
  assign n22475 = n22474 ^ n21931;
  assign n22476 = n21869 & n22475;
  assign n22477 = ~n21867 & n21953;
  assign n22478 = n22477 ^ n21958;
  assign n22479 = n21987 & n22478;
  assign n22480 = n22479 ^ n21958;
  assign n22481 = ~n22476 & ~n22480;
  assign n22482 = ~n21866 & n22001;
  assign n22483 = n22482 ^ n21975;
  assign n22484 = n21867 & n22483;
  assign n22485 = n22484 ^ n21975;
  assign n22486 = n22481 & ~n22485;
  assign n22487 = ~n21972 & n22486;
  assign n22488 = ~n22011 & n22487;
  assign n22492 = ~n21866 & n21931;
  assign n22489 = n21960 ^ n21936;
  assign n22490 = ~n21866 & n22489;
  assign n22491 = n22490 ^ n21960;
  assign n22493 = n22492 ^ n22491;
  assign n22494 = ~n21867 & n22493;
  assign n22495 = n22494 ^ n22491;
  assign n22496 = n22488 & ~n22495;
  assign n22499 = n21867 & n21945;
  assign n22497 = n21867 & ~n21957;
  assign n22498 = n22497 ^ n21948;
  assign n22500 = n22499 ^ n22498;
  assign n22501 = ~n21987 & ~n22500;
  assign n22502 = n22501 ^ n22498;
  assign n22503 = n22496 & n22502;
  assign n22504 = n21976 ^ n21934;
  assign n22505 = n21867 & n22504;
  assign n22506 = n22505 ^ n21934;
  assign n22507 = n21987 & n22506;
  assign n22508 = n22503 & ~n22507;
  assign n22509 = ~n22473 & n22508;
  assign n22510 = n21966 & n22509;
  assign n22511 = n22510 ^ n20680;
  assign n22512 = n22135 ^ x790;
  assign n22513 = n21296 ^ x795;
  assign n22514 = ~n22512 & ~n22513;
  assign n22515 = n22514 ^ n22512;
  assign n22516 = n22515 ^ n22513;
  assign n22517 = n22178 ^ x791;
  assign n22518 = n21774 ^ x793;
  assign n22520 = n22311 ^ x792;
  assign n22521 = n22518 & n22520;
  assign n22522 = ~n22517 & n22521;
  assign n22523 = n22522 ^ n22517;
  assign n22519 = ~n22517 & ~n22518;
  assign n22524 = n22523 ^ n22519;
  assign n22525 = n19551 ^ x794;
  assign n22526 = ~n22524 & ~n22525;
  assign n22527 = n22526 ^ n22524;
  assign n22528 = ~n22516 & ~n22527;
  assign n22534 = n22519 ^ n22518;
  assign n22530 = n22517 & n22525;
  assign n22533 = ~n22518 & n22530;
  assign n22535 = n22534 ^ n22533;
  assign n22536 = ~n22520 & ~n22535;
  assign n22537 = n22536 ^ n22535;
  assign n22529 = n22521 ^ n22518;
  assign n22531 = n22530 ^ n22517;
  assign n22532 = n22529 & n22531;
  assign n22538 = n22537 ^ n22532;
  assign n22539 = ~n22515 & ~n22538;
  assign n22540 = ~n22515 & ~n22524;
  assign n22554 = n22522 & n22525;
  assign n22555 = n22554 ^ n22522;
  assign n22550 = n22519 & ~n22520;
  assign n22551 = ~n22525 & n22550;
  assign n22552 = n22551 ^ n22550;
  assign n22547 = n22525 ^ n22520;
  assign n22548 = n22519 & ~n22547;
  assign n22549 = n22548 ^ n22519;
  assign n22553 = n22552 ^ n22549;
  assign n22556 = n22555 ^ n22553;
  assign n22543 = n22522 ^ n22521;
  assign n22542 = n22521 & n22530;
  assign n22544 = n22543 ^ n22542;
  assign n22541 = n22529 & n22530;
  assign n22545 = n22544 ^ n22541;
  assign n22546 = n22545 ^ n22536;
  assign n22557 = n22556 ^ n22546;
  assign n22558 = n22557 ^ n22546;
  assign n22559 = n22515 & n22558;
  assign n22560 = n22559 ^ n22546;
  assign n22561 = n22514 ^ n22513;
  assign n22562 = n22560 & n22561;
  assign n22563 = n22562 ^ n22546;
  assign n22564 = ~n22540 & ~n22563;
  assign n22565 = n22513 ^ n22512;
  assign n22566 = ~n22520 & n22533;
  assign n22567 = n22566 ^ n22533;
  assign n22574 = n22567 ^ n22548;
  assign n22575 = ~n22513 & n22574;
  assign n22576 = n22575 ^ n22548;
  assign n22571 = n22544 ^ n22537;
  assign n22572 = n22513 & ~n22571;
  assign n22568 = n22567 ^ n22532;
  assign n22569 = n22568 ^ n22566;
  assign n22570 = n22569 ^ n22544;
  assign n22573 = n22572 ^ n22570;
  assign n22577 = n22576 ^ n22573;
  assign n22578 = n22565 & n22577;
  assign n22579 = n22578 ^ n22573;
  assign n22580 = n22564 & ~n22579;
  assign n22581 = ~n22539 & n22580;
  assign n22582 = ~n22528 & n22581;
  assign n22583 = n22554 ^ n22526;
  assign n22584 = n22583 ^ n22552;
  assign n22585 = n22512 & n22584;
  assign n22586 = n22585 ^ n22552;
  assign n22587 = ~n22513 & n22586;
  assign n22588 = n22582 & ~n22587;
  assign n22592 = ~n22512 & n22542;
  assign n22589 = n22554 ^ n22548;
  assign n22590 = n22512 & n22589;
  assign n22591 = n22590 ^ n22554;
  assign n22593 = n22592 ^ n22591;
  assign n22594 = n22513 & n22593;
  assign n22595 = n22594 ^ n22591;
  assign n22596 = n22588 & ~n22595;
  assign n22597 = n22566 ^ n22554;
  assign n22598 = n22512 & n22597;
  assign n22599 = n22598 ^ n22566;
  assign n22600 = n22513 & n22599;
  assign n22601 = n22596 & ~n22600;
  assign n22602 = n22601 ^ n19802;
  assign n22603 = n21936 ^ n21869;
  assign n22604 = n21971 ^ n21952;
  assign n22605 = n21936 & n22604;
  assign n22606 = n22605 ^ n21952;
  assign n22607 = n22603 & ~n22606;
  assign n22608 = n22607 ^ n21869;
  assign n22610 = n21951 ^ n21939;
  assign n22609 = n21976 ^ n21967;
  assign n22611 = n22610 ^ n22609;
  assign n22612 = n21867 & n22611;
  assign n22613 = n22612 ^ n22609;
  assign n22614 = n21987 & n22613;
  assign n22615 = ~n22608 & ~n22614;
  assign n22617 = ~n21971 & n22474;
  assign n22616 = ~n21867 & n21956;
  assign n22618 = n22617 ^ n22616;
  assign n22619 = n22615 & ~n22618;
  assign n22620 = ~n22005 & n22619;
  assign n22621 = ~n22016 & n22620;
  assign n22622 = ~n22495 & n22621;
  assign n22623 = n21978 ^ n21939;
  assign n22624 = n22623 ^ n21969;
  assign n22625 = n21866 & n22624;
  assign n22626 = n22625 ^ n21969;
  assign n22627 = n21867 & n22626;
  assign n22628 = n22622 & ~n22627;
  assign n22629 = ~n22473 & n22628;
  assign n22630 = n21966 & n22629;
  assign n22631 = n22630 ^ n19506;
  assign n22632 = n20853 ^ x814;
  assign n22633 = n21656 ^ x819;
  assign n22636 = n21458 ^ x818;
  assign n22634 = n20290 ^ x815;
  assign n22641 = n22038 ^ x817;
  assign n22642 = ~n22634 & ~n22641;
  assign n22650 = n22642 ^ n22641;
  assign n22653 = n22636 & ~n22650;
  assign n22654 = n22653 ^ n22650;
  assign n22635 = n22425 ^ x816;
  assign n22640 = ~n22635 & ~n22636;
  assign n22651 = n22640 ^ n22636;
  assign n22652 = ~n22650 & ~n22651;
  assign n22655 = n22654 ^ n22652;
  assign n22643 = n22642 ^ n22634;
  assign n22644 = n22643 ^ n22641;
  assign n22646 = n22636 & ~n22644;
  assign n22647 = ~n22635 & n22646;
  assign n22648 = n22647 ^ n22646;
  assign n22645 = n22640 & ~n22644;
  assign n22649 = n22648 ^ n22645;
  assign n22656 = n22655 ^ n22649;
  assign n22666 = ~n22633 & ~n22656;
  assign n22658 = n22646 ^ n22644;
  assign n22659 = n22658 ^ n22645;
  assign n22637 = n22636 ^ n22635;
  assign n22638 = n22634 & n22637;
  assign n22639 = n22638 ^ n22634;
  assign n22657 = n22656 ^ n22639;
  assign n22660 = n22659 ^ n22657;
  assign n22661 = n22660 ^ n22655;
  assign n22662 = n22661 ^ n22645;
  assign n22663 = n22662 ^ n22638;
  assign n22664 = n22633 & ~n22663;
  assign n22665 = n22664 ^ n22638;
  assign n22667 = n22666 ^ n22665;
  assign n22668 = ~n22632 & n22667;
  assign n22669 = n22668 ^ n22665;
  assign n22670 = n22633 ^ n22632;
  assign n22677 = n22645 ^ n22640;
  assign n22676 = n22640 & ~n22643;
  assign n22678 = n22677 ^ n22676;
  assign n22679 = n22678 ^ n22655;
  assign n22674 = n22636 & n22642;
  assign n22675 = n22674 ^ n22642;
  assign n22680 = n22679 ^ n22675;
  assign n22671 = n22636 & ~n22643;
  assign n22672 = ~n22635 & n22671;
  assign n22673 = n22672 ^ n22671;
  assign n22681 = n22680 ^ n22673;
  assign n22682 = ~n22670 & ~n22681;
  assign n22683 = ~n22669 & ~n22682;
  assign n22687 = ~n22635 & n22674;
  assign n22688 = n22687 ^ n22674;
  assign n22684 = n22671 ^ n22643;
  assign n22685 = n22684 ^ n22676;
  assign n22686 = n22685 ^ n22648;
  assign n22689 = n22688 ^ n22686;
  assign n22690 = n22689 ^ n22688;
  assign n22691 = ~n22632 & ~n22690;
  assign n22692 = n22691 ^ n22688;
  assign n22693 = n22633 & n22692;
  assign n22694 = n22693 ^ n22688;
  assign n22695 = n22683 & ~n22694;
  assign n22696 = n22657 ^ n22652;
  assign n22697 = n22696 ^ n22653;
  assign n22698 = n22697 ^ n22681;
  assign n22699 = ~n22633 & n22698;
  assign n22700 = n22699 ^ n22697;
  assign n22701 = n22670 & ~n22700;
  assign n22702 = n22695 & ~n22701;
  assign n22703 = n22679 ^ n22672;
  assign n22704 = n22703 ^ n22676;
  assign n22705 = n22704 ^ n22676;
  assign n22706 = n22633 & ~n22705;
  assign n22707 = n22706 ^ n22676;
  assign n22708 = n22670 & n22707;
  assign n22709 = n22708 ^ n22676;
  assign n22710 = n22702 & ~n22709;
  assign n22711 = n22679 ^ n22660;
  assign n22712 = n22633 & ~n22711;
  assign n22713 = n22712 ^ n22679;
  assign n22714 = n22713 ^ n22687;
  assign n22715 = n22670 & ~n22714;
  assign n22716 = n22715 ^ n22687;
  assign n22717 = n22710 & ~n22716;
  assign n22718 = n22717 ^ n20148;
  assign n22719 = ~n22633 & ~n22659;
  assign n22720 = n22719 ^ n22659;
  assign n22721 = n22720 ^ n22674;
  assign n22722 = n22670 & ~n22721;
  assign n22723 = n22722 ^ n22674;
  assign n22724 = n22685 ^ n22672;
  assign n22725 = n22632 & ~n22724;
  assign n22726 = n22725 ^ n22685;
  assign n22727 = ~n22633 & ~n22726;
  assign n22728 = ~n22723 & ~n22727;
  assign n22729 = n22632 & ~n22633;
  assign n22730 = n22729 ^ n22632;
  assign n22731 = n22730 ^ n22633;
  assign n22732 = n22731 ^ n22632;
  assign n22733 = n22660 & ~n22732;
  assign n22734 = n22647 ^ n22645;
  assign n22735 = n22734 ^ n22730;
  assign n22736 = n22732 ^ n22696;
  assign n22737 = ~n22734 & ~n22736;
  assign n22738 = n22737 ^ n22732;
  assign n22739 = n22735 & ~n22738;
  assign n22740 = n22739 ^ n22730;
  assign n22741 = ~n22733 & ~n22740;
  assign n22743 = n22681 ^ n22676;
  assign n22744 = n22743 ^ n22672;
  assign n22742 = n22697 ^ n22649;
  assign n22745 = n22744 ^ n22742;
  assign n22746 = n22633 & n22745;
  assign n22747 = n22746 ^ n22742;
  assign n22748 = n22670 & ~n22747;
  assign n22749 = n22741 & ~n22748;
  assign n22750 = n22677 & n22730;
  assign n22751 = n22750 ^ n22655;
  assign n22752 = n22749 & n22751;
  assign n22753 = n22728 & n22752;
  assign n22754 = ~n22701 & n22753;
  assign n22755 = n22754 ^ n20557;
  assign n22761 = n21712 ^ n21686;
  assign n22757 = n21775 ^ n21661;
  assign n22756 = n21709 ^ n21675;
  assign n22758 = n22757 ^ n22756;
  assign n22759 = ~n21543 & ~n22758;
  assign n22760 = n22759 ^ n22756;
  assign n22762 = n22761 ^ n22760;
  assign n22763 = n22762 ^ n22760;
  assign n22764 = ~n21543 & ~n22763;
  assign n22765 = n22764 ^ n22760;
  assign n22766 = n21544 & n22765;
  assign n22767 = n22766 ^ n22760;
  assign n22768 = n21729 ^ n21699;
  assign n22769 = n21707 ^ n21695;
  assign n22770 = n21699 & n22769;
  assign n22771 = n22770 ^ n21695;
  assign n22772 = n22768 & ~n22771;
  assign n22773 = n22772 ^ n21729;
  assign n22774 = ~n22767 & ~n22773;
  assign n22775 = ~n21722 & n22774;
  assign n22776 = ~n21731 & n22775;
  assign n22777 = n21783 & n22776;
  assign n22778 = n22777 ^ n19731;
  assign n22779 = n21188 ^ x802;
  assign n22784 = n21359 ^ x803;
  assign n22781 = n21853 ^ x805;
  assign n22782 = n20029 ^ x806;
  assign n22783 = ~n22781 & ~n22782;
  assign n22803 = n22783 ^ n22781;
  assign n22785 = n22354 ^ x804;
  assign n22804 = n22803 ^ n22785;
  assign n22791 = n22782 ^ n22781;
  assign n22805 = n22804 ^ n22791;
  assign n22838 = ~n22784 & n22805;
  assign n22839 = n22838 ^ n22791;
  assign n22780 = n20751 ^ x807;
  assign n22843 = n22839 ^ n22780;
  assign n22786 = n22784 & n22785;
  assign n22798 = n22786 ^ n22784;
  assign n22799 = n22798 ^ n22785;
  assign n22800 = n22799 ^ n22784;
  assign n22801 = n22783 ^ n22782;
  assign n22802 = n22800 & n22801;
  assign n22806 = n22805 ^ n22802;
  assign n22826 = n22806 ^ n22785;
  assign n22820 = ~n22800 & n22803;
  assign n22821 = n22820 ^ n22801;
  assign n22808 = n22784 ^ n22781;
  assign n22809 = n22808 ^ n22785;
  assign n22810 = ~n22782 & n22809;
  assign n22818 = n22785 & n22810;
  assign n22790 = n22785 ^ n22781;
  assign n22792 = n22791 ^ n22785;
  assign n22793 = n22791 ^ n22784;
  assign n22794 = n22792 & ~n22793;
  assign n22795 = n22794 ^ n22791;
  assign n22796 = ~n22790 & n22795;
  assign n22815 = n22796 ^ n22791;
  assign n22819 = n22818 ^ n22815;
  assign n22822 = n22821 ^ n22819;
  assign n22811 = n22810 ^ n22785;
  assign n22823 = ~n22791 & ~n22811;
  assign n22824 = ~n22822 & ~n22823;
  assign n22788 = n22782 & n22786;
  assign n22825 = n22824 ^ n22788;
  assign n22827 = n22826 ^ n22825;
  assign n22812 = n22784 ^ n22782;
  assign n22817 = n22812 ^ n22785;
  assign n22828 = n22827 ^ n22817;
  assign n22840 = n22839 ^ n22828;
  assign n22841 = n22780 & ~n22840;
  assign n22842 = n22841 ^ n22828;
  assign n22844 = n22843 ^ n22842;
  assign n22845 = n22844 ^ n22828;
  assign n22829 = n22828 ^ n22791;
  assign n22813 = n22811 & n22812;
  assign n22814 = n22813 ^ n22809;
  assign n22816 = n22815 ^ n22814;
  assign n22830 = n22829 ^ n22816;
  assign n22831 = n22830 ^ n22808;
  assign n22787 = ~n22783 & n22786;
  assign n22789 = n22788 ^ n22787;
  assign n22797 = n22796 ^ n22789;
  assign n22807 = n22806 ^ n22797;
  assign n22832 = n22831 ^ n22807;
  assign n22833 = n22780 & ~n22832;
  assign n22834 = n22833 ^ n22807;
  assign n22835 = n22834 ^ n22780;
  assign n22836 = n22835 ^ n22831;
  assign n22837 = n22836 ^ n22807;
  assign n22846 = n22845 ^ n22837;
  assign n22847 = n22779 & ~n22846;
  assign n22848 = n22847 ^ n22837;
  assign n22849 = n22848 ^ n18622;
  assign n22850 = n22565 & n22576;
  assign n22852 = n22553 ^ n22527;
  assign n22851 = n22552 ^ n22526;
  assign n22853 = n22852 ^ n22851;
  assign n22854 = ~n22516 & ~n22853;
  assign n22855 = n22542 ^ n22536;
  assign n22856 = ~n22565 & n22855;
  assign n22857 = ~n22854 & ~n22856;
  assign n22861 = n22568 ^ n22545;
  assign n22858 = n22525 ^ n22518;
  assign n22859 = n22858 ^ n22512;
  assign n22860 = ~n22517 & n22859;
  assign n22862 = n22861 ^ n22860;
  assign n22863 = n22862 ^ n22860;
  assign n22864 = ~n22512 & n22863;
  assign n22865 = n22864 ^ n22860;
  assign n22866 = n22513 & n22865;
  assign n22867 = n22866 ^ n22860;
  assign n22868 = n22514 & ~n22571;
  assign n22869 = n22868 ^ n22571;
  assign n22870 = n22869 ^ n22572;
  assign n22871 = ~n22867 & n22870;
  assign n22872 = n22857 & n22871;
  assign n22880 = n22514 & n22568;
  assign n22876 = n22513 & ~n22537;
  assign n22873 = n22566 ^ n22555;
  assign n22874 = n22513 & n22873;
  assign n22875 = n22874 ^ n22566;
  assign n22877 = n22876 ^ n22875;
  assign n22878 = ~n22565 & n22877;
  assign n22879 = n22878 ^ n22875;
  assign n22881 = n22880 ^ n22879;
  assign n22882 = n22872 & ~n22881;
  assign n22883 = ~n22850 & n22882;
  assign n22884 = ~n22600 & n22883;
  assign n22885 = n22884 ^ n20230;
  assign n22886 = n20030 & n20997;
  assign n22887 = n22886 ^ n20992;
  assign n22888 = n20291 & n22887;
  assign n22889 = n22888 ^ n20992;
  assign n22890 = ~n21010 & ~n22889;
  assign n22897 = n21022 ^ n20996;
  assign n22898 = n22897 ^ n21001;
  assign n22896 = n21012 ^ n21006;
  assign n22899 = n22898 ^ n22896;
  assign n22900 = ~n20030 & ~n22899;
  assign n22901 = n22900 ^ n22896;
  assign n22902 = n22901 ^ n21009;
  assign n22903 = ~n22901 & n22902;
  assign n22892 = n21023 ^ n20999;
  assign n22891 = n21015 ^ n21007;
  assign n22893 = n22892 ^ n22891;
  assign n22894 = n20030 & ~n22893;
  assign n22895 = n22894 ^ n22891;
  assign n22904 = n22903 ^ n22895;
  assign n22905 = n20291 & n22904;
  assign n22906 = n22905 ^ n22903;
  assign n22907 = ~n21059 & n22906;
  assign n22908 = ~n21041 & n22907;
  assign n22909 = ~n21046 & n22908;
  assign n22910 = n22890 & n22909;
  assign n22911 = ~n22384 & n22910;
  assign n22912 = ~n21070 & n22911;
  assign n22913 = n22912 ^ n20619;
  assign n22914 = n22687 ^ n22680;
  assign n22915 = n22731 & ~n22914;
  assign n22916 = n22632 & n22687;
  assign n22917 = n22655 ^ n22647;
  assign n22918 = n22917 ^ n22673;
  assign n22919 = n22918 ^ n22697;
  assign n22920 = n22730 & n22919;
  assign n22921 = ~n22916 & ~n22920;
  assign n22922 = ~n22633 & ~n22743;
  assign n22923 = n22922 ^ n22685;
  assign n22924 = n22670 & ~n22923;
  assign n22925 = n22924 ^ n22685;
  assign n22926 = n22921 & n22925;
  assign n22940 = ~n22633 & ~n22917;
  assign n22941 = n22940 ^ n22719;
  assign n22938 = n22917 ^ n22660;
  assign n22939 = n22731 & ~n22938;
  assign n22942 = n22941 ^ n22939;
  assign n22928 = ~n22732 & ~n22917;
  assign n22936 = n22928 ^ n22733;
  assign n22934 = n22688 ^ n22649;
  assign n22935 = ~n22732 & n22934;
  assign n22937 = n22936 ^ n22935;
  assign n22943 = n22942 ^ n22937;
  assign n22932 = n22648 & n22729;
  assign n22927 = n22917 ^ n22732;
  assign n22929 = n22928 ^ n22927;
  assign n22930 = n22672 ^ n22652;
  assign n22931 = n22929 & n22930;
  assign n22933 = n22932 ^ n22931;
  assign n22944 = n22943 ^ n22933;
  assign n22945 = n22926 & ~n22944;
  assign n22946 = ~n22709 & n22945;
  assign n22947 = ~n22915 & n22946;
  assign n22948 = n22947 ^ n19760;
  assign n22949 = ~n22633 & n22672;
  assign n22950 = n22676 ^ n22673;
  assign n22951 = n22729 & n22950;
  assign n22952 = ~n22949 & ~n22951;
  assign n22953 = n22633 & n22645;
  assign n22954 = n22953 ^ n22680;
  assign n22955 = n22670 & ~n22954;
  assign n22956 = n22955 ^ n22680;
  assign n22957 = n22952 & n22956;
  assign n22958 = ~n22632 & n22653;
  assign n22959 = n22688 ^ n22685;
  assign n22960 = n22730 & ~n22959;
  assign n22961 = n22685 ^ n22673;
  assign n22962 = n22731 & ~n22961;
  assign n22966 = n22661 ^ n22652;
  assign n22963 = n22730 & n22929;
  assign n22964 = n22963 ^ n22649;
  assign n22965 = n22964 ^ n22733;
  assign n22967 = n22966 ^ n22965;
  assign n22968 = n22967 ^ n22965;
  assign n22969 = ~n22633 & ~n22968;
  assign n22970 = n22969 ^ n22965;
  assign n22971 = n22670 & n22970;
  assign n22972 = n22971 ^ n22965;
  assign n22973 = ~n22962 & ~n22972;
  assign n22974 = ~n22915 & n22973;
  assign n22975 = ~n22960 & n22974;
  assign n22976 = ~n22958 & n22975;
  assign n22977 = n22957 & n22976;
  assign n22978 = ~n22716 & n22977;
  assign n22979 = n22978 ^ n19103;
  assign n22980 = n21971 ^ n21967;
  assign n22983 = n21952 ^ n21935;
  assign n22981 = n21959 ^ n21927;
  assign n22982 = n22981 ^ n21941;
  assign n22984 = n22983 ^ n22982;
  assign n22985 = n22984 ^ n21869;
  assign n22986 = ~n21971 & ~n22985;
  assign n22987 = n22986 ^ n21869;
  assign n22988 = ~n22980 & ~n22987;
  assign n22989 = n22988 ^ n21967;
  assign n22990 = n22475 ^ n21961;
  assign n22991 = ~n21867 & n22990;
  assign n22992 = n22991 ^ n21961;
  assign n22993 = n21987 & n22992;
  assign n22994 = ~n22989 & ~n22993;
  assign n22995 = ~n21949 & n22994;
  assign n22996 = ~n22019 & n22995;
  assign n22997 = n22502 & n22996;
  assign n22998 = ~n22627 & n22997;
  assign n22999 = ~n22507 & n22998;
  assign n23000 = ~n22473 & n22999;
  assign n23001 = n23000 ^ n21097;
  assign n23002 = ~n22516 & n22542;
  assign n23003 = ~n22538 & ~n22561;
  assign n23014 = ~n22513 & n22522;
  assign n23005 = n22551 ^ n22527;
  assign n23006 = n23005 ^ n22555;
  assign n23004 = n22536 ^ n22526;
  assign n23007 = n23006 ^ n23004;
  assign n23008 = n23006 ^ n22513;
  assign n23009 = n22565 & n23008;
  assign n23010 = n23009 ^ n22513;
  assign n23011 = ~n23007 & n23010;
  assign n23012 = n23011 ^ n23004;
  assign n23013 = ~n22552 & ~n23012;
  assign n23015 = n23014 ^ n23013;
  assign n23016 = n22565 & ~n23015;
  assign n23017 = n23016 ^ n23013;
  assign n23018 = ~n22868 & n23017;
  assign n23019 = n22567 ^ n22541;
  assign n23020 = n23019 ^ n22569;
  assign n23021 = n23020 ^ n22569;
  assign n23022 = n22561 & n23021;
  assign n23023 = n23022 ^ n22569;
  assign n23024 = n22515 & n23023;
  assign n23025 = n23024 ^ n22569;
  assign n23026 = n23018 & ~n23025;
  assign n23027 = ~n22595 & n23026;
  assign n23028 = ~n23003 & n23027;
  assign n23029 = ~n23002 & n23028;
  assign n23030 = n22536 ^ n22515;
  assign n23031 = n22851 ^ n22561;
  assign n23032 = ~n22536 & n23031;
  assign n23033 = n23032 ^ n22561;
  assign n23034 = ~n23030 & ~n23033;
  assign n23035 = n23034 ^ n22515;
  assign n23036 = n23029 & n23035;
  assign n23037 = ~n22879 & n23036;
  assign n23038 = n23037 ^ n20582;
  assign n23045 = n22824 ^ n22787;
  assign n23046 = n23045 ^ n22819;
  assign n23047 = n22779 & ~n23046;
  assign n23048 = n23047 ^ n22819;
  assign n23040 = n22818 ^ n22798;
  assign n23039 = n22820 ^ n22802;
  assign n23041 = n23040 ^ n23039;
  assign n23042 = n23041 ^ n22814;
  assign n23043 = n22779 & ~n23042;
  assign n23044 = n23043 ^ n23041;
  assign n23049 = n23048 ^ n23044;
  assign n23050 = ~n22780 & n23049;
  assign n23051 = n23050 ^ n23048;
  assign n23052 = n23051 ^ n19563;
  assign n23053 = n22545 ^ n22532;
  assign n23054 = ~n22561 & n23053;
  assign n23068 = n22851 ^ n22555;
  assign n23069 = n23068 ^ n22519;
  assign n23070 = n22513 & n23069;
  assign n23071 = n23070 ^ n22519;
  assign n23056 = n22518 ^ n22517;
  assign n23057 = n22858 & ~n23056;
  assign n23058 = n23057 ^ n22518;
  assign n23059 = n22547 ^ n22517;
  assign n23060 = n23059 ^ n22518;
  assign n23061 = n23060 ^ n22525;
  assign n23062 = n23061 ^ n22517;
  assign n23063 = ~n23058 & ~n23062;
  assign n23064 = n23063 ^ n23059;
  assign n23055 = n22852 ^ n22583;
  assign n23065 = n23064 ^ n23055;
  assign n23066 = n22513 & n23065;
  assign n23067 = n23066 ^ n23055;
  assign n23072 = n23071 ^ n23067;
  assign n23073 = ~n22512 & ~n23072;
  assign n23074 = n23073 ^ n23071;
  assign n23075 = ~n22600 & ~n23074;
  assign n23076 = ~n23054 & n23075;
  assign n23078 = n22566 ^ n22545;
  assign n23077 = n22542 ^ n22537;
  assign n23079 = n23078 ^ n23077;
  assign n23080 = n22513 & ~n23079;
  assign n23081 = n23080 ^ n23077;
  assign n23082 = ~n22565 & ~n23081;
  assign n23083 = n23076 & ~n23082;
  assign n23084 = ~n22881 & n23083;
  assign n23085 = n23084 ^ n18856;
  assign n23086 = n22842 ^ n22834;
  assign n23087 = n22779 & ~n23086;
  assign n23088 = n23087 ^ n22834;
  assign n23089 = n23088 ^ n21104;
  assign n23090 = n22780 ^ n22779;
  assign n23093 = n23041 ^ n22825;
  assign n23094 = ~n22780 & n23093;
  assign n23095 = n23094 ^ n23041;
  assign n23091 = ~n22780 & n22816;
  assign n23092 = n23091 ^ n22814;
  assign n23096 = n23095 ^ n23092;
  assign n23097 = ~n23090 & ~n23096;
  assign n23098 = n23097 ^ n23095;
  assign n23099 = ~n22818 & n23098;
  assign n23100 = n23099 ^ n20195;
  assign n23101 = n22222 ^ n22150;
  assign n23102 = ~n22181 & n23101;
  assign n23103 = n22180 & n22268;
  assign n23104 = n22149 ^ n22144;
  assign n23105 = n22210 & ~n23104;
  assign n23106 = n22196 ^ n22149;
  assign n23107 = n23106 ^ n22223;
  assign n23108 = ~n22180 & ~n23107;
  assign n23109 = n22222 ^ n22148;
  assign n23110 = ~n23108 & ~n23109;
  assign n23111 = ~n23105 & ~n23110;
  assign n23113 = ~n22152 & n22200;
  assign n23112 = n22182 & n22219;
  assign n23114 = n23113 ^ n23112;
  assign n23115 = n23111 & ~n23114;
  assign n23116 = ~n23103 & n23115;
  assign n23117 = ~n23102 & n23116;
  assign n23118 = ~n22242 & n23117;
  assign n23119 = ~n22290 & n23118;
  assign n23120 = n22204 ^ n22201;
  assign n23121 = ~n22179 & n23120;
  assign n23122 = n23121 ^ n22201;
  assign n23123 = ~n22255 & n23122;
  assign n23124 = n23119 & ~n23123;
  assign n23125 = n22182 & n22267;
  assign n23126 = n23125 ^ n22285;
  assign n23127 = n23124 & ~n23126;
  assign n23128 = n23127 ^ n19602;
  assign n23129 = n22180 & n22203;
  assign n23130 = n22182 & n22217;
  assign n23131 = ~n22179 & n22202;
  assign n23132 = n22143 & n22180;
  assign n23133 = n23132 ^ n22210;
  assign n23134 = ~n22220 & n23133;
  assign n23135 = ~n23131 & ~n23134;
  assign n23136 = n23107 ^ n22219;
  assign n23137 = ~n22181 & n23136;
  assign n23138 = n22222 ^ n22180;
  assign n23139 = n22210 ^ n22150;
  assign n23140 = n22222 & n23139;
  assign n23141 = n23140 ^ n22210;
  assign n23142 = ~n23138 & n23141;
  assign n23143 = n23142 ^ n22180;
  assign n23144 = ~n23137 & ~n23143;
  assign n23145 = n23135 & n23144;
  assign n23146 = ~n23130 & n23145;
  assign n23147 = ~n23129 & n23146;
  assign n23148 = ~n23123 & n23147;
  assign n23149 = ~n22248 & n23148;
  assign n23150 = ~n23126 & n23149;
  assign n23151 = n23150 ^ n18133;
  assign n23152 = n21035 ^ n20997;
  assign n23153 = n23152 ^ n21011;
  assign n23154 = n23153 ^ n21012;
  assign n23155 = n23154 ^ n21012;
  assign n23156 = ~n20291 & n23155;
  assign n23157 = n23156 ^ n21012;
  assign n23158 = n21034 & n23157;
  assign n23159 = n23158 ^ n21012;
  assign n23165 = ~n20030 & n21006;
  assign n23161 = n21024 ^ n21018;
  assign n23160 = n22358 ^ n21001;
  assign n23162 = n23161 ^ n23160;
  assign n23163 = ~n20030 & ~n23162;
  assign n23164 = n23163 ^ n23160;
  assign n23166 = n23165 ^ n23164;
  assign n23167 = ~n20291 & ~n23166;
  assign n23168 = n23167 ^ n23164;
  assign n23169 = ~n23159 & n23168;
  assign n23170 = ~n22355 & n23169;
  assign n23171 = ~n21063 & n23170;
  assign n23172 = n22890 & n23171;
  assign n23173 = n23172 ^ n20460;
  assign y0 = n19551;
  assign y1 = n21072;
  assign y2 = n20029;
  assign y3 = n21418;
  assign y4 = n21458;
  assign y5 = n21489;
  assign y6 = n21511;
  assign y7 = n21740;
  assign y8 = n21774;
  assign y9 = n21820;
  assign y10 = n21853;
  assign y11 = n22022;
  assign y12 = n22038;
  assign y13 = n22250;
  assign y14 = n21926;
  assign y15 = n22292;
  assign y16 = n22311;
  assign y17 = n22332;
  assign y18 = n22354;
  assign y19 = n22388;
  assign y20 = n22425;
  assign y21 = n22448;
  assign y22 = n21897;
  assign y23 = n22472;
  assign y24 = n22178;
  assign y25 = n22511;
  assign y26 = n21359;
  assign y27 = n22602;
  assign y28 = n20290;
  assign y29 = n22631;
  assign y30 = n21542;
  assign y31 = n22718;
  assign y32 = n22135;
  assign y33 = n22755;
  assign y34 = n21188;
  assign y35 = n22778;
  assign y36 = n20853;
  assign y37 = ~n22849;
  assign y38 = n21614;
  assign y39 = n22885;
  assign y40 = n22074;
  assign y41 = n22913;
  assign y42 = n21223;
  assign y43 = n22948;
  assign y44 = n20524;
  assign y45 = n22979;
  assign y46 = n21577;
  assign y47 = n23001;
  assign y48 = n22109;
  assign y49 = n23038;
  assign y50 = n21260;
  assign y51 = n23052;
  assign y52 = n20981;
  assign y53 = n23085;
  assign y54 = n21617;
  assign y55 = n23089;
  assign y56 = n21865;
  assign y57 = n23100;
  assign y58 = n21296;
  assign y59 = n23128;
  assign y60 = n20751;
  assign y61 = n23151;
  assign y62 = n21656;
  assign y63 = n23173;
endmodule
