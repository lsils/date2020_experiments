module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 ;
  assign n66 = ~x15 & ~x31 ;
  assign n65 = ~x47 & ~x63 ;
  assign n67 = n66 ^ n65 ;
  assign n138 = x30 ^ x14 ;
  assign n139 = x31 ^ x15 ;
  assign n141 = x28 ^ x12 ;
  assign n143 = x26 ^ x10 ;
  assign n145 = x24 ^ x8 ;
  assign n147 = x22 ^ x6 ;
  assign n149 = x20 ^ x4 ;
  assign n151 = x18 ^ x2 ;
  assign n153 = x0 & ~x16 ;
  assign n154 = n153 ^ x18 ;
  assign n152 = x18 ^ x1 ;
  assign n155 = n154 ^ n152 ;
  assign n156 = x17 ^ x1 ;
  assign n157 = n155 & ~n156 ;
  assign n158 = n157 ^ n152 ;
  assign n159 = ~n151 & n158 ;
  assign n160 = n159 ^ x2 ;
  assign n161 = n160 ^ x20 ;
  assign n150 = x20 ^ x3 ;
  assign n162 = n161 ^ n150 ;
  assign n163 = x19 ^ x3 ;
  assign n164 = n162 & ~n163 ;
  assign n165 = n164 ^ n150 ;
  assign n166 = ~n149 & n165 ;
  assign n167 = n166 ^ x4 ;
  assign n168 = n167 ^ x22 ;
  assign n148 = x22 ^ x5 ;
  assign n169 = n168 ^ n148 ;
  assign n170 = x21 ^ x5 ;
  assign n171 = n169 & ~n170 ;
  assign n172 = n171 ^ n148 ;
  assign n173 = ~n147 & n172 ;
  assign n174 = n173 ^ x6 ;
  assign n175 = n174 ^ x24 ;
  assign n146 = x24 ^ x7 ;
  assign n176 = n175 ^ n146 ;
  assign n177 = x23 ^ x7 ;
  assign n178 = n176 & ~n177 ;
  assign n179 = n178 ^ n146 ;
  assign n180 = ~n145 & n179 ;
  assign n181 = n180 ^ x8 ;
  assign n182 = n181 ^ x26 ;
  assign n144 = x26 ^ x9 ;
  assign n183 = n182 ^ n144 ;
  assign n184 = x25 ^ x9 ;
  assign n185 = n183 & ~n184 ;
  assign n186 = n185 ^ n144 ;
  assign n187 = ~n143 & n186 ;
  assign n188 = n187 ^ x10 ;
  assign n189 = n188 ^ x28 ;
  assign n142 = x28 ^ x11 ;
  assign n190 = n189 ^ n142 ;
  assign n191 = x27 ^ x11 ;
  assign n192 = n190 & ~n191 ;
  assign n193 = n192 ^ n142 ;
  assign n194 = ~n141 & n193 ;
  assign n195 = n194 ^ x12 ;
  assign n196 = n195 ^ x30 ;
  assign n140 = x30 ^ x13 ;
  assign n197 = n196 ^ n140 ;
  assign n198 = x29 ^ x13 ;
  assign n199 = n197 & ~n198 ;
  assign n200 = n199 ^ n140 ;
  assign n201 = ~n138 & n200 ;
  assign n202 = n201 ^ x14 ;
  assign n203 = n202 ^ x31 ;
  assign n204 = ~n139 & n203 ;
  assign n205 = n204 ^ x15 ;
  assign n206 = n138 & ~n205 ;
  assign n207 = n206 ^ x14 ;
  assign n68 = x62 ^ x46 ;
  assign n69 = x63 ^ x47 ;
  assign n71 = x60 ^ x44 ;
  assign n73 = x58 ^ x42 ;
  assign n75 = x56 ^ x40 ;
  assign n77 = x54 ^ x38 ;
  assign n79 = x52 ^ x36 ;
  assign n81 = x50 ^ x34 ;
  assign n83 = x32 & ~x48 ;
  assign n84 = n83 ^ x50 ;
  assign n82 = x50 ^ x33 ;
  assign n85 = n84 ^ n82 ;
  assign n86 = x49 ^ x33 ;
  assign n87 = n85 & ~n86 ;
  assign n88 = n87 ^ n82 ;
  assign n89 = ~n81 & n88 ;
  assign n90 = n89 ^ x34 ;
  assign n91 = n90 ^ x52 ;
  assign n80 = x52 ^ x35 ;
  assign n92 = n91 ^ n80 ;
  assign n93 = x51 ^ x35 ;
  assign n94 = n92 & ~n93 ;
  assign n95 = n94 ^ n80 ;
  assign n96 = ~n79 & n95 ;
  assign n97 = n96 ^ x36 ;
  assign n98 = n97 ^ x54 ;
  assign n78 = x54 ^ x37 ;
  assign n99 = n98 ^ n78 ;
  assign n100 = x53 ^ x37 ;
  assign n101 = n99 & ~n100 ;
  assign n102 = n101 ^ n78 ;
  assign n103 = ~n77 & n102 ;
  assign n104 = n103 ^ x38 ;
  assign n105 = n104 ^ x56 ;
  assign n76 = x56 ^ x39 ;
  assign n106 = n105 ^ n76 ;
  assign n107 = x55 ^ x39 ;
  assign n108 = n106 & ~n107 ;
  assign n109 = n108 ^ n76 ;
  assign n110 = ~n75 & n109 ;
  assign n111 = n110 ^ x40 ;
  assign n112 = n111 ^ x58 ;
  assign n74 = x58 ^ x41 ;
  assign n113 = n112 ^ n74 ;
  assign n114 = x57 ^ x41 ;
  assign n115 = n113 & ~n114 ;
  assign n116 = n115 ^ n74 ;
  assign n117 = ~n73 & n116 ;
  assign n118 = n117 ^ x42 ;
  assign n119 = n118 ^ x60 ;
  assign n72 = x60 ^ x43 ;
  assign n120 = n119 ^ n72 ;
  assign n121 = x59 ^ x43 ;
  assign n122 = n120 & ~n121 ;
  assign n123 = n122 ^ n72 ;
  assign n124 = ~n71 & n123 ;
  assign n125 = n124 ^ x44 ;
  assign n126 = n125 ^ x62 ;
  assign n70 = x62 ^ x45 ;
  assign n127 = n126 ^ n70 ;
  assign n128 = x61 ^ x45 ;
  assign n129 = n127 & ~n128 ;
  assign n130 = n129 ^ n70 ;
  assign n131 = ~n68 & n130 ;
  assign n132 = n131 ^ x46 ;
  assign n133 = n132 ^ x63 ;
  assign n134 = ~n69 & n133 ;
  assign n135 = n134 ^ x47 ;
  assign n136 = n68 & ~n135 ;
  assign n137 = n136 ^ x46 ;
  assign n208 = n207 ^ n137 ;
  assign n211 = n128 & ~n135 ;
  assign n212 = n211 ^ x45 ;
  assign n209 = n198 & ~n205 ;
  assign n210 = n209 ^ x13 ;
  assign n213 = n212 ^ n210 ;
  assign n216 = n71 & ~n135 ;
  assign n217 = n216 ^ x44 ;
  assign n214 = n141 & ~n205 ;
  assign n215 = n214 ^ x12 ;
  assign n218 = n217 ^ n215 ;
  assign n221 = n191 & ~n205 ;
  assign n222 = n221 ^ x11 ;
  assign n219 = n121 & ~n135 ;
  assign n220 = n219 ^ x43 ;
  assign n223 = n222 ^ n220 ;
  assign n226 = n73 & ~n135 ;
  assign n227 = n226 ^ x42 ;
  assign n224 = n143 & ~n205 ;
  assign n225 = n224 ^ x10 ;
  assign n228 = n227 ^ n225 ;
  assign n231 = n184 & ~n205 ;
  assign n232 = n231 ^ x9 ;
  assign n229 = n114 & ~n135 ;
  assign n230 = n229 ^ x41 ;
  assign n233 = n232 ^ n230 ;
  assign n236 = n75 & ~n135 ;
  assign n237 = n236 ^ x40 ;
  assign n234 = n145 & ~n205 ;
  assign n235 = n234 ^ x8 ;
  assign n238 = n237 ^ n235 ;
  assign n241 = n177 & ~n205 ;
  assign n242 = n241 ^ x7 ;
  assign n239 = n107 & ~n135 ;
  assign n240 = n239 ^ x39 ;
  assign n243 = n242 ^ n240 ;
  assign n246 = n147 & ~n205 ;
  assign n247 = n246 ^ x6 ;
  assign n244 = n77 & ~n135 ;
  assign n245 = n244 ^ x38 ;
  assign n248 = n247 ^ n245 ;
  assign n251 = n170 & ~n205 ;
  assign n252 = n251 ^ x5 ;
  assign n249 = n100 & ~n135 ;
  assign n250 = n249 ^ x37 ;
  assign n253 = n252 ^ n250 ;
  assign n256 = n79 & ~n135 ;
  assign n257 = n256 ^ x36 ;
  assign n254 = n149 & ~n205 ;
  assign n255 = n254 ^ x4 ;
  assign n258 = n257 ^ n255 ;
  assign n261 = n93 & ~n135 ;
  assign n262 = n261 ^ x35 ;
  assign n259 = n163 & ~n205 ;
  assign n260 = n259 ^ x3 ;
  assign n263 = n262 ^ n260 ;
  assign n266 = n151 & ~n205 ;
  assign n267 = n266 ^ x2 ;
  assign n264 = n81 & ~n135 ;
  assign n265 = n264 ^ x34 ;
  assign n268 = n267 ^ n265 ;
  assign n271 = n156 & ~n205 ;
  assign n272 = n271 ^ x1 ;
  assign n269 = n86 & ~n135 ;
  assign n270 = n269 ^ x33 ;
  assign n273 = n272 ^ n270 ;
  assign n274 = x48 ^ x32 ;
  assign n275 = ~n135 & n274 ;
  assign n276 = n275 ^ x32 ;
  assign n277 = x16 ^ x0 ;
  assign n278 = ~n205 & n277 ;
  assign n279 = n278 ^ x0 ;
  assign n280 = ~n276 & n279 ;
  assign n281 = n280 ^ n272 ;
  assign n282 = ~n273 & n281 ;
  assign n283 = n282 ^ n272 ;
  assign n284 = n283 ^ n267 ;
  assign n285 = ~n268 & n284 ;
  assign n286 = n285 ^ n267 ;
  assign n287 = n286 ^ n262 ;
  assign n288 = ~n263 & ~n287 ;
  assign n289 = n288 ^ n262 ;
  assign n290 = n289 ^ n255 ;
  assign n291 = ~n258 & ~n290 ;
  assign n292 = n291 ^ n255 ;
  assign n293 = n292 ^ n252 ;
  assign n294 = ~n253 & n293 ;
  assign n295 = n294 ^ n252 ;
  assign n296 = n295 ^ n245 ;
  assign n297 = ~n248 & ~n296 ;
  assign n298 = n297 ^ n245 ;
  assign n299 = n298 ^ n242 ;
  assign n300 = ~n243 & ~n299 ;
  assign n301 = n300 ^ n242 ;
  assign n302 = n301 ^ n235 ;
  assign n303 = ~n238 & n302 ;
  assign n304 = n303 ^ n235 ;
  assign n305 = n304 ^ n232 ;
  assign n306 = ~n233 & n305 ;
  assign n307 = n306 ^ n232 ;
  assign n308 = n307 ^ n225 ;
  assign n309 = ~n228 & n308 ;
  assign n310 = n309 ^ n225 ;
  assign n311 = n310 ^ n222 ;
  assign n312 = ~n223 & n311 ;
  assign n313 = n312 ^ n222 ;
  assign n314 = n313 ^ n217 ;
  assign n315 = ~n218 & ~n314 ;
  assign n316 = n315 ^ n217 ;
  assign n317 = n316 ^ n212 ;
  assign n318 = ~n213 & ~n317 ;
  assign n319 = n318 ^ n210 ;
  assign n320 = n319 ^ n207 ;
  assign n321 = ~n208 & ~n320 ;
  assign n322 = n321 ^ n137 ;
  assign n323 = n322 ^ n66 ;
  assign n324 = ~n67 & ~n323 ;
  assign n325 = n324 ^ n65 ;
  assign n326 = n205 ^ n135 ;
  assign n327 = n325 & n326 ;
  assign n328 = n327 ^ n135 ;
  assign n329 = n279 ^ n276 ;
  assign n330 = n325 & n329 ;
  assign n331 = n330 ^ n276 ;
  assign n332 = n273 & n325 ;
  assign n333 = n332 ^ n270 ;
  assign n334 = n268 & n325 ;
  assign n335 = n334 ^ n265 ;
  assign n336 = n263 & n325 ;
  assign n337 = n336 ^ n262 ;
  assign n338 = n258 & n325 ;
  assign n339 = n338 ^ n257 ;
  assign n340 = n253 & n325 ;
  assign n341 = n340 ^ n250 ;
  assign n342 = n248 & n325 ;
  assign n343 = n342 ^ n245 ;
  assign n344 = n243 & ~n325 ;
  assign n345 = n344 ^ n242 ;
  assign n346 = n238 & n325 ;
  assign n347 = n346 ^ n237 ;
  assign n348 = n233 & n325 ;
  assign n349 = n348 ^ n230 ;
  assign n350 = n228 & ~n325 ;
  assign n351 = n350 ^ n225 ;
  assign n352 = n223 & ~n325 ;
  assign n353 = n352 ^ n222 ;
  assign n354 = n218 & n325 ;
  assign n355 = n354 ^ n217 ;
  assign n356 = n213 & n325 ;
  assign n357 = n356 ^ n212 ;
  assign n358 = n208 & n325 ;
  assign n359 = n358 ^ n137 ;
  assign n360 = n65 & n66 ;
  assign y0 = ~n328 ;
  assign y1 = ~n325 ;
  assign y2 = n331 ;
  assign y3 = n333 ;
  assign y4 = n335 ;
  assign y5 = n337 ;
  assign y6 = n339 ;
  assign y7 = n341 ;
  assign y8 = n343 ;
  assign y9 = n345 ;
  assign y10 = n347 ;
  assign y11 = n349 ;
  assign y12 = n351 ;
  assign y13 = n353 ;
  assign y14 = n355 ;
  assign y15 = n357 ;
  assign y16 = n359 ;
  assign y17 = ~n360 ;
endmodule
