module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128;
  wire n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437;
  assign n257 = x125 & ~x253;
  assign n258 = ~x126 & ~n257;
  assign n259 = ~x254 & ~n258;
  assign n260 = ~x127 & ~n259;
  assign n261 = ~x252 & ~x253;
  assign n262 = ~x254 & n261;
  assign n263 = x121 & ~x249;
  assign n264 = ~x122 & ~n263;
  assign n265 = ~x250 & ~n264;
  assign n266 = ~x123 & ~n265;
  assign n267 = ~x248 & ~x250;
  assign n268 = ~x249 & n267;
  assign n269 = x120 & n268;
  assign n270 = n266 & ~n269;
  assign n271 = ~x251 & ~n270;
  assign n272 = ~x124 & ~n271;
  assign n273 = ~x247 & ~x251;
  assign n274 = n268 & n273;
  assign n275 = x119 & n274;
  assign n276 = n272 & ~n275;
  assign n277 = ~x246 & n274;
  assign n278 = x118 & n277;
  assign n279 = n276 & ~n278;
  assign n280 = ~x245 & n277;
  assign n281 = x114 & ~x242;
  assign n282 = ~x115 & ~n281;
  assign n283 = ~x241 & ~x242;
  assign n284 = x113 & n283;
  assign n285 = n282 & ~n284;
  assign n286 = ~x243 & ~n285;
  assign n287 = ~x116 & ~n286;
  assign n288 = ~x244 & ~n287;
  assign n289 = ~x117 & ~n288;
  assign n290 = n280 & ~n289;
  assign n291 = n279 & ~n290;
  assign n292 = ~x240 & n283;
  assign n293 = ~x243 & n292;
  assign n294 = ~x244 & n293;
  assign n295 = n280 & n294;
  assign n296 = x111 & ~x239;
  assign n297 = ~x112 & ~n296;
  assign n298 = n295 & ~n297;
  assign n299 = n291 & ~n298;
  assign n300 = x102 & ~x230;
  assign n301 = ~x103 & ~n300;
  assign n302 = ~x229 & ~x230;
  assign n303 = x101 & n302;
  assign n304 = n301 & ~n303;
  assign n305 = ~x231 & ~n304;
  assign n306 = ~x104 & ~n305;
  assign n307 = ~x228 & n302;
  assign n308 = ~x231 & n307;
  assign n309 = x100 & n308;
  assign n310 = n306 & ~n309;
  assign n311 = ~x232 & ~n310;
  assign n312 = ~x105 & ~n311;
  assign n313 = ~x227 & ~x232;
  assign n314 = n308 & n313;
  assign n315 = x99 & n314;
  assign n316 = n312 & ~n315;
  assign n317 = ~x233 & ~n316;
  assign n318 = ~x106 & ~n317;
  assign n319 = ~x234 & ~n318;
  assign n320 = ~x107 & ~n319;
  assign n321 = ~x235 & ~x237;
  assign n322 = ~x236 & n321;
  assign n323 = ~n320 & n322;
  assign n324 = x108 & ~x236;
  assign n325 = ~x109 & ~n324;
  assign n326 = ~x237 & ~n325;
  assign n327 = ~x110 & ~n326;
  assign n328 = ~n323 & n327;
  assign n329 = ~x238 & ~x239;
  assign n330 = n295 & n329;
  assign n331 = ~n328 & n330;
  assign n332 = n299 & ~n331;
  assign n333 = ~x221 & ~x222;
  assign n334 = x93 & n333;
  assign n335 = ~x96 & ~n334;
  assign n336 = x94 & ~x222;
  assign n337 = ~x95 & ~n336;
  assign n338 = ~x97 & ~x98;
  assign n339 = n337 & n338;
  assign n340 = n335 & n339;
  assign n341 = ~x226 & ~x233;
  assign n342 = n314 & n341;
  assign n343 = ~x234 & n342;
  assign n344 = n322 & n343;
  assign n345 = n330 & n344;
  assign n346 = ~x224 & ~x225;
  assign n347 = ~x223 & n346;
  assign n348 = x96 & n346;
  assign n349 = x97 & ~x225;
  assign n350 = ~x98 & ~n349;
  assign n351 = ~n348 & n350;
  assign n352 = ~n347 & n351;
  assign n353 = n345 & ~n352;
  assign n354 = ~n340 & n353;
  assign n355 = n332 & ~n354;
  assign n356 = n345 & n347;
  assign n357 = n333 & n356;
  assign n358 = x89 & ~x217;
  assign n359 = ~x90 & ~n358;
  assign n360 = ~x218 & ~n359;
  assign n361 = ~x91 & ~n360;
  assign n362 = ~x219 & ~n361;
  assign n363 = ~x92 & ~n362;
  assign n364 = ~x216 & ~x217;
  assign n365 = ~x218 & n364;
  assign n366 = ~x219 & n365;
  assign n367 = x85 & ~x213;
  assign n368 = ~x86 & ~n367;
  assign n369 = ~x214 & ~n368;
  assign n370 = ~x87 & ~n369;
  assign n371 = ~x215 & ~n370;
  assign n372 = ~x88 & ~n371;
  assign n373 = ~x212 & ~x213;
  assign n374 = ~x214 & n373;
  assign n375 = ~x215 & n374;
  assign n376 = x82 & ~x210;
  assign n377 = ~x83 & ~n376;
  assign n378 = ~x209 & ~x210;
  assign n379 = x81 & n378;
  assign n380 = n377 & ~n379;
  assign n381 = ~x211 & ~n380;
  assign n382 = ~x84 & ~n381;
  assign n383 = n375 & ~n382;
  assign n384 = n372 & ~n383;
  assign n385 = n366 & ~n384;
  assign n386 = n363 & ~n385;
  assign n387 = x78 & ~x206;
  assign n388 = ~x79 & ~n387;
  assign n389 = ~x207 & ~n388;
  assign n390 = ~x80 & ~n389;
  assign n391 = ~x205 & ~x206;
  assign n392 = ~x207 & n391;
  assign n393 = x76 & ~x204;
  assign n394 = ~x77 & ~n393;
  assign n395 = n392 & ~n394;
  assign n396 = n390 & ~n395;
  assign n397 = ~x203 & ~x204;
  assign n398 = n392 & n397;
  assign n399 = x73 & ~x201;
  assign n400 = ~x74 & ~n399;
  assign n401 = ~x202 & ~n400;
  assign n402 = ~x75 & ~n401;
  assign n403 = n398 & ~n402;
  assign n404 = n396 & ~n403;
  assign n405 = ~x208 & n378;
  assign n406 = ~x211 & n405;
  assign n407 = n375 & n406;
  assign n408 = n366 & n407;
  assign n409 = ~n404 & n408;
  assign n410 = n386 & ~n409;
  assign n411 = ~x220 & ~n410;
  assign n412 = n357 & n411;
  assign n413 = n355 & ~n412;
  assign n414 = x70 & ~x198;
  assign n415 = ~x71 & ~n414;
  assign n416 = ~x197 & ~x198;
  assign n417 = x69 & n416;
  assign n418 = n415 & ~n417;
  assign n419 = ~x199 & ~n418;
  assign n420 = ~x72 & ~n419;
  assign n421 = ~x196 & n416;
  assign n422 = ~x199 & n421;
  assign n423 = x66 & ~x194;
  assign n424 = ~x67 & ~n423;
  assign n425 = ~x193 & ~x194;
  assign n426 = x65 & n425;
  assign n427 = n424 & ~n426;
  assign n428 = ~x195 & ~n427;
  assign n429 = ~x68 & ~n428;
  assign n430 = n422 & ~n429;
  assign n431 = n420 & ~n430;
  assign n432 = ~x192 & n425;
  assign n433 = ~x195 & n432;
  assign n434 = n422 & n433;
  assign n435 = x61 & ~x189;
  assign n436 = ~x62 & ~n435;
  assign n437 = ~x190 & ~n436;
  assign n438 = ~x63 & ~n437;
  assign n439 = ~x191 & ~n438;
  assign n440 = ~x64 & ~n439;
  assign n441 = ~x188 & ~x189;
  assign n442 = ~x190 & n441;
  assign n443 = ~x191 & n442;
  assign n444 = x57 & ~x185;
  assign n445 = ~x58 & ~n444;
  assign n446 = ~x186 & ~n445;
  assign n447 = ~x59 & ~n446;
  assign n448 = ~x187 & ~n447;
  assign n449 = ~x60 & ~n448;
  assign n450 = n443 & ~n449;
  assign n451 = n440 & ~n450;
  assign n452 = n434 & ~n451;
  assign n453 = n431 & ~n452;
  assign n454 = ~x200 & ~x202;
  assign n455 = ~x201 & n454;
  assign n456 = n398 & n455;
  assign n457 = n408 & n456;
  assign n458 = ~x220 & n457;
  assign n459 = n357 & n458;
  assign n460 = ~n453 & n459;
  assign n461 = n413 & ~n460;
  assign n462 = ~x184 & ~x185;
  assign n463 = ~x186 & n462;
  assign n464 = ~x187 & n463;
  assign n465 = n443 & n464;
  assign n466 = n434 & n465;
  assign n467 = n459 & n466;
  assign n468 = x53 & ~x181;
  assign n469 = ~x54 & ~n468;
  assign n470 = ~x182 & ~n469;
  assign n471 = ~x55 & ~n470;
  assign n472 = ~x183 & ~n471;
  assign n473 = ~x56 & ~n472;
  assign n474 = ~x180 & ~x181;
  assign n475 = ~x182 & n474;
  assign n476 = ~x183 & n475;
  assign n477 = x49 & ~x177;
  assign n478 = ~x50 & ~n477;
  assign n479 = ~x178 & ~n478;
  assign n480 = ~x51 & ~n479;
  assign n481 = ~x179 & ~n480;
  assign n482 = ~x52 & ~n481;
  assign n483 = n476 & ~n482;
  assign n484 = n473 & ~n483;
  assign n485 = n467 & ~n484;
  assign n486 = n461 & ~n485;
  assign n487 = n262 & ~n486;
  assign n488 = n260 & ~n487;
  assign n489 = ~x176 & ~x178;
  assign n490 = ~x177 & n489;
  assign n491 = ~x179 & n490;
  assign n492 = n476 & n491;
  assign n493 = n467 & n492;
  assign n494 = n262 & n493;
  assign n495 = x46 & ~x174;
  assign n496 = ~x47 & ~n495;
  assign n497 = ~x173 & ~x174;
  assign n498 = x45 & n497;
  assign n499 = n496 & ~n498;
  assign n500 = ~x172 & n497;
  assign n501 = x44 & n500;
  assign n502 = n499 & ~n501;
  assign n503 = ~x175 & ~n502;
  assign n504 = ~x171 & ~x175;
  assign n505 = n500 & n504;
  assign n506 = x43 & n505;
  assign n507 = ~x48 & ~n506;
  assign n508 = ~n503 & n507;
  assign n509 = ~x170 & n505;
  assign n510 = x41 & ~x169;
  assign n511 = ~x42 & ~n510;
  assign n512 = n509 & ~n511;
  assign n513 = n508 & ~n512;
  assign n514 = n494 & ~n513;
  assign n515 = n488 & ~n514;
  assign n516 = ~x168 & ~x169;
  assign n517 = n509 & n516;
  assign n518 = n494 & n517;
  assign n519 = x38 & ~x166;
  assign n520 = ~x39 & ~n519;
  assign n521 = ~x165 & ~x166;
  assign n522 = x37 & n521;
  assign n523 = n520 & ~n522;
  assign n524 = ~x167 & ~n523;
  assign n525 = ~x40 & ~n524;
  assign n526 = n518 & ~n525;
  assign n527 = n515 & ~n526;
  assign n528 = x34 & ~x162;
  assign n529 = ~x35 & ~n528;
  assign n530 = ~x161 & ~x162;
  assign n531 = x33 & n530;
  assign n532 = n529 & ~n531;
  assign n533 = ~x163 & ~n532;
  assign n534 = ~x36 & ~n533;
  assign n535 = ~x164 & n521;
  assign n536 = ~x167 & n535;
  assign n537 = n518 & n536;
  assign n538 = ~n534 & n537;
  assign n539 = n527 & ~n538;
  assign n540 = ~x160 & n530;
  assign n541 = ~x163 & n540;
  assign n542 = n537 & n541;
  assign n543 = x30 & ~x158;
  assign n544 = ~x31 & ~n543;
  assign n545 = ~x157 & ~x158;
  assign n546 = x29 & n545;
  assign n547 = n544 & ~n546;
  assign n548 = ~x159 & ~n547;
  assign n549 = ~x32 & ~n548;
  assign n550 = n542 & ~n549;
  assign n551 = n539 & ~n550;
  assign n552 = ~x156 & n545;
  assign n553 = ~x159 & n552;
  assign n554 = n542 & n553;
  assign n555 = x27 & ~x155;
  assign n556 = ~x28 & ~n555;
  assign n557 = n554 & ~n556;
  assign n558 = n551 & ~n557;
  assign n559 = ~x154 & ~x155;
  assign n560 = n554 & n559;
  assign n561 = x26 & n560;
  assign n562 = n558 & ~n561;
  assign n563 = ~x153 & n560;
  assign n564 = ~x150 & ~x151;
  assign n565 = ~x149 & n564;
  assign n566 = x20 & ~x148;
  assign n567 = n565 & n566;
  assign n568 = x23 & ~x151;
  assign n569 = ~x24 & ~n568;
  assign n570 = x22 & n564;
  assign n571 = n569 & ~n570;
  assign n572 = x21 & n565;
  assign n573 = n571 & ~n572;
  assign n574 = ~x147 & ~x148;
  assign n575 = n565 & n574;
  assign n576 = x19 & n575;
  assign n577 = n573 & ~n576;
  assign n578 = ~n567 & n577;
  assign n579 = ~x152 & ~n578;
  assign n580 = ~x25 & ~n579;
  assign n581 = n563 & ~n580;
  assign n582 = n562 & ~n581;
  assign n583 = x15 & ~x143;
  assign n584 = ~x16 & ~n583;
  assign n585 = ~x144 & ~n584;
  assign n586 = ~x17 & ~n585;
  assign n587 = ~x145 & ~n586;
  assign n588 = ~x18 & ~n587;
  assign n589 = ~x142 & ~x144;
  assign n590 = ~x143 & n589;
  assign n591 = ~x145 & n590;
  assign n592 = x14 & n591;
  assign n593 = n588 & ~n592;
  assign n594 = ~x146 & ~x152;
  assign n595 = n575 & n594;
  assign n596 = n563 & n595;
  assign n597 = ~n593 & n596;
  assign n598 = n582 & ~n597;
  assign n599 = ~x141 & n591;
  assign n600 = n596 & n599;
  assign n601 = ~x139 & ~x140;
  assign n602 = x11 & n601;
  assign n603 = x12 & ~x140;
  assign n604 = ~x13 & ~n603;
  assign n605 = ~n602 & n604;
  assign n606 = n600 & ~n605;
  assign n607 = n598 & ~n606;
  assign n608 = x7 & ~x135;
  assign n609 = ~x8 & ~n608;
  assign n610 = ~x136 & ~n609;
  assign n611 = ~x9 & ~n610;
  assign n612 = ~x134 & ~x135;
  assign n613 = ~x136 & n612;
  assign n614 = x6 & n613;
  assign n615 = n611 & ~n614;
  assign n616 = ~x137 & ~n615;
  assign n617 = ~x10 & ~n616;
  assign n618 = ~x138 & n601;
  assign n619 = n600 & n618;
  assign n620 = ~n617 & n619;
  assign n621 = n607 & ~n620;
  assign n622 = ~x255 & ~n621;
  assign n623 = ~x0 & ~n622;
  assign n624 = ~x133 & ~x137;
  assign n625 = n613 & n624;
  assign n626 = ~x255 & n625;
  assign n627 = n619 & n626;
  assign n628 = x4 & ~x132;
  assign n629 = ~x5 & ~n628;
  assign n630 = ~x129 & ~x130;
  assign n631 = x1 & n630;
  assign n632 = x2 & ~x130;
  assign n633 = ~x3 & ~n632;
  assign n634 = ~n631 & n633;
  assign n635 = ~x131 & ~x132;
  assign n636 = ~n634 & n635;
  assign n637 = n629 & ~n636;
  assign n638 = n627 & ~n637;
  assign n639 = n623 & ~n638;
  assign n640 = x128 & ~n639;
  assign n641 = ~n633 & n635;
  assign n642 = n629 & ~n641;
  assign n643 = n627 & ~n642;
  assign n644 = n623 & ~n643;
  assign n645 = ~x128 & ~n644;
  assign n646 = ~x1 & ~n645;
  assign n647 = x129 & ~n646;
  assign n648 = x3 & n635;
  assign n649 = n629 & ~n648;
  assign n650 = n627 & ~n649;
  assign n651 = n623 & ~n650;
  assign n652 = ~x128 & ~n651;
  assign n653 = ~x1 & ~n652;
  assign n654 = ~x129 & ~n653;
  assign n655 = ~x2 & ~n654;
  assign n656 = x130 & ~n655;
  assign n657 = ~x128 & n630;
  assign n658 = ~n653 & n657;
  assign n659 = n634 & ~n658;
  assign n660 = x131 & ~n659;
  assign n661 = x5 & n627;
  assign n662 = n623 & ~n661;
  assign n663 = n657 & ~n662;
  assign n664 = n634 & ~n663;
  assign n665 = ~x131 & ~n664;
  assign n666 = ~x4 & ~n665;
  assign n667 = x132 & ~n666;
  assign n668 = n635 & n657;
  assign n669 = ~n623 & n668;
  assign n670 = n637 & ~n669;
  assign n671 = ~x133 & ~n670;
  assign n672 = n671 ^ n670;
  assign n673 = ~x6 & ~n671;
  assign n674 = ~x134 & ~n673;
  assign n675 = n674 ^ n673;
  assign n676 = ~x7 & ~n674;
  assign n677 = ~x135 & ~n676;
  assign n678 = n677 ^ n676;
  assign n679 = ~x8 & ~n677;
  assign n680 = x136 & ~n679;
  assign n681 = n613 & ~n673;
  assign n682 = n611 & ~n681;
  assign n683 = x137 & ~n682;
  assign n684 = x0 & n668;
  assign n685 = n637 & ~n684;
  assign n686 = n625 & ~n685;
  assign n687 = n617 & ~n686;
  assign n688 = n626 & n668;
  assign n689 = ~n607 & n688;
  assign n690 = n687 & ~n689;
  assign n691 = x138 & ~n690;
  assign n692 = x13 & n600;
  assign n693 = n598 & ~n692;
  assign n694 = ~x138 & n688;
  assign n695 = ~n693 & n694;
  assign n696 = ~x138 & ~n687;
  assign n697 = ~x11 & ~n696;
  assign n698 = ~n695 & n697;
  assign n699 = n603 & n694;
  assign n700 = n600 & n699;
  assign n701 = n698 & ~n700;
  assign n702 = x139 & ~n701;
  assign n703 = ~x139 & ~n698;
  assign n704 = ~x12 & ~n703;
  assign n705 = x140 & ~n704;
  assign n706 = n618 & ~n687;
  assign n707 = n605 & ~n706;
  assign n708 = n618 & n688;
  assign n709 = ~n598 & n708;
  assign n710 = n707 & ~n709;
  assign n711 = x141 & ~n710;
  assign n712 = ~x141 & n708;
  assign n713 = ~n582 & n712;
  assign n714 = ~x141 & ~n707;
  assign n715 = ~x14 & ~n714;
  assign n716 = ~n713 & n715;
  assign n717 = n596 & n712;
  assign n718 = ~n588 & n717;
  assign n719 = n716 & ~n718;
  assign n720 = x142 & ~n719;
  assign n721 = x18 & n717;
  assign n722 = n716 & ~n721;
  assign n723 = ~x145 & n717;
  assign n724 = x17 & n723;
  assign n725 = n722 & ~n724;
  assign n726 = ~x142 & ~n725;
  assign n727 = ~x15 & ~n726;
  assign n728 = x16 & n589;
  assign n729 = n723 & n728;
  assign n730 = n727 & ~n729;
  assign n731 = x143 & ~n730;
  assign n732 = ~x143 & ~n727;
  assign n733 = ~x16 & ~n732;
  assign n734 = x144 & ~n733;
  assign n735 = n590 & ~n722;
  assign n736 = n586 & ~n735;
  assign n737 = x145 & ~n736;
  assign n738 = n591 & ~n716;
  assign n739 = n588 & ~n738;
  assign n740 = x146 & ~n739;
  assign n741 = n599 & ~n707;
  assign n742 = n593 & ~n741;
  assign n743 = n599 & n708;
  assign n744 = x25 & n563;
  assign n745 = n562 & ~n744;
  assign n746 = n743 & ~n745;
  assign n747 = n742 & ~n746;
  assign n748 = ~x146 & ~n747;
  assign n749 = ~x19 & ~n748;
  assign n750 = n594 & n743;
  assign n751 = n563 & n750;
  assign n752 = ~n573 & n751;
  assign n753 = n749 & ~n752;
  assign n754 = n567 & n751;
  assign n755 = n753 & ~n754;
  assign n756 = x147 & ~n755;
  assign n757 = ~x147 & ~n753;
  assign n758 = ~x20 & ~n757;
  assign n759 = x148 & ~n758;
  assign n760 = n574 & ~n749;
  assign n761 = ~x21 & ~n566;
  assign n762 = ~n760 & n761;
  assign n763 = n574 & n751;
  assign n764 = ~n571 & n763;
  assign n765 = n762 & ~n764;
  assign n766 = x149 & ~n765;
  assign n767 = ~n569 & n763;
  assign n768 = n762 & ~n767;
  assign n769 = ~x149 & ~n768;
  assign n770 = ~x22 & ~n769;
  assign n771 = x150 & ~n770;
  assign n772 = x24 & n763;
  assign n773 = n762 & ~n772;
  assign n774 = ~x149 & ~n773;
  assign n775 = ~x22 & ~n774;
  assign n776 = ~x150 & ~n775;
  assign n777 = ~x23 & ~n776;
  assign n778 = x151 & ~n777;
  assign n779 = n565 & ~n762;
  assign n780 = n571 & ~n779;
  assign n781 = x152 & ~n780;
  assign n782 = n595 & ~n742;
  assign n783 = n580 & ~n782;
  assign n784 = n595 & n743;
  assign n785 = ~n562 & n784;
  assign n786 = n783 & ~n785;
  assign n787 = x153 & ~n786;
  assign n788 = ~x153 & ~n783;
  assign n789 = ~x26 & ~n788;
  assign n790 = ~x153 & n784;
  assign n791 = ~n558 & n790;
  assign n792 = n789 & ~n791;
  assign n793 = x154 & ~n792;
  assign n794 = x28 & n554;
  assign n795 = n551 & ~n794;
  assign n796 = n790 & ~n795;
  assign n797 = n789 & ~n796;
  assign n798 = ~x154 & ~n797;
  assign n799 = ~x27 & ~n798;
  assign n800 = x155 & ~n799;
  assign n801 = n559 & ~n789;
  assign n802 = n556 & ~n801;
  assign n803 = n559 & n790;
  assign n804 = ~n551 & n803;
  assign n805 = n802 & ~n804;
  assign n806 = x156 & ~n805;
  assign n807 = x32 & n542;
  assign n808 = n539 & ~n807;
  assign n809 = n803 & ~n808;
  assign n810 = n802 & ~n809;
  assign n811 = ~x159 & n803;
  assign n812 = n542 & n811;
  assign n813 = ~n544 & n812;
  assign n814 = n810 & ~n813;
  assign n815 = ~x156 & ~n814;
  assign n816 = ~x29 & ~n815;
  assign n817 = x157 & ~n816;
  assign n818 = x31 & n812;
  assign n819 = n810 & ~n818;
  assign n820 = ~x156 & ~n819;
  assign n821 = ~x29 & ~n820;
  assign n822 = ~x157 & ~n821;
  assign n823 = ~x30 & ~n822;
  assign n824 = x158 & ~n823;
  assign n825 = n552 & ~n810;
  assign n826 = n547 & ~n825;
  assign n827 = x159 & ~n826;
  assign n828 = n553 & ~n802;
  assign n829 = n549 & ~n828;
  assign n830 = n553 & n803;
  assign n831 = ~n539 & n830;
  assign n832 = n829 & ~n831;
  assign n833 = x160 & ~n832;
  assign n834 = x36 & n537;
  assign n835 = n527 & ~n834;
  assign n836 = n830 & ~n835;
  assign n837 = n829 & ~n836;
  assign n838 = ~x163 & n830;
  assign n839 = n537 & n838;
  assign n840 = ~n529 & n839;
  assign n841 = n837 & ~n840;
  assign n842 = ~x160 & ~n841;
  assign n843 = ~x33 & ~n842;
  assign n844 = x161 & ~n843;
  assign n845 = x35 & n839;
  assign n846 = n837 & ~n845;
  assign n847 = ~x160 & ~n846;
  assign n848 = ~x33 & ~n847;
  assign n849 = ~x161 & ~n848;
  assign n850 = ~x34 & ~n849;
  assign n851 = x162 & ~n850;
  assign n852 = n540 & ~n837;
  assign n853 = n532 & ~n852;
  assign n854 = x163 & ~n853;
  assign n855 = n541 & ~n829;
  assign n856 = n534 & ~n855;
  assign n857 = n541 & n830;
  assign n858 = ~n527 & n857;
  assign n859 = n856 & ~n858;
  assign n860 = x164 & ~n859;
  assign n861 = x40 & n518;
  assign n862 = n515 & ~n861;
  assign n863 = n857 & ~n862;
  assign n864 = n856 & ~n863;
  assign n865 = ~x167 & n857;
  assign n866 = n518 & n865;
  assign n867 = ~n520 & n866;
  assign n868 = n864 & ~n867;
  assign n869 = ~x164 & ~n868;
  assign n870 = ~x37 & ~n869;
  assign n871 = x165 & ~n870;
  assign n872 = x39 & n866;
  assign n873 = n864 & ~n872;
  assign n874 = ~x164 & ~n873;
  assign n875 = ~x37 & ~n874;
  assign n876 = ~x165 & ~n875;
  assign n877 = ~x38 & ~n876;
  assign n878 = x166 & ~n877;
  assign n879 = n535 & ~n864;
  assign n880 = n523 & ~n879;
  assign n881 = x167 & ~n880;
  assign n882 = n536 & ~n856;
  assign n883 = n525 & ~n882;
  assign n884 = n536 & n857;
  assign n885 = ~n515 & n884;
  assign n886 = n883 & ~n885;
  assign n887 = x168 & ~n886;
  assign n888 = ~n488 & n884;
  assign n889 = n883 & ~n888;
  assign n890 = n494 & n884;
  assign n891 = x42 & n509;
  assign n892 = n508 & ~n891;
  assign n893 = n890 & ~n892;
  assign n894 = n889 & ~n893;
  assign n895 = ~x168 & ~n894;
  assign n896 = ~x41 & ~n895;
  assign n897 = x169 & ~n896;
  assign n898 = n516 & ~n889;
  assign n899 = n511 & ~n898;
  assign n900 = n516 & n890;
  assign n901 = ~n508 & n900;
  assign n902 = n899 & ~n901;
  assign n903 = x170 & ~n902;
  assign n904 = ~x170 & ~n899;
  assign n905 = ~x170 & n900;
  assign n906 = x48 & n905;
  assign n907 = ~x43 & ~n906;
  assign n908 = ~n904 & n907;
  assign n909 = n503 & n905;
  assign n910 = n908 & ~n909;
  assign n911 = x171 & ~n910;
  assign n912 = ~x171 & ~n908;
  assign n913 = ~x44 & ~n912;
  assign n914 = n504 & n905;
  assign n915 = ~n499 & n914;
  assign n916 = n913 & ~n915;
  assign n917 = x172 & ~n916;
  assign n918 = ~n496 & n914;
  assign n919 = n913 & ~n918;
  assign n920 = ~x172 & ~n919;
  assign n921 = ~x45 & ~n920;
  assign n922 = x173 & ~n921;
  assign n923 = x47 & n914;
  assign n924 = n913 & ~n923;
  assign n925 = ~x172 & ~n924;
  assign n926 = ~x45 & ~n925;
  assign n927 = ~x173 & ~n926;
  assign n928 = ~x46 & ~n927;
  assign n929 = x174 & ~n928;
  assign n930 = n500 & ~n913;
  assign n931 = n499 & ~n930;
  assign n932 = x175 & ~n931;
  assign n933 = n517 & ~n889;
  assign n934 = n513 & ~n933;
  assign n935 = x176 & ~n934;
  assign n936 = n517 & n884;
  assign n937 = ~n260 & n936;
  assign n938 = n517 & ~n883;
  assign n939 = n513 & ~n938;
  assign n940 = ~n937 & n939;
  assign n941 = n262 & n936;
  assign n942 = ~n461 & n941;
  assign n943 = n940 & ~n942;
  assign n944 = n467 & n941;
  assign n945 = x52 & n476;
  assign n946 = n473 & ~n945;
  assign n947 = n944 & ~n946;
  assign n948 = n943 & ~n947;
  assign n949 = ~x179 & n476;
  assign n950 = n944 & n949;
  assign n951 = x51 & n950;
  assign n952 = n948 & ~n951;
  assign n953 = ~x176 & ~n952;
  assign n954 = ~x49 & ~n953;
  assign n955 = x50 & n489;
  assign n956 = n950 & n955;
  assign n957 = n954 & ~n956;
  assign n958 = x177 & ~n957;
  assign n959 = ~x177 & ~n954;
  assign n960 = ~x50 & ~n959;
  assign n961 = x178 & ~n960;
  assign n962 = n490 & ~n948;
  assign n963 = n480 & ~n962;
  assign n964 = x179 & ~n963;
  assign n965 = n491 & ~n943;
  assign n966 = n482 & ~n965;
  assign n967 = n491 & n944;
  assign n968 = ~n473 & n967;
  assign n969 = n966 & ~n968;
  assign n970 = x180 & ~n969;
  assign n971 = x56 & n967;
  assign n972 = n966 & ~n971;
  assign n973 = ~x183 & n967;
  assign n974 = x55 & n973;
  assign n975 = n972 & ~n974;
  assign n976 = x54 & ~x182;
  assign n977 = n973 & n976;
  assign n978 = n975 & ~n977;
  assign n979 = ~x180 & ~n978;
  assign n980 = ~x53 & ~n979;
  assign n981 = x181 & ~n980;
  assign n982 = n474 & ~n975;
  assign n983 = n469 & ~n982;
  assign n984 = x182 & ~n983;
  assign n985 = n475 & ~n972;
  assign n986 = n471 & ~n985;
  assign n987 = x183 & ~n986;
  assign n988 = n476 & ~n966;
  assign n989 = n473 & ~n988;
  assign n990 = x184 & ~n989;
  assign n991 = n492 & ~n940;
  assign n992 = n484 & ~n991;
  assign n993 = n492 & n941;
  assign n994 = ~n413 & n993;
  assign n995 = n992 & ~n994;
  assign n996 = n459 & n993;
  assign n997 = ~n431 & n996;
  assign n998 = n995 & ~n997;
  assign n999 = n434 & n996;
  assign n1000 = ~n440 & n999;
  assign n1001 = n998 & ~n1000;
  assign n1002 = n443 & n999;
  assign n1003 = x60 & n1002;
  assign n1004 = n1001 & ~n1003;
  assign n1005 = ~x187 & n1002;
  assign n1006 = x59 & n1005;
  assign n1007 = n1004 & ~n1006;
  assign n1008 = x58 & ~x186;
  assign n1009 = n1005 & n1008;
  assign n1010 = n1007 & ~n1009;
  assign n1011 = ~x184 & ~n1010;
  assign n1012 = ~x57 & ~n1011;
  assign n1013 = x185 & ~n1012;
  assign n1014 = n462 & ~n1007;
  assign n1015 = n445 & ~n1014;
  assign n1016 = x186 & ~n1015;
  assign n1017 = n463 & ~n1004;
  assign n1018 = n447 & ~n1017;
  assign n1019 = x187 & ~n1018;
  assign n1020 = n464 & ~n1001;
  assign n1021 = n449 & ~n1020;
  assign n1022 = x188 & ~n1021;
  assign n1023 = x64 & n999;
  assign n1024 = n998 & ~n1023;
  assign n1025 = n464 & ~n1024;
  assign n1026 = n449 & ~n1025;
  assign n1027 = ~x191 & n464;
  assign n1028 = n999 & n1027;
  assign n1029 = x63 & n1028;
  assign n1030 = n1026 & ~n1029;
  assign n1031 = x62 & ~x190;
  assign n1032 = n1028 & n1031;
  assign n1033 = n1030 & ~n1032;
  assign n1034 = ~x188 & ~n1033;
  assign n1035 = ~x61 & ~n1034;
  assign n1036 = x189 & ~n1035;
  assign n1037 = n441 & ~n1030;
  assign n1038 = n436 & ~n1037;
  assign n1039 = x190 & ~n1038;
  assign n1040 = n442 & ~n1026;
  assign n1041 = n438 & ~n1040;
  assign n1042 = x191 & ~n1041;
  assign n1043 = n465 & ~n998;
  assign n1044 = n451 & ~n1043;
  assign n1045 = x192 & ~n1044;
  assign n1046 = n465 & ~n995;
  assign n1047 = n451 & ~n1046;
  assign n1048 = n465 & n996;
  assign n1049 = ~n420 & n1048;
  assign n1050 = n1047 & ~n1049;
  assign n1051 = n422 & n1048;
  assign n1052 = x68 & n1051;
  assign n1053 = n1050 & ~n1052;
  assign n1054 = ~x195 & n1051;
  assign n1055 = ~n424 & n1054;
  assign n1056 = n1053 & ~n1055;
  assign n1057 = ~x192 & ~n1056;
  assign n1058 = ~x65 & ~n1057;
  assign n1059 = x193 & ~n1058;
  assign n1060 = x67 & n1054;
  assign n1061 = n1053 & ~n1060;
  assign n1062 = ~x192 & ~n1061;
  assign n1063 = ~x65 & ~n1062;
  assign n1064 = ~x193 & ~n1063;
  assign n1065 = ~x66 & ~n1064;
  assign n1066 = x194 & ~n1065;
  assign n1067 = n432 & ~n1053;
  assign n1068 = n427 & ~n1067;
  assign n1069 = x195 & ~n1068;
  assign n1070 = n433 & ~n1050;
  assign n1071 = n429 & ~n1070;
  assign n1072 = x196 & ~n1071;
  assign n1073 = x72 & n1048;
  assign n1074 = n1047 & ~n1073;
  assign n1075 = n433 & ~n1074;
  assign n1076 = n429 & ~n1075;
  assign n1077 = ~x199 & n433;
  assign n1078 = n1048 & n1077;
  assign n1079 = ~n415 & n1078;
  assign n1080 = n1076 & ~n1079;
  assign n1081 = ~x196 & ~n1080;
  assign n1082 = ~x69 & ~n1081;
  assign n1083 = x197 & ~n1082;
  assign n1084 = x71 & n1078;
  assign n1085 = n1076 & ~n1084;
  assign n1086 = ~x196 & ~n1085;
  assign n1087 = ~x69 & ~n1086;
  assign n1088 = ~x197 & ~n1087;
  assign n1089 = ~x70 & ~n1088;
  assign n1090 = x198 & ~n1089;
  assign n1091 = n421 & ~n1076;
  assign n1092 = n418 & ~n1091;
  assign n1093 = x199 & ~n1092;
  assign n1094 = n434 & ~n1047;
  assign n1095 = n431 & ~n1094;
  assign n1096 = x200 & ~n1095;
  assign n1097 = n466 & ~n992;
  assign n1098 = n453 & ~n1097;
  assign n1099 = n466 & n993;
  assign n1100 = ~n355 & n1099;
  assign n1101 = n1098 & ~n1100;
  assign n1102 = ~x220 & n357;
  assign n1103 = n1099 & n1102;
  assign n1104 = ~n386 & n1103;
  assign n1105 = n1101 & ~n1104;
  assign n1106 = n408 & n1103;
  assign n1107 = x75 & n398;
  assign n1108 = n396 & ~n1107;
  assign n1109 = n1106 & ~n1108;
  assign n1110 = n1105 & ~n1109;
  assign n1111 = ~x200 & ~n1110;
  assign n1112 = ~x73 & ~n1111;
  assign n1113 = x74 & n454;
  assign n1114 = n398 & n1113;
  assign n1115 = n1106 & n1114;
  assign n1116 = n1112 & ~n1115;
  assign n1117 = x201 & ~n1116;
  assign n1118 = ~x201 & ~n1112;
  assign n1119 = ~x74 & ~n1118;
  assign n1120 = x202 & ~n1119;
  assign n1121 = n455 & ~n1105;
  assign n1122 = n402 & ~n1121;
  assign n1123 = n455 & n1106;
  assign n1124 = ~n396 & n1123;
  assign n1125 = n1122 & ~n1124;
  assign n1126 = x203 & ~n1125;
  assign n1127 = x77 & n392;
  assign n1128 = n390 & ~n1127;
  assign n1129 = n1123 & ~n1128;
  assign n1130 = n1122 & ~n1129;
  assign n1131 = ~x203 & ~n1130;
  assign n1132 = ~x76 & ~n1131;
  assign n1133 = x204 & ~n1132;
  assign n1134 = n397 & ~n1122;
  assign n1135 = n394 & ~n1134;
  assign n1136 = n397 & n1123;
  assign n1137 = ~n390 & n1136;
  assign n1138 = n1135 & ~n1137;
  assign n1139 = x205 & ~n1138;
  assign n1140 = x80 & n1136;
  assign n1141 = n1135 & ~n1140;
  assign n1142 = x79 & ~x207;
  assign n1143 = n1136 & n1142;
  assign n1144 = n1141 & ~n1143;
  assign n1145 = ~x205 & ~n1144;
  assign n1146 = ~x78 & ~n1145;
  assign n1147 = x206 & ~n1146;
  assign n1148 = n391 & ~n1141;
  assign n1149 = n388 & ~n1148;
  assign n1150 = x207 & ~n1149;
  assign n1151 = n392 & ~n1135;
  assign n1152 = n390 & ~n1151;
  assign n1153 = x208 & ~n1152;
  assign n1154 = n456 & ~n1101;
  assign n1155 = n404 & ~n1154;
  assign n1156 = n456 & n1103;
  assign n1157 = ~n363 & n1156;
  assign n1158 = n1155 & ~n1157;
  assign n1159 = n366 & n1156;
  assign n1160 = x84 & n375;
  assign n1161 = n372 & ~n1160;
  assign n1162 = n1159 & ~n1161;
  assign n1163 = n1158 & ~n1162;
  assign n1164 = ~x211 & n375;
  assign n1165 = n1159 & n1164;
  assign n1166 = ~n377 & n1165;
  assign n1167 = n1163 & ~n1166;
  assign n1168 = ~x208 & ~n1167;
  assign n1169 = ~x81 & ~n1168;
  assign n1170 = x209 & ~n1169;
  assign n1171 = x83 & n1165;
  assign n1172 = n1163 & ~n1171;
  assign n1173 = ~x208 & ~n1172;
  assign n1174 = ~x81 & ~n1173;
  assign n1175 = ~x209 & ~n1174;
  assign n1176 = ~x82 & ~n1175;
  assign n1177 = x210 & ~n1176;
  assign n1178 = n405 & ~n1163;
  assign n1179 = n380 & ~n1178;
  assign n1180 = x211 & ~n1179;
  assign n1181 = n406 & ~n1158;
  assign n1182 = n382 & ~n1181;
  assign n1183 = n406 & n1159;
  assign n1184 = ~n372 & n1183;
  assign n1185 = n1182 & ~n1184;
  assign n1186 = x212 & ~n1185;
  assign n1187 = x88 & n1183;
  assign n1188 = n1182 & ~n1187;
  assign n1189 = ~x215 & n1183;
  assign n1190 = x87 & n1189;
  assign n1191 = n1188 & ~n1190;
  assign n1192 = x86 & ~x214;
  assign n1193 = n1189 & n1192;
  assign n1194 = n1191 & ~n1193;
  assign n1195 = ~x212 & ~n1194;
  assign n1196 = ~x85 & ~n1195;
  assign n1197 = x213 & ~n1196;
  assign n1198 = n373 & ~n1191;
  assign n1199 = n368 & ~n1198;
  assign n1200 = x214 & ~n1199;
  assign n1201 = n374 & ~n1188;
  assign n1202 = n370 & ~n1201;
  assign n1203 = x215 & ~n1202;
  assign n1204 = n375 & ~n1182;
  assign n1205 = n372 & ~n1204;
  assign n1206 = x216 & ~n1205;
  assign n1207 = x92 & n1156;
  assign n1208 = n1155 & ~n1207;
  assign n1209 = n407 & ~n1208;
  assign n1210 = n384 & ~n1209;
  assign n1211 = ~x219 & n407;
  assign n1212 = n1156 & n1211;
  assign n1213 = x91 & n1212;
  assign n1214 = n1210 & ~n1213;
  assign n1215 = x90 & ~x218;
  assign n1216 = n1212 & n1215;
  assign n1217 = n1214 & ~n1216;
  assign n1218 = ~x216 & ~n1217;
  assign n1219 = ~x89 & ~n1218;
  assign n1220 = x217 & ~n1219;
  assign n1221 = n364 & ~n1214;
  assign n1222 = n359 & ~n1221;
  assign n1223 = x218 & ~n1222;
  assign n1224 = n365 & ~n1210;
  assign n1225 = n361 & ~n1224;
  assign n1226 = x219 & ~n1225;
  assign n1227 = n457 & ~n1101;
  assign n1228 = n410 & ~n1227;
  assign n1229 = x220 & ~n1228;
  assign n1230 = n458 & ~n1098;
  assign n1231 = ~x93 & ~n411;
  assign n1232 = ~n1230 & n1231;
  assign n1233 = n458 & n1099;
  assign n1234 = n345 & ~n351;
  assign n1235 = n332 & ~n1234;
  assign n1236 = x95 & n356;
  assign n1237 = n1235 & ~n1236;
  assign n1238 = n1233 & ~n1237;
  assign n1239 = n1232 & ~n1238;
  assign n1240 = n336 & n356;
  assign n1241 = n1233 & n1240;
  assign n1242 = n1239 & ~n1241;
  assign n1243 = x221 & ~n1242;
  assign n1244 = ~x221 & ~n1239;
  assign n1245 = ~x94 & ~n1244;
  assign n1246 = x222 & ~n1245;
  assign n1247 = n333 & ~n1232;
  assign n1248 = n337 & ~n1247;
  assign n1249 = n333 & n1233;
  assign n1250 = ~n1235 & n1249;
  assign n1251 = n1248 & ~n1250;
  assign n1252 = x223 & ~n1251;
  assign n1253 = ~n332 & n1249;
  assign n1254 = n1248 & ~n1253;
  assign n1255 = n345 & n1249;
  assign n1256 = ~n350 & n1255;
  assign n1257 = n1254 & ~n1256;
  assign n1258 = ~x223 & ~n1257;
  assign n1259 = ~x96 & ~n1258;
  assign n1260 = x224 & ~n1259;
  assign n1261 = x98 & n1255;
  assign n1262 = n1254 & ~n1261;
  assign n1263 = ~x223 & ~n1262;
  assign n1264 = ~x96 & ~n1263;
  assign n1265 = ~x224 & ~n1264;
  assign n1266 = ~x97 & ~n1265;
  assign n1267 = x225 & ~n1266;
  assign n1268 = n340 & ~n1247;
  assign n1269 = ~n1253 & n1268;
  assign n1270 = x226 & ~n352;
  assign n1271 = ~n1269 & n1270;
  assign n1272 = ~n352 & ~n1268;
  assign n1273 = n347 & n1249;
  assign n1274 = x110 & n330;
  assign n1275 = n299 & ~n1274;
  assign n1276 = n1273 & ~n1275;
  assign n1277 = ~n1272 & ~n1276;
  assign n1278 = n330 & n1273;
  assign n1279 = n322 & n1278;
  assign n1280 = x107 & n1279;
  assign n1281 = n326 & n1278;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = n1277 & n1282;
  assign n1284 = ~x234 & n1279;
  assign n1285 = x106 & n1284;
  assign n1286 = n1283 & ~n1285;
  assign n1287 = ~x226 & ~n1286;
  assign n1288 = ~x99 & ~n1287;
  assign n1289 = n341 & n1284;
  assign n1290 = ~n312 & n1289;
  assign n1291 = n1288 & ~n1290;
  assign n1292 = x227 & ~n1291;
  assign n1293 = ~x231 & ~n301;
  assign n1294 = ~x104 & ~n1293;
  assign n1295 = ~x232 & ~n1294;
  assign n1296 = ~x105 & ~n1295;
  assign n1297 = n1289 & ~n1296;
  assign n1298 = n1288 & ~n1297;
  assign n1299 = ~x227 & ~n1298;
  assign n1300 = ~x100 & ~n1299;
  assign n1301 = ~n306 & n313;
  assign n1302 = n1289 & n1301;
  assign n1303 = n1300 & ~n1302;
  assign n1304 = x228 & ~n1303;
  assign n1305 = ~x228 & ~n1300;
  assign n1306 = ~x101 & ~n1305;
  assign n1307 = ~x229 & ~n1306;
  assign n1308 = n1307 ^ n1306;
  assign n1309 = ~x102 & ~n1307;
  assign n1310 = x230 & ~n1309;
  assign n1311 = n307 & ~n1300;
  assign n1312 = n304 & ~n1311;
  assign n1313 = ~x231 & ~n1312;
  assign n1314 = n1313 ^ n1312;
  assign n1315 = ~x104 & ~n1313;
  assign n1316 = x232 & ~n1315;
  assign n1317 = n314 & ~n1288;
  assign n1318 = n312 & ~n1317;
  assign n1319 = x233 & ~n1318;
  assign n1320 = n342 & ~n1283;
  assign n1321 = n318 & ~n1320;
  assign n1322 = x234 & ~n1321;
  assign n1323 = n343 & ~n1277;
  assign n1324 = n320 & ~n1323;
  assign n1325 = n343 & n1281;
  assign n1326 = n1324 & ~n1325;
  assign n1327 = x235 & ~n1326;
  assign n1328 = ~x235 & ~n1324;
  assign n1329 = ~x108 & ~n1328;
  assign n1330 = x109 & n321;
  assign n1331 = n343 & n1330;
  assign n1332 = n1278 & n1331;
  assign n1333 = n1329 & ~n1332;
  assign n1334 = x236 & ~n1333;
  assign n1335 = ~x236 & ~n1329;
  assign n1336 = ~x109 & ~n1335;
  assign n1337 = x237 & ~n1336;
  assign n1338 = n344 & ~n1277;
  assign n1339 = n328 & ~n1338;
  assign n1340 = ~x238 & ~n1339;
  assign n1341 = n1340 ^ n1339;
  assign n1342 = ~x111 & ~n1340;
  assign n1343 = x239 & ~n1342;
  assign n1344 = ~n328 & n329;
  assign n1345 = n297 & ~n1344;
  assign n1346 = n329 & n344;
  assign n1347 = n1272 & n1346;
  assign n1348 = n1345 & ~n1347;
  assign n1349 = n1273 & n1346;
  assign n1350 = ~n291 & n1349;
  assign n1351 = n1348 & ~n1350;
  assign n1352 = x240 & ~n1351;
  assign n1353 = ~n279 & n1349;
  assign n1354 = n1348 & ~n1353;
  assign n1355 = n280 & n1349;
  assign n1356 = x117 & n1355;
  assign n1357 = n1354 & ~n1356;
  assign n1358 = ~x244 & n1355;
  assign n1359 = x116 & n1358;
  assign n1360 = n1357 & ~n1359;
  assign n1361 = ~x243 & n1358;
  assign n1362 = ~n282 & n1361;
  assign n1363 = n1360 & ~n1362;
  assign n1364 = ~x240 & ~n1363;
  assign n1365 = ~x113 & ~n1364;
  assign n1366 = x241 & ~n1365;
  assign n1367 = x115 & n1361;
  assign n1368 = n1360 & ~n1367;
  assign n1369 = ~x240 & ~n1368;
  assign n1370 = ~x113 & ~n1369;
  assign n1371 = ~x241 & ~n1370;
  assign n1372 = ~x114 & ~n1371;
  assign n1373 = x242 & ~n1372;
  assign n1374 = n292 & ~n1360;
  assign n1375 = n285 & ~n1374;
  assign n1376 = x243 & ~n1375;
  assign n1377 = n293 & ~n1357;
  assign n1378 = n287 & ~n1377;
  assign n1379 = x244 & ~n1378;
  assign n1380 = n294 & ~n1354;
  assign n1381 = n289 & ~n1380;
  assign n1382 = x245 & ~n1381;
  assign n1383 = ~x245 & n294;
  assign n1384 = ~n1348 & n1383;
  assign n1385 = ~x245 & ~n289;
  assign n1386 = ~x118 & ~n1385;
  assign n1387 = ~n1384 & n1386;
  assign n1388 = n1349 & n1383;
  assign n1389 = ~n276 & n1388;
  assign n1390 = n1387 & ~n1389;
  assign n1391 = x246 & ~n1390;
  assign n1392 = ~x246 & ~n1387;
  assign n1393 = ~x246 & n1388;
  assign n1394 = ~n272 & n1393;
  assign n1395 = ~x119 & ~n1394;
  assign n1396 = ~n1392 & n1395;
  assign n1397 = x247 & ~n1396;
  assign n1398 = x124 & n1393;
  assign n1399 = ~x119 & ~n1398;
  assign n1400 = ~n1392 & n1399;
  assign n1401 = ~x247 & ~n1400;
  assign n1402 = ~x120 & ~n1401;
  assign n1403 = n273 & n1393;
  assign n1404 = ~n266 & n1403;
  assign n1405 = n1402 & ~n1404;
  assign n1406 = x248 & ~n1405;
  assign n1407 = x123 & n1403;
  assign n1408 = n1402 & ~n1407;
  assign n1409 = ~x248 & ~n1408;
  assign n1410 = ~x121 & ~n1409;
  assign n1411 = x122 & n267;
  assign n1412 = n1403 & n1411;
  assign n1413 = n1410 & ~n1412;
  assign n1414 = x249 & ~n1413;
  assign n1415 = ~x249 & ~n1410;
  assign n1416 = ~x122 & ~n1415;
  assign n1417 = x250 & ~n1416;
  assign n1418 = n268 & ~n1402;
  assign n1419 = n266 & ~n1418;
  assign n1420 = x251 & ~n1419;
  assign n1421 = n493 & ~n992;
  assign n1422 = n486 & ~n1421;
  assign n1423 = ~x252 & ~n1422;
  assign n1424 = n1423 ^ n1422;
  assign n1425 = ~x125 & ~n1423;
  assign n1426 = x253 & ~n1425;
  assign n1427 = x127 & n936;
  assign n1428 = n939 & ~n1427;
  assign n1429 = n493 & ~n1428;
  assign n1430 = n486 & ~n1429;
  assign n1431 = n261 & ~n1430;
  assign n1432 = n258 & ~n1431;
  assign n1433 = x254 & ~n1432;
  assign n1434 = n494 & ~n939;
  assign n1435 = n488 & ~n1434;
  assign n1436 = x255 & ~n1435;
  assign n1437 = n494 & n936;
  assign y0 = n640;
  assign y1 = n647;
  assign y2 = n656;
  assign y3 = n660;
  assign y4 = n667;
  assign y5 = ~n672;
  assign y6 = ~n675;
  assign y7 = ~n678;
  assign y8 = n680;
  assign y9 = n683;
  assign y10 = n691;
  assign y11 = n702;
  assign y12 = n705;
  assign y13 = n711;
  assign y14 = n720;
  assign y15 = n731;
  assign y16 = n734;
  assign y17 = n737;
  assign y18 = n740;
  assign y19 = n756;
  assign y20 = n759;
  assign y21 = n766;
  assign y22 = n771;
  assign y23 = n778;
  assign y24 = n781;
  assign y25 = n787;
  assign y26 = n793;
  assign y27 = n800;
  assign y28 = n806;
  assign y29 = n817;
  assign y30 = n824;
  assign y31 = n827;
  assign y32 = n833;
  assign y33 = n844;
  assign y34 = n851;
  assign y35 = n854;
  assign y36 = n860;
  assign y37 = n871;
  assign y38 = n878;
  assign y39 = n881;
  assign y40 = n887;
  assign y41 = n897;
  assign y42 = n903;
  assign y43 = n911;
  assign y44 = n917;
  assign y45 = n922;
  assign y46 = n929;
  assign y47 = n932;
  assign y48 = n935;
  assign y49 = n958;
  assign y50 = n961;
  assign y51 = n964;
  assign y52 = n970;
  assign y53 = n981;
  assign y54 = n984;
  assign y55 = n987;
  assign y56 = n990;
  assign y57 = n1013;
  assign y58 = n1016;
  assign y59 = n1019;
  assign y60 = n1022;
  assign y61 = n1036;
  assign y62 = n1039;
  assign y63 = n1042;
  assign y64 = n1045;
  assign y65 = n1059;
  assign y66 = n1066;
  assign y67 = n1069;
  assign y68 = n1072;
  assign y69 = n1083;
  assign y70 = n1090;
  assign y71 = n1093;
  assign y72 = n1096;
  assign y73 = n1117;
  assign y74 = n1120;
  assign y75 = n1126;
  assign y76 = n1133;
  assign y77 = n1139;
  assign y78 = n1147;
  assign y79 = n1150;
  assign y80 = n1153;
  assign y81 = n1170;
  assign y82 = n1177;
  assign y83 = n1180;
  assign y84 = n1186;
  assign y85 = n1197;
  assign y86 = n1200;
  assign y87 = n1203;
  assign y88 = n1206;
  assign y89 = n1220;
  assign y90 = n1223;
  assign y91 = n1226;
  assign y92 = n1229;
  assign y93 = n1243;
  assign y94 = n1246;
  assign y95 = n1252;
  assign y96 = n1260;
  assign y97 = n1267;
  assign y98 = n1271;
  assign y99 = n1292;
  assign y100 = n1304;
  assign y101 = ~n1308;
  assign y102 = n1310;
  assign y103 = ~n1314;
  assign y104 = n1316;
  assign y105 = n1319;
  assign y106 = n1322;
  assign y107 = n1327;
  assign y108 = n1334;
  assign y109 = n1337;
  assign y110 = ~n1341;
  assign y111 = n1343;
  assign y112 = n1352;
  assign y113 = n1366;
  assign y114 = n1373;
  assign y115 = n1376;
  assign y116 = n1379;
  assign y117 = n1382;
  assign y118 = n1391;
  assign y119 = n1397;
  assign y120 = n1406;
  assign y121 = n1414;
  assign y122 = n1417;
  assign y123 = n1420;
  assign y124 = ~n1424;
  assign y125 = n1426;
  assign y126 = n1433;
  assign y127 = n1436;
  assign y128 = ~n1437;
endmodule
