module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127;
  wire n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180;
  assign n1160 = x245 ^ x241;
  assign n1149 = x246 ^ x244;
  assign n1161 = n1160 ^ n1149;
  assign n1150 = x243 ^ x240;
  assign n1145 = x242 ^ x241;
  assign n1146 = n1145 ^ x247;
  assign n1147 = n1146 ^ x243;
  assign n1188 = n1150 ^ n1147;
  assign n1172 = x245 ^ x242;
  assign n1179 = n1172 ^ n1149;
  assign n1187 = n1179 ^ n1146;
  assign n1192 = n1188 ^ n1187;
  assign n1189 = n1187 & n1188;
  assign n1152 = x246 ^ x240;
  assign n1183 = n1152 & n1179;
  assign n1190 = n1189 ^ n1183;
  assign n1151 = n1150 ^ n1149;
  assign n1156 = n1151 ^ n1145;
  assign n1157 = x245 ^ x240;
  assign n1163 = n1156 & n1157;
  assign n1162 = n1150 & n1161;
  assign n1164 = n1163 ^ n1162;
  assign n1191 = n1190 ^ n1164;
  assign n1193 = n1192 ^ n1191;
  assign n1182 = ~x246 & n1146;
  assign n1184 = n1183 ^ n1182;
  assign n1180 = n1179 ^ n1152;
  assign n1144 = x245 ^ x243;
  assign n1173 = n1172 ^ n1150;
  assign n1174 = n1144 & n1173;
  assign n1175 = n1174 ^ n1162;
  assign n1181 = n1180 ^ n1175;
  assign n1185 = n1184 ^ n1181;
  assign n1197 = n1193 ^ n1185;
  assign n1171 = n1160 ^ n1151;
  assign n1176 = n1175 ^ n1171;
  assign n1166 = n1151 ^ x247;
  assign n1167 = n1146 ^ x246;
  assign n1168 = n1167 ^ n1157;
  assign n1169 = n1166 & n1168;
  assign n1153 = n1152 ^ n1144;
  assign n1154 = n1151 & n1153;
  assign n1170 = n1169 ^ n1154;
  assign n1177 = n1176 ^ n1170;
  assign n1186 = n1177 & n1185;
  assign n1158 = n1157 ^ n1156;
  assign n1148 = x247 & n1147;
  assign n1155 = n1154 ^ n1148;
  assign n1159 = n1158 ^ n1155;
  assign n1165 = n1164 ^ n1159;
  assign n1198 = n1186 ^ n1165;
  assign n1199 = n1197 & n1198;
  assign n1200 = n1199 ^ n1193;
  assign n1178 = n1177 ^ n1165;
  assign n1194 = n1193 ^ n1186;
  assign n1195 = n1178 & n1194;
  assign n1196 = n1195 ^ n1165;
  assign n1201 = n1200 ^ n1196;
  assign n1655 = n1161 & n1201;
  assign n1208 = n1197 ^ n1186;
  assign n1206 = n1165 & n1185;
  assign n1207 = ~n1193 & n1206;
  assign n1209 = n1208 ^ n1207;
  assign n1204 = n1186 ^ n1178;
  assign n1202 = ~n1165 & n1177;
  assign n1203 = n1193 & n1202;
  assign n1205 = n1204 ^ n1203;
  assign n1210 = n1209 ^ n1205;
  assign n1211 = n1210 ^ n1201;
  assign n1250 = n1173 & n1211;
  assign n1656 = n1655 ^ n1250;
  assign n1219 = n1209 ^ n1200;
  assign n1641 = n1151 & n1219;
  assign n1221 = n1166 & n1209;
  assign n1220 = n1153 & n1219;
  assign n1222 = n1221 ^ n1220;
  assign n1642 = n1641 ^ n1222;
  assign n1738 = n1656 ^ n1642;
  assign n1217 = n1168 & n1209;
  assign n1213 = n1150 & n1201;
  assign n1212 = n1144 & n1211;
  assign n1214 = n1213 ^ n1212;
  assign n1737 = n1217 ^ n1214;
  assign n1739 = n1738 ^ n1737;
  assign n1740 = n1739 ^ x137;
  assign n1741 = n1740 ^ x169;
  assign n1742 = n1741 ^ x201;
  assign n1743 = n1742 ^ x233;
  assign n1716 = n1655 ^ n1213;
  assign n1713 = n1157 & n1210;
  assign n1714 = n1713 ^ x138;
  assign n1710 = n1188 & n1196;
  assign n1226 = x247 & n1200;
  assign n1709 = n1641 ^ n1226;
  assign n1711 = n1710 ^ n1709;
  assign n1248 = n1156 & n1210;
  assign n1246 = n1205 ^ n1196;
  assign n1247 = n1152 & n1246;
  assign n1249 = n1248 ^ n1247;
  assign n1712 = n1711 ^ n1249;
  assign n1715 = n1714 ^ n1712;
  assign n1717 = n1716 ^ n1715;
  assign n1718 = n1717 ^ x170;
  assign n1719 = n1718 ^ x202;
  assign n1720 = n1719 ^ x234;
  assign n5055 = n1743 ^ n1720;
  assign n1244 = n1167 & n1205;
  assign n1225 = n1187 & n1196;
  assign n1245 = n1244 ^ n1225;
  assign n1751 = n1709 ^ n1245;
  assign n1638 = n1179 & n1246;
  assign n1639 = n1638 ^ n1214;
  assign n1750 = n1639 ^ n1247;
  assign n1752 = n1751 ^ n1750;
  assign n1753 = n1752 ^ x143;
  assign n1754 = n1753 ^ x175;
  assign n1755 = n1754 ^ x207;
  assign n1756 = n1755 ^ x239;
  assign n5056 = n5055 ^ n1756;
  assign n1787 = n1147 & n1200;
  assign n1216 = n1146 & n1205;
  assign n1218 = n1217 ^ n1216;
  assign n1788 = n1787 ^ n1218;
  assign n1251 = n1250 ^ n1249;
  assign n1785 = n1711 ^ n1251;
  assign n1784 = n1639 ^ x141;
  assign n1786 = n1785 ^ n1784;
  assign n1789 = n1788 ^ n1786;
  assign n1790 = n1789 ^ x173;
  assign n1791 = n1790 ^ x205;
  assign n1792 = n1791 ^ x237;
  assign n5059 = n1792 ^ n1720;
  assign n1253 = n1216 ^ n1214;
  assign n1252 = n1251 ^ n1245;
  assign n1254 = n1253 ^ n1252;
  assign n1255 = n1254 ^ x142;
  assign n1256 = n1255 ^ x174;
  assign n1257 = n1256 ^ x206;
  assign n1258 = n1257 ^ x238;
  assign n1227 = n1226 ^ n1225;
  assign n1223 = n1222 ^ n1218;
  assign n1215 = n1214 ^ x140;
  assign n1224 = n1223 ^ n1215;
  assign n1228 = n1227 ^ n1224;
  assign n1229 = n1228 ^ x172;
  assign n1230 = n1229 ^ x204;
  assign n1231 = n1230 ^ x236;
  assign n5051 = n1258 ^ n1231;
  assign n5060 = n5059 ^ n5051;
  assign n5061 = n5060 ^ n5056;
  assign n1643 = n1642 ^ n1218;
  assign n1640 = n1639 ^ x139;
  assign n1644 = n1643 ^ n1640;
  assign n1645 = n1644 ^ x171;
  assign n1646 = n1645 ^ x203;
  assign n1647 = n1646 ^ x235;
  assign n5057 = n5056 ^ n1647;
  assign n1657 = n1656 ^ n1218;
  assign n1654 = n1639 ^ n1220;
  assign n1658 = n1657 ^ n1654;
  assign n1659 = n1658 ^ x136;
  assign n1660 = n1659 ^ x168;
  assign n1661 = n1660 ^ x200;
  assign n1662 = n1661 ^ x232;
  assign n5052 = n1662 ^ n1647;
  assign n5058 = n5057 ^ n5052;
  assign n5074 = n5061 ^ n5058;
  assign n5069 = n1792 ^ n1743;
  assign n5070 = n5069 ^ n5051;
  assign n5071 = n5052 & n5070;
  assign n5066 = n1792 ^ n1662;
  assign n5053 = n5052 ^ n5051;
  assign n5067 = n5055 ^ n5053;
  assign n5068 = n5066 & ~n5067;
  assign n5072 = n5071 ^ n5068;
  assign n5063 = n1662 ^ n1258;
  assign n5064 = n5060 & ~n5063;
  assign n5062 = ~n5058 & ~n5061;
  assign n5065 = n5064 ^ n5062;
  assign n5073 = n5072 ^ n5065;
  assign n5075 = n5074 ^ n5073;
  assign n5089 = n5067 ^ n5066;
  assign n5076 = n1792 ^ n1647;
  assign n5086 = n5076 ^ n5063;
  assign n5087 = ~n5053 & ~n5086;
  assign n5085 = ~n1756 & ~n5057;
  assign n5088 = n5087 ^ n5085;
  assign n5090 = n5089 ^ n5088;
  assign n5091 = n5090 ^ n5072;
  assign n5099 = n5069 ^ n5053;
  assign n5077 = n5059 ^ n5052;
  assign n5078 = n5076 & ~n5077;
  assign n5079 = n5078 ^ n5071;
  assign n5100 = n5099 ^ n5079;
  assign n5054 = n5053 ^ n1756;
  assign n5095 = n5056 ^ n1258;
  assign n5096 = n5095 ^ n5066;
  assign n5097 = n5054 & n5096;
  assign n5098 = n5097 ^ n5087;
  assign n5101 = n5100 ^ n5098;
  assign n5116 = n5091 & n5101;
  assign n5117 = n5075 & n5116;
  assign n5114 = n5101 ^ n5091;
  assign n5082 = n1258 & ~n5056;
  assign n5083 = n5082 ^ n5064;
  assign n5080 = n5063 ^ n5060;
  assign n5081 = n5080 ^ n5079;
  assign n5084 = n5083 ^ n5081;
  assign n5102 = ~n5084 & n5101;
  assign n5115 = n5114 ^ n5102;
  assign n5118 = n5117 ^ n5115;
  assign n5635 = ~n5056 & ~n5118;
  assign n5094 = n5084 ^ n5075;
  assign n5103 = n5102 ^ n5094;
  assign n5092 = ~n5084 & ~n5091;
  assign n5093 = ~n5075 & n5092;
  assign n5104 = n5103 ^ n5093;
  assign n5132 = n5096 & ~n5104;
  assign n5636 = n5635 ^ n5132;
  assign n5120 = n5102 ^ n5075;
  assign n5121 = ~n5114 & n5120;
  assign n5122 = n5121 ^ n5091;
  assign n5106 = n5102 ^ n5091;
  assign n5107 = ~n5094 & ~n5106;
  assign n5108 = n5107 ^ n5075;
  assign n5123 = n5122 ^ n5108;
  assign n5126 = n5070 & ~n5123;
  assign n5119 = n5118 ^ n5104;
  assign n5124 = n5123 ^ n5119;
  assign n5125 = ~n5077 & ~n5124;
  assign n5127 = n5126 ^ n5125;
  assign n5673 = n5636 ^ n5127;
  assign n5527 = n5122 ^ n5118;
  assign n5584 = n5060 & n5527;
  assign n5130 = n5052 & ~n5123;
  assign n5129 = n5076 & ~n5124;
  assign n5131 = n5130 ^ n5129;
  assign n5585 = n5584 ^ n5131;
  assign n5109 = n5108 ^ n5104;
  assign n5110 = ~n5086 & ~n5109;
  assign n5672 = n5585 ^ n5110;
  assign n5674 = n5673 ^ n5672;
  assign n2798 = x234 ^ x233;
  assign n2799 = n2798 ^ x239;
  assign n2811 = x237 ^ x233;
  assign n2801 = x235 ^ x232;
  assign n2796 = x238 ^ x236;
  assign n2807 = n2801 ^ n2796;
  assign n2839 = n2811 ^ n2807;
  assign n2792 = x237 ^ x235;
  assign n2795 = x237 ^ x234;
  assign n2818 = n2801 ^ n2795;
  assign n2819 = n2792 & n2818;
  assign n2812 = n2811 ^ n2796;
  assign n2813 = n2801 & n2812;
  assign n2820 = n2819 ^ n2813;
  assign n2840 = n2839 ^ n2820;
  assign n2834 = n2807 ^ x239;
  assign n2835 = n2799 ^ x238;
  assign n2809 = x237 ^ x232;
  assign n2836 = n2835 ^ n2809;
  assign n2837 = n2834 & n2836;
  assign n2793 = x238 ^ x232;
  assign n2794 = n2793 ^ n2792;
  assign n2827 = n2794 & n2807;
  assign n2838 = n2837 ^ n2827;
  assign n2841 = n2840 ^ n2838;
  assign n2808 = n2807 ^ n2798;
  assign n2829 = n2809 ^ n2808;
  assign n2802 = n2799 ^ x235;
  assign n2826 = x239 & n2802;
  assign n2828 = n2827 ^ n2826;
  assign n2830 = n2829 ^ n2828;
  assign n2810 = n2808 & n2809;
  assign n2814 = n2813 ^ n2810;
  assign n2831 = n2830 ^ n2814;
  assign n2853 = n2841 ^ n2831;
  assign n2823 = ~x238 & n2799;
  assign n2797 = n2796 ^ n2795;
  assign n2805 = n2793 & n2797;
  assign n2824 = n2823 ^ n2805;
  assign n2821 = n2797 ^ n2793;
  assign n2822 = n2821 ^ n2820;
  assign n2825 = n2824 ^ n2822;
  assign n2842 = n2825 & n2841;
  assign n2854 = n2853 ^ n2842;
  assign n2803 = n2802 ^ n2801;
  assign n2800 = n2799 ^ n2797;
  assign n2816 = n2803 ^ n2800;
  assign n2804 = n2800 & n2803;
  assign n2806 = n2805 ^ n2804;
  assign n2815 = n2814 ^ n2806;
  assign n2817 = n2816 ^ n2815;
  assign n2851 = ~n2831 & n2841;
  assign n2852 = n2817 & n2851;
  assign n2855 = n2854 ^ n2852;
  assign n2873 = n2799 & n2855;
  assign n2843 = n2825 ^ n2817;
  assign n2844 = n2843 ^ n2842;
  assign n2832 = n2825 & n2831;
  assign n2833 = ~n2817 & n2832;
  assign n2845 = n2844 ^ n2833;
  assign n2872 = n2836 & n2845;
  assign n2874 = n2873 ^ n2872;
  assign n2857 = n2842 ^ n2817;
  assign n2858 = n2853 & n2857;
  assign n2859 = n2858 ^ n2831;
  assign n2846 = n2842 ^ n2831;
  assign n2847 = n2843 & n2846;
  assign n2848 = n2847 ^ n2817;
  assign n2860 = n2859 ^ n2848;
  assign n2856 = n2855 ^ n2845;
  assign n2861 = n2860 ^ n2856;
  assign n2870 = n2818 & n2861;
  assign n2869 = n2812 & n2860;
  assign n2871 = n2870 ^ n2869;
  assign n2875 = n2874 ^ n2871;
  assign n2865 = n2859 ^ n2855;
  assign n2866 = n2797 & n2865;
  assign n2863 = n2801 & n2860;
  assign n2862 = n2792 & n2861;
  assign n2864 = n2863 ^ n2862;
  assign n2867 = n2866 ^ n2864;
  assign n2849 = n2848 ^ n2845;
  assign n2850 = n2794 & n2849;
  assign n2868 = n2867 ^ n2850;
  assign n2876 = n2875 ^ n2868;
  assign n2877 = n2876 ^ x128;
  assign n5675 = n5674 ^ n2877;
  assign n2878 = n2877 ^ x160;
  assign n5676 = n5675 ^ n2878;
  assign n2879 = n2878 ^ x192;
  assign n7570 = n5676 ^ n2879;
  assign n4460 = n2879 ^ x224;
  assign n8250 = n7570 ^ n4460;
  assign n5112 = ~n5053 & ~n5109;
  assign n5105 = n5054 & ~n5104;
  assign n5111 = n5110 ^ n5105;
  assign n5113 = n5112 ^ n5111;
  assign n5707 = n5636 ^ n5113;
  assign n3301 = n2834 & n2845;
  assign n3302 = n3301 ^ n2850;
  assign n3254 = n2807 & n2849;
  assign n3303 = n3302 ^ n3254;
  assign n3304 = n3303 ^ n2874;
  assign n3300 = n2867 ^ x131;
  assign n3305 = n3304 ^ n3300;
  assign n5706 = n5585 ^ n3305;
  assign n5708 = n5707 ^ n5706;
  assign n3306 = n3305 ^ x163;
  assign n5709 = n5708 ^ n3306;
  assign n3307 = n3306 ^ x195;
  assign n7579 = n5709 ^ n3307;
  assign n4454 = n3307 ^ x227;
  assign n8249 = n7579 ^ n4454;
  assign n8251 = n8250 ^ n8249;
  assign n5133 = n5132 ^ n5131;
  assign n5128 = n5127 ^ n5113;
  assign n5134 = n5133 ^ n5128;
  assign n3396 = n2872 ^ n2864;
  assign n3395 = n3303 ^ n2871;
  assign n3397 = n3396 ^ n3395;
  assign n3398 = n3397 ^ x129;
  assign n5135 = n5134 ^ n3398;
  assign n3399 = n3398 ^ x161;
  assign n5136 = n5135 ^ n3399;
  assign n3400 = n3399 ^ x193;
  assign n7596 = n5136 ^ n3400;
  assign n4488 = n3400 ^ x225;
  assign n8262 = n7596 ^ n4488;
  assign n5534 = n5130 ^ n5126;
  assign n5531 = n5066 & n5119;
  assign n3371 = n2869 ^ n2863;
  assign n3368 = n2809 & n2856;
  assign n3369 = n3368 ^ x130;
  assign n3257 = n2803 & n2859;
  assign n3255 = x239 & n2848;
  assign n3256 = n3255 ^ n3254;
  assign n3258 = n3257 ^ n3256;
  assign n3231 = n2808 & n2856;
  assign n3230 = n2793 & n2865;
  assign n3232 = n3231 ^ n3230;
  assign n3367 = n3258 ^ n3232;
  assign n3370 = n3369 ^ n3367;
  assign n3372 = n3371 ^ n3370;
  assign n5532 = n5531 ^ n3372;
  assign n5528 = ~n5063 & n5527;
  assign n5526 = ~n5067 & n5119;
  assign n5529 = n5528 ^ n5526;
  assign n5524 = ~n5058 & ~n5122;
  assign n5522 = ~n1756 & n5108;
  assign n5523 = n5522 ^ n5112;
  assign n5525 = n5524 ^ n5523;
  assign n5530 = n5529 ^ n5525;
  assign n5533 = n5532 ^ n5530;
  assign n5535 = n5534 ^ n5533;
  assign n3373 = n3372 ^ x162;
  assign n5536 = n5535 ^ n3373;
  assign n3374 = n3373 ^ x194;
  assign n7591 = n5536 ^ n3374;
  assign n4483 = n3374 ^ x226;
  assign n8258 = n7591 ^ n4483;
  assign n8272 = n8262 ^ n8258;
  assign n5631 = n5529 ^ n5125;
  assign n5588 = ~n5061 & ~n5122;
  assign n5587 = n5095 & ~n5118;
  assign n5589 = n5588 ^ n5587;
  assign n5728 = n5631 ^ n5589;
  assign n5727 = n5635 ^ n5131;
  assign n5729 = n5728 ^ n5727;
  assign n3235 = n2873 ^ n2864;
  assign n3233 = n3232 ^ n2870;
  assign n3228 = n2800 & n2859;
  assign n3227 = n2835 & n2855;
  assign n3229 = n3228 ^ n3227;
  assign n3234 = n3233 ^ n3229;
  assign n3236 = n3235 ^ n3234;
  assign n3237 = n3236 ^ x134;
  assign n5730 = n5729 ^ n3237;
  assign n3238 = n3237 ^ x166;
  assign n5731 = n5730 ^ n3238;
  assign n3239 = n3238 ^ x198;
  assign n7559 = n5731 ^ n3239;
  assign n4467 = n3239 ^ x230;
  assign n8253 = n7559 ^ n4467;
  assign n5747 = n5588 ^ n5522;
  assign n5745 = n5636 ^ n5111;
  assign n3344 = n3255 ^ n3228;
  assign n3342 = n3302 ^ n2874;
  assign n3341 = n2864 ^ x132;
  assign n3343 = n3342 ^ n3341;
  assign n3345 = n3344 ^ n3343;
  assign n5744 = n5131 ^ n3345;
  assign n5746 = n5745 ^ n5744;
  assign n5748 = n5747 ^ n5746;
  assign n3346 = n3345 ^ x164;
  assign n5749 = n5748 ^ n3346;
  assign n3347 = n3346 ^ x196;
  assign n7564 = n5749 ^ n3347;
  assign n4475 = n3347 ^ x228;
  assign n8252 = n7564 ^ n4475;
  assign n8254 = n8253 ^ n8252;
  assign n8255 = n8254 ^ n8251;
  assign n8279 = n8272 ^ n8255;
  assign n5634 = ~n5057 & n5108;
  assign n5637 = n5636 ^ n5634;
  assign n5632 = n5631 ^ n5525;
  assign n3261 = n2802 & n2848;
  assign n3262 = n3261 ^ n2874;
  assign n3259 = n3258 ^ n3233;
  assign n3253 = n2867 ^ x133;
  assign n3260 = n3259 ^ n3253;
  assign n3263 = n3262 ^ n3260;
  assign n5630 = n5585 ^ n3263;
  assign n5633 = n5632 ^ n5630;
  assign n5638 = n5637 ^ n5633;
  assign n3264 = n3263 ^ x165;
  assign n5639 = n5638 ^ n3264;
  assign n3265 = n3264 ^ x197;
  assign n7604 = n5639 ^ n3265;
  assign n4498 = n3265 ^ x229;
  assign n8256 = n7604 ^ n4498;
  assign n8278 = n8256 ^ n8250;
  assign n8304 = n8279 ^ n8278;
  assign n5590 = n5589 ^ n5523;
  assign n5586 = n5585 ^ n5528;
  assign n5591 = n5590 ^ n5586;
  assign n3427 = n3256 ^ n3229;
  assign n3426 = n3230 ^ n2867;
  assign n3428 = n3427 ^ n3426;
  assign n3429 = n3428 ^ x135;
  assign n5592 = n5591 ^ n3429;
  assign n3430 = n3429 ^ x167;
  assign n5593 = n5592 ^ n3430;
  assign n3431 = n3430 ^ x199;
  assign n7584 = n5593 ^ n3431;
  assign n4448 = n3431 ^ x231;
  assign n8271 = n7584 ^ n4448;
  assign n8273 = n8272 ^ n8271;
  assign n8283 = n8273 ^ n8249;
  assign n8302 = ~n8271 & ~n8283;
  assign n8267 = n8253 ^ n8250;
  assign n8257 = n8256 ^ n8249;
  assign n8295 = n8267 ^ n8257;
  assign n8296 = n8255 & n8295;
  assign n8303 = n8302 ^ n8296;
  assign n8305 = n8304 ^ n8303;
  assign n8280 = n8278 & n8279;
  assign n8263 = n8262 ^ n8256;
  assign n8264 = n8263 ^ n8254;
  assign n8265 = n8251 & ~n8264;
  assign n8281 = n8280 ^ n8265;
  assign n8306 = n8305 ^ n8281;
  assign n8298 = n8263 ^ n8255;
  assign n8259 = n8258 ^ n8256;
  assign n8260 = n8259 ^ n8251;
  assign n8261 = n8257 & ~n8260;
  assign n8266 = n8265 ^ n8261;
  assign n8299 = n8298 ^ n8266;
  assign n8291 = n8273 ^ n8253;
  assign n8292 = n8291 ^ n8278;
  assign n8293 = n8271 ^ n8255;
  assign n8294 = ~n8292 & ~n8293;
  assign n8297 = n8296 ^ n8294;
  assign n8300 = n8299 ^ n8297;
  assign n8320 = n8306 ^ n8300;
  assign n8268 = n8259 ^ n8254;
  assign n8275 = n8267 & ~n8268;
  assign n8274 = ~n8253 & ~n8273;
  assign n8276 = n8275 ^ n8274;
  assign n8269 = n8268 ^ n8267;
  assign n8270 = n8269 ^ n8266;
  assign n8277 = n8276 ^ n8270;
  assign n8301 = ~n8277 & ~n8300;
  assign n8284 = n8283 ^ n8251;
  assign n8282 = n8273 ^ n8268;
  assign n8288 = n8284 ^ n8282;
  assign n8285 = n8282 & ~n8284;
  assign n8286 = n8285 ^ n8275;
  assign n8287 = n8286 ^ n8281;
  assign n8289 = n8288 ^ n8287;
  assign n8321 = n8301 ^ n8289;
  assign n8322 = ~n8320 & ~n8321;
  assign n8323 = n8322 ^ n8306;
  assign n8290 = n8289 ^ n8277;
  assign n8307 = n8306 ^ n8301;
  assign n8308 = n8290 & n8307;
  assign n8309 = n8308 ^ n8289;
  assign n8324 = n8323 ^ n8309;
  assign n8335 = n8251 & ~n8324;
  assign n8332 = ~n8264 & ~n8324;
  assign n8741 = n8335 ^ n8332;
  assign n8327 = n8320 ^ n8301;
  assign n8325 = ~n8300 & ~n8306;
  assign n8326 = ~n8289 & n8325;
  assign n8328 = n8327 ^ n8326;
  assign n8311 = ~n8277 & n8306;
  assign n8312 = n8289 & n8311;
  assign n8310 = n8301 ^ n8290;
  assign n8313 = n8312 ^ n8310;
  assign n8329 = n8328 ^ n8313;
  assign n8738 = n8278 & ~n8329;
  assign n5978 = n4498 ^ n4488;
  assign n5960 = n4475 ^ n4467;
  assign n5979 = n5978 ^ n5960;
  assign n5962 = n4488 ^ n4483;
  assign n5963 = n5962 ^ n4448;
  assign n5959 = n4498 ^ n4483;
  assign n5961 = n5960 ^ n5959;
  assign n6004 = n5963 ^ n5961;
  assign n5966 = n4460 ^ n4454;
  assign n5964 = n5963 ^ n4454;
  assign n6003 = n5966 ^ n5964;
  assign n6008 = n6004 ^ n6003;
  assign n6005 = n6003 & n6004;
  assign n5969 = n4467 ^ n4460;
  assign n5998 = n5961 & ~n5969;
  assign n6006 = n6005 ^ n5998;
  assign n5980 = n5966 & n5979;
  assign n5973 = n4498 ^ n4460;
  assign n5967 = n5966 ^ n5960;
  assign n5974 = n5967 ^ n5962;
  assign n5977 = n5973 & ~n5974;
  assign n5981 = n5980 ^ n5977;
  assign n6007 = n6006 ^ n5981;
  assign n6009 = n6008 ^ n6007;
  assign n5997 = n4467 & n5963;
  assign n5999 = n5998 ^ n5997;
  assign n5995 = n5969 ^ n5961;
  assign n5968 = n4498 ^ n4454;
  assign n5984 = n5966 ^ n5959;
  assign n5985 = n5968 & ~n5984;
  assign n5986 = n5985 ^ n5980;
  assign n5996 = n5995 ^ n5986;
  assign n6000 = n5999 ^ n5996;
  assign n6018 = n6009 ^ n6000;
  assign n5988 = n5967 ^ n4448;
  assign n5989 = n5963 ^ n4467;
  assign n5990 = n5989 ^ n5973;
  assign n5991 = ~n5988 & ~n5990;
  assign n5970 = n5969 ^ n5968;
  assign n5971 = ~n5967 & ~n5970;
  assign n5992 = n5991 ^ n5971;
  assign n5983 = n5978 ^ n5967;
  assign n5987 = n5986 ^ n5983;
  assign n5993 = n5992 ^ n5987;
  assign n6001 = n5993 & ~n6000;
  assign n5975 = n5974 ^ n5973;
  assign n5965 = n4448 & n5964;
  assign n5972 = n5971 ^ n5965;
  assign n5976 = n5975 ^ n5972;
  assign n5982 = n5981 ^ n5976;
  assign n6019 = n6001 ^ n5982;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = n6020 ^ n6009;
  assign n5994 = n5993 ^ n5982;
  assign n6013 = n6009 ^ n6001;
  assign n6014 = ~n5994 & n6013;
  assign n6015 = n6014 ^ n5982;
  assign n6022 = n6021 ^ n6015;
  assign n6482 = n5979 & ~n6022;
  assign n6023 = n5966 & ~n6022;
  assign n6575 = n6482 ^ n6023;
  assign n6026 = n6018 ^ n6001;
  assign n6024 = ~n5982 & ~n6000;
  assign n6025 = ~n6009 & n6024;
  assign n6027 = n6026 ^ n6025;
  assign n6010 = n5982 & n5993;
  assign n6011 = n6009 & n6010;
  assign n6002 = n6001 ^ n5994;
  assign n6012 = n6011 ^ n6002;
  assign n6028 = n6027 ^ n6012;
  assign n6572 = n5973 & n6028;
  assign n1963 = x227 ^ x224;
  assign n1980 = x229 ^ x225;
  assign n1964 = x230 ^ x228;
  assign n1965 = n1964 ^ n1963;
  assign n2009 = n1980 ^ n1965;
  assign n1987 = x229 ^ x227;
  assign n1970 = x229 ^ x226;
  assign n1988 = n1970 ^ n1963;
  assign n1989 = n1987 & n1988;
  assign n1981 = n1980 ^ n1964;
  assign n1982 = n1963 & n1981;
  assign n1990 = n1989 ^ n1982;
  assign n2010 = n2009 ^ n1990;
  assign n1966 = x226 ^ x225;
  assign n1967 = n1966 ^ x231;
  assign n2004 = n1967 ^ x230;
  assign n1977 = x229 ^ x224;
  assign n2005 = n2004 ^ n1977;
  assign n2006 = n1965 ^ x231;
  assign n2007 = n2005 & n2006;
  assign n1974 = x230 ^ x224;
  assign n1998 = n1987 ^ n1974;
  assign n1999 = n1965 & n1998;
  assign n2008 = n2007 ^ n1999;
  assign n2011 = n2010 ^ n2008;
  assign n1978 = n1966 ^ n1965;
  assign n2001 = n1978 ^ n1977;
  assign n1968 = n1967 ^ x227;
  assign n1997 = x231 & n1968;
  assign n2000 = n1999 ^ n1997;
  assign n2002 = n2001 ^ n2000;
  assign n1979 = n1977 & n1978;
  assign n1983 = n1982 ^ n1979;
  assign n2003 = n2002 ^ n1983;
  assign n2026 = n2011 ^ n2003;
  assign n1993 = ~x230 & n1967;
  assign n1971 = n1970 ^ n1964;
  assign n1975 = n1971 & n1974;
  assign n1994 = n1993 ^ n1975;
  assign n1991 = n1974 ^ n1971;
  assign n1992 = n1991 ^ n1990;
  assign n1995 = n1994 ^ n1992;
  assign n2012 = n1995 & n2011;
  assign n1972 = n1971 ^ n1967;
  assign n1969 = n1968 ^ n1963;
  assign n1985 = n1972 ^ n1969;
  assign n1973 = n1969 & n1972;
  assign n1976 = n1975 ^ n1973;
  assign n1984 = n1983 ^ n1976;
  assign n1986 = n1985 ^ n1984;
  assign n2027 = n2012 ^ n1986;
  assign n2028 = n2026 & n2027;
  assign n2029 = n2028 ^ n2003;
  assign n1996 = n1995 ^ n1986;
  assign n2013 = n2012 ^ n2003;
  assign n2014 = n1996 & n2013;
  assign n2015 = n2014 ^ n1986;
  assign n2030 = n2029 ^ n2015;
  assign n2042 = n1963 & n2030;
  assign n2031 = n1981 & n2030;
  assign n2404 = n2042 ^ n2031;
  assign n2034 = n2026 ^ n2012;
  assign n2032 = ~n2003 & n2011;
  assign n2033 = n1986 & n2032;
  assign n2035 = n2034 ^ n2033;
  assign n2018 = n2012 ^ n1996;
  assign n2016 = n1995 & n2003;
  assign n2017 = ~n1986 & n2016;
  assign n2019 = n2018 ^ n2017;
  assign n2036 = n2035 ^ n2019;
  assign n2401 = n1977 & n2036;
  assign n2402 = n2401 ^ x154;
  assign n2398 = n1978 & n2036;
  assign n2396 = n2035 ^ n2029;
  assign n2397 = n1974 & n2396;
  assign n2399 = n2398 ^ n2397;
  assign n2394 = n1969 & n2029;
  assign n2392 = x231 & n2015;
  assign n2020 = n2019 ^ n2015;
  assign n2021 = n1965 & n2020;
  assign n2393 = n2392 ^ n2021;
  assign n2395 = n2394 ^ n2393;
  assign n2400 = n2399 ^ n2395;
  assign n2403 = n2402 ^ n2400;
  assign n2405 = n2404 ^ n2403;
  assign n6573 = n6572 ^ n2405;
  assign n6569 = n6003 & ~n6015;
  assign n6039 = n6027 ^ n6021;
  assign n6040 = ~n5967 & ~n6039;
  assign n6038 = n4448 & n6021;
  assign n6041 = n6040 ^ n6038;
  assign n6570 = n6569 ^ n6041;
  assign n6499 = ~n5974 & n6028;
  assign n6016 = n6015 ^ n6012;
  assign n6033 = ~n5969 & n6016;
  assign n6500 = n6499 ^ n6033;
  assign n6571 = n6570 ^ n6500;
  assign n6574 = n6573 ^ n6571;
  assign n6576 = n6575 ^ n6574;
  assign n8739 = n8738 ^ n6576;
  assign n8735 = n8279 & ~n8329;
  assign n8733 = n8328 ^ n8323;
  assign n8734 = n8267 & ~n8733;
  assign n8736 = n8735 ^ n8734;
  assign n8730 = ~n8271 & ~n8309;
  assign n8314 = n8313 ^ n8309;
  assign n8315 = n8255 & ~n8314;
  assign n8731 = n8730 ^ n8315;
  assign n8729 = ~n8284 & n8323;
  assign n8732 = n8731 ^ n8729;
  assign n8737 = n8736 ^ n8732;
  assign n8740 = n8739 ^ n8737;
  assign n8742 = n8741 ^ n8740;
  assign n2406 = n2405 ^ x186;
  assign n7189 = n6576 ^ n2406;
  assign n10768 = n8742 ^ n7189;
  assign n3986 = n2406 ^ x218;
  assign n8148 = n7189 ^ n3986;
  assign n10769 = n10768 ^ n8148;
  assign n4079 = n3986 ^ x250;
  assign n8149 = n8148 ^ n4079;
  assign n10770 = n10769 ^ n8149;
  assign n8338 = ~n8292 & n8313;
  assign n8330 = n8329 ^ n8324;
  assign n8336 = n8257 & n8330;
  assign n8337 = n8336 ^ n8335;
  assign n8339 = n8338 ^ n8337;
  assign n8331 = ~n8260 & n8330;
  assign n8333 = n8332 ^ n8331;
  assign n8317 = ~n8293 & n8313;
  assign n8316 = n8295 & ~n8314;
  assign n8318 = n8317 ^ n8316;
  assign n8319 = n8318 ^ n8315;
  assign n8334 = n8333 ^ n8319;
  assign n8340 = n8339 ^ n8334;
  assign n6029 = n6028 ^ n6022;
  assign n6481 = ~n5984 & ~n6029;
  assign n6483 = n6482 ^ n6481;
  assign n6419 = ~n5988 & ~n6027;
  assign n6418 = ~n5970 & ~n6039;
  assign n6420 = n6419 ^ n6418;
  assign n6421 = n6420 ^ n6040;
  assign n6607 = n6483 ^ n6421;
  assign n6416 = ~n5990 & ~n6027;
  assign n6030 = n5968 & ~n6029;
  assign n6031 = n6030 ^ n6023;
  assign n6606 = n6416 ^ n6031;
  assign n6608 = n6607 ^ n6606;
  assign n2044 = n2005 & n2019;
  assign n2037 = n2036 ^ n2030;
  assign n2041 = n1987 & n2037;
  assign n2043 = n2042 ^ n2041;
  assign n2045 = n2044 ^ n2043;
  assign n2038 = n1988 & n2037;
  assign n2039 = n2038 ^ n2031;
  assign n2023 = n2006 & n2019;
  assign n2022 = n1998 & n2020;
  assign n2024 = n2023 ^ n2022;
  assign n2025 = n2024 ^ n2021;
  assign n2040 = n2039 ^ n2025;
  assign n2046 = n2045 ^ n2040;
  assign n2047 = n2046 ^ x153;
  assign n6609 = n6608 ^ n2047;
  assign n8341 = n8340 ^ n6609;
  assign n2048 = n2047 ^ x185;
  assign n7184 = n6609 ^ n2048;
  assign n10760 = n8341 ^ n7184;
  assign n3991 = n2048 ^ x217;
  assign n8111 = n7184 ^ n3991;
  assign n10761 = n10760 ^ n8111;
  assign n4086 = n3991 ^ x249;
  assign n8112 = n8111 ^ n4086;
  assign n10762 = n10761 ^ n8112;
  assign n11438 = n10770 ^ n10762;
  assign n8790 = n8282 & n8323;
  assign n8789 = ~n8291 & ~n8328;
  assign n8791 = n8790 ^ n8789;
  assign n8792 = n8791 ^ n8731;
  assign n8786 = ~n8268 & ~n8733;
  assign n8787 = n8786 ^ n8337;
  assign n8788 = n8787 ^ n8734;
  assign n8793 = n8792 ^ n8788;
  assign n6036 = n6004 & ~n6015;
  assign n6035 = ~n5989 & ~n6012;
  assign n6037 = n6036 ^ n6035;
  assign n6042 = n6041 ^ n6037;
  assign n6017 = n5961 & n6016;
  assign n6032 = n6031 ^ n6017;
  assign n6034 = n6033 ^ n6032;
  assign n6043 = n6042 ^ n6034;
  assign n2467 = n1972 & n2029;
  assign n2466 = n2004 & n2035;
  assign n2468 = n2467 ^ n2466;
  assign n2555 = n2468 ^ n2393;
  assign n2524 = n1971 & n2396;
  assign n2525 = n2524 ^ n2043;
  assign n2554 = n2525 ^ n2397;
  assign n2556 = n2555 ^ n2554;
  assign n2557 = n2556 ^ x159;
  assign n6044 = n6043 ^ n2557;
  assign n8794 = n8793 ^ n6044;
  assign n2558 = n2557 ^ x191;
  assign n7179 = n6044 ^ n2558;
  assign n10834 = n8794 ^ n7179;
  assign n3975 = n2558 ^ x223;
  assign n8142 = n7179 ^ n3975;
  assign n10835 = n10834 ^ n8142;
  assign n4088 = n3975 ^ x255;
  assign n8143 = n8142 ^ n4088;
  assign n10836 = n10835 ^ n8143;
  assign n11439 = n11438 ^ n10836;
  assign n8834 = n8736 ^ n8331;
  assign n8928 = n8834 ^ n8791;
  assign n8838 = ~n8273 & ~n8328;
  assign n8927 = n8838 ^ n8337;
  assign n8929 = n8928 ^ n8927;
  assign n6501 = n6500 ^ n6481;
  assign n6502 = n6501 ^ n6037;
  assign n6415 = n5963 & ~n6012;
  assign n6498 = n6415 ^ n6031;
  assign n6503 = n6502 ^ n6498;
  assign n2471 = n1967 & n2035;
  assign n2472 = n2471 ^ n2043;
  assign n2469 = n2399 ^ n2038;
  assign n2470 = n2469 ^ n2468;
  assign n2473 = n2472 ^ n2470;
  assign n2474 = n2473 ^ x158;
  assign n6504 = n6503 ^ n2474;
  assign n8930 = n8929 ^ n6504;
  assign n2475 = n2474 ^ x190;
  assign n7167 = n6504 ^ n2475;
  assign n10777 = n8930 ^ n7167;
  assign n3964 = n2475 ^ x222;
  assign n8125 = n7167 ^ n3964;
  assign n10778 = n10777 ^ n8125;
  assign n4082 = n3964 ^ x254;
  assign n8126 = n8125 ^ n4082;
  assign n10779 = n10778 ^ n8126;
  assign n11459 = n11439 ^ n10779;
  assign n8839 = n8838 ^ n8338;
  assign n8837 = ~n8283 & ~n8309;
  assign n8840 = n8839 ^ n8837;
  assign n8835 = n8834 ^ n8732;
  assign n6642 = n5964 & n6021;
  assign n6417 = n6416 ^ n6415;
  assign n6643 = n6642 ^ n6417;
  assign n6640 = n6570 ^ n6501;
  assign n2578 = n1968 & n2015;
  assign n2487 = n2471 ^ n2044;
  assign n2579 = n2578 ^ n2487;
  assign n2576 = n2469 ^ n2395;
  assign n2575 = n2525 ^ x157;
  assign n2577 = n2576 ^ n2575;
  assign n2580 = n2579 ^ n2577;
  assign n6639 = n6032 ^ n2580;
  assign n6641 = n6640 ^ n6639;
  assign n6644 = n6643 ^ n6641;
  assign n8833 = n8787 ^ n6644;
  assign n8836 = n8835 ^ n8833;
  assign n8841 = n8840 ^ n8836;
  assign n2581 = n2580 ^ x189;
  assign n7198 = n6644 ^ n2581;
  assign n10816 = n8841 ^ n7198;
  assign n3980 = n2581 ^ x221;
  assign n8117 = n7198 ^ n3980;
  assign n10817 = n10816 ^ n8117;
  assign n4080 = n3980 ^ x253;
  assign n8118 = n8117 ^ n4080;
  assign n10818 = n10817 ^ n8118;
  assign n8876 = n8839 ^ n8333;
  assign n8875 = n8787 ^ n8316;
  assign n8877 = n8876 ^ n8875;
  assign n6484 = n6483 ^ n6417;
  assign n6480 = n6418 ^ n6032;
  assign n6485 = n6484 ^ n6480;
  assign n2545 = n2487 ^ n2039;
  assign n2544 = n2525 ^ n2022;
  assign n2546 = n2545 ^ n2544;
  assign n2547 = n2546 ^ x152;
  assign n6486 = n6485 ^ n2547;
  assign n8878 = n8877 ^ n6486;
  assign n2548 = n2547 ^ x184;
  assign n7160 = n6486 ^ n2548;
  assign n10805 = n8878 ^ n7160;
  assign n3955 = n2548 ^ x216;
  assign n8165 = n7160 ^ n3955;
  assign n10806 = n10805 ^ n8165;
  assign n4077 = n3955 ^ x248;
  assign n8166 = n8165 ^ n4077;
  assign n10807 = n10806 ^ n8166;
  assign n11449 = n10818 ^ n10807;
  assign n11460 = n11459 ^ n11449;
  assign n8909 = n8839 ^ n8319;
  assign n6422 = n6421 ^ n6417;
  assign n2527 = n2487 ^ n2025;
  assign n2526 = n2525 ^ x155;
  assign n2528 = n2527 ^ n2526;
  assign n6414 = n6032 ^ n2528;
  assign n6423 = n6422 ^ n6414;
  assign n8908 = n8787 ^ n6423;
  assign n8910 = n8909 ^ n8908;
  assign n2529 = n2528 ^ x187;
  assign n7155 = n6423 ^ n2529;
  assign n10796 = n8910 ^ n7155;
  assign n3952 = n2529 ^ x219;
  assign n8156 = n7155 ^ n3952;
  assign n10797 = n10796 ^ n8156;
  assign n4076 = n3952 ^ x251;
  assign n8157 = n8156 ^ n4076;
  assign n10798 = n10797 ^ n8157;
  assign n11440 = n11439 ^ n10798;
  assign n11437 = n10807 ^ n10798;
  assign n11481 = n11440 ^ n11437;
  assign n11465 = n10818 ^ n10770;
  assign n8952 = n8790 ^ n8730;
  assign n8950 = n8839 ^ n8318;
  assign n6552 = n6038 ^ n6036;
  assign n6550 = n6420 ^ n6417;
  assign n2490 = n2467 ^ n2392;
  assign n2488 = n2487 ^ n2024;
  assign n2486 = n2043 ^ x156;
  assign n2489 = n2488 ^ n2486;
  assign n2491 = n2490 ^ n2489;
  assign n6549 = n6031 ^ n2491;
  assign n6551 = n6550 ^ n6549;
  assign n6553 = n6552 ^ n6551;
  assign n8949 = n8337 ^ n6553;
  assign n8951 = n8950 ^ n8949;
  assign n8953 = n8952 ^ n8951;
  assign n2492 = n2491 ^ x188;
  assign n7172 = n6553 ^ n2492;
  assign n10788 = n8953 ^ n7172;
  assign n3970 = n2492 ^ x220;
  assign n8134 = n7172 ^ n3970;
  assign n10789 = n10788 ^ n8134;
  assign n4083 = n3970 ^ x252;
  assign n8135 = n8134 ^ n4083;
  assign n10790 = n10789 ^ n8135;
  assign n11442 = n10790 ^ n10779;
  assign n11472 = n11465 ^ n11442;
  assign n11480 = n11472 ^ n11439;
  assign n11485 = n11481 ^ n11480;
  assign n11482 = ~n11480 & ~n11481;
  assign n11445 = n10807 ^ n10779;
  assign n11475 = ~n11445 & n11472;
  assign n11483 = n11482 ^ n11475;
  assign n11454 = n10818 ^ n10762;
  assign n11455 = n11454 ^ n11442;
  assign n11456 = n11437 & n11455;
  assign n11443 = n11442 ^ n11437;
  assign n11450 = n11443 ^ n11438;
  assign n11453 = n11449 & ~n11450;
  assign n11457 = n11456 ^ n11453;
  assign n11484 = n11483 ^ n11457;
  assign n11486 = n11485 ^ n11484;
  assign n11476 = n10779 & ~n11439;
  assign n11477 = n11476 ^ n11475;
  assign n11473 = n11472 ^ n11445;
  assign n11444 = n10818 ^ n10798;
  assign n11466 = n11465 ^ n11437;
  assign n11467 = n11444 & ~n11466;
  assign n11468 = n11467 ^ n11456;
  assign n11474 = n11473 ^ n11468;
  assign n11478 = n11477 ^ n11474;
  assign n11490 = n11486 ^ n11478;
  assign n11464 = n11454 ^ n11443;
  assign n11469 = n11468 ^ n11464;
  assign n11461 = n11443 ^ n10836;
  assign n11462 = n11460 & n11461;
  assign n11446 = n11445 ^ n11444;
  assign n11447 = ~n11443 & ~n11446;
  assign n11463 = n11462 ^ n11447;
  assign n11470 = n11469 ^ n11463;
  assign n11479 = n11470 & ~n11478;
  assign n11502 = n11490 ^ n11479;
  assign n11451 = n11450 ^ n11449;
  assign n11441 = ~n10836 & ~n11440;
  assign n11448 = n11447 ^ n11441;
  assign n11452 = n11451 ^ n11448;
  assign n11458 = n11457 ^ n11452;
  assign n11500 = ~n11458 & ~n11478;
  assign n11501 = ~n11486 & n11500;
  assign n11503 = n11502 ^ n11501;
  assign n11514 = n11460 & ~n11503;
  assign n11497 = n11458 & n11470;
  assign n11498 = n11486 & n11497;
  assign n11471 = n11470 ^ n11458;
  assign n11496 = n11479 ^ n11471;
  assign n11499 = n11498 ^ n11496;
  assign n11504 = n11503 ^ n11499;
  assign n11491 = n11479 ^ n11458;
  assign n11492 = ~n11490 & ~n11491;
  assign n11493 = n11492 ^ n11486;
  assign n11487 = n11486 ^ n11479;
  assign n11488 = ~n11471 & n11487;
  assign n11489 = n11488 ^ n11458;
  assign n11494 = n11493 ^ n11489;
  assign n11505 = n11504 ^ n11494;
  assign n11506 = n11444 & ~n11505;
  assign n11495 = n11437 & ~n11494;
  assign n11507 = n11506 ^ n11495;
  assign n12124 = n11514 ^ n11507;
  assign n12048 = n11455 & ~n11494;
  assign n11936 = ~n11466 & ~n11505;
  assign n12122 = n12048 ^ n11936;
  assign n11510 = n11503 ^ n11493;
  assign n11998 = ~n11443 & ~n11510;
  assign n11511 = ~n11446 & ~n11510;
  assign n11509 = n11461 & ~n11503;
  assign n11512 = n11511 ^ n11509;
  assign n12112 = n11998 ^ n11512;
  assign n12123 = n12122 ^ n12112;
  assign n12125 = n12124 ^ n12123;
  assign n9544 = n8118 ^ n8112;
  assign n9526 = n8135 ^ n8126;
  assign n9545 = n9544 ^ n9526;
  assign n9528 = n8149 ^ n8112;
  assign n9529 = n9528 ^ n8143;
  assign n9525 = n8149 ^ n8118;
  assign n9527 = n9526 ^ n9525;
  assign n9570 = n9529 ^ n9527;
  assign n9532 = n8166 ^ n8157;
  assign n9530 = n9529 ^ n8157;
  assign n9569 = n9532 ^ n9530;
  assign n9574 = n9570 ^ n9569;
  assign n9571 = ~n9569 & ~n9570;
  assign n9535 = n8166 ^ n8126;
  assign n9564 = n9527 & ~n9535;
  assign n9572 = n9571 ^ n9564;
  assign n9546 = n9532 & n9545;
  assign n9539 = n8166 ^ n8118;
  assign n9533 = n9532 ^ n9526;
  assign n9540 = n9533 ^ n9528;
  assign n9543 = n9539 & ~n9540;
  assign n9547 = n9546 ^ n9543;
  assign n9573 = n9572 ^ n9547;
  assign n9575 = n9574 ^ n9573;
  assign n9563 = n8126 & ~n9529;
  assign n9565 = n9564 ^ n9563;
  assign n9561 = n9535 ^ n9527;
  assign n9534 = n8157 ^ n8118;
  assign n9550 = n9532 ^ n9525;
  assign n9551 = n9534 & ~n9550;
  assign n9552 = n9551 ^ n9546;
  assign n9562 = n9561 ^ n9552;
  assign n9566 = n9565 ^ n9562;
  assign n9584 = n9575 ^ n9566;
  assign n9554 = n9533 ^ n8143;
  assign n9555 = n9529 ^ n8126;
  assign n9556 = n9555 ^ n9539;
  assign n9557 = n9554 & n9556;
  assign n9536 = n9535 ^ n9534;
  assign n9537 = ~n9533 & ~n9536;
  assign n9558 = n9557 ^ n9537;
  assign n9549 = n9544 ^ n9533;
  assign n9553 = n9552 ^ n9549;
  assign n9559 = n9558 ^ n9553;
  assign n9567 = n9559 & ~n9566;
  assign n9541 = n9540 ^ n9539;
  assign n9531 = ~n8143 & ~n9530;
  assign n9538 = n9537 ^ n9531;
  assign n9542 = n9541 ^ n9538;
  assign n9548 = n9547 ^ n9542;
  assign n9585 = n9567 ^ n9548;
  assign n9586 = ~n9584 & ~n9585;
  assign n9587 = n9586 ^ n9575;
  assign n9560 = n9559 ^ n9548;
  assign n9579 = n9575 ^ n9567;
  assign n9580 = ~n9560 & n9579;
  assign n9581 = n9580 ^ n9548;
  assign n9588 = n9587 ^ n9581;
  assign n9641 = n9545 & ~n9588;
  assign n9592 = n9584 ^ n9567;
  assign n9590 = ~n9548 & ~n9566;
  assign n9591 = ~n9575 & n9590;
  assign n9593 = n9592 ^ n9591;
  assign n9576 = n9548 & n9559;
  assign n9577 = n9575 & n9576;
  assign n9568 = n9567 ^ n9560;
  assign n9578 = n9577 ^ n9568;
  assign n9594 = n9593 ^ n9578;
  assign n9595 = n9594 ^ n9588;
  assign n9640 = ~n9550 & ~n9595;
  assign n9642 = n9641 ^ n9640;
  assign n9601 = n9593 ^ n9587;
  assign n9604 = ~n9533 & ~n9601;
  assign n9602 = ~n9536 & ~n9601;
  assign n9600 = n9554 & ~n9593;
  assign n9603 = n9602 ^ n9600;
  assign n9605 = n9604 ^ n9603;
  assign n9859 = n9642 ^ n9605;
  assign n9607 = n9556 & ~n9593;
  assign n9596 = n9534 & ~n9595;
  assign n9589 = n9532 & ~n9588;
  assign n9597 = n9596 ^ n9589;
  assign n9858 = n9607 ^ n9597;
  assign n9860 = n9859 ^ n9858;
  assign n4087 = n4086 ^ n4079;
  assign n4089 = n4088 ^ n4087;
  assign n4120 = n4089 ^ n4082;
  assign n4097 = n4080 ^ n4077;
  assign n4121 = n4120 ^ n4097;
  assign n4114 = n4082 & ~n4089;
  assign n4084 = n4083 ^ n4082;
  assign n4081 = n4080 ^ n4079;
  assign n4085 = n4084 ^ n4081;
  assign n4094 = n4082 ^ n4077;
  assign n4095 = n4085 & ~n4094;
  assign n4115 = n4114 ^ n4095;
  assign n4109 = n4080 ^ n4076;
  assign n4078 = n4077 ^ n4076;
  assign n4110 = n4081 ^ n4078;
  assign n4111 = n4109 & ~n4110;
  assign n4101 = n4086 ^ n4080;
  assign n4102 = n4101 ^ n4084;
  assign n4103 = n4078 & n4102;
  assign n4112 = n4111 ^ n4103;
  assign n4108 = n4094 ^ n4085;
  assign n4113 = n4112 ^ n4108;
  assign n4116 = n4115 ^ n4113;
  assign n4098 = n4084 ^ n4078;
  assign n4125 = n4101 ^ n4098;
  assign n4126 = n4125 ^ n4112;
  assign n4122 = n4098 ^ n4088;
  assign n4123 = n4121 & n4122;
  assign n4118 = n4109 ^ n4094;
  assign n4119 = ~n4098 & ~n4118;
  assign n4124 = n4123 ^ n4119;
  assign n4127 = n4126 ^ n4124;
  assign n4128 = ~n4116 & n4127;
  assign n4091 = n4089 ^ n4076;
  assign n4092 = n4091 ^ n4078;
  assign n4090 = n4089 ^ n4085;
  assign n4106 = n4092 ^ n4090;
  assign n4099 = n4098 ^ n4087;
  assign n4100 = n4097 & ~n4099;
  assign n4104 = n4103 ^ n4100;
  assign n4093 = ~n4090 & ~n4092;
  assign n4096 = n4095 ^ n4093;
  assign n4105 = n4104 ^ n4096;
  assign n4107 = n4106 ^ n4105;
  assign n4117 = n4116 ^ n4107;
  assign n4149 = n4128 ^ n4117;
  assign n4131 = n4099 ^ n4097;
  assign n4129 = ~n4088 & ~n4091;
  assign n4130 = n4129 ^ n4119;
  assign n4132 = n4131 ^ n4130;
  assign n4133 = n4132 ^ n4104;
  assign n4147 = ~n4116 & ~n4133;
  assign n4148 = ~n4107 & n4147;
  assign n4150 = n4149 ^ n4148;
  assign n4166 = n4121 & ~n4150;
  assign n4144 = n4127 & n4133;
  assign n4145 = n4107 & n4144;
  assign n4137 = n4133 ^ n4127;
  assign n4143 = n4137 ^ n4128;
  assign n4146 = n4145 ^ n4143;
  assign n4151 = n4150 ^ n4146;
  assign n4138 = n4128 ^ n4107;
  assign n4139 = ~n4137 & n4138;
  assign n4140 = n4139 ^ n4133;
  assign n4134 = n4133 ^ n4128;
  assign n4135 = ~n4117 & ~n4134;
  assign n4136 = n4135 ^ n4107;
  assign n4141 = n4140 ^ n4136;
  assign n4152 = n4151 ^ n4141;
  assign n4153 = n4109 & ~n4152;
  assign n4142 = n4078 & ~n4141;
  assign n4154 = n4153 ^ n4142;
  assign n4795 = n4166 ^ n4154;
  assign n4586 = n4102 & ~n4141;
  assign n4585 = ~n4110 & ~n4152;
  assign n4587 = n4586 ^ n4585;
  assign n4160 = n4150 ^ n4136;
  assign n4163 = ~n4098 & ~n4160;
  assign n4161 = ~n4118 & ~n4160;
  assign n4159 = n4122 & ~n4150;
  assign n4162 = n4161 ^ n4159;
  assign n4164 = n4163 ^ n4162;
  assign n4794 = n4587 ^ n4164;
  assign n4796 = n4795 ^ n4794;
  assign n352 = x254 ^ x252;
  assign n351 = x251 ^ x248;
  assign n353 = n352 ^ n351;
  assign n354 = x250 ^ x249;
  assign n363 = n354 ^ x255;
  assign n397 = ~x254 & n363;
  assign n361 = x253 ^ x250;
  assign n362 = n361 ^ n352;
  assign n368 = x254 ^ x248;
  assign n369 = n362 & n368;
  assign n398 = n397 ^ n369;
  assign n395 = n368 ^ n362;
  assign n349 = x253 ^ x251;
  assign n382 = n361 ^ n351;
  assign n383 = n349 & n382;
  assign n357 = x253 ^ x249;
  assign n358 = n357 ^ n352;
  assign n359 = n351 & n358;
  assign n384 = n383 ^ n359;
  assign n396 = n395 ^ n384;
  assign n399 = n398 ^ n396;
  assign n365 = n363 ^ x251;
  assign n366 = n365 ^ n351;
  assign n364 = n363 ^ n362;
  assign n372 = n366 ^ n364;
  assign n367 = n364 & n366;
  assign n370 = n369 ^ n367;
  assign n350 = x253 ^ x248;
  assign n355 = n354 ^ n353;
  assign n356 = n350 & n355;
  assign n360 = n359 ^ n356;
  assign n371 = n370 ^ n360;
  assign n373 = n372 ^ n371;
  assign n405 = n399 ^ n373;
  assign n381 = n357 ^ n353;
  assign n385 = n384 ^ n381;
  assign n378 = n368 ^ n349;
  assign n379 = n353 & n378;
  assign n374 = n353 ^ x255;
  assign n375 = n363 ^ x254;
  assign n376 = n375 ^ n350;
  assign n377 = n374 & n376;
  assign n380 = n379 ^ n377;
  assign n386 = n385 ^ n380;
  assign n400 = n386 & n399;
  assign n389 = n355 ^ n350;
  assign n387 = x255 & n365;
  assign n388 = n387 ^ n379;
  assign n390 = n389 ^ n388;
  assign n391 = n390 ^ n360;
  assign n412 = n400 ^ n391;
  assign n413 = n405 & n412;
  assign n414 = n413 ^ n373;
  assign n406 = n405 ^ n400;
  assign n403 = n391 & n399;
  assign n404 = ~n373 & n403;
  assign n407 = n406 ^ n404;
  assign n422 = n414 ^ n407;
  assign n867 = n353 & n422;
  assign n423 = n378 & n422;
  assign n421 = n374 & n407;
  assign n424 = n423 ^ n421;
  assign n868 = n867 ^ n424;
  assign n394 = n391 ^ n386;
  assign n409 = n400 ^ n373;
  assign n410 = n394 & n409;
  assign n411 = n410 ^ n391;
  assign n415 = n414 ^ n411;
  assign n840 = n358 & n415;
  assign n401 = n400 ^ n394;
  assign n392 = n386 & ~n391;
  assign n393 = n373 & n392;
  assign n402 = n401 ^ n393;
  assign n408 = n407 ^ n402;
  assign n416 = n415 ^ n408;
  assign n756 = n382 & n416;
  assign n841 = n840 ^ n756;
  assign n913 = n868 ^ n841;
  assign n426 = n376 & n407;
  assign n418 = n351 & n415;
  assign n417 = n349 & n416;
  assign n419 = n418 ^ n417;
  assign n912 = n426 ^ n419;
  assign n914 = n913 ^ n912;
  assign n915 = n914 ^ x145;
  assign n4797 = n4796 ^ n915;
  assign n9861 = n9860 ^ n4797;
  assign n12126 = n12125 ^ n9861;
  assign n3538 = n915 ^ x177;
  assign n4798 = n4797 ^ n3538;
  assign n9862 = n9861 ^ n4798;
  assign n12127 = n12126 ^ n9862;
  assign n3539 = n3538 ^ x209;
  assign n4799 = n4798 ^ n3539;
  assign n9863 = n9862 ^ n4799;
  assign n12128 = n12127 ^ n9863;
  assign n3540 = n3539 ^ x241;
  assign n4800 = n4799 ^ n3540;
  assign n9864 = n9863 ^ n4800;
  assign n13634 = n12128 ^ n9864;
  assign n12049 = n12048 ^ n11495;
  assign n12045 = n11449 & n11504;
  assign n9837 = n9641 ^ n9589;
  assign n9834 = n9539 & n9594;
  assign n4772 = n4586 ^ n4142;
  assign n4769 = n4097 & n4151;
  assign n908 = n840 ^ n418;
  assign n905 = n350 & n408;
  assign n906 = n905 ^ x146;
  assign n902 = n366 & n411;
  assign n431 = x255 & n414;
  assign n901 = n867 ^ n431;
  assign n903 = n902 ^ n901;
  assign n754 = n355 & n408;
  assign n752 = n411 ^ n402;
  assign n753 = n368 & n752;
  assign n755 = n754 ^ n753;
  assign n904 = n903 ^ n755;
  assign n907 = n906 ^ n904;
  assign n909 = n908 ^ n907;
  assign n4770 = n4769 ^ n909;
  assign n4728 = ~n4092 & ~n4140;
  assign n4624 = ~n4088 & n4136;
  assign n4727 = n4624 ^ n4163;
  assign n4729 = n4728 ^ n4727;
  assign n4155 = n4146 ^ n4140;
  assign n4644 = ~n4094 & n4155;
  assign n4643 = ~n4099 & n4151;
  assign n4645 = n4644 ^ n4643;
  assign n4768 = n4729 ^ n4645;
  assign n4771 = n4770 ^ n4768;
  assign n4773 = n4772 ^ n4771;
  assign n9835 = n9834 ^ n4773;
  assign n9800 = ~n9569 & ~n9581;
  assign n9716 = ~n8143 & n9587;
  assign n9770 = n9716 ^ n9604;
  assign n9801 = n9800 ^ n9770;
  assign n9582 = n9581 ^ n9578;
  assign n9702 = ~n9535 & n9582;
  assign n9701 = ~n9540 & n9594;
  assign n9703 = n9702 ^ n9701;
  assign n9833 = n9801 ^ n9703;
  assign n9836 = n9835 ^ n9833;
  assign n9838 = n9837 ^ n9836;
  assign n12046 = n12045 ^ n9838;
  assign n12000 = ~n11481 & ~n11489;
  assign n11519 = ~n10836 & n11493;
  assign n11999 = n11998 ^ n11519;
  assign n12001 = n12000 ^ n11999;
  assign n11938 = n11499 ^ n11489;
  assign n11939 = ~n11445 & n11938;
  assign n11937 = ~n11450 & n11504;
  assign n11940 = n11939 ^ n11937;
  assign n12044 = n12001 ^ n11940;
  assign n12047 = n12046 ^ n12044;
  assign n12050 = n12049 ^ n12047;
  assign n3527 = n909 ^ x178;
  assign n4774 = n4773 ^ n3527;
  assign n9839 = n9838 ^ n4774;
  assign n12051 = n12050 ^ n9839;
  assign n3528 = n3527 ^ x210;
  assign n4775 = n4774 ^ n3528;
  assign n9840 = n9839 ^ n4775;
  assign n12052 = n12051 ^ n9840;
  assign n3529 = n3528 ^ x242;
  assign n4776 = n4775 ^ n3529;
  assign n9841 = n9840 ^ n4776;
  assign n13611 = n12052 ^ n9841;
  assign n14144 = n13634 ^ n13611;
  assign n11934 = n11459 & ~n11499;
  assign n11518 = ~n11480 & ~n11489;
  assign n11935 = n11934 ^ n11518;
  assign n12090 = n11999 ^ n11935;
  assign n11995 = n11472 & n11938;
  assign n11996 = n11995 ^ n11507;
  assign n12089 = n11996 ^ n11939;
  assign n12091 = n12090 ^ n12089;
  assign n9699 = ~n9570 & ~n9581;
  assign n9698 = n9555 & ~n9578;
  assign n9700 = n9699 ^ n9698;
  assign n9771 = n9770 ^ n9700;
  assign n9583 = n9527 & n9582;
  assign n9598 = n9597 ^ n9583;
  assign n9769 = n9702 ^ n9598;
  assign n9772 = n9771 ^ n9769;
  assign n4641 = n4120 & ~n4146;
  assign n4623 = ~n4090 & ~n4140;
  assign n4642 = n4641 ^ n4623;
  assign n4836 = n4727 ^ n4642;
  assign n4156 = n4085 & n4155;
  assign n4157 = n4156 ^ n4154;
  assign n4835 = n4644 ^ n4157;
  assign n4837 = n4836 ^ n4835;
  assign n750 = n375 & n402;
  assign n430 = n364 & n411;
  assign n751 = n750 ^ n430;
  assign n944 = n901 ^ n751;
  assign n837 = n362 & n752;
  assign n838 = n837 ^ n419;
  assign n943 = n838 ^ n753;
  assign n945 = n944 ^ n943;
  assign n946 = n945 ^ x151;
  assign n4838 = n4837 ^ n946;
  assign n9773 = n9772 ^ n4838;
  assign n12092 = n12091 ^ n9773;
  assign n3535 = n946 ^ x183;
  assign n4839 = n4838 ^ n3535;
  assign n9774 = n9773 ^ n4839;
  assign n12093 = n12092 ^ n9774;
  assign n3536 = n3535 ^ x215;
  assign n4840 = n4839 ^ n3536;
  assign n9775 = n9774 ^ n4840;
  assign n12094 = n12093 ^ n9775;
  assign n3537 = n3536 ^ x247;
  assign n4841 = n4840 ^ n3537;
  assign n9776 = n9775 ^ n4841;
  assign n13667 = n12094 ^ n9776;
  assign n14145 = n14144 ^ n13667;
  assign n11513 = ~n11439 & ~n11499;
  assign n11515 = n11514 ^ n11513;
  assign n12113 = n12112 ^ n11515;
  assign n9606 = ~n9529 & ~n9578;
  assign n9608 = n9607 ^ n9606;
  assign n9609 = n9608 ^ n9605;
  assign n4165 = ~n4089 & ~n4146;
  assign n4167 = n4166 ^ n4165;
  assign n4168 = n4167 ^ n4164;
  assign n425 = n363 & n402;
  assign n427 = n426 ^ n425;
  assign n869 = n868 ^ n427;
  assign n866 = n838 ^ x147;
  assign n870 = n869 ^ n866;
  assign n4158 = n4157 ^ n870;
  assign n4169 = n4168 ^ n4158;
  assign n9599 = n9598 ^ n4169;
  assign n9610 = n9609 ^ n9599;
  assign n12111 = n11996 ^ n9610;
  assign n12114 = n12113 ^ n12111;
  assign n3543 = n870 ^ x179;
  assign n4170 = n4169 ^ n3543;
  assign n9611 = n9610 ^ n4170;
  assign n12115 = n12114 ^ n9611;
  assign n3544 = n3543 ^ x211;
  assign n4171 = n4170 ^ n3544;
  assign n9612 = n9611 ^ n4171;
  assign n12116 = n12115 ^ n9612;
  assign n3545 = n3544 ^ x243;
  assign n4172 = n4171 ^ n3545;
  assign n9613 = n9612 ^ n4172;
  assign n13624 = n12116 ^ n9613;
  assign n14155 = n14145 ^ n13624;
  assign n12152 = n12122 ^ n11515;
  assign n12151 = n11996 ^ n11511;
  assign n12153 = n12152 ^ n12151;
  assign n9643 = n9642 ^ n9608;
  assign n9639 = n9602 ^ n9598;
  assign n9644 = n9643 ^ n9639;
  assign n4588 = n4587 ^ n4167;
  assign n4584 = n4161 ^ n4157;
  assign n4589 = n4588 ^ n4584;
  assign n842 = n841 ^ n427;
  assign n839 = n838 ^ n423;
  assign n843 = n842 ^ n839;
  assign n844 = n843 ^ x144;
  assign n4590 = n4589 ^ n844;
  assign n9645 = n9644 ^ n4590;
  assign n12154 = n12153 ^ n9645;
  assign n3548 = n844 ^ x176;
  assign n4591 = n4590 ^ n3548;
  assign n9646 = n9645 ^ n4591;
  assign n12155 = n12154 ^ n9646;
  assign n3549 = n3548 ^ x208;
  assign n4592 = n4591 ^ n3549;
  assign n9647 = n9646 ^ n4592;
  assign n12156 = n12155 ^ n9647;
  assign n3550 = n3549 ^ x240;
  assign n4593 = n4592 ^ n3550;
  assign n9648 = n9647 ^ n4593;
  assign n13618 = n12156 ^ n9648;
  assign n14129 = n13624 ^ n13618;
  assign n14156 = n14155 ^ n14129;
  assign n12004 = ~n11440 & n11493;
  assign n12005 = n12004 ^ n11515;
  assign n11941 = n11940 ^ n11936;
  assign n12002 = n12001 ^ n11941;
  assign n9804 = ~n9530 & n9587;
  assign n9805 = n9804 ^ n9608;
  assign n9704 = n9703 ^ n9640;
  assign n9802 = n9801 ^ n9704;
  assign n4732 = ~n4091 & n4136;
  assign n4733 = n4732 ^ n4167;
  assign n4646 = n4645 ^ n4585;
  assign n4730 = n4729 ^ n4646;
  assign n971 = n365 & n414;
  assign n972 = n971 ^ n427;
  assign n757 = n756 ^ n755;
  assign n969 = n903 ^ n757;
  assign n968 = n838 ^ x149;
  assign n970 = n969 ^ n968;
  assign n973 = n972 ^ n970;
  assign n4726 = n4157 ^ n973;
  assign n4731 = n4730 ^ n4726;
  assign n4734 = n4733 ^ n4731;
  assign n9799 = n9598 ^ n4734;
  assign n9803 = n9802 ^ n9799;
  assign n9806 = n9805 ^ n9803;
  assign n11997 = n11996 ^ n9806;
  assign n12003 = n12002 ^ n11997;
  assign n12006 = n12005 ^ n12003;
  assign n3530 = n973 ^ x181;
  assign n4735 = n4734 ^ n3530;
  assign n9807 = n9806 ^ n4735;
  assign n12007 = n12006 ^ n9807;
  assign n3531 = n3530 ^ x213;
  assign n4736 = n4735 ^ n3531;
  assign n9808 = n9807 ^ n4736;
  assign n12008 = n12007 ^ n9808;
  assign n3532 = n3531 ^ x245;
  assign n4737 = n4736 ^ n3532;
  assign n9809 = n9808 ^ n4737;
  assign n13605 = n12008 ^ n9809;
  assign n14133 = n13611 ^ n13605;
  assign n11942 = n11941 ^ n11935;
  assign n11933 = n11513 ^ n11507;
  assign n11943 = n11942 ^ n11933;
  assign n9705 = n9704 ^ n9700;
  assign n9697 = n9606 ^ n9597;
  assign n9706 = n9705 ^ n9697;
  assign n4647 = n4646 ^ n4642;
  assign n4640 = n4165 ^ n4154;
  assign n4648 = n4647 ^ n4640;
  assign n759 = n425 ^ n419;
  assign n758 = n757 ^ n751;
  assign n760 = n759 ^ n758;
  assign n761 = n760 ^ x150;
  assign n4649 = n4648 ^ n761;
  assign n9707 = n9706 ^ n4649;
  assign n11944 = n11943 ^ n9707;
  assign n3523 = n761 ^ x182;
  assign n4650 = n4649 ^ n3523;
  assign n9708 = n9707 ^ n4650;
  assign n11945 = n11944 ^ n9708;
  assign n3524 = n3523 ^ x214;
  assign n4651 = n4650 ^ n3524;
  assign n9709 = n9708 ^ n4651;
  assign n11946 = n11945 ^ n9709;
  assign n3525 = n3524 ^ x246;
  assign n4652 = n4651 ^ n3525;
  assign n9710 = n9709 ^ n4652;
  assign n13643 = n11946 ^ n9710;
  assign n11520 = n11519 ^ n11518;
  assign n11516 = n11515 ^ n11512;
  assign n9717 = n9716 ^ n9699;
  assign n9714 = n9608 ^ n9603;
  assign n4625 = n4624 ^ n4623;
  assign n4621 = n4167 ^ n4162;
  assign n432 = n431 ^ n430;
  assign n428 = n427 ^ n424;
  assign n420 = n419 ^ x148;
  assign n429 = n428 ^ n420;
  assign n433 = n432 ^ n429;
  assign n4620 = n4154 ^ n433;
  assign n4622 = n4621 ^ n4620;
  assign n4626 = n4625 ^ n4622;
  assign n9713 = n9597 ^ n4626;
  assign n9715 = n9714 ^ n9713;
  assign n9718 = n9717 ^ n9715;
  assign n11508 = n11507 ^ n9718;
  assign n11517 = n11516 ^ n11508;
  assign n11521 = n11520 ^ n11517;
  assign n3520 = n433 ^ x180;
  assign n4627 = n4626 ^ n3520;
  assign n9719 = n9718 ^ n4627;
  assign n11522 = n11521 ^ n9719;
  assign n3521 = n3520 ^ x212;
  assign n4628 = n4627 ^ n3521;
  assign n9720 = n9719 ^ n4628;
  assign n11523 = n11522 ^ n9720;
  assign n3522 = n3521 ^ x244;
  assign n4629 = n4628 ^ n3522;
  assign n9721 = n9720 ^ n4629;
  assign n13641 = n11523 ^ n9721;
  assign n14130 = n13643 ^ n13641;
  assign n14141 = n14133 ^ n14130;
  assign n14154 = n14145 ^ n14141;
  assign n14160 = n14156 ^ n14154;
  assign n14157 = ~n14154 & ~n14156;
  assign n14140 = n13643 ^ n13618;
  assign n14147 = ~n14140 & n14141;
  assign n14158 = n14157 ^ n14147;
  assign n14150 = n13618 ^ n13605;
  assign n14131 = n14130 ^ n14129;
  assign n14151 = n14144 ^ n14131;
  assign n14152 = n14150 & ~n14151;
  assign n14136 = n13634 ^ n13605;
  assign n14137 = n14136 ^ n14130;
  assign n14138 = n14129 & n14137;
  assign n14153 = n14152 ^ n14138;
  assign n14159 = n14158 ^ n14153;
  assign n14161 = n14160 ^ n14159;
  assign n14146 = n13643 & ~n14145;
  assign n14148 = n14147 ^ n14146;
  assign n14142 = n14141 ^ n14140;
  assign n14132 = n13624 ^ n13605;
  assign n14134 = n14133 ^ n14129;
  assign n14135 = n14132 & ~n14134;
  assign n14139 = n14138 ^ n14135;
  assign n14143 = n14142 ^ n14139;
  assign n14149 = n14148 ^ n14143;
  assign n14162 = n14161 ^ n14149;
  assign n14175 = n14136 ^ n14131;
  assign n14176 = n14175 ^ n14139;
  assign n14170 = n14145 ^ n13643;
  assign n14171 = n14170 ^ n14150;
  assign n14172 = n14131 ^ n13667;
  assign n14173 = n14171 & n14172;
  assign n14164 = n14140 ^ n14132;
  assign n14165 = ~n14131 & ~n14164;
  assign n14174 = n14173 ^ n14165;
  assign n14177 = n14176 ^ n14174;
  assign n14178 = ~n14149 & n14177;
  assign n14167 = n14151 ^ n14150;
  assign n14163 = ~n13667 & ~n14155;
  assign n14166 = n14165 ^ n14163;
  assign n14168 = n14167 ^ n14166;
  assign n14169 = n14168 ^ n14153;
  assign n14179 = n14178 ^ n14169;
  assign n14180 = ~n14162 & ~n14179;
  assign n14181 = n14180 ^ n14161;
  assign n14392 = ~n14155 & n14181;
  assign n14199 = n14169 & n14177;
  assign n14200 = n14161 & n14199;
  assign n14192 = n14177 ^ n14169;
  assign n14198 = n14192 ^ n14178;
  assign n14201 = n14200 ^ n14198;
  assign n14353 = ~n14145 & ~n14201;
  assign n14184 = n14178 ^ n14162;
  assign n14182 = ~n14149 & ~n14169;
  assign n14183 = ~n14161 & n14182;
  assign n14185 = n14184 ^ n14183;
  assign n14210 = n14171 & ~n14185;
  assign n14391 = n14353 ^ n14210;
  assign n14393 = n14392 ^ n14391;
  assign n14202 = n14201 ^ n14185;
  assign n14272 = ~n14151 & n14202;
  assign n14193 = n14178 ^ n14161;
  assign n14194 = ~n14192 & n14193;
  assign n14195 = n14194 ^ n14169;
  assign n14270 = n14201 ^ n14195;
  assign n14271 = ~n14140 & n14270;
  assign n14273 = n14272 ^ n14271;
  assign n14196 = n14195 ^ n14181;
  assign n14203 = n14202 ^ n14196;
  assign n14204 = ~n14134 & ~n14203;
  assign n14355 = n14273 ^ n14204;
  assign n14268 = ~n14156 & ~n14195;
  assign n14266 = ~n13667 & n14181;
  assign n14186 = n14185 ^ n14181;
  assign n14187 = ~n14131 & ~n14186;
  assign n14267 = n14266 ^ n14187;
  assign n14269 = n14268 ^ n14267;
  assign n14389 = n14355 ^ n14269;
  assign n14291 = n14141 & n14270;
  assign n14208 = n14132 & ~n14203;
  assign n14207 = n14129 & ~n14196;
  assign n14209 = n14208 ^ n14207;
  assign n14292 = n14291 ^ n14209;
  assign n9967 = n9864 ^ n9841;
  assign n9968 = n9967 ^ n9776;
  assign n9969 = n9968 ^ n9613;
  assign n9971 = n9648 ^ n9613;
  assign n10008 = n9971 ^ n9969;
  assign n9965 = n9841 ^ n9809;
  assign n9964 = n9721 ^ n9710;
  assign n9966 = n9965 ^ n9964;
  assign n10007 = n9968 ^ n9966;
  assign n10012 = n10008 ^ n10007;
  assign n10009 = ~n10007 & ~n10008;
  assign n9974 = n9710 ^ n9648;
  assign n10003 = n9966 & ~n9974;
  assign n10010 = n10009 ^ n10003;
  assign n9972 = n9971 ^ n9964;
  assign n9978 = n9972 ^ n9967;
  assign n9979 = n9809 ^ n9648;
  assign n9985 = ~n9978 & n9979;
  assign n9982 = n9864 ^ n9809;
  assign n9983 = n9982 ^ n9964;
  assign n9984 = n9971 & n9983;
  assign n9986 = n9985 ^ n9984;
  assign n10011 = n10010 ^ n9986;
  assign n10013 = n10012 ^ n10011;
  assign n10002 = n9710 & ~n9968;
  assign n10004 = n10003 ^ n10002;
  assign n10000 = n9974 ^ n9966;
  assign n9973 = n9809 ^ n9613;
  assign n9994 = n9971 ^ n9965;
  assign n9995 = n9973 & ~n9994;
  assign n9996 = n9995 ^ n9984;
  assign n10001 = n10000 ^ n9996;
  assign n10005 = n10004 ^ n10001;
  assign n10023 = n10013 ^ n10005;
  assign n9993 = n9982 ^ n9972;
  assign n9997 = n9996 ^ n9993;
  assign n9988 = n9968 ^ n9710;
  assign n9989 = n9988 ^ n9979;
  assign n9990 = n9972 ^ n9776;
  assign n9991 = n9989 & n9990;
  assign n9975 = n9974 ^ n9973;
  assign n9976 = ~n9972 & ~n9975;
  assign n9992 = n9991 ^ n9976;
  assign n9998 = n9997 ^ n9992;
  assign n10006 = n9998 & ~n10005;
  assign n9980 = n9979 ^ n9978;
  assign n9970 = ~n9776 & ~n9969;
  assign n9977 = n9976 ^ n9970;
  assign n9981 = n9980 ^ n9977;
  assign n9987 = n9986 ^ n9981;
  assign n10024 = n10006 ^ n9987;
  assign n10025 = ~n10023 & ~n10024;
  assign n10026 = n10025 ^ n10013;
  assign n10287 = ~n9969 & n10026;
  assign n10031 = n10023 ^ n10006;
  assign n10029 = ~n9987 & ~n10005;
  assign n10030 = ~n10013 & n10029;
  assign n10032 = n10031 ^ n10030;
  assign n10040 = n9989 & ~n10032;
  assign n10018 = n9987 & n9998;
  assign n10019 = n10013 & n10018;
  assign n9999 = n9998 ^ n9987;
  assign n10017 = n10006 ^ n9999;
  assign n10020 = n10019 ^ n10017;
  assign n10039 = ~n9968 & ~n10020;
  assign n10041 = n10040 ^ n10039;
  assign n10288 = n10287 ^ n10041;
  assign n10014 = n10013 ^ n10006;
  assign n10015 = ~n9999 & n10014;
  assign n10016 = n10015 ^ n9987;
  assign n10232 = ~n10008 & ~n10016;
  assign n10096 = ~n9776 & n10026;
  assign n10042 = n10032 ^ n10026;
  assign n10043 = ~n9972 & ~n10042;
  assign n10199 = n10096 ^ n10043;
  assign n10233 = n10232 ^ n10199;
  assign n10033 = n10032 ^ n10020;
  assign n10149 = ~n9978 & n10033;
  assign n10021 = n10020 ^ n10016;
  assign n10148 = ~n9974 & n10021;
  assign n10150 = n10149 ^ n10148;
  assign n10027 = n10026 ^ n10016;
  assign n10034 = n10033 ^ n10027;
  assign n10076 = ~n9994 & ~n10034;
  assign n10151 = n10150 ^ n10076;
  assign n10285 = n10233 ^ n10151;
  assign n10035 = n9973 & ~n10034;
  assign n10028 = n9971 & ~n10027;
  assign n10036 = n10035 ^ n10028;
  assign n10022 = n9966 & n10021;
  assign n10037 = n10036 ^ n10022;
  assign n7692 = n4800 ^ n4776;
  assign n7693 = n7692 ^ n4841;
  assign n7694 = n7693 ^ n4172;
  assign n7696 = n4593 ^ n4172;
  assign n7733 = n7696 ^ n7694;
  assign n7690 = n4776 ^ n4737;
  assign n7689 = n4652 ^ n4629;
  assign n7691 = n7690 ^ n7689;
  assign n7732 = n7693 ^ n7691;
  assign n7737 = n7733 ^ n7732;
  assign n7734 = ~n7732 & ~n7733;
  assign n7699 = n4652 ^ n4593;
  assign n7728 = n7691 & ~n7699;
  assign n7735 = n7734 ^ n7728;
  assign n7697 = n7696 ^ n7689;
  assign n7703 = n7697 ^ n7692;
  assign n7704 = n4737 ^ n4593;
  assign n7710 = ~n7703 & n7704;
  assign n7707 = n4800 ^ n4737;
  assign n7708 = n7707 ^ n7689;
  assign n7709 = n7696 & n7708;
  assign n7711 = n7710 ^ n7709;
  assign n7736 = n7735 ^ n7711;
  assign n7738 = n7737 ^ n7736;
  assign n7727 = n4652 & ~n7693;
  assign n7729 = n7728 ^ n7727;
  assign n7725 = n7699 ^ n7691;
  assign n7698 = n4737 ^ n4172;
  assign n7719 = n7696 ^ n7690;
  assign n7720 = n7698 & ~n7719;
  assign n7721 = n7720 ^ n7709;
  assign n7726 = n7725 ^ n7721;
  assign n7730 = n7729 ^ n7726;
  assign n7748 = n7738 ^ n7730;
  assign n7718 = n7707 ^ n7697;
  assign n7722 = n7721 ^ n7718;
  assign n7713 = n7697 ^ n4841;
  assign n7714 = n7693 ^ n4652;
  assign n7715 = n7714 ^ n7704;
  assign n7716 = n7713 & n7715;
  assign n7700 = n7699 ^ n7698;
  assign n7701 = ~n7697 & ~n7700;
  assign n7717 = n7716 ^ n7701;
  assign n7723 = n7722 ^ n7717;
  assign n7731 = n7723 & ~n7730;
  assign n7705 = n7704 ^ n7703;
  assign n7695 = ~n4841 & ~n7694;
  assign n7702 = n7701 ^ n7695;
  assign n7706 = n7705 ^ n7702;
  assign n7712 = n7711 ^ n7706;
  assign n7749 = n7731 ^ n7712;
  assign n7750 = ~n7748 & ~n7749;
  assign n7751 = n7750 ^ n7738;
  assign n7910 = ~n7694 & n7751;
  assign n7756 = n7748 ^ n7731;
  assign n7754 = ~n7712 & ~n7730;
  assign n7755 = ~n7738 & n7754;
  assign n7757 = n7756 ^ n7755;
  assign n7765 = n7715 & ~n7757;
  assign n7743 = n7712 & n7723;
  assign n7744 = n7738 & n7743;
  assign n7724 = n7723 ^ n7712;
  assign n7742 = n7731 ^ n7724;
  assign n7745 = n7744 ^ n7742;
  assign n7764 = ~n7693 & ~n7745;
  assign n7766 = n7765 ^ n7764;
  assign n7911 = n7910 ^ n7766;
  assign n7739 = n7738 ^ n7731;
  assign n7740 = ~n7724 & n7739;
  assign n7741 = n7740 ^ n7712;
  assign n7746 = n7745 ^ n7741;
  assign n7855 = ~n7699 & n7746;
  assign n7758 = n7757 ^ n7745;
  assign n7854 = ~n7703 & n7758;
  assign n7856 = n7855 ^ n7854;
  assign n7752 = n7751 ^ n7741;
  assign n7759 = n7758 ^ n7752;
  assign n7803 = ~n7719 & ~n7759;
  assign n7907 = n7856 ^ n7803;
  assign n7859 = ~n7733 & ~n7741;
  assign n7857 = ~n4841 & n7751;
  assign n7768 = n7757 ^ n7751;
  assign n7771 = ~n7697 & ~n7768;
  assign n7858 = n7857 ^ n7771;
  assign n7860 = n7859 ^ n7858;
  assign n7908 = n7907 ^ n7860;
  assign n7760 = n7698 & ~n7759;
  assign n7753 = n7696 & ~n7752;
  assign n7761 = n7760 ^ n7753;
  assign n7747 = n7691 & n7746;
  assign n7762 = n7761 ^ n7747;
  assign n3541 = n3540 ^ n3529;
  assign n3542 = n3541 ^ n3537;
  assign n3546 = n3545 ^ n3542;
  assign n3551 = n3550 ^ n3545;
  assign n3588 = n3551 ^ n3546;
  assign n3533 = n3532 ^ n3529;
  assign n3526 = n3525 ^ n3522;
  assign n3534 = n3533 ^ n3526;
  assign n3587 = n3542 ^ n3534;
  assign n3592 = n3588 ^ n3587;
  assign n3589 = ~n3587 & ~n3588;
  assign n3554 = n3550 ^ n3525;
  assign n3583 = n3534 & ~n3554;
  assign n3590 = n3589 ^ n3583;
  assign n3552 = n3551 ^ n3526;
  assign n3558 = n3552 ^ n3541;
  assign n3559 = n3550 ^ n3532;
  assign n3565 = ~n3558 & n3559;
  assign n3562 = n3540 ^ n3532;
  assign n3563 = n3562 ^ n3526;
  assign n3564 = n3551 & n3563;
  assign n3566 = n3565 ^ n3564;
  assign n3591 = n3590 ^ n3566;
  assign n3593 = n3592 ^ n3591;
  assign n3582 = n3525 & ~n3542;
  assign n3584 = n3583 ^ n3582;
  assign n3580 = n3554 ^ n3534;
  assign n3553 = n3545 ^ n3532;
  assign n3574 = n3551 ^ n3533;
  assign n3575 = n3553 & ~n3574;
  assign n3576 = n3575 ^ n3564;
  assign n3581 = n3580 ^ n3576;
  assign n3585 = n3584 ^ n3581;
  assign n3603 = n3593 ^ n3585;
  assign n3573 = n3562 ^ n3552;
  assign n3577 = n3576 ^ n3573;
  assign n3568 = n3542 ^ n3525;
  assign n3569 = n3568 ^ n3559;
  assign n3570 = n3552 ^ n3537;
  assign n3571 = n3569 & n3570;
  assign n3555 = n3554 ^ n3553;
  assign n3556 = ~n3552 & ~n3555;
  assign n3572 = n3571 ^ n3556;
  assign n3578 = n3577 ^ n3572;
  assign n3586 = n3578 & ~n3585;
  assign n3560 = n3559 ^ n3558;
  assign n3547 = ~n3537 & ~n3546;
  assign n3557 = n3556 ^ n3547;
  assign n3561 = n3560 ^ n3557;
  assign n3567 = n3566 ^ n3561;
  assign n3604 = n3586 ^ n3567;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = n3605 ^ n3593;
  assign n3635 = ~n3546 & n3606;
  assign n3611 = n3603 ^ n3586;
  assign n3609 = ~n3567 & ~n3585;
  assign n3610 = ~n3593 & n3609;
  assign n3612 = n3611 ^ n3610;
  assign n3633 = n3569 & ~n3612;
  assign n3598 = n3567 & n3578;
  assign n3599 = n3593 & n3598;
  assign n3579 = n3578 ^ n3567;
  assign n3597 = n3586 ^ n3579;
  assign n3600 = n3599 ^ n3597;
  assign n3632 = ~n3542 & ~n3600;
  assign n3634 = n3633 ^ n3632;
  assign n3636 = n3635 ^ n3634;
  assign n3594 = n3593 ^ n3586;
  assign n3595 = ~n3579 & n3594;
  assign n3596 = n3595 ^ n3567;
  assign n3628 = ~n3588 & ~n3596;
  assign n3625 = n3612 ^ n3606;
  assign n3626 = ~n3552 & ~n3625;
  assign n3624 = ~n3537 & n3606;
  assign n3627 = n3626 ^ n3624;
  assign n3629 = n3628 ^ n3627;
  assign n3613 = n3612 ^ n3600;
  assign n3607 = n3606 ^ n3596;
  assign n3614 = n3613 ^ n3607;
  assign n3622 = ~n3574 & ~n3614;
  assign n3601 = n3600 ^ n3596;
  assign n3620 = ~n3554 & n3601;
  assign n3619 = ~n3558 & n3613;
  assign n3621 = n3620 ^ n3619;
  assign n3623 = n3622 ^ n3621;
  assign n3630 = n3629 ^ n3623;
  assign n3615 = n3553 & ~n3614;
  assign n3608 = n3551 & ~n3607;
  assign n3616 = n3615 ^ n3608;
  assign n3602 = n3534 & n3601;
  assign n3617 = n3616 ^ n3602;
  assign n3618 = n3617 ^ n1789;
  assign n3631 = n3630 ^ n3618;
  assign n3637 = n3636 ^ n3631;
  assign n7906 = n7762 ^ n3637;
  assign n7909 = n7908 ^ n7906;
  assign n7912 = n7911 ^ n7909;
  assign n10284 = n10037 ^ n7912;
  assign n10286 = n10285 ^ n10284;
  assign n10289 = n10288 ^ n10286;
  assign n14388 = n14292 ^ n10289;
  assign n14390 = n14389 ^ n14388;
  assign n14394 = n14393 ^ n14390;
  assign n3638 = n3637 ^ n1790;
  assign n7913 = n7912 ^ n3638;
  assign n10290 = n10289 ^ n7913;
  assign n14395 = n14394 ^ n10290;
  assign n3639 = n3638 ^ n1791;
  assign n7914 = n7913 ^ n3639;
  assign n13177 = n10290 ^ n7914;
  assign n16848 = n14395 ^ n13177;
  assign n6741 = n3639 ^ n1792;
  assign n10920 = n7914 ^ n6741;
  assign n13178 = n13177 ^ n10920;
  assign n18662 = n16848 ^ n13178;
  assign n14211 = n14210 ^ n14209;
  assign n14197 = n14137 & ~n14196;
  assign n14205 = n14204 ^ n14197;
  assign n14189 = ~n14164 & ~n14186;
  assign n14188 = n14172 & ~n14185;
  assign n14190 = n14189 ^ n14188;
  assign n14191 = n14190 ^ n14187;
  assign n14206 = n14205 ^ n14191;
  assign n14212 = n14211 ^ n14206;
  assign n10258 = n10040 ^ n10036;
  assign n10077 = n9983 & ~n10027;
  assign n10078 = n10077 ^ n10076;
  assign n10045 = ~n9975 & ~n10042;
  assign n10044 = n9990 & ~n10032;
  assign n10046 = n10045 ^ n10044;
  assign n10047 = n10046 ^ n10043;
  assign n10257 = n10078 ^ n10047;
  assign n10259 = n10258 ^ n10257;
  assign n7802 = n7708 & ~n7752;
  assign n7804 = n7803 ^ n7802;
  assign n7769 = ~n7700 & ~n7768;
  assign n7767 = n7713 & ~n7757;
  assign n7770 = n7769 ^ n7767;
  assign n7772 = n7771 ^ n7770;
  assign n8015 = n7804 ^ n7772;
  assign n8014 = n7765 ^ n7761;
  assign n8016 = n8015 ^ n8014;
  assign n3696 = n3633 ^ n3616;
  assign n3693 = n3563 & ~n3607;
  assign n3694 = n3693 ^ n3622;
  assign n3690 = ~n3555 & ~n3625;
  assign n3689 = n3570 & ~n3612;
  assign n3691 = n3690 ^ n3689;
  assign n3692 = n3691 ^ n3626;
  assign n3695 = n3694 ^ n3692;
  assign n3697 = n3696 ^ n3695;
  assign n3698 = n3697 ^ n1740;
  assign n8017 = n8016 ^ n3698;
  assign n10260 = n10259 ^ n8017;
  assign n14213 = n14212 ^ n10260;
  assign n3699 = n3698 ^ n1741;
  assign n8018 = n8017 ^ n3699;
  assign n10261 = n10260 ^ n8018;
  assign n14214 = n14213 ^ n10261;
  assign n3700 = n3699 ^ n1742;
  assign n8019 = n8018 ^ n3700;
  assign n13199 = n10261 ^ n8019;
  assign n16875 = n14214 ^ n13199;
  assign n6734 = n3700 ^ n1743;
  assign n10935 = n8019 ^ n6734;
  assign n13200 = n13199 ^ n10935;
  assign n18388 = n16875 ^ n13200;
  assign n19226 = n18662 ^ n18388;
  assign n14295 = ~n14154 & ~n14195;
  assign n14424 = n14295 ^ n14266;
  assign n14422 = n14391 ^ n14190;
  assign n10095 = ~n10007 & ~n10016;
  assign n10097 = n10096 ^ n10095;
  assign n10093 = n10046 ^ n10041;
  assign n7925 = ~n7732 & ~n7741;
  assign n7926 = n7925 ^ n7857;
  assign n7923 = n7770 ^ n7766;
  assign n3711 = ~n3587 & ~n3596;
  assign n3712 = n3711 ^ n3624;
  assign n3709 = n3691 ^ n3634;
  assign n3708 = n3616 ^ n1228;
  assign n3710 = n3709 ^ n3708;
  assign n3713 = n3712 ^ n3710;
  assign n7922 = n7761 ^ n3713;
  assign n7924 = n7923 ^ n7922;
  assign n7927 = n7926 ^ n7924;
  assign n10092 = n10036 ^ n7927;
  assign n10094 = n10093 ^ n10092;
  assign n10098 = n10097 ^ n10094;
  assign n14421 = n14209 ^ n10098;
  assign n14423 = n14422 ^ n14421;
  assign n14425 = n14424 ^ n14423;
  assign n3714 = n3713 ^ n1229;
  assign n7928 = n7927 ^ n3714;
  assign n10099 = n10098 ^ n7928;
  assign n14426 = n14425 ^ n10099;
  assign n3715 = n3714 ^ n1230;
  assign n7929 = n7928 ^ n3715;
  assign n13182 = n10099 ^ n7929;
  assign n16836 = n14426 ^ n13182;
  assign n6730 = n3715 ^ n1231;
  assign n10923 = n7929 ^ n6730;
  assign n13183 = n13182 ^ n10923;
  assign n18588 = n16836 ^ n13183;
  assign n14294 = n14170 & ~n14201;
  assign n14296 = n14295 ^ n14294;
  assign n14356 = n14355 ^ n14296;
  assign n14354 = n14353 ^ n14209;
  assign n14357 = n14356 ^ n14354;
  assign n10146 = n9988 & ~n10020;
  assign n10147 = n10146 ^ n10095;
  assign n10152 = n10151 ^ n10147;
  assign n10145 = n10039 ^ n10036;
  assign n10153 = n10152 ^ n10145;
  assign n7955 = n7714 & ~n7745;
  assign n7956 = n7955 ^ n7925;
  assign n7957 = n7956 ^ n7907;
  assign n7954 = n7764 ^ n7761;
  assign n7958 = n7957 ^ n7954;
  assign n3752 = n3568 & ~n3600;
  assign n3753 = n3752 ^ n3711;
  assign n3754 = n3753 ^ n3623;
  assign n3751 = n3632 ^ n3616;
  assign n3755 = n3754 ^ n3751;
  assign n3756 = n3755 ^ n1255;
  assign n7959 = n7958 ^ n3756;
  assign n10154 = n10153 ^ n7959;
  assign n14358 = n14357 ^ n10154;
  assign n3757 = n3756 ^ n1256;
  assign n7960 = n7959 ^ n3757;
  assign n10155 = n10154 ^ n7960;
  assign n14359 = n14358 ^ n10155;
  assign n3758 = n3757 ^ n1257;
  assign n7961 = n7960 ^ n3758;
  assign n13180 = n10155 ^ n7961;
  assign n16833 = n14359 ^ n13180;
  assign n6729 = n3758 ^ n1258;
  assign n10922 = n7961 ^ n6729;
  assign n13181 = n13180 ^ n10922;
  assign n18573 = n16833 ^ n13181;
  assign n19221 = n18588 ^ n18573;
  assign n19227 = n19226 ^ n19221;
  assign n14278 = n14207 ^ n14197;
  assign n14275 = n14150 & n14202;
  assign n10238 = n10077 ^ n10028;
  assign n10235 = n9979 & n10033;
  assign n7865 = n7802 ^ n7753;
  assign n7862 = n7704 & n7758;
  assign n3843 = n3693 ^ n3608;
  assign n3840 = n3559 & n3613;
  assign n3841 = n3840 ^ n1717;
  assign n3839 = n3629 ^ n3621;
  assign n3842 = n3841 ^ n3839;
  assign n3844 = n3843 ^ n3842;
  assign n7863 = n7862 ^ n3844;
  assign n7861 = n7860 ^ n7856;
  assign n7864 = n7863 ^ n7861;
  assign n7866 = n7865 ^ n7864;
  assign n10236 = n10235 ^ n7866;
  assign n10234 = n10233 ^ n10150;
  assign n10237 = n10236 ^ n10234;
  assign n10239 = n10238 ^ n10237;
  assign n14276 = n14275 ^ n10239;
  assign n14274 = n14273 ^ n14269;
  assign n14277 = n14276 ^ n14274;
  assign n14279 = n14278 ^ n14277;
  assign n3845 = n3844 ^ n1718;
  assign n7867 = n7866 ^ n3845;
  assign n10240 = n10239 ^ n7867;
  assign n14280 = n14279 ^ n10240;
  assign n3846 = n3845 ^ n1719;
  assign n7868 = n7867 ^ n3846;
  assign n13175 = n10240 ^ n7868;
  assign n16853 = n14280 ^ n13175;
  assign n6733 = n3846 ^ n1720;
  assign n10919 = n7868 ^ n6733;
  assign n13176 = n13175 ^ n10919;
  assign n18457 = n16853 ^ n13176;
  assign n19223 = n18457 ^ n18388;
  assign n14297 = n14296 ^ n14267;
  assign n14293 = n14292 ^ n14271;
  assign n14298 = n14297 ^ n14293;
  assign n10200 = n10199 ^ n10147;
  assign n10198 = n10148 ^ n10037;
  assign n10201 = n10200 ^ n10198;
  assign n7992 = n7956 ^ n7858;
  assign n7991 = n7855 ^ n7762;
  assign n7993 = n7992 ^ n7991;
  assign n3786 = n3753 ^ n3627;
  assign n3785 = n3620 ^ n3617;
  assign n3787 = n3786 ^ n3785;
  assign n3788 = n3787 ^ n1753;
  assign n7994 = n7993 ^ n3788;
  assign n10202 = n10201 ^ n7994;
  assign n14299 = n14298 ^ n10202;
  assign n3789 = n3788 ^ n1754;
  assign n7995 = n7994 ^ n3789;
  assign n10203 = n10202 ^ n7995;
  assign n14300 = n14299 ^ n10203;
  assign n3790 = n3789 ^ n1755;
  assign n7996 = n7995 ^ n3790;
  assign n13197 = n10203 ^ n7996;
  assign n16884 = n14300 ^ n13197;
  assign n6737 = n3790 ^ n1756;
  assign n10937 = n7996 ^ n6737;
  assign n13198 = n13197 ^ n10937;
  assign n18505 = n16884 ^ n13198;
  assign n19232 = n19223 ^ n18505;
  assign n19266 = ~n18573 & n19232;
  assign n14410 = n14391 ^ n14205;
  assign n14409 = n14292 ^ n14189;
  assign n14411 = n14410 ^ n14409;
  assign n10079 = n10078 ^ n10041;
  assign n10075 = n10045 ^ n10037;
  assign n10080 = n10079 ^ n10075;
  assign n7805 = n7804 ^ n7766;
  assign n7801 = n7769 ^ n7762;
  assign n7806 = n7805 ^ n7801;
  assign n3856 = n3694 ^ n3634;
  assign n3855 = n3690 ^ n3617;
  assign n3857 = n3856 ^ n3855;
  assign n3858 = n3857 ^ n1659;
  assign n7807 = n7806 ^ n3858;
  assign n10081 = n10080 ^ n7807;
  assign n14412 = n14411 ^ n10081;
  assign n3859 = n3858 ^ n1660;
  assign n7808 = n7807 ^ n3859;
  assign n10082 = n10081 ^ n7808;
  assign n14413 = n14412 ^ n10082;
  assign n3860 = n3859 ^ n1661;
  assign n7809 = n7808 ^ n3860;
  assign n13186 = n10082 ^ n7809;
  assign n16860 = n14413 ^ n13186;
  assign n6726 = n3860 ^ n1662;
  assign n10926 = n7809 ^ n6726;
  assign n13187 = n13186 ^ n10926;
  assign n18631 = n16860 ^ n13187;
  assign n19218 = n18631 ^ n18573;
  assign n19230 = n18662 ^ n18457;
  assign n19231 = n19230 ^ n19221;
  assign n19237 = n19218 & n19231;
  assign n19267 = n19266 ^ n19237;
  assign n19264 = n19231 ^ n19218;
  assign n14463 = n14391 ^ n14191;
  assign n10048 = n10047 ^ n10041;
  assign n7773 = n7772 ^ n7766;
  assign n3817 = n3692 ^ n3634;
  assign n3816 = n3617 ^ n1644;
  assign n3818 = n3817 ^ n3816;
  assign n7763 = n7762 ^ n3818;
  assign n7774 = n7773 ^ n7763;
  assign n10038 = n10037 ^ n7774;
  assign n10049 = n10048 ^ n10038;
  assign n14462 = n14292 ^ n10049;
  assign n14464 = n14463 ^ n14462;
  assign n3819 = n3818 ^ n1645;
  assign n7775 = n7774 ^ n3819;
  assign n10050 = n10049 ^ n7775;
  assign n14465 = n14464 ^ n10050;
  assign n3820 = n3819 ^ n1646;
  assign n7776 = n7775 ^ n3820;
  assign n13188 = n10050 ^ n7776;
  assign n16868 = n14465 ^ n13188;
  assign n6727 = n3820 ^ n1647;
  assign n10927 = n7776 ^ n6727;
  assign n13189 = n13188 ^ n10927;
  assign n18540 = n16868 ^ n13189;
  assign n19246 = n18662 ^ n18540;
  assign n19220 = n18631 ^ n18540;
  assign n19251 = n19230 ^ n19220;
  assign n19252 = n19246 & n19251;
  assign n19228 = n19220 & n19227;
  assign n19253 = n19252 ^ n19228;
  assign n19265 = n19264 ^ n19253;
  assign n19268 = n19267 ^ n19265;
  assign n19234 = n19232 ^ n18540;
  assign n19235 = n19234 ^ n19220;
  assign n19233 = n19232 ^ n19231;
  assign n19240 = n19235 ^ n19233;
  assign n19236 = n19233 & n19235;
  assign n19238 = n19237 ^ n19236;
  assign n19219 = n18662 ^ n18631;
  assign n19222 = n19221 ^ n19220;
  assign n19224 = n19223 ^ n19222;
  assign n19225 = n19219 & n19224;
  assign n19229 = n19228 ^ n19225;
  assign n19239 = n19238 ^ n19229;
  assign n19241 = n19240 ^ n19239;
  assign n19279 = n19268 ^ n19241;
  assign n19250 = n19226 ^ n19222;
  assign n19254 = n19253 ^ n19250;
  assign n19247 = n19246 ^ n19218;
  assign n19248 = n19222 & n19247;
  assign n19242 = n19232 ^ n18573;
  assign n19243 = n19242 ^ n19219;
  assign n19244 = n19222 ^ n18505;
  assign n19245 = n19243 & n19244;
  assign n19249 = n19248 ^ n19245;
  assign n19255 = n19254 ^ n19249;
  assign n19269 = n19255 & n19268;
  assign n19258 = n19224 ^ n19219;
  assign n19256 = n18505 & n19234;
  assign n19257 = n19256 ^ n19248;
  assign n19259 = n19258 ^ n19257;
  assign n19260 = n19259 ^ n19229;
  assign n19285 = n19269 ^ n19260;
  assign n19286 = n19279 & n19285;
  assign n19287 = n19286 ^ n19241;
  assign n19263 = n19260 ^ n19255;
  assign n19272 = n19269 ^ n19241;
  assign n19273 = n19263 & n19272;
  assign n19274 = n19273 ^ n19260;
  assign n19298 = n19287 ^ n19274;
  assign n19300 = n19227 & n19298;
  assign n19299 = n19220 & n19298;
  assign n19301 = n19300 ^ n19299;
  assign n19280 = n19279 ^ n19269;
  assign n19277 = n19260 & n19268;
  assign n19278 = ~n19241 & n19277;
  assign n19281 = n19280 ^ n19278;
  assign n19270 = n19269 ^ n19263;
  assign n19261 = n19255 & ~n19260;
  assign n19262 = n19241 & n19261;
  assign n19271 = n19270 ^ n19262;
  assign n19282 = n19281 ^ n19271;
  assign n19295 = n19219 & n19282;
  assign n13208 = n13200 ^ n13178;
  assign n13184 = n13183 ^ n13181;
  assign n13210 = n13208 ^ n13184;
  assign n13201 = n13200 ^ n13176;
  assign n13202 = n13201 ^ n13198;
  assign n13224 = n13202 ^ n13189;
  assign n13190 = n13189 ^ n13187;
  assign n13236 = n13224 ^ n13190;
  assign n13179 = n13178 ^ n13176;
  assign n13185 = n13184 ^ n13179;
  assign n13235 = n13202 ^ n13185;
  assign n13240 = n13236 ^ n13235;
  assign n13237 = ~n13235 & ~n13236;
  assign n13192 = n13187 ^ n13181;
  assign n13220 = n13185 & ~n13192;
  assign n13238 = n13237 ^ n13220;
  assign n13196 = n13187 ^ n13178;
  assign n13191 = n13190 ^ n13184;
  assign n13227 = n13201 ^ n13191;
  assign n13230 = n13196 & ~n13227;
  assign n13211 = n13190 & n13210;
  assign n13231 = n13230 ^ n13211;
  assign n13239 = n13238 ^ n13231;
  assign n13241 = n13240 ^ n13239;
  assign n13219 = n13181 & ~n13202;
  assign n13221 = n13220 ^ n13219;
  assign n13217 = n13192 ^ n13185;
  assign n13193 = n13189 ^ n13178;
  assign n13212 = n13190 ^ n13179;
  assign n13213 = n13193 & ~n13212;
  assign n13214 = n13213 ^ n13211;
  assign n13218 = n13217 ^ n13214;
  assign n13222 = n13221 ^ n13218;
  assign n13252 = n13241 ^ n13222;
  assign n13228 = n13227 ^ n13196;
  assign n13225 = ~n13198 & ~n13224;
  assign n13194 = n13193 ^ n13192;
  assign n13195 = ~n13191 & ~n13194;
  assign n13226 = n13225 ^ n13195;
  assign n13229 = n13228 ^ n13226;
  assign n13232 = n13231 ^ n13229;
  assign n13209 = n13208 ^ n13191;
  assign n13215 = n13214 ^ n13209;
  assign n13203 = n13202 ^ n13181;
  assign n13204 = n13203 ^ n13196;
  assign n13205 = n13198 ^ n13191;
  assign n13206 = n13204 & n13205;
  assign n13207 = n13206 ^ n13195;
  assign n13216 = n13215 ^ n13207;
  assign n13223 = n13216 & ~n13222;
  assign n13256 = n13232 ^ n13223;
  assign n13257 = ~n13252 & ~n13256;
  assign n13258 = n13257 ^ n13241;
  assign n13233 = n13232 ^ n13216;
  assign n13245 = n13241 ^ n13223;
  assign n13246 = ~n13233 & n13245;
  assign n13247 = n13246 ^ n13232;
  assign n13259 = n13258 ^ n13247;
  assign n13272 = n13210 & ~n13259;
  assign n13262 = n13190 & ~n13259;
  assign n13497 = n13272 ^ n13262;
  assign n13253 = n13252 ^ n13223;
  assign n13250 = ~n13222 & ~n13232;
  assign n13251 = ~n13241 & n13250;
  assign n13254 = n13253 ^ n13251;
  assign n13242 = n13216 & n13232;
  assign n13243 = n13241 & n13242;
  assign n13234 = n13233 ^ n13223;
  assign n13244 = n13243 ^ n13234;
  assign n13255 = n13254 ^ n13244;
  assign n13494 = n13196 & n13255;
  assign n10944 = n10935 ^ n10920;
  assign n10924 = n10923 ^ n10922;
  assign n10946 = n10944 ^ n10924;
  assign n10936 = n10935 ^ n10919;
  assign n10938 = n10937 ^ n10936;
  assign n10960 = n10938 ^ n10927;
  assign n10928 = n10927 ^ n10926;
  assign n10972 = n10960 ^ n10928;
  assign n10921 = n10920 ^ n10919;
  assign n10925 = n10924 ^ n10921;
  assign n10971 = n10938 ^ n10925;
  assign n10976 = n10972 ^ n10971;
  assign n10973 = ~n10971 & ~n10972;
  assign n10930 = n10926 ^ n10922;
  assign n10956 = n10925 & ~n10930;
  assign n10974 = n10973 ^ n10956;
  assign n10934 = n10926 ^ n10920;
  assign n10929 = n10928 ^ n10924;
  assign n10963 = n10936 ^ n10929;
  assign n10966 = n10934 & ~n10963;
  assign n10947 = n10928 & n10946;
  assign n10967 = n10966 ^ n10947;
  assign n10975 = n10974 ^ n10967;
  assign n10977 = n10976 ^ n10975;
  assign n10955 = n10922 & ~n10938;
  assign n10957 = n10956 ^ n10955;
  assign n10953 = n10930 ^ n10925;
  assign n10931 = n10927 ^ n10920;
  assign n10948 = n10928 ^ n10921;
  assign n10949 = n10931 & ~n10948;
  assign n10950 = n10949 ^ n10947;
  assign n10954 = n10953 ^ n10950;
  assign n10958 = n10957 ^ n10954;
  assign n10988 = n10977 ^ n10958;
  assign n10964 = n10963 ^ n10934;
  assign n10961 = ~n10937 & ~n10960;
  assign n10932 = n10931 ^ n10930;
  assign n10933 = ~n10929 & ~n10932;
  assign n10962 = n10961 ^ n10933;
  assign n10965 = n10964 ^ n10962;
  assign n10968 = n10967 ^ n10965;
  assign n10945 = n10944 ^ n10929;
  assign n10951 = n10950 ^ n10945;
  assign n10939 = n10938 ^ n10922;
  assign n10940 = n10939 ^ n10934;
  assign n10941 = n10937 ^ n10929;
  assign n10942 = n10940 & n10941;
  assign n10943 = n10942 ^ n10933;
  assign n10952 = n10951 ^ n10943;
  assign n10959 = n10952 & ~n10958;
  assign n10992 = n10968 ^ n10959;
  assign n10993 = ~n10988 & ~n10992;
  assign n10994 = n10993 ^ n10977;
  assign n10969 = n10968 ^ n10952;
  assign n10981 = n10977 ^ n10959;
  assign n10982 = ~n10969 & n10981;
  assign n10983 = n10982 ^ n10968;
  assign n10995 = n10994 ^ n10983;
  assign n11066 = n10946 & ~n10995;
  assign n10998 = n10928 & ~n10995;
  assign n11067 = n11066 ^ n10998;
  assign n10989 = n10988 ^ n10959;
  assign n10986 = ~n10958 & ~n10968;
  assign n10987 = ~n10977 & n10986;
  assign n10990 = n10989 ^ n10987;
  assign n10978 = n10952 & n10968;
  assign n10979 = n10977 & n10978;
  assign n10970 = n10969 ^ n10959;
  assign n10980 = n10979 ^ n10970;
  assign n10991 = n10990 ^ n10980;
  assign n11063 = n10934 & n10991;
  assign n6751 = n6741 ^ n6734;
  assign n6731 = n6730 ^ n6729;
  assign n6752 = n6751 ^ n6731;
  assign n6735 = n6734 ^ n6733;
  assign n6738 = n6737 ^ n6735;
  assign n6739 = n6738 ^ n6727;
  assign n6728 = n6727 ^ n6726;
  assign n6779 = n6739 ^ n6728;
  assign n6762 = n6741 ^ n6733;
  assign n6769 = n6762 ^ n6731;
  assign n6778 = n6769 ^ n6738;
  assign n6783 = n6779 ^ n6778;
  assign n6780 = ~n6778 & ~n6779;
  assign n6743 = n6729 ^ n6726;
  assign n6772 = ~n6743 & n6769;
  assign n6781 = n6780 ^ n6772;
  assign n6753 = n6728 & n6752;
  assign n6732 = n6731 ^ n6728;
  assign n6736 = n6735 ^ n6732;
  assign n6747 = n6741 ^ n6726;
  assign n6750 = ~n6736 & n6747;
  assign n6754 = n6753 ^ n6750;
  assign n6782 = n6781 ^ n6754;
  assign n6784 = n6783 ^ n6782;
  assign n6773 = n6729 & ~n6738;
  assign n6774 = n6773 ^ n6772;
  assign n6770 = n6769 ^ n6743;
  assign n6742 = n6741 ^ n6727;
  assign n6763 = n6762 ^ n6728;
  assign n6764 = n6742 & ~n6763;
  assign n6765 = n6764 ^ n6753;
  assign n6771 = n6770 ^ n6765;
  assign n6775 = n6774 ^ n6771;
  assign n6790 = n6784 ^ n6775;
  assign n6761 = n6751 ^ n6732;
  assign n6766 = n6765 ^ n6761;
  assign n6756 = n6738 ^ n6729;
  assign n6757 = n6756 ^ n6747;
  assign n6758 = n6737 ^ n6732;
  assign n6759 = n6757 & n6758;
  assign n6744 = n6743 ^ n6742;
  assign n6745 = ~n6732 & ~n6744;
  assign n6760 = n6759 ^ n6745;
  assign n6767 = n6766 ^ n6760;
  assign n6776 = n6767 & ~n6775;
  assign n6748 = n6747 ^ n6736;
  assign n6740 = ~n6737 & ~n6739;
  assign n6746 = n6745 ^ n6740;
  assign n6749 = n6748 ^ n6746;
  assign n6755 = n6754 ^ n6749;
  assign n6801 = n6776 ^ n6755;
  assign n6802 = ~n6790 & ~n6801;
  assign n6803 = n6802 ^ n6784;
  assign n6768 = n6767 ^ n6755;
  assign n6795 = n6784 ^ n6776;
  assign n6796 = ~n6768 & n6795;
  assign n6797 = n6796 ^ n6755;
  assign n6814 = n6803 ^ n6797;
  assign n6816 = n6752 & ~n6814;
  assign n6815 = n6728 & ~n6814;
  assign n6817 = n6816 ^ n6815;
  assign n6791 = n6790 ^ n6776;
  assign n6788 = ~n6755 & ~n6775;
  assign n6789 = ~n6784 & n6788;
  assign n6792 = n6791 ^ n6789;
  assign n6785 = n6755 & n6767;
  assign n6786 = n6784 & n6785;
  assign n6777 = n6776 ^ n6768;
  assign n6787 = n6786 ^ n6777;
  assign n6793 = n6792 ^ n6787;
  assign n6811 = n6747 & n6793;
  assign n6812 = n6811 ^ n5535;
  assign n6808 = ~n6779 & ~n6797;
  assign n6805 = n6803 ^ n6792;
  assign n6806 = ~n6732 & ~n6805;
  assign n6804 = ~n6737 & n6803;
  assign n6807 = n6806 ^ n6804;
  assign n6809 = n6808 ^ n6807;
  assign n6798 = n6797 ^ n6787;
  assign n6799 = ~n6743 & n6798;
  assign n6794 = ~n6736 & n6793;
  assign n6800 = n6799 ^ n6794;
  assign n6810 = n6809 ^ n6800;
  assign n6813 = n6812 ^ n6810;
  assign n6818 = n6817 ^ n6813;
  assign n11064 = n11063 ^ n6818;
  assign n11011 = ~n10972 & ~n10983;
  assign n11008 = n10994 ^ n10990;
  assign n11009 = ~n10929 & ~n11008;
  assign n11007 = ~n10937 & n10994;
  assign n11010 = n11009 ^ n11007;
  assign n11012 = n11011 ^ n11010;
  assign n10984 = n10983 ^ n10980;
  assign n11004 = ~n10930 & n10984;
  assign n11003 = ~n10963 & n10991;
  assign n11005 = n11004 ^ n11003;
  assign n11062 = n11012 ^ n11005;
  assign n11065 = n11064 ^ n11062;
  assign n11068 = n11067 ^ n11065;
  assign n13495 = n13494 ^ n11068;
  assign n13491 = ~n13236 & ~n13247;
  assign n13421 = ~n13198 & n13258;
  assign n13265 = n13258 ^ n13254;
  assign n13321 = ~n13191 & ~n13265;
  assign n13440 = n13421 ^ n13321;
  assign n13492 = n13491 ^ n13440;
  assign n13248 = n13247 ^ n13244;
  assign n13375 = ~n13192 & n13248;
  assign n13374 = ~n13227 & n13255;
  assign n13376 = n13375 ^ n13374;
  assign n13493 = n13492 ^ n13376;
  assign n13496 = n13495 ^ n13493;
  assign n13498 = n13497 ^ n13496;
  assign n19296 = n19295 ^ n13498;
  assign n19292 = n19235 & n19274;
  assign n19289 = n19287 ^ n19281;
  assign n19290 = n19222 & n19289;
  assign n19288 = n18505 & n19287;
  assign n19291 = n19290 ^ n19288;
  assign n19293 = n19292 ^ n19291;
  assign n19283 = n19224 & n19282;
  assign n19275 = n19274 ^ n19271;
  assign n19276 = n19218 & n19275;
  assign n19284 = n19283 ^ n19276;
  assign n19294 = n19293 ^ n19284;
  assign n19297 = n19296 ^ n19294;
  assign n19302 = n19301 ^ n19297;
  assign n6819 = n6818 ^ n5536;
  assign n14032 = n11068 ^ n6819;
  assign n17134 = n14032 ^ n13498;
  assign n19303 = n19302 ^ n17134;
  assign n11651 = n7591 ^ n6819;
  assign n14702 = n14032 ^ n11651;
  assign n17359 = n17134 ^ n14702;
  assign n19304 = n19303 ^ n17359;
  assign n12502 = n11651 ^ n8258;
  assign n14703 = n14702 ^ n12502;
  assign n17360 = n17359 ^ n14703;
  assign n21965 = n19304 ^ n17360;
  assign n19376 = n19243 & n19281;
  assign n19365 = n19298 ^ n19282;
  assign n19366 = n19246 & n19365;
  assign n19367 = n19366 ^ n19299;
  assign n19477 = n19376 ^ n19367;
  assign n19370 = n19251 & n19365;
  assign n19449 = n19370 ^ n19300;
  assign n19422 = n19244 & n19281;
  assign n19421 = n19247 & n19289;
  assign n19423 = n19422 ^ n19421;
  assign n19424 = n19423 ^ n19290;
  assign n19476 = n19449 ^ n19424;
  assign n19478 = n19477 ^ n19476;
  assign n13269 = n13204 & ~n13254;
  assign n13260 = n13259 ^ n13255;
  assign n13261 = n13193 & ~n13260;
  assign n13263 = n13262 ^ n13261;
  assign n13467 = n13269 ^ n13263;
  assign n13319 = n13205 & ~n13254;
  assign n13266 = ~n13194 & ~n13265;
  assign n13320 = n13319 ^ n13266;
  assign n13322 = n13321 ^ n13320;
  assign n13271 = ~n13212 & ~n13260;
  assign n13273 = n13272 ^ n13271;
  assign n13466 = n13322 ^ n13273;
  assign n13468 = n13467 ^ n13466;
  assign n11017 = n10940 & ~n10990;
  assign n10996 = n10995 ^ n10991;
  assign n10997 = n10931 & ~n10996;
  assign n10999 = n10998 ^ n10997;
  assign n11193 = n11017 ^ n10999;
  assign n11002 = ~n10948 & ~n10996;
  assign n11134 = n11066 ^ n11002;
  assign n11109 = n10941 & ~n10990;
  assign n11108 = ~n10932 & ~n11008;
  assign n11110 = n11109 ^ n11108;
  assign n11111 = n11110 ^ n11009;
  assign n11192 = n11134 ^ n11111;
  assign n11194 = n11193 ^ n11192;
  assign n6879 = n6757 & ~n6792;
  assign n6873 = n6814 ^ n6793;
  assign n6877 = n6742 & ~n6873;
  assign n6878 = n6877 ^ n6815;
  assign n6880 = n6879 ^ n6878;
  assign n6874 = ~n6763 & ~n6873;
  assign n6875 = n6874 ^ n6816;
  assign n6870 = n6758 & ~n6792;
  assign n6869 = ~n6744 & ~n6805;
  assign n6871 = n6870 ^ n6869;
  assign n6872 = n6871 ^ n6806;
  assign n6876 = n6875 ^ n6872;
  assign n6881 = n6880 ^ n6876;
  assign n6882 = n6881 ^ n5135;
  assign n11195 = n11194 ^ n6882;
  assign n13469 = n13468 ^ n11195;
  assign n19479 = n19478 ^ n13469;
  assign n6883 = n6882 ^ n5136;
  assign n14027 = n11195 ^ n6883;
  assign n17140 = n14027 ^ n13469;
  assign n19480 = n19479 ^ n17140;
  assign n11656 = n7596 ^ n6883;
  assign n14692 = n14027 ^ n11656;
  assign n17368 = n17140 ^ n14692;
  assign n19481 = n19480 ^ n17368;
  assign n12498 = n11656 ^ n8262;
  assign n14693 = n14692 ^ n12498;
  assign n17369 = n17368 ^ n14693;
  assign n21961 = n19481 ^ n17369;
  assign n22457 = n21965 ^ n21961;
  assign n19505 = n19233 & n19274;
  assign n19504 = n19242 & n19271;
  assign n19506 = n19505 ^ n19504;
  assign n19507 = n19506 ^ n19291;
  assign n19364 = n19231 & n19275;
  assign n19368 = n19367 ^ n19364;
  assign n19503 = n19368 ^ n19276;
  assign n19508 = n19507 ^ n19503;
  assign n13379 = ~n13235 & ~n13247;
  assign n13378 = n13203 & ~n13244;
  assign n13380 = n13379 ^ n13378;
  assign n13441 = n13440 ^ n13380;
  assign n13249 = n13185 & n13248;
  assign n13264 = n13263 ^ n13249;
  assign n13439 = n13375 ^ n13264;
  assign n13442 = n13441 ^ n13439;
  assign n11169 = ~n10971 & ~n10983;
  assign n11168 = n10939 & ~n10980;
  assign n11170 = n11169 ^ n11168;
  assign n11209 = n11170 ^ n11010;
  assign n10985 = n10925 & n10984;
  assign n11000 = n10999 ^ n10985;
  assign n11208 = n11004 ^ n11000;
  assign n11210 = n11209 ^ n11208;
  assign n6924 = ~n6778 & ~n6797;
  assign n6923 = n6756 & ~n6787;
  assign n6925 = n6924 ^ n6923;
  assign n6926 = n6925 ^ n6807;
  assign n6920 = n6769 & n6798;
  assign n6921 = n6920 ^ n6878;
  assign n6922 = n6921 ^ n6799;
  assign n6927 = n6926 ^ n6922;
  assign n6928 = n6927 ^ n5592;
  assign n11211 = n11210 ^ n6928;
  assign n13443 = n13442 ^ n11211;
  assign n19509 = n19508 ^ n13443;
  assign n6929 = n6928 ^ n5593;
  assign n14052 = n11211 ^ n6929;
  assign n17128 = n14052 ^ n13443;
  assign n19510 = n19509 ^ n17128;
  assign n11647 = n7584 ^ n6929;
  assign n14711 = n14052 ^ n11647;
  assign n17371 = n17128 ^ n14711;
  assign n19511 = n19510 ^ n17371;
  assign n12494 = n11647 ^ n8271;
  assign n14712 = n14711 ^ n12494;
  assign n17372 = n17371 ^ n14712;
  assign n21969 = n19511 ^ n17372;
  assign n22458 = n22457 ^ n21969;
  assign n19375 = n19232 & n19271;
  assign n19532 = n19375 ^ n19367;
  assign n19371 = n19370 ^ n19284;
  assign n19531 = n19506 ^ n19371;
  assign n19533 = n19532 ^ n19531;
  assign n13377 = n13376 ^ n13271;
  assign n13381 = n13380 ^ n13377;
  assign n13268 = ~n13202 & ~n13244;
  assign n13373 = n13268 ^ n13263;
  assign n13382 = n13381 ^ n13373;
  assign n11006 = n11005 ^ n11002;
  assign n11171 = n11170 ^ n11006;
  assign n11016 = ~n10938 & ~n10980;
  assign n11167 = n11016 ^ n10999;
  assign n11172 = n11171 ^ n11167;
  assign n7014 = n6874 ^ n6800;
  assign n7039 = n7014 ^ n6925;
  assign n6950 = ~n6738 & ~n6787;
  assign n7038 = n6950 ^ n6878;
  assign n7040 = n7039 ^ n7038;
  assign n7041 = n7040 ^ n5730;
  assign n11173 = n11172 ^ n7041;
  assign n13383 = n13382 ^ n11173;
  assign n19534 = n19533 ^ n13383;
  assign n7042 = n7041 ^ n5731;
  assign n14013 = n11173 ^ n7042;
  assign n17101 = n14013 ^ n13383;
  assign n19535 = n19534 ^ n17101;
  assign n11678 = n7559 ^ n7042;
  assign n14684 = n14013 ^ n11678;
  assign n17364 = n17101 ^ n14684;
  assign n19536 = n19535 ^ n17364;
  assign n12521 = n11678 ^ n8253;
  assign n14685 = n14684 ^ n12521;
  assign n17365 = n17364 ^ n14685;
  assign n21957 = n19536 ^ n17365;
  assign n22480 = n22458 ^ n21957;
  assign n19377 = n19376 ^ n19375;
  assign n19450 = n19449 ^ n19377;
  assign n19448 = n19421 ^ n19368;
  assign n19451 = n19450 ^ n19448;
  assign n13270 = n13269 ^ n13268;
  assign n13274 = n13273 ^ n13270;
  assign n13267 = n13266 ^ n13264;
  assign n13275 = n13274 ^ n13267;
  assign n11018 = n11017 ^ n11016;
  assign n11135 = n11134 ^ n11018;
  assign n11133 = n11108 ^ n11000;
  assign n11136 = n11135 ^ n11133;
  assign n6951 = n6950 ^ n6879;
  assign n6952 = n6951 ^ n6875;
  assign n6949 = n6921 ^ n6869;
  assign n6953 = n6952 ^ n6949;
  assign n6954 = n6953 ^ n5675;
  assign n11137 = n11136 ^ n6954;
  assign n13276 = n13275 ^ n11137;
  assign n19452 = n19451 ^ n13276;
  assign n6955 = n6954 ^ n5676;
  assign n14005 = n11137 ^ n6955;
  assign n17114 = n14005 ^ n13276;
  assign n19453 = n19452 ^ n17114;
  assign n11671 = n7570 ^ n6955;
  assign n14682 = n14005 ^ n11671;
  assign n17378 = n17114 ^ n14682;
  assign n19454 = n19453 ^ n17378;
  assign n12514 = n11671 ^ n8250;
  assign n14683 = n14682 ^ n12514;
  assign n17379 = n17378 ^ n14683;
  assign n21988 = n19454 ^ n17379;
  assign n19374 = n19234 & n19287;
  assign n19378 = n19377 ^ n19374;
  assign n19372 = n19371 ^ n19293;
  assign n13523 = ~n13224 & n13258;
  assign n13524 = n13523 ^ n13270;
  assign n13521 = n13492 ^ n13377;
  assign n11015 = ~n10960 & n10994;
  assign n11019 = n11018 ^ n11015;
  assign n11013 = n11012 ^ n11006;
  assign n7017 = ~n6739 & n6803;
  assign n7018 = n7017 ^ n6951;
  assign n7015 = n7014 ^ n6809;
  assign n7013 = n6921 ^ n5638;
  assign n7016 = n7015 ^ n7013;
  assign n7019 = n7018 ^ n7016;
  assign n11001 = n11000 ^ n7019;
  assign n11014 = n11013 ^ n11001;
  assign n11020 = n11019 ^ n11014;
  assign n13520 = n13264 ^ n11020;
  assign n13522 = n13521 ^ n13520;
  assign n13525 = n13524 ^ n13522;
  assign n19369 = n19368 ^ n13525;
  assign n19373 = n19372 ^ n19369;
  assign n19379 = n19378 ^ n19373;
  assign n7020 = n7019 ^ n5639;
  assign n14040 = n11020 ^ n7020;
  assign n17146 = n14040 ^ n13525;
  assign n19380 = n19379 ^ n17146;
  assign n11692 = n7604 ^ n7020;
  assign n14690 = n14040 ^ n11692;
  assign n17357 = n17146 ^ n14690;
  assign n19381 = n19380 ^ n17357;
  assign n12531 = n11692 ^ n8256;
  assign n14691 = n14690 ^ n12531;
  assign n17358 = n17357 ^ n14691;
  assign n21982 = n19381 ^ n17358;
  assign n22466 = n21988 ^ n21982;
  assign n22481 = n22480 ^ n22466;
  assign n22501 = n21957 & ~n22458;
  assign n22453 = n21988 ^ n21957;
  assign n19560 = n19505 ^ n19288;
  assign n19558 = n19423 ^ n19377;
  assign n13422 = n13421 ^ n13379;
  assign n13419 = n13320 ^ n13270;
  assign n11238 = n11169 ^ n11007;
  assign n11236 = n11110 ^ n11018;
  assign n7066 = n6924 ^ n6804;
  assign n7064 = n6951 ^ n6871;
  assign n7063 = n6878 ^ n5748;
  assign n7065 = n7064 ^ n7063;
  assign n7067 = n7066 ^ n7065;
  assign n11235 = n10999 ^ n7067;
  assign n11237 = n11236 ^ n11235;
  assign n11239 = n11238 ^ n11237;
  assign n13418 = n13263 ^ n11239;
  assign n13420 = n13419 ^ n13418;
  assign n13423 = n13422 ^ n13420;
  assign n19557 = n19367 ^ n13423;
  assign n19559 = n19558 ^ n19557;
  assign n19561 = n19560 ^ n19559;
  assign n7068 = n7067 ^ n5749;
  assign n14019 = n11239 ^ n7068;
  assign n17107 = n14019 ^ n13423;
  assign n19562 = n19561 ^ n17107;
  assign n11685 = n7564 ^ n7068;
  assign n14695 = n14019 ^ n11685;
  assign n17362 = n17107 ^ n14695;
  assign n19563 = n19562 ^ n17362;
  assign n12526 = n11685 ^ n8252;
  assign n14696 = n14695 ^ n12526;
  assign n17363 = n17362 ^ n14696;
  assign n21977 = n19563 ^ n17363;
  assign n22455 = n21977 ^ n21957;
  assign n22454 = n21982 ^ n21965;
  assign n22456 = n22455 ^ n22454;
  assign n22464 = ~n22453 & n22456;
  assign n22502 = n22501 ^ n22464;
  assign n22499 = n22456 ^ n22453;
  assign n19425 = n19424 ^ n19377;
  assign n13323 = n13322 ^ n13270;
  assign n11112 = n11111 ^ n11018;
  assign n6977 = n6951 ^ n6872;
  assign n6976 = n6921 ^ n5708;
  assign n6978 = n6977 ^ n6976;
  assign n11107 = n11000 ^ n6978;
  assign n11113 = n11112 ^ n11107;
  assign n13318 = n13264 ^ n11113;
  assign n13324 = n13323 ^ n13318;
  assign n19420 = n19368 ^ n13324;
  assign n19426 = n19425 ^ n19420;
  assign n6979 = n6978 ^ n5709;
  assign n13999 = n11113 ^ n6979;
  assign n17120 = n13999 ^ n13324;
  assign n19427 = n19426 ^ n17120;
  assign n11664 = n7579 ^ n6979;
  assign n14687 = n13999 ^ n11664;
  assign n17375 = n17120 ^ n14687;
  assign n19428 = n19427 ^ n17375;
  assign n12509 = n11664 ^ n8249;
  assign n14688 = n14687 ^ n12509;
  assign n17376 = n17375 ^ n14688;
  assign n21995 = n19428 ^ n17376;
  assign n22477 = n21995 ^ n21982;
  assign n22461 = n21995 ^ n21988;
  assign n22486 = n22461 ^ n22454;
  assign n22487 = n22477 & ~n22486;
  assign n22470 = n21982 ^ n21961;
  assign n22471 = n22470 ^ n22455;
  assign n22472 = n22461 & ~n22471;
  assign n22488 = n22487 ^ n22472;
  assign n22500 = n22499 ^ n22488;
  assign n22503 = n22502 ^ n22500;
  assign n22460 = n22458 ^ n21995;
  assign n22462 = n22461 ^ n22460;
  assign n22459 = n22458 ^ n22456;
  assign n22475 = n22462 ^ n22459;
  assign n22467 = n22461 ^ n22455;
  assign n22468 = n22467 ^ n22457;
  assign n22469 = n22466 & n22468;
  assign n22473 = n22472 ^ n22469;
  assign n22463 = ~n22459 & ~n22462;
  assign n22465 = n22464 ^ n22463;
  assign n22474 = n22473 ^ n22465;
  assign n22476 = n22475 ^ n22474;
  assign n22514 = n22503 ^ n22476;
  assign n22485 = n22470 ^ n22467;
  assign n22489 = n22488 ^ n22485;
  assign n22482 = n22467 ^ n21969;
  assign n22483 = n22481 & ~n22482;
  assign n22478 = n22477 ^ n22453;
  assign n22479 = ~n22467 & ~n22478;
  assign n22484 = n22483 ^ n22479;
  assign n22490 = n22489 ^ n22484;
  assign n22504 = ~n22490 & ~n22503;
  assign n22515 = n22514 ^ n22504;
  assign n22493 = n22468 ^ n22466;
  assign n22491 = n21969 & ~n22460;
  assign n22492 = n22491 ^ n22479;
  assign n22494 = n22493 ^ n22492;
  assign n22495 = n22494 ^ n22473;
  assign n22512 = n22495 & ~n22503;
  assign n22513 = ~n22476 & n22512;
  assign n22516 = n22515 ^ n22513;
  assign n22594 = n22481 & ~n22516;
  assign n22520 = n22504 ^ n22495;
  assign n22521 = ~n22514 & n22520;
  assign n22522 = n22521 ^ n22476;
  assign n22498 = n22495 ^ n22490;
  assign n22507 = n22504 ^ n22476;
  assign n22508 = ~n22498 & n22507;
  assign n22509 = n22508 ^ n22495;
  assign n22523 = n22522 ^ n22509;
  assign n22533 = n22461 & n22523;
  assign n22505 = n22504 ^ n22498;
  assign n22496 = ~n22490 & ~n22495;
  assign n22497 = n22476 & n22496;
  assign n22506 = n22505 ^ n22497;
  assign n22517 = n22516 ^ n22506;
  assign n22524 = n22523 ^ n22517;
  assign n22532 = n22477 & n22524;
  assign n22534 = n22533 ^ n22532;
  assign n22789 = n22594 ^ n22534;
  assign n22688 = ~n22471 & n22523;
  assign n22525 = ~n22486 & n22524;
  assign n22740 = n22688 ^ n22525;
  assign n22596 = n22522 ^ n22516;
  assign n22642 = ~n22467 & ~n22596;
  assign n22598 = ~n22482 & ~n22516;
  assign n22597 = ~n22478 & ~n22596;
  assign n22599 = n22598 ^ n22597;
  assign n22714 = n22642 ^ n22599;
  assign n22788 = n22740 ^ n22714;
  assign n22790 = n22789 ^ n22788;
  assign n17370 = n17369 ^ n17360;
  assign n17373 = n17372 ^ n17370;
  assign n17400 = n17373 ^ n17365;
  assign n17386 = n17379 ^ n17358;
  assign n17401 = n17400 ^ n17386;
  assign n17421 = ~n17365 & ~n17373;
  assign n17366 = n17365 ^ n17363;
  assign n17361 = n17360 ^ n17358;
  assign n17367 = n17366 ^ n17361;
  assign n17383 = n17379 ^ n17365;
  assign n17384 = n17367 & n17383;
  assign n17422 = n17421 ^ n17384;
  assign n17419 = n17383 ^ n17367;
  assign n17397 = n17376 ^ n17358;
  assign n17380 = n17379 ^ n17376;
  assign n17406 = n17380 ^ n17361;
  assign n17407 = ~n17397 & ~n17406;
  assign n17390 = n17369 ^ n17358;
  assign n17391 = n17390 ^ n17366;
  assign n17392 = ~n17380 & n17391;
  assign n17408 = n17407 ^ n17392;
  assign n17420 = n17419 ^ n17408;
  assign n17423 = n17422 ^ n17420;
  assign n17377 = n17376 ^ n17373;
  assign n17381 = n17380 ^ n17377;
  assign n17374 = n17373 ^ n17367;
  assign n17395 = n17381 ^ n17374;
  assign n17387 = n17380 ^ n17366;
  assign n17388 = n17387 ^ n17370;
  assign n17389 = n17386 & ~n17388;
  assign n17393 = n17392 ^ n17389;
  assign n17382 = ~n17374 & ~n17381;
  assign n17385 = n17384 ^ n17382;
  assign n17394 = n17393 ^ n17385;
  assign n17396 = n17395 ^ n17394;
  assign n17434 = n17423 ^ n17396;
  assign n17405 = n17390 ^ n17387;
  assign n17409 = n17408 ^ n17405;
  assign n17402 = n17387 ^ n17372;
  assign n17403 = ~n17401 & n17402;
  assign n17398 = n17397 ^ n17383;
  assign n17399 = ~n17387 & ~n17398;
  assign n17404 = n17403 ^ n17399;
  assign n17410 = n17409 ^ n17404;
  assign n17424 = ~n17410 & n17423;
  assign n17435 = n17434 ^ n17424;
  assign n17413 = n17388 ^ n17386;
  assign n17411 = ~n17372 & n17377;
  assign n17412 = n17411 ^ n17399;
  assign n17414 = n17413 ^ n17412;
  assign n17415 = n17414 ^ n17393;
  assign n17432 = ~n17415 & n17423;
  assign n17433 = ~n17396 & n17432;
  assign n17436 = n17435 ^ n17433;
  assign n17451 = ~n17401 & n17436;
  assign n17438 = n17424 ^ n17415;
  assign n17439 = n17434 & ~n17438;
  assign n17440 = n17439 ^ n17396;
  assign n17418 = n17415 ^ n17410;
  assign n17427 = n17424 ^ n17396;
  assign n17428 = n17418 & n17427;
  assign n17429 = n17428 ^ n17415;
  assign n17441 = n17440 ^ n17429;
  assign n17444 = ~n17380 & ~n17441;
  assign n17425 = n17424 ^ n17418;
  assign n17416 = ~n17410 & n17415;
  assign n17417 = n17396 & n17416;
  assign n17426 = n17425 ^ n17417;
  assign n17437 = n17436 ^ n17426;
  assign n17442 = n17441 ^ n17437;
  assign n17443 = ~n17397 & ~n17442;
  assign n17445 = n17444 ^ n17443;
  assign n17593 = n17451 ^ n17445;
  assign n17589 = n17402 & n17436;
  assign n17447 = n17440 ^ n17436;
  assign n17448 = ~n17398 & n17447;
  assign n17590 = n17589 ^ n17448;
  assign n17550 = ~n17387 & n17447;
  assign n17591 = n17590 ^ n17550;
  assign n17454 = n17391 & ~n17441;
  assign n17453 = ~n17406 & ~n17442;
  assign n17455 = n17454 ^ n17453;
  assign n17592 = n17591 ^ n17455;
  assign n17594 = n17593 ^ n17592;
  assign n14704 = n14703 ^ n14693;
  assign n14713 = n14712 ^ n14704;
  assign n14730 = n14713 ^ n14685;
  assign n14700 = n14691 ^ n14683;
  assign n14731 = n14730 ^ n14700;
  assign n14708 = n14703 ^ n14691;
  assign n14697 = n14696 ^ n14685;
  assign n14709 = n14708 ^ n14697;
  assign n14716 = n14713 ^ n14709;
  assign n14714 = n14713 ^ n14688;
  assign n14689 = n14688 ^ n14683;
  assign n14715 = n14714 ^ n14689;
  assign n14720 = n14716 ^ n14715;
  assign n14717 = ~n14715 & n14716;
  assign n14686 = n14685 ^ n14683;
  assign n14710 = ~n14686 & ~n14709;
  assign n14718 = n14717 ^ n14710;
  assign n14701 = n14697 ^ n14689;
  assign n14705 = n14704 ^ n14701;
  assign n14706 = n14700 & n14705;
  assign n14694 = n14693 ^ n14691;
  assign n14698 = n14697 ^ n14694;
  assign n14699 = n14689 & ~n14698;
  assign n14707 = n14706 ^ n14699;
  assign n14719 = n14718 ^ n14707;
  assign n14721 = n14720 ^ n14719;
  assign n14727 = n14705 ^ n14700;
  assign n14725 = ~n14712 & ~n14714;
  assign n14722 = n14691 ^ n14688;
  assign n14723 = n14722 ^ n14686;
  assign n14724 = n14701 & ~n14723;
  assign n14726 = n14725 ^ n14724;
  assign n14728 = n14727 ^ n14726;
  assign n14729 = n14728 ^ n14707;
  assign n14746 = n14685 & ~n14713;
  assign n14747 = n14746 ^ n14710;
  assign n14744 = n14709 ^ n14686;
  assign n14736 = n14708 ^ n14689;
  assign n14737 = n14722 & ~n14736;
  assign n14738 = n14737 ^ n14699;
  assign n14745 = n14744 ^ n14738;
  assign n14748 = n14747 ^ n14745;
  assign n14759 = n14729 & n14748;
  assign n14760 = n14721 & n14759;
  assign n14757 = n14748 ^ n14721;
  assign n14735 = n14701 ^ n14694;
  assign n14739 = n14738 ^ n14735;
  assign n14732 = n14712 ^ n14701;
  assign n14733 = n14731 & ~n14732;
  assign n14734 = n14733 ^ n14724;
  assign n14740 = n14739 ^ n14734;
  assign n14749 = ~n14740 & n14748;
  assign n14758 = n14757 ^ n14749;
  assign n14761 = n14760 ^ n14758;
  assign n15205 = n14731 & ~n14761;
  assign n14765 = n14749 ^ n14729;
  assign n14766 = ~n14757 & n14765;
  assign n14767 = n14766 ^ n14721;
  assign n14743 = n14740 ^ n14729;
  assign n14752 = n14749 ^ n14721;
  assign n14753 = ~n14743 & ~n14752;
  assign n14754 = n14753 ^ n14729;
  assign n14768 = n14767 ^ n14754;
  assign n14778 = n14689 & ~n14768;
  assign n14750 = n14749 ^ n14743;
  assign n14741 = ~n14729 & ~n14740;
  assign n14742 = ~n14721 & n14741;
  assign n14751 = n14750 ^ n14742;
  assign n14762 = n14761 ^ n14751;
  assign n14769 = n14768 ^ n14762;
  assign n14777 = n14722 & ~n14769;
  assign n14779 = n14778 ^ n14777;
  assign n15367 = n15205 ^ n14779;
  assign n15202 = n14767 ^ n14761;
  assign n15278 = n14701 & n15202;
  assign n15246 = ~n14732 & ~n14761;
  assign n15203 = ~n14723 & n15202;
  assign n15247 = n15246 ^ n15203;
  assign n15279 = n15278 ^ n15247;
  assign n15207 = ~n14698 & ~n14768;
  assign n14770 = ~n14736 & ~n14769;
  assign n15208 = n15207 ^ n14770;
  assign n15366 = n15279 ^ n15208;
  assign n15368 = n15367 ^ n15366;
  assign n12762 = n12502 ^ n12498;
  assign n12768 = n12762 ^ n12494;
  assign n12785 = n12768 ^ n12521;
  assign n12760 = n12531 ^ n12514;
  assign n12786 = n12785 ^ n12760;
  assign n12770 = n12768 ^ n12509;
  assign n12756 = n12514 ^ n12509;
  assign n12771 = n12770 ^ n12756;
  assign n12754 = n12526 ^ n12521;
  assign n12753 = n12531 ^ n12502;
  assign n12755 = n12754 ^ n12753;
  assign n12769 = n12768 ^ n12755;
  assign n12775 = n12771 ^ n12769;
  assign n12772 = n12769 & ~n12771;
  assign n12766 = n12521 ^ n12514;
  assign n12767 = ~n12755 & ~n12766;
  assign n12773 = n12772 ^ n12767;
  assign n12761 = n12756 ^ n12754;
  assign n12763 = n12762 ^ n12761;
  assign n12764 = ~n12760 & ~n12763;
  assign n12757 = n12531 ^ n12498;
  assign n12758 = n12757 ^ n12754;
  assign n12759 = n12756 & ~n12758;
  assign n12765 = n12764 ^ n12759;
  assign n12774 = n12773 ^ n12765;
  assign n12776 = n12775 ^ n12774;
  assign n12782 = n12763 ^ n12760;
  assign n12780 = ~n12494 & ~n12770;
  assign n12777 = n12531 ^ n12509;
  assign n12778 = n12777 ^ n12766;
  assign n12779 = ~n12761 & n12778;
  assign n12781 = n12780 ^ n12779;
  assign n12783 = n12782 ^ n12781;
  assign n12784 = n12783 ^ n12765;
  assign n12801 = n12521 & ~n12768;
  assign n12802 = n12801 ^ n12767;
  assign n12799 = n12766 ^ n12755;
  assign n12791 = n12756 ^ n12753;
  assign n12792 = ~n12777 & n12791;
  assign n12793 = n12792 ^ n12759;
  assign n12800 = n12799 ^ n12793;
  assign n12803 = n12802 ^ n12800;
  assign n12814 = n12784 & n12803;
  assign n12815 = n12776 & n12814;
  assign n12812 = n12803 ^ n12776;
  assign n12790 = n12761 ^ n12757;
  assign n12794 = n12793 ^ n12790;
  assign n12787 = n12761 ^ n12494;
  assign n12788 = ~n12786 & n12787;
  assign n12789 = n12788 ^ n12779;
  assign n12795 = n12794 ^ n12789;
  assign n12804 = ~n12795 & n12803;
  assign n12813 = n12812 ^ n12804;
  assign n12816 = n12815 ^ n12813;
  assign n12829 = ~n12786 & ~n12816;
  assign n12818 = n12804 ^ n12784;
  assign n12819 = ~n12812 & n12818;
  assign n12820 = n12819 ^ n12776;
  assign n12798 = n12795 ^ n12784;
  assign n12807 = n12804 ^ n12776;
  assign n12808 = ~n12798 & ~n12807;
  assign n12809 = n12808 ^ n12784;
  assign n12821 = n12820 ^ n12809;
  assign n12824 = n12756 & ~n12821;
  assign n12805 = n12804 ^ n12798;
  assign n12796 = ~n12784 & ~n12795;
  assign n12797 = ~n12776 & n12796;
  assign n12806 = n12805 ^ n12797;
  assign n12817 = n12816 ^ n12806;
  assign n12822 = n12821 ^ n12817;
  assign n12823 = ~n12777 & ~n12822;
  assign n12825 = n12824 ^ n12823;
  assign n13072 = n12829 ^ n12825;
  assign n12980 = ~n12758 & ~n12821;
  assign n12904 = n12791 & ~n12822;
  assign n12981 = n12980 ^ n12904;
  assign n12831 = n12820 ^ n12816;
  assign n12835 = ~n12761 & n12831;
  assign n12833 = n12787 & ~n12816;
  assign n12832 = n12778 & n12831;
  assign n12834 = n12833 ^ n12832;
  assign n12836 = n12835 ^ n12834;
  assign n13071 = n12981 ^ n12836;
  assign n13073 = n13072 ^ n13071;
  assign n13074 = n13073 ^ n8341;
  assign n15369 = n15368 ^ n13074;
  assign n17595 = n17594 ^ n15369;
  assign n22791 = n22790 ^ n17595;
  assign n13075 = n13074 ^ n10760;
  assign n15370 = n15369 ^ n13075;
  assign n17596 = n17595 ^ n15370;
  assign n22792 = n22791 ^ n17596;
  assign n13076 = n13075 ^ n10761;
  assign n15371 = n15370 ^ n13076;
  assign n19667 = n17596 ^ n15371;
  assign n22793 = n22792 ^ n19667;
  assign n13077 = n13076 ^ n10762;
  assign n15372 = n15371 ^ n13077;
  assign n19668 = n19667 ^ n15372;
  assign n22794 = n22793 ^ n19668;
  assign n22689 = n22688 ^ n22533;
  assign n22685 = n22466 & n22517;
  assign n17626 = n17454 ^ n17444;
  assign n17623 = n17386 & n17437;
  assign n15332 = n15207 ^ n14778;
  assign n15329 = n14700 & n14762;
  assign n13050 = n12980 ^ n12824;
  assign n13047 = ~n12760 & n12817;
  assign n13048 = n13047 ^ n8742;
  assign n12908 = ~n12771 & n12809;
  assign n12906 = ~n12494 & ~n12820;
  assign n12907 = n12906 ^ n12835;
  assign n12909 = n12908 ^ n12907;
  assign n12902 = ~n12763 & n12817;
  assign n12810 = n12809 ^ n12806;
  assign n12901 = ~n12766 & ~n12810;
  assign n12903 = n12902 ^ n12901;
  assign n13046 = n12909 ^ n12903;
  assign n13049 = n13048 ^ n13046;
  assign n13051 = n13050 ^ n13049;
  assign n15330 = n15329 ^ n13051;
  assign n15326 = ~n14715 & n14754;
  assign n15250 = ~n14712 & ~n14767;
  assign n15314 = n15278 ^ n15250;
  assign n15327 = n15326 ^ n15314;
  assign n14763 = n14705 & n14762;
  assign n14755 = n14754 ^ n14751;
  assign n14756 = ~n14686 & ~n14755;
  assign n14764 = n14763 ^ n14756;
  assign n15328 = n15327 ^ n14764;
  assign n15331 = n15330 ^ n15328;
  assign n15333 = n15332 ^ n15331;
  assign n17624 = n17623 ^ n15333;
  assign n17620 = ~n17381 & ~n17429;
  assign n17549 = ~n17372 & n17440;
  assign n17551 = n17550 ^ n17549;
  assign n17621 = n17620 ^ n17551;
  assign n17520 = ~n17388 & n17437;
  assign n17430 = n17429 ^ n17426;
  assign n17519 = n17383 & ~n17430;
  assign n17521 = n17520 ^ n17519;
  assign n17622 = n17621 ^ n17521;
  assign n17625 = n17624 ^ n17622;
  assign n17627 = n17626 ^ n17625;
  assign n22686 = n22685 ^ n17627;
  assign n22644 = ~n22462 & n22509;
  assign n22602 = n21969 & n22522;
  assign n22643 = n22642 ^ n22602;
  assign n22645 = n22644 ^ n22643;
  assign n22518 = n22468 & n22517;
  assign n22510 = n22509 ^ n22506;
  assign n22511 = ~n22453 & ~n22510;
  assign n22519 = n22518 ^ n22511;
  assign n22684 = n22645 ^ n22519;
  assign n22687 = n22686 ^ n22684;
  assign n22690 = n22689 ^ n22687;
  assign n13052 = n13051 ^ n10768;
  assign n15334 = n15333 ^ n13052;
  assign n17628 = n17627 ^ n15334;
  assign n22691 = n22690 ^ n17628;
  assign n13053 = n13052 ^ n10769;
  assign n15335 = n15334 ^ n13053;
  assign n19660 = n17628 ^ n15335;
  assign n22692 = n22691 ^ n19660;
  assign n13054 = n13053 ^ n10770;
  assign n15336 = n15335 ^ n13054;
  assign n19661 = n19660 ^ n15336;
  assign n22693 = n22692 ^ n19661;
  assign n24750 = n22794 ^ n22693;
  assign n22528 = ~n22459 & n22509;
  assign n22527 = n22480 & ~n22506;
  assign n22529 = n22528 ^ n22527;
  assign n22764 = n22643 ^ n22529;
  assign n22639 = n22456 & ~n22510;
  assign n22640 = n22639 ^ n22534;
  assign n22763 = n22640 ^ n22511;
  assign n22765 = n22764 ^ n22763;
  assign n17524 = ~n17400 & n17426;
  assign n17523 = ~n17374 & ~n17429;
  assign n17525 = n17524 ^ n17523;
  assign n17552 = n17551 ^ n17525;
  assign n17431 = n17367 & ~n17430;
  assign n17446 = n17445 ^ n17431;
  assign n17548 = n17519 ^ n17446;
  assign n17553 = n17552 ^ n17548;
  assign n14773 = n14730 & ~n14751;
  assign n14772 = n14716 & n14754;
  assign n14774 = n14773 ^ n14772;
  assign n15315 = n15314 ^ n14774;
  assign n15200 = ~n14709 & ~n14755;
  assign n15201 = n15200 ^ n14779;
  assign n15313 = n15201 ^ n14756;
  assign n15316 = n15315 ^ n15313;
  assign n12948 = n12769 & n12809;
  assign n12947 = n12785 & ~n12806;
  assign n12949 = n12948 ^ n12947;
  assign n13096 = n12949 ^ n12907;
  assign n12811 = ~n12755 & ~n12810;
  assign n12826 = n12825 ^ n12811;
  assign n13095 = n12901 ^ n12826;
  assign n13097 = n13096 ^ n13095;
  assign n13098 = n13097 ^ n8794;
  assign n15317 = n15316 ^ n13098;
  assign n17554 = n17553 ^ n15317;
  assign n22766 = n22765 ^ n17554;
  assign n13099 = n13098 ^ n10834;
  assign n15318 = n15317 ^ n13099;
  assign n17555 = n17554 ^ n15318;
  assign n22767 = n22766 ^ n17555;
  assign n13100 = n13099 ^ n10835;
  assign n15319 = n15318 ^ n13100;
  assign n19670 = n17555 ^ n15319;
  assign n22768 = n22767 ^ n19670;
  assign n13101 = n13100 ^ n10836;
  assign n15320 = n15319 ^ n13101;
  assign n19671 = n19670 ^ n15320;
  assign n22769 = n22768 ^ n19671;
  assign n24751 = n24750 ^ n22769;
  assign n22603 = n22602 ^ n22528;
  assign n22531 = ~n22458 & ~n22506;
  assign n22595 = n22594 ^ n22531;
  assign n22600 = n22599 ^ n22595;
  assign n17686 = n17549 ^ n17523;
  assign n17450 = ~n17373 & n17426;
  assign n17452 = n17451 ^ n17450;
  assign n17684 = n17590 ^ n17452;
  assign n15251 = n15250 ^ n14772;
  assign n14776 = ~n14713 & ~n14751;
  assign n15206 = n15205 ^ n14776;
  assign n15248 = n15247 ^ n15206;
  assign n13017 = n12948 ^ n12906;
  assign n12828 = ~n12768 & ~n12806;
  assign n12830 = n12829 ^ n12828;
  assign n13015 = n12834 ^ n12830;
  assign n13014 = n12825 ^ n8953;
  assign n13016 = n13015 ^ n13014;
  assign n13018 = n13017 ^ n13016;
  assign n15245 = n14779 ^ n13018;
  assign n15249 = n15248 ^ n15245;
  assign n15252 = n15251 ^ n15249;
  assign n17683 = n17445 ^ n15252;
  assign n17685 = n17684 ^ n17683;
  assign n17687 = n17686 ^ n17685;
  assign n22593 = n22534 ^ n17687;
  assign n22601 = n22600 ^ n22593;
  assign n22604 = n22603 ^ n22601;
  assign n13019 = n13018 ^ n10788;
  assign n15253 = n15252 ^ n13019;
  assign n17688 = n17687 ^ n15253;
  assign n22605 = n22604 ^ n17688;
  assign n13020 = n13019 ^ n10789;
  assign n15254 = n15253 ^ n13020;
  assign n19663 = n17688 ^ n15254;
  assign n22606 = n22605 ^ n19663;
  assign n13021 = n13020 ^ n10790;
  assign n15255 = n15254 ^ n13021;
  assign n19664 = n19663 ^ n15255;
  assign n22607 = n22606 ^ n19664;
  assign n22535 = n22534 ^ n22531;
  assign n22526 = n22525 ^ n22519;
  assign n22530 = n22529 ^ n22526;
  assign n22536 = n22535 ^ n22530;
  assign n17527 = n17450 ^ n17445;
  assign n17522 = n17521 ^ n17453;
  assign n17526 = n17525 ^ n17522;
  assign n17528 = n17527 ^ n17526;
  assign n14780 = n14779 ^ n14776;
  assign n14771 = n14770 ^ n14764;
  assign n14775 = n14774 ^ n14771;
  assign n14781 = n14780 ^ n14775;
  assign n12951 = n12828 ^ n12825;
  assign n12905 = n12904 ^ n12903;
  assign n12950 = n12949 ^ n12905;
  assign n12952 = n12951 ^ n12950;
  assign n12953 = n12952 ^ n8930;
  assign n14782 = n14781 ^ n12953;
  assign n17529 = n17528 ^ n14782;
  assign n22537 = n22536 ^ n17529;
  assign n12954 = n12953 ^ n10777;
  assign n14783 = n14782 ^ n12954;
  assign n17530 = n17529 ^ n14783;
  assign n22538 = n22537 ^ n17530;
  assign n12955 = n12954 ^ n10778;
  assign n14784 = n14783 ^ n12955;
  assign n19655 = n17530 ^ n14784;
  assign n22539 = n22538 ^ n19655;
  assign n12956 = n12955 ^ n10779;
  assign n14785 = n14784 ^ n12956;
  assign n19656 = n19655 ^ n14785;
  assign n22540 = n22539 ^ n19656;
  assign n24748 = n22607 ^ n22540;
  assign n22648 = ~n22460 & n22522;
  assign n22649 = n22648 ^ n22595;
  assign n22646 = n22645 ^ n22526;
  assign n17712 = n17377 & n17440;
  assign n17713 = n17712 ^ n17452;
  assign n17710 = n17621 ^ n17522;
  assign n15406 = ~n14714 & ~n14767;
  assign n15407 = n15406 ^ n15206;
  assign n12913 = ~n12770 & ~n12820;
  assign n12914 = n12913 ^ n12830;
  assign n12911 = n12826 ^ n8841;
  assign n12910 = n12909 ^ n12905;
  assign n12912 = n12911 ^ n12910;
  assign n12915 = n12914 ^ n12912;
  assign n15404 = n15201 ^ n12915;
  assign n15403 = n15327 ^ n14771;
  assign n15405 = n15404 ^ n15403;
  assign n15408 = n15407 ^ n15405;
  assign n17709 = n17446 ^ n15408;
  assign n17711 = n17710 ^ n17709;
  assign n17714 = n17713 ^ n17711;
  assign n22641 = n22640 ^ n17714;
  assign n22647 = n22646 ^ n22641;
  assign n22650 = n22649 ^ n22647;
  assign n12916 = n12915 ^ n10816;
  assign n15409 = n15408 ^ n12916;
  assign n17715 = n17714 ^ n15409;
  assign n22651 = n22650 ^ n17715;
  assign n12917 = n12916 ^ n10817;
  assign n15410 = n15409 ^ n12917;
  assign n19658 = n17715 ^ n15410;
  assign n22652 = n22651 ^ n19658;
  assign n12918 = n12917 ^ n10818;
  assign n15411 = n15410 ^ n12918;
  assign n19659 = n19658 ^ n15411;
  assign n22653 = n22652 ^ n19659;
  assign n24747 = n22693 ^ n22653;
  assign n24749 = n24748 ^ n24747;
  assign n24752 = n24751 ^ n24749;
  assign n22741 = n22740 ^ n22595;
  assign n22739 = n22640 ^ n22597;
  assign n22742 = n22741 ^ n22739;
  assign n17456 = n17455 ^ n17452;
  assign n17449 = n17448 ^ n17446;
  assign n17457 = n17456 ^ n17449;
  assign n15209 = n15208 ^ n15206;
  assign n15204 = n15203 ^ n15201;
  assign n15210 = n15209 ^ n15204;
  assign n12982 = n12981 ^ n12830;
  assign n12979 = n12832 ^ n12826;
  assign n12983 = n12982 ^ n12979;
  assign n12984 = n12983 ^ n8878;
  assign n15211 = n15210 ^ n12984;
  assign n17458 = n17457 ^ n15211;
  assign n22743 = n22742 ^ n17458;
  assign n12985 = n12984 ^ n10805;
  assign n15212 = n15211 ^ n12985;
  assign n17459 = n17458 ^ n15212;
  assign n22744 = n22743 ^ n17459;
  assign n12986 = n12985 ^ n10806;
  assign n15213 = n15212 ^ n12986;
  assign n19653 = n17459 ^ n15213;
  assign n22745 = n22744 ^ n19653;
  assign n12987 = n12986 ^ n10807;
  assign n15214 = n15213 ^ n12987;
  assign n19654 = n19653 ^ n15214;
  assign n22746 = n22745 ^ n19654;
  assign n22715 = n22714 ^ n22595;
  assign n17651 = n17591 ^ n17452;
  assign n15280 = n15279 ^ n15206;
  assign n12837 = n12836 ^ n12830;
  assign n12827 = n12826 ^ n8910;
  assign n12838 = n12837 ^ n12827;
  assign n15277 = n15201 ^ n12838;
  assign n15281 = n15280 ^ n15277;
  assign n17650 = n17446 ^ n15281;
  assign n17652 = n17651 ^ n17650;
  assign n22713 = n22640 ^ n17652;
  assign n22716 = n22715 ^ n22713;
  assign n12839 = n12838 ^ n10796;
  assign n15282 = n15281 ^ n12839;
  assign n17653 = n17652 ^ n15282;
  assign n22717 = n22716 ^ n17653;
  assign n12840 = n12839 ^ n10797;
  assign n15283 = n15282 ^ n12840;
  assign n19674 = n17653 ^ n15283;
  assign n22718 = n22717 ^ n19674;
  assign n12841 = n12840 ^ n10798;
  assign n15284 = n15283 ^ n12841;
  assign n19675 = n19674 ^ n15284;
  assign n22719 = n22718 ^ n19675;
  assign n24754 = n22746 ^ n22719;
  assign n24760 = n24754 ^ n24748;
  assign n24761 = n24760 ^ n24750;
  assign n24759 = n22746 ^ n22653;
  assign n24786 = n24761 ^ n24759;
  assign n24753 = n24751 ^ n22719;
  assign n24784 = n22769 & n24753;
  assign n24774 = n22719 ^ n22653;
  assign n24746 = n22746 ^ n22540;
  assign n24775 = n24774 ^ n24746;
  assign n24776 = n24760 & n24775;
  assign n24785 = n24784 ^ n24776;
  assign n24787 = n24786 ^ n24785;
  assign n24763 = n22794 ^ n22653;
  assign n24764 = n24763 ^ n24748;
  assign n24765 = n24754 & n24764;
  assign n24762 = n24759 & n24761;
  assign n24766 = n24765 ^ n24762;
  assign n24788 = n24787 ^ n24766;
  assign n24779 = n24754 ^ n24747;
  assign n24780 = n24774 & n24779;
  assign n24781 = n24780 ^ n24765;
  assign n24778 = n24763 ^ n24760;
  assign n24782 = n24781 ^ n24778;
  assign n24770 = n24751 ^ n22540;
  assign n24771 = n24770 ^ n24759;
  assign n24772 = n24760 ^ n22769;
  assign n24773 = n24771 & n24772;
  assign n24777 = n24776 ^ n24773;
  assign n24783 = n24782 ^ n24777;
  assign n24791 = n24788 ^ n24783;
  assign n24794 = ~n22540 & n24751;
  assign n24757 = n24746 & n24749;
  assign n24795 = n24794 ^ n24757;
  assign n24792 = n24749 ^ n24746;
  assign n24793 = n24792 ^ n24781;
  assign n24796 = n24795 ^ n24793;
  assign n24797 = n24783 & n24796;
  assign n24755 = n24754 ^ n24753;
  assign n24768 = n24755 ^ n24752;
  assign n24756 = n24752 & n24755;
  assign n24758 = n24757 ^ n24756;
  assign n24767 = n24766 ^ n24758;
  assign n24769 = n24768 ^ n24767;
  assign n24800 = n24797 ^ n24769;
  assign n24801 = n24791 & n24800;
  assign n24802 = n24801 ^ n24788;
  assign n25039 = n24752 & n24802;
  assign n24798 = n24797 ^ n24791;
  assign n24789 = n24783 & ~n24788;
  assign n24790 = n24769 & n24789;
  assign n24799 = n24798 ^ n24790;
  assign n25038 = n24770 & n24799;
  assign n25040 = n25039 ^ n25038;
  assign n24807 = n24796 ^ n24769;
  assign n24813 = n24797 ^ n24788;
  assign n24814 = n24807 & n24813;
  assign n24815 = n24814 ^ n24769;
  assign n24808 = n24807 ^ n24797;
  assign n24805 = n24788 & n24796;
  assign n24806 = ~n24769 & n24805;
  assign n24809 = n24808 ^ n24806;
  assign n24817 = n24815 ^ n24809;
  assign n24818 = n24760 & n24817;
  assign n24816 = n22769 & n24815;
  assign n24819 = n24818 ^ n24816;
  assign n25095 = n25040 ^ n24819;
  assign n24826 = n24815 ^ n24802;
  assign n24810 = n24809 ^ n24799;
  assign n24893 = n24826 ^ n24810;
  assign n24894 = n24774 & n24893;
  assign n24828 = n24754 & n24826;
  assign n24895 = n24894 ^ n24828;
  assign n24803 = n24802 ^ n24799;
  assign n24892 = n24749 & n24803;
  assign n24896 = n24895 ^ n24892;
  assign n24804 = n24746 & n24803;
  assign n25094 = n24896 ^ n24804;
  assign n25096 = n25095 ^ n25094;
  assign n19677 = n19675 ^ n19654;
  assign n19665 = n19664 ^ n19656;
  assign n19683 = n19677 ^ n19665;
  assign n19669 = n19668 ^ n19661;
  assign n19672 = n19671 ^ n19669;
  assign n19717 = ~n19656 & n19672;
  assign n19657 = n19656 ^ n19654;
  assign n19662 = n19661 ^ n19659;
  assign n19666 = n19665 ^ n19662;
  assign n19680 = n19657 & n19666;
  assign n19718 = n19717 ^ n19680;
  assign n19715 = n19666 ^ n19657;
  assign n19697 = n19675 ^ n19659;
  assign n19702 = n19677 ^ n19662;
  assign n19703 = n19697 & n19702;
  assign n19686 = n19668 ^ n19659;
  assign n19687 = n19686 ^ n19665;
  assign n19688 = n19677 & n19687;
  assign n19704 = n19703 ^ n19688;
  assign n19716 = n19715 ^ n19704;
  assign n19719 = n19718 ^ n19716;
  assign n19676 = n19675 ^ n19672;
  assign n19678 = n19677 ^ n19676;
  assign n19673 = n19672 ^ n19666;
  assign n19691 = n19678 ^ n19673;
  assign n19682 = n19659 ^ n19654;
  assign n19684 = n19683 ^ n19669;
  assign n19685 = n19682 & n19684;
  assign n19689 = n19688 ^ n19685;
  assign n19679 = n19673 & n19678;
  assign n19681 = n19680 ^ n19679;
  assign n19690 = n19689 ^ n19681;
  assign n19692 = n19691 ^ n19690;
  assign n19730 = n19719 ^ n19692;
  assign n19701 = n19686 ^ n19683;
  assign n19705 = n19704 ^ n19701;
  assign n19698 = n19697 ^ n19657;
  assign n19699 = n19683 & n19698;
  assign n19693 = n19672 ^ n19656;
  assign n19694 = n19693 ^ n19682;
  assign n19695 = n19683 ^ n19671;
  assign n19696 = n19694 & n19695;
  assign n19700 = n19699 ^ n19696;
  assign n19706 = n19705 ^ n19700;
  assign n19720 = n19706 & n19719;
  assign n19709 = n19684 ^ n19682;
  assign n19707 = n19671 & n19676;
  assign n19708 = n19707 ^ n19699;
  assign n19710 = n19709 ^ n19708;
  assign n19711 = n19710 ^ n19689;
  assign n19736 = n19720 ^ n19711;
  assign n19737 = n19730 & n19736;
  assign n19738 = n19737 ^ n19692;
  assign n19731 = n19730 ^ n19720;
  assign n19728 = n19711 & n19719;
  assign n19729 = ~n19692 & n19728;
  assign n19732 = n19731 ^ n19729;
  assign n19769 = n19738 ^ n19732;
  assign n19860 = n19683 & n19769;
  assign n19775 = n19671 & n19738;
  assign n19861 = n19860 ^ n19775;
  assign n19714 = n19711 ^ n19706;
  assign n19723 = n19720 ^ n19692;
  assign n19724 = n19714 & n19723;
  assign n19725 = n19724 ^ n19711;
  assign n19744 = n19673 & n19725;
  assign n19721 = n19720 ^ n19714;
  assign n19712 = n19706 & ~n19711;
  assign n19713 = n19692 & n19712;
  assign n19722 = n19721 ^ n19713;
  assign n19743 = n19693 & n19722;
  assign n19745 = n19744 ^ n19743;
  assign n19987 = n19861 ^ n19745;
  assign n19726 = n19725 ^ n19722;
  assign n19857 = n19666 & n19726;
  assign n19739 = n19738 ^ n19725;
  assign n19749 = n19677 & n19739;
  assign n19733 = n19732 ^ n19722;
  assign n19740 = n19739 ^ n19733;
  assign n19748 = n19697 & n19740;
  assign n19750 = n19749 ^ n19748;
  assign n19858 = n19857 ^ n19750;
  assign n19727 = n19657 & n19726;
  assign n19986 = n19858 ^ n19727;
  assign n19988 = n19987 ^ n19986;
  assign n16431 = n15284 ^ n15214;
  assign n16424 = n15255 ^ n14785;
  assign n16437 = n16431 ^ n16424;
  assign n16427 = n15372 ^ n15336;
  assign n16428 = n16427 ^ n15320;
  assign n16471 = ~n14785 & n16428;
  assign n16423 = n15214 ^ n14785;
  assign n16425 = n15411 ^ n15336;
  assign n16426 = n16425 ^ n16424;
  assign n16434 = n16423 & n16426;
  assign n16472 = n16471 ^ n16434;
  assign n16469 = n16426 ^ n16423;
  assign n16447 = n15411 ^ n15284;
  assign n16456 = n16431 ^ n16425;
  assign n16457 = n16447 & n16456;
  assign n16440 = n15411 ^ n15372;
  assign n16441 = n16440 ^ n16424;
  assign n16442 = n16431 & n16441;
  assign n16458 = n16457 ^ n16442;
  assign n16470 = n16469 ^ n16458;
  assign n16473 = n16472 ^ n16470;
  assign n16430 = n16428 ^ n15284;
  assign n16432 = n16431 ^ n16430;
  assign n16429 = n16428 ^ n16426;
  assign n16445 = n16432 ^ n16429;
  assign n16436 = n15411 ^ n15214;
  assign n16438 = n16437 ^ n16427;
  assign n16439 = n16436 & n16438;
  assign n16443 = n16442 ^ n16439;
  assign n16433 = n16429 & n16432;
  assign n16435 = n16434 ^ n16433;
  assign n16444 = n16443 ^ n16435;
  assign n16446 = n16445 ^ n16444;
  assign n16484 = n16473 ^ n16446;
  assign n16455 = n16440 ^ n16437;
  assign n16459 = n16458 ^ n16455;
  assign n16450 = n16428 ^ n14785;
  assign n16451 = n16450 ^ n16436;
  assign n16452 = n16437 ^ n15320;
  assign n16453 = n16451 & n16452;
  assign n16448 = n16447 ^ n16423;
  assign n16449 = n16437 & n16448;
  assign n16454 = n16453 ^ n16449;
  assign n16460 = n16459 ^ n16454;
  assign n16474 = n16460 & n16473;
  assign n16463 = n16438 ^ n16436;
  assign n16461 = n15320 & n16430;
  assign n16462 = n16461 ^ n16449;
  assign n16464 = n16463 ^ n16462;
  assign n16465 = n16464 ^ n16443;
  assign n16490 = n16474 ^ n16465;
  assign n16491 = n16484 & n16490;
  assign n16492 = n16491 ^ n16446;
  assign n16485 = n16484 ^ n16474;
  assign n16482 = n16465 & n16473;
  assign n16483 = ~n16446 & n16482;
  assign n16486 = n16485 ^ n16483;
  assign n16519 = n16492 ^ n16486;
  assign n16611 = n16437 & n16519;
  assign n16525 = n15320 & n16492;
  assign n16612 = n16611 ^ n16525;
  assign n16468 = n16465 ^ n16460;
  assign n16475 = n16474 ^ n16468;
  assign n16466 = n16460 & ~n16465;
  assign n16467 = n16446 & n16466;
  assign n16476 = n16475 ^ n16467;
  assign n16498 = n16450 & n16476;
  assign n16477 = n16474 ^ n16446;
  assign n16478 = n16468 & n16477;
  assign n16479 = n16478 ^ n16465;
  assign n16497 = n16429 & n16479;
  assign n16499 = n16498 ^ n16497;
  assign n16666 = n16612 ^ n16499;
  assign n16480 = n16479 ^ n16476;
  assign n16644 = n16426 & n16480;
  assign n16493 = n16492 ^ n16479;
  assign n16503 = n16431 & n16493;
  assign n16487 = n16486 ^ n16476;
  assign n16494 = n16493 ^ n16487;
  assign n16502 = n16447 & n16494;
  assign n16504 = n16503 ^ n16502;
  assign n16645 = n16644 ^ n16504;
  assign n16481 = n16423 & n16480;
  assign n16665 = n16645 ^ n16481;
  assign n16667 = n16666 ^ n16665;
  assign n15622 = n13021 ^ n12956;
  assign n15617 = n12987 ^ n12841;
  assign n15623 = n15622 ^ n15617;
  assign n15618 = n13077 ^ n13054;
  assign n15619 = n15618 ^ n13101;
  assign n15620 = n15619 ^ n12841;
  assign n15661 = n15620 ^ n15617;
  assign n15645 = n13054 ^ n12918;
  assign n15652 = n15645 ^ n15622;
  assign n15660 = n15652 ^ n15619;
  assign n15665 = n15661 ^ n15660;
  assign n15662 = ~n15660 & ~n15661;
  assign n15625 = n12987 ^ n12956;
  assign n15655 = ~n15625 & n15652;
  assign n15663 = n15662 ^ n15655;
  assign n15634 = n13077 ^ n12918;
  assign n15635 = n15634 ^ n15622;
  assign n15636 = n15617 & n15635;
  assign n15629 = n15623 ^ n15618;
  assign n15630 = n12987 ^ n12918;
  assign n15633 = ~n15629 & n15630;
  assign n15637 = n15636 ^ n15633;
  assign n15664 = n15663 ^ n15637;
  assign n15666 = n15665 ^ n15664;
  assign n15656 = n12956 & ~n15619;
  assign n15657 = n15656 ^ n15655;
  assign n15653 = n15652 ^ n15625;
  assign n15624 = n12918 ^ n12841;
  assign n15646 = n15645 ^ n15617;
  assign n15647 = n15624 & ~n15646;
  assign n15648 = n15647 ^ n15636;
  assign n15654 = n15653 ^ n15648;
  assign n15658 = n15657 ^ n15654;
  assign n15670 = n15666 ^ n15658;
  assign n15644 = n15634 ^ n15623;
  assign n15649 = n15648 ^ n15644;
  assign n15639 = n15619 ^ n12956;
  assign n15640 = n15639 ^ n15630;
  assign n15641 = n15623 ^ n13101;
  assign n15642 = n15640 & n15641;
  assign n15626 = n15625 ^ n15624;
  assign n15627 = ~n15623 & ~n15626;
  assign n15643 = n15642 ^ n15627;
  assign n15650 = n15649 ^ n15643;
  assign n15659 = n15650 & ~n15658;
  assign n15682 = n15670 ^ n15659;
  assign n15631 = n15630 ^ n15629;
  assign n15621 = ~n13101 & ~n15620;
  assign n15628 = n15627 ^ n15621;
  assign n15632 = n15631 ^ n15628;
  assign n15638 = n15637 ^ n15632;
  assign n15680 = ~n15638 & ~n15658;
  assign n15681 = ~n15666 & n15680;
  assign n15683 = n15682 ^ n15681;
  assign n15671 = n15659 ^ n15638;
  assign n15672 = ~n15670 & ~n15671;
  assign n15673 = n15672 ^ n15666;
  assign n15692 = n15683 ^ n15673;
  assign n16181 = ~n15623 & ~n15692;
  assign n15699 = ~n13101 & n15673;
  assign n16182 = n16181 ^ n15699;
  assign n15677 = n15638 & n15650;
  assign n15678 = n15666 & n15677;
  assign n15651 = n15650 ^ n15638;
  assign n15676 = n15659 ^ n15651;
  assign n15679 = n15678 ^ n15676;
  assign n16095 = n15639 & ~n15679;
  assign n15667 = n15666 ^ n15659;
  assign n15668 = ~n15651 & n15667;
  assign n15669 = n15668 ^ n15638;
  assign n15698 = ~n15660 & ~n15669;
  assign n16096 = n16095 ^ n15698;
  assign n16268 = n16182 ^ n16096;
  assign n16090 = n15679 ^ n15669;
  assign n16178 = n15652 & n16090;
  assign n15684 = n15683 ^ n15679;
  assign n15674 = n15673 ^ n15669;
  assign n15685 = n15684 ^ n15674;
  assign n15686 = n15624 & ~n15685;
  assign n15675 = n15617 & ~n15674;
  assign n15687 = n15686 ^ n15675;
  assign n16179 = n16178 ^ n15687;
  assign n16091 = ~n15625 & n16090;
  assign n16267 = n16179 ^ n16091;
  assign n16269 = n16268 ^ n16267;
  assign n16270 = n16269 ^ n12092;
  assign n16668 = n16667 ^ n16270;
  assign n19989 = n19988 ^ n16668;
  assign n25097 = n25096 ^ n19989;
  assign n16271 = n16270 ^ n12093;
  assign n19984 = n16668 ^ n16271;
  assign n19990 = n19989 ^ n19984;
  assign n25098 = n25097 ^ n19990;
  assign n16272 = n16271 ^ n12094;
  assign n19985 = n19984 ^ n16272;
  assign n19991 = n19990 ^ n19985;
  assign n25099 = n25098 ^ n19991;
  assign n17020 = n16272 ^ n13667;
  assign n20376 = n19985 ^ n17020;
  assign n23442 = n20376 ^ n19991;
  assign n26533 = n25099 ^ n23442;
  assign n24903 = n24771 & n24809;
  assign n25007 = n24903 ^ n24895;
  assign n24898 = n24779 & n24893;
  assign n24827 = n24764 & n24826;
  assign n24977 = n24898 ^ n24827;
  assign n24950 = n24772 & n24809;
  assign n24949 = n24775 & n24817;
  assign n24951 = n24950 ^ n24949;
  assign n24952 = n24951 ^ n24818;
  assign n25006 = n24977 ^ n24952;
  assign n25008 = n25007 ^ n25006;
  assign n19767 = n19694 & n19732;
  assign n20012 = n19767 ^ n19750;
  assign n19907 = n19687 & n19739;
  assign n19741 = n19702 & n19740;
  assign n19961 = n19907 ^ n19741;
  assign n19771 = n19695 & n19732;
  assign n19770 = n19698 & n19769;
  assign n19772 = n19771 ^ n19770;
  assign n19934 = n19860 ^ n19772;
  assign n20011 = n19961 ^ n19934;
  assign n20013 = n20012 ^ n20011;
  assign n16517 = n16451 & n16486;
  assign n16713 = n16517 ^ n16504;
  assign n16619 = n16441 & n16493;
  assign n16495 = n16456 & n16494;
  assign n16711 = n16619 ^ n16495;
  assign n16521 = n16452 & n16486;
  assign n16520 = n16448 & n16519;
  assign n16522 = n16521 ^ n16520;
  assign n16687 = n16611 ^ n16522;
  assign n16712 = n16711 ^ n16687;
  assign n16714 = n16713 ^ n16712;
  assign n15690 = n15640 & ~n15683;
  assign n16295 = n15690 ^ n15687;
  assign n16226 = n15635 & ~n15674;
  assign n16093 = ~n15646 & ~n15685;
  assign n16293 = n16226 ^ n16093;
  assign n15694 = n15641 & ~n15683;
  assign n15693 = ~n15626 & ~n15692;
  assign n15695 = n15694 ^ n15693;
  assign n16251 = n16181 ^ n15695;
  assign n16294 = n16293 ^ n16251;
  assign n16296 = n16295 ^ n16294;
  assign n16297 = n16296 ^ n12126;
  assign n16715 = n16714 ^ n16297;
  assign n20014 = n20013 ^ n16715;
  assign n25009 = n25008 ^ n20014;
  assign n16298 = n16297 ^ n12127;
  assign n20009 = n16715 ^ n16298;
  assign n20015 = n20014 ^ n20009;
  assign n25010 = n25009 ^ n20015;
  assign n16299 = n16298 ^ n12128;
  assign n20010 = n20009 ^ n16299;
  assign n20016 = n20015 ^ n20010;
  assign n25011 = n25010 ^ n20016;
  assign n17013 = n16299 ^ n13634;
  assign n20380 = n20010 ^ n17013;
  assign n23429 = n20380 ^ n20016;
  assign n26525 = n25011 ^ n23429;
  assign n24829 = n24828 ^ n24827;
  assign n24823 = n24759 & n24810;
  assign n19908 = n19907 ^ n19749;
  assign n19904 = n19682 & n19733;
  assign n16620 = n16619 ^ n16503;
  assign n16616 = n16436 & n16487;
  assign n16227 = n16226 ^ n15675;
  assign n16223 = n15630 & n15684;
  assign n16224 = n16223 ^ n12050;
  assign n16183 = ~n15661 & ~n15669;
  assign n16184 = n16183 ^ n16182;
  assign n16089 = ~n15629 & n15684;
  assign n16092 = n16091 ^ n16089;
  assign n16222 = n16184 ^ n16092;
  assign n16225 = n16224 ^ n16222;
  assign n16228 = n16227 ^ n16225;
  assign n16617 = n16616 ^ n16228;
  assign n16613 = n16432 & n16479;
  assign n16614 = n16613 ^ n16612;
  assign n16488 = n16438 & n16487;
  assign n16489 = n16488 ^ n16481;
  assign n16615 = n16614 ^ n16489;
  assign n16618 = n16617 ^ n16615;
  assign n16621 = n16620 ^ n16618;
  assign n19905 = n19904 ^ n16621;
  assign n19862 = n19678 & n19725;
  assign n19863 = n19862 ^ n19861;
  assign n19734 = n19684 & n19733;
  assign n19735 = n19734 ^ n19727;
  assign n19903 = n19863 ^ n19735;
  assign n19906 = n19905 ^ n19903;
  assign n19909 = n19908 ^ n19906;
  assign n24824 = n24823 ^ n19909;
  assign n24820 = n24755 & n24802;
  assign n24821 = n24820 ^ n24819;
  assign n24811 = n24761 & n24810;
  assign n24812 = n24811 ^ n24804;
  assign n24822 = n24821 ^ n24812;
  assign n24825 = n24824 ^ n24822;
  assign n24830 = n24829 ^ n24825;
  assign n16229 = n16228 ^ n12051;
  assign n19901 = n16621 ^ n16229;
  assign n19910 = n19909 ^ n19901;
  assign n24831 = n24830 ^ n19910;
  assign n16230 = n16229 ^ n12052;
  assign n19902 = n19901 ^ n16230;
  assign n19911 = n19910 ^ n19902;
  assign n24832 = n24831 ^ n19911;
  assign n16976 = n16230 ^ n13611;
  assign n20362 = n19902 ^ n16976;
  assign n23435 = n20362 ^ n19911;
  assign n26514 = n24832 ^ n23435;
  assign n26526 = n26525 ^ n26514;
  assign n26534 = n26533 ^ n26526;
  assign n24905 = n24753 & n24815;
  assign n24902 = n24751 & n24799;
  assign n24904 = n24903 ^ n24902;
  assign n24906 = n24905 ^ n24904;
  assign n24899 = n24898 ^ n24812;
  assign n24900 = n24899 ^ n24821;
  assign n19866 = n19676 & n19738;
  assign n19747 = n19672 & n19722;
  assign n19768 = n19767 ^ n19747;
  assign n19867 = n19866 ^ n19768;
  assign n19742 = n19741 ^ n19735;
  assign n19864 = n19863 ^ n19742;
  assign n16649 = n16430 & n16492;
  assign n16501 = n16428 & n16476;
  assign n16518 = n16517 ^ n16501;
  assign n16650 = n16649 ^ n16518;
  assign n16496 = n16495 ^ n16489;
  assign n16647 = n16614 ^ n16496;
  assign n16187 = ~n15620 & n15673;
  assign n15689 = ~n15619 & ~n15679;
  assign n15691 = n15690 ^ n15689;
  assign n16188 = n16187 ^ n15691;
  assign n16094 = n16093 ^ n16092;
  assign n16185 = n16184 ^ n16094;
  assign n16180 = n16179 ^ n12006;
  assign n16186 = n16185 ^ n16180;
  assign n16189 = n16188 ^ n16186;
  assign n16646 = n16645 ^ n16189;
  assign n16648 = n16647 ^ n16646;
  assign n16651 = n16650 ^ n16648;
  assign n19859 = n19858 ^ n16651;
  assign n19865 = n19864 ^ n19859;
  assign n19868 = n19867 ^ n19865;
  assign n24897 = n24896 ^ n19868;
  assign n24901 = n24900 ^ n24897;
  assign n24907 = n24906 ^ n24901;
  assign n16190 = n16189 ^ n12007;
  assign n19855 = n16651 ^ n16190;
  assign n19869 = n19868 ^ n19855;
  assign n24908 = n24907 ^ n19869;
  assign n16191 = n16190 ^ n12008;
  assign n19856 = n19855 ^ n16191;
  assign n19870 = n19869 ^ n19856;
  assign n24909 = n24908 ^ n19870;
  assign n16985 = n16191 ^ n13605;
  assign n20368 = n19856 ^ n16985;
  assign n23455 = n20368 ^ n19870;
  assign n26513 = n24909 ^ n23455;
  assign n26529 = n26525 ^ n26513;
  assign n24953 = n24952 ^ n24904;
  assign n19935 = n19934 ^ n19768;
  assign n16688 = n16687 ^ n16518;
  assign n16252 = n16251 ^ n15691;
  assign n16250 = n16179 ^ n12114;
  assign n16253 = n16252 ^ n16250;
  assign n16686 = n16645 ^ n16253;
  assign n16689 = n16688 ^ n16686;
  assign n19933 = n19858 ^ n16689;
  assign n19936 = n19935 ^ n19933;
  assign n24948 = n24896 ^ n19936;
  assign n24954 = n24953 ^ n24948;
  assign n16254 = n16253 ^ n12115;
  assign n19931 = n16689 ^ n16254;
  assign n19937 = n19936 ^ n19931;
  assign n24955 = n24954 ^ n19937;
  assign n16255 = n16254 ^ n12116;
  assign n19932 = n19931 ^ n16255;
  assign n19938 = n19937 ^ n19932;
  assign n24956 = n24955 ^ n19938;
  assign n17000 = n16255 ^ n13624;
  assign n20389 = n19932 ^ n17000;
  assign n23464 = n20389 ^ n19938;
  assign n26522 = n24956 ^ n23464;
  assign n24978 = n24977 ^ n24904;
  assign n24976 = n24949 ^ n24896;
  assign n24979 = n24978 ^ n24976;
  assign n19962 = n19961 ^ n19768;
  assign n19960 = n19858 ^ n19770;
  assign n19963 = n19962 ^ n19960;
  assign n16735 = n16711 ^ n16518;
  assign n16734 = n16645 ^ n16520;
  assign n16736 = n16735 ^ n16734;
  assign n16318 = n16293 ^ n15691;
  assign n16317 = n16179 ^ n15693;
  assign n16319 = n16318 ^ n16317;
  assign n16320 = n16319 ^ n12154;
  assign n16737 = n16736 ^ n16320;
  assign n19964 = n19963 ^ n16737;
  assign n24980 = n24979 ^ n19964;
  assign n16321 = n16320 ^ n12155;
  assign n19958 = n16737 ^ n16321;
  assign n19965 = n19964 ^ n19958;
  assign n24981 = n24980 ^ n19965;
  assign n16322 = n16321 ^ n12156;
  assign n19959 = n19958 ^ n16322;
  assign n19966 = n19965 ^ n19959;
  assign n24982 = n24981 ^ n19966;
  assign n16993 = n16322 ^ n13618;
  assign n20396 = n19959 ^ n16993;
  assign n23449 = n20396 ^ n19966;
  assign n26520 = n24982 ^ n23449;
  assign n26523 = n26522 ^ n26520;
  assign n25042 = n24902 ^ n24895;
  assign n25041 = n25040 ^ n24899;
  assign n25043 = n25042 ^ n25041;
  assign n19751 = n19750 ^ n19747;
  assign n19746 = n19745 ^ n19742;
  assign n19752 = n19751 ^ n19746;
  assign n16505 = n16504 ^ n16501;
  assign n16500 = n16499 ^ n16496;
  assign n16506 = n16505 ^ n16500;
  assign n16097 = n16096 ^ n16094;
  assign n16088 = n15689 ^ n15687;
  assign n16098 = n16097 ^ n16088;
  assign n16099 = n16098 ^ n11944;
  assign n16507 = n16506 ^ n16099;
  assign n19753 = n19752 ^ n16507;
  assign n25044 = n25043 ^ n19753;
  assign n16100 = n16099 ^ n11945;
  assign n19651 = n16507 ^ n16100;
  assign n19754 = n19753 ^ n19651;
  assign n25045 = n25044 ^ n19754;
  assign n16101 = n16100 ^ n11946;
  assign n19652 = n19651 ^ n16101;
  assign n19755 = n19754 ^ n19652;
  assign n25046 = n25045 ^ n19755;
  assign n16965 = n16101 ^ n13643;
  assign n20351 = n19652 ^ n16965;
  assign n23423 = n20351 ^ n19755;
  assign n26517 = n25046 ^ n23423;
  assign n25052 = n25039 ^ n24816;
  assign n25050 = n24951 ^ n24904;
  assign n19776 = n19775 ^ n19744;
  assign n19773 = n19772 ^ n19768;
  assign n16526 = n16525 ^ n16497;
  assign n16523 = n16522 ^ n16518;
  assign n15700 = n15699 ^ n15698;
  assign n15696 = n15695 ^ n15691;
  assign n15688 = n15687 ^ n11521;
  assign n15697 = n15696 ^ n15688;
  assign n15701 = n15700 ^ n15697;
  assign n16516 = n16504 ^ n15701;
  assign n16524 = n16523 ^ n16516;
  assign n16527 = n16526 ^ n16524;
  assign n19766 = n19750 ^ n16527;
  assign n19774 = n19773 ^ n19766;
  assign n19777 = n19776 ^ n19774;
  assign n25049 = n24895 ^ n19777;
  assign n25051 = n25050 ^ n25049;
  assign n25053 = n25052 ^ n25051;
  assign n15702 = n15701 ^ n11522;
  assign n19764 = n16527 ^ n15702;
  assign n19778 = n19777 ^ n19764;
  assign n25054 = n25053 ^ n19778;
  assign n15703 = n15702 ^ n11523;
  assign n19765 = n19764 ^ n15703;
  assign n19779 = n19778 ^ n19765;
  assign n25055 = n25054 ^ n19779;
  assign n16968 = n15703 ^ n13641;
  assign n20345 = n19765 ^ n16968;
  assign n23469 = n20345 ^ n19779;
  assign n26516 = n25055 ^ n23469;
  assign n26518 = n26517 ^ n26516;
  assign n26524 = n26523 ^ n26518;
  assign n26553 = n26529 ^ n26524;
  assign n26538 = n26522 ^ n26513;
  assign n26515 = n26514 ^ n26513;
  assign n26550 = n26523 ^ n26515;
  assign n26551 = n26538 & n26550;
  assign n26530 = n26529 ^ n26518;
  assign n26531 = n26523 & n26530;
  assign n26552 = n26551 ^ n26531;
  assign n26554 = n26553 ^ n26552;
  assign n26545 = n26534 ^ n26517;
  assign n26521 = n26520 ^ n26513;
  assign n26546 = n26545 ^ n26521;
  assign n26547 = n26533 ^ n26524;
  assign n26548 = n26546 & n26547;
  assign n26537 = n26520 ^ n26517;
  assign n26539 = n26538 ^ n26537;
  assign n26540 = n26524 & n26539;
  assign n26549 = n26548 ^ n26540;
  assign n26555 = n26554 ^ n26549;
  assign n26567 = ~n26517 & n26534;
  assign n26519 = n26518 ^ n26515;
  assign n26560 = n26519 & n26537;
  assign n26568 = n26567 ^ n26560;
  assign n26565 = n26537 ^ n26519;
  assign n26566 = n26565 ^ n26552;
  assign n26569 = n26568 ^ n26566;
  assign n26570 = n26555 & n26569;
  assign n26527 = n26526 ^ n26524;
  assign n26542 = n26527 ^ n26521;
  assign n26535 = n26534 ^ n26522;
  assign n26536 = n26533 & n26535;
  assign n26541 = n26540 ^ n26536;
  assign n26543 = n26542 ^ n26541;
  assign n26528 = n26521 & n26527;
  assign n26532 = n26531 ^ n26528;
  assign n26544 = n26543 ^ n26532;
  assign n26556 = n26555 ^ n26544;
  assign n26576 = n26570 ^ n26556;
  assign n26558 = n26535 ^ n26523;
  assign n26557 = n26534 ^ n26519;
  assign n26563 = n26558 ^ n26557;
  assign n26559 = n26557 & n26558;
  assign n26561 = n26560 ^ n26559;
  assign n26562 = n26561 ^ n26532;
  assign n26564 = n26563 ^ n26562;
  assign n26574 = ~n26544 & n26555;
  assign n26575 = n26564 & n26574;
  assign n26577 = n26576 ^ n26575;
  assign n26596 = n26534 & n26577;
  assign n26582 = n26569 ^ n26564;
  assign n26586 = n26570 ^ n26544;
  assign n26587 = n26582 & n26586;
  assign n26588 = n26587 ^ n26564;
  assign n26571 = n26570 ^ n26564;
  assign n26572 = n26556 & n26571;
  assign n26573 = n26572 ^ n26544;
  assign n26589 = n26588 ^ n26573;
  assign n26592 = n26523 & n26589;
  assign n26583 = n26582 ^ n26570;
  assign n26580 = n26544 & n26569;
  assign n26581 = ~n26564 & n26580;
  assign n26584 = n26583 ^ n26581;
  assign n26585 = n26584 ^ n26577;
  assign n26590 = n26589 ^ n26585;
  assign n26591 = n26538 & n26590;
  assign n26593 = n26592 ^ n26591;
  assign n26678 = n26596 ^ n26593;
  assign n26578 = n26577 ^ n26573;
  assign n26626 = n26537 & n26578;
  assign n26625 = n26527 & n26585;
  assign n26627 = n26626 ^ n26625;
  assign n26612 = n26550 & n26590;
  assign n26659 = n26627 ^ n26612;
  assign n26647 = n26545 & n26577;
  assign n26646 = n26557 & n26573;
  assign n26648 = n26647 ^ n26646;
  assign n26677 = n26659 ^ n26648;
  assign n26679 = n26678 ^ n26677;
  assign n23826 = n23455 ^ n23435;
  assign n23825 = n23469 ^ n23423;
  assign n23827 = n23826 ^ n23825;
  assign n23823 = n23435 ^ n23429;
  assign n23824 = n23823 ^ n23442;
  assign n23828 = n23827 ^ n23824;
  assign n23840 = n23455 ^ n23449;
  assign n23822 = n23464 ^ n23449;
  assign n23838 = n23825 ^ n23822;
  assign n23839 = n23838 ^ n23823;
  assign n23869 = n23840 ^ n23839;
  assign n23829 = n23824 ^ n23464;
  assign n23867 = n23442 & n23829;
  assign n23847 = n23464 ^ n23455;
  assign n23832 = n23449 ^ n23423;
  assign n23860 = n23847 ^ n23832;
  assign n23861 = n23838 & n23860;
  assign n23868 = n23867 ^ n23861;
  assign n23870 = n23869 ^ n23868;
  assign n23841 = n23839 & n23840;
  assign n23835 = n23455 ^ n23429;
  assign n23836 = n23835 ^ n23825;
  assign n23837 = n23822 & n23836;
  assign n23842 = n23841 ^ n23837;
  assign n23871 = n23870 ^ n23842;
  assign n23863 = n23838 ^ n23835;
  assign n23848 = n23826 ^ n23822;
  assign n23849 = n23847 & n23848;
  assign n23850 = n23849 ^ n23837;
  assign n23864 = n23863 ^ n23850;
  assign n23856 = n23838 ^ n23442;
  assign n23857 = n23824 ^ n23423;
  assign n23858 = n23857 ^ n23840;
  assign n23859 = n23856 & n23858;
  assign n23862 = n23861 ^ n23859;
  assign n23865 = n23864 ^ n23862;
  assign n23875 = n23871 ^ n23865;
  assign n23852 = ~n23423 & n23824;
  assign n23833 = n23827 & n23832;
  assign n23853 = n23852 ^ n23833;
  assign n23846 = n23832 ^ n23827;
  assign n23851 = n23850 ^ n23846;
  assign n23854 = n23853 ^ n23851;
  assign n23866 = n23854 & n23865;
  assign n23830 = n23829 ^ n23822;
  assign n23844 = n23830 ^ n23828;
  assign n23831 = n23828 & n23830;
  assign n23834 = n23833 ^ n23831;
  assign n23843 = n23842 ^ n23834;
  assign n23845 = n23844 ^ n23843;
  assign n23876 = n23866 ^ n23845;
  assign n23877 = n23875 & n23876;
  assign n23878 = n23877 ^ n23871;
  assign n24099 = n23828 & n23878;
  assign n23887 = n23875 ^ n23866;
  assign n23885 = n23865 & ~n23871;
  assign n23886 = n23845 & n23885;
  assign n23888 = n23887 ^ n23886;
  assign n24098 = n23857 & n23888;
  assign n24100 = n24099 ^ n24098;
  assign n23855 = n23854 ^ n23845;
  assign n23883 = n23866 ^ n23855;
  assign n23881 = n23854 & n23871;
  assign n23882 = ~n23845 & n23881;
  assign n23884 = n23883 ^ n23882;
  assign n23889 = n23888 ^ n23884;
  assign n23872 = n23871 ^ n23866;
  assign n23873 = n23855 & n23872;
  assign n23874 = n23873 ^ n23845;
  assign n23879 = n23878 ^ n23874;
  assign n23890 = n23889 ^ n23879;
  assign n23972 = n23848 & n23890;
  assign n23893 = n23888 ^ n23878;
  assign n23970 = n23832 & n23893;
  assign n23969 = n23839 & n23889;
  assign n23971 = n23970 ^ n23969;
  assign n23973 = n23972 ^ n23971;
  assign n24101 = n24100 ^ n23973;
  assign n23897 = n23824 & n23888;
  assign n23891 = n23847 & n23890;
  assign n23880 = n23822 & n23879;
  assign n23892 = n23891 ^ n23880;
  assign n24097 = n23897 ^ n23892;
  assign n24102 = n24101 ^ n24097;
  assign n20619 = n20380 ^ n20362;
  assign n20620 = n20619 ^ n20376;
  assign n20623 = n20396 ^ n20389;
  assign n20617 = n20351 ^ n20345;
  assign n20632 = n20623 ^ n20617;
  assign n20629 = n20380 ^ n20368;
  assign n20656 = n20632 ^ n20629;
  assign n20640 = n20389 ^ n20368;
  assign n20616 = n20368 ^ n20362;
  assign n20653 = n20623 ^ n20616;
  assign n20654 = n20640 & n20653;
  assign n20630 = n20629 ^ n20617;
  assign n20631 = n20623 & n20630;
  assign n20655 = n20654 ^ n20631;
  assign n20657 = n20656 ^ n20655;
  assign n20648 = n20620 ^ n20351;
  assign n20634 = n20396 ^ n20368;
  assign n20649 = n20648 ^ n20634;
  assign n20650 = n20632 ^ n20376;
  assign n20651 = n20649 & n20650;
  assign n20626 = n20396 ^ n20351;
  assign n20641 = n20640 ^ n20626;
  assign n20642 = n20632 & n20641;
  assign n20652 = n20651 ^ n20642;
  assign n20658 = n20657 ^ n20652;
  assign n20633 = n20632 ^ n20619;
  assign n20645 = n20634 ^ n20633;
  assign n20622 = n20620 ^ n20389;
  assign n20643 = n20376 & n20622;
  assign n20644 = n20643 ^ n20642;
  assign n20646 = n20645 ^ n20644;
  assign n20635 = n20633 & n20634;
  assign n20636 = n20635 ^ n20631;
  assign n20647 = n20646 ^ n20636;
  assign n20667 = n20658 ^ n20647;
  assign n20663 = ~n20351 & n20620;
  assign n20618 = n20617 ^ n20616;
  assign n20627 = n20618 & n20626;
  assign n20664 = n20663 ^ n20627;
  assign n20661 = n20626 ^ n20618;
  assign n20662 = n20661 ^ n20655;
  assign n20665 = n20664 ^ n20662;
  assign n20666 = n20658 & n20665;
  assign n20668 = n20667 ^ n20666;
  assign n20624 = n20623 ^ n20622;
  assign n20621 = n20620 ^ n20618;
  assign n20638 = n20624 ^ n20621;
  assign n20625 = n20621 & n20624;
  assign n20628 = n20627 ^ n20625;
  assign n20637 = n20636 ^ n20628;
  assign n20639 = n20638 ^ n20637;
  assign n20659 = ~n20647 & n20658;
  assign n20660 = n20639 & n20659;
  assign n20669 = n20668 ^ n20660;
  assign n20746 = n20620 & n20669;
  assign n20677 = n20665 ^ n20639;
  assign n20681 = n20666 ^ n20647;
  assign n20682 = n20677 & n20681;
  assign n20683 = n20682 ^ n20639;
  assign n20670 = n20666 ^ n20639;
  assign n20671 = n20667 & n20670;
  assign n20672 = n20671 ^ n20647;
  assign n20684 = n20683 ^ n20672;
  assign n20687 = n20623 & n20684;
  assign n20678 = n20677 ^ n20666;
  assign n20675 = n20647 & n20665;
  assign n20676 = ~n20639 & n20675;
  assign n20679 = n20678 ^ n20676;
  assign n20680 = n20679 ^ n20669;
  assign n20685 = n20684 ^ n20680;
  assign n20686 = n20640 & n20685;
  assign n20688 = n20687 ^ n20686;
  assign n20747 = n20746 ^ n20688;
  assign n20743 = n20653 & n20685;
  assign n20741 = n20633 & n20680;
  assign n20673 = n20672 ^ n20669;
  assign n20690 = n20626 & n20673;
  assign n20742 = n20741 ^ n20690;
  assign n20744 = n20743 ^ n20742;
  assign n20697 = n20621 & n20672;
  assign n20696 = n20648 & n20669;
  assign n20698 = n20697 ^ n20696;
  assign n20745 = n20744 ^ n20698;
  assign n20748 = n20747 ^ n20745;
  assign n18307 = n17013 ^ n16976;
  assign n18308 = n18307 ^ n17020;
  assign n18320 = n17013 ^ n16985;
  assign n18311 = n17000 ^ n16993;
  assign n18305 = n16968 ^ n16965;
  assign n18317 = n18311 ^ n18305;
  assign n18349 = n18320 ^ n18317;
  assign n18302 = n17000 ^ n16985;
  assign n18304 = n16985 ^ n16976;
  assign n18334 = n18311 ^ n18304;
  assign n18335 = n18302 & n18334;
  assign n18321 = n18320 ^ n18305;
  assign n18322 = n18311 & n18321;
  assign n18336 = n18335 ^ n18322;
  assign n18350 = n18349 ^ n18336;
  assign n18344 = n18317 ^ n17020;
  assign n18345 = n18308 ^ n16965;
  assign n18316 = n16993 ^ n16985;
  assign n18346 = n18345 ^ n18316;
  assign n18347 = n18344 & n18346;
  assign n18301 = n16993 ^ n16965;
  assign n18303 = n18302 ^ n18301;
  assign n18328 = n18303 & n18317;
  assign n18348 = n18347 ^ n18328;
  assign n18351 = n18350 ^ n18348;
  assign n18318 = n18317 ^ n18307;
  assign n18330 = n18318 ^ n18316;
  assign n18310 = n18308 ^ n17000;
  assign n18327 = n17020 & n18310;
  assign n18329 = n18328 ^ n18327;
  assign n18331 = n18330 ^ n18329;
  assign n18319 = n18316 & n18318;
  assign n18323 = n18322 ^ n18319;
  assign n18332 = n18331 ^ n18323;
  assign n18366 = n18351 ^ n18332;
  assign n18338 = ~n16965 & n18308;
  assign n18306 = n18305 ^ n18304;
  assign n18314 = n18301 & n18306;
  assign n18339 = n18338 ^ n18314;
  assign n18333 = n18306 ^ n18301;
  assign n18337 = n18336 ^ n18333;
  assign n18340 = n18339 ^ n18337;
  assign n18352 = n18340 & n18351;
  assign n18367 = n18366 ^ n18352;
  assign n18312 = n18311 ^ n18310;
  assign n18309 = n18308 ^ n18306;
  assign n18325 = n18312 ^ n18309;
  assign n18313 = n18309 & n18312;
  assign n18315 = n18314 ^ n18313;
  assign n18324 = n18323 ^ n18315;
  assign n18326 = n18325 ^ n18324;
  assign n18364 = ~n18332 & n18351;
  assign n18365 = n18326 & n18364;
  assign n18368 = n18367 ^ n18365;
  assign n18534 = n18308 & n18368;
  assign n18370 = n18352 ^ n18326;
  assign n18371 = n18366 & n18370;
  assign n18372 = n18371 ^ n18332;
  assign n18343 = n18340 ^ n18326;
  assign n18355 = n18352 ^ n18332;
  assign n18356 = n18343 & n18355;
  assign n18357 = n18356 ^ n18326;
  assign n18373 = n18372 ^ n18357;
  assign n18381 = n18311 & n18373;
  assign n18353 = n18352 ^ n18343;
  assign n18341 = n18332 & n18340;
  assign n18342 = ~n18326 & n18341;
  assign n18354 = n18353 ^ n18342;
  assign n18369 = n18368 ^ n18354;
  assign n18374 = n18373 ^ n18369;
  assign n18380 = n18302 & n18374;
  assign n18382 = n18381 ^ n18380;
  assign n18568 = n18534 ^ n18382;
  assign n18446 = n18372 ^ n18368;
  assign n18447 = n18301 & n18446;
  assign n18445 = n18318 & n18369;
  assign n18448 = n18447 ^ n18445;
  assign n18375 = n18334 & n18374;
  assign n18566 = n18448 ^ n18375;
  assign n18498 = n18309 & n18372;
  assign n18497 = n18345 & n18368;
  assign n18499 = n18498 ^ n18497;
  assign n18567 = n18566 ^ n18499;
  assign n18569 = n18568 ^ n18567;
  assign n18570 = n18569 ^ n14358;
  assign n20749 = n20748 ^ n18570;
  assign n24103 = n24102 ^ n20749;
  assign n26680 = n26679 ^ n24103;
  assign n18571 = n18570 ^ n14359;
  assign n20750 = n20749 ^ n18571;
  assign n24104 = n24103 ^ n20750;
  assign n26681 = n26680 ^ n24104;
  assign n18572 = n18571 ^ n16833;
  assign n22889 = n20750 ^ n18572;
  assign n26115 = n24104 ^ n22889;
  assign n26682 = n26681 ^ n26115;
  assign n18574 = n18573 ^ n18572;
  assign n22890 = n22889 ^ n18574;
  assign n26116 = n26115 ^ n22890;
  assign n26683 = n26682 ^ n26116;
  assign n26622 = n26533 & n26588;
  assign n26599 = n26588 ^ n26584;
  assign n26603 = n26524 & n26599;
  assign n26623 = n26622 ^ n26603;
  assign n26649 = n26648 ^ n26623;
  assign n26579 = n26519 & n26578;
  assign n26594 = n26593 ^ n26579;
  assign n26645 = n26626 ^ n26594;
  assign n26650 = n26649 ^ n26645;
  assign n23975 = n23442 & n23874;
  assign n23900 = n23884 ^ n23874;
  assign n23904 = n23838 & n23900;
  assign n23976 = n23975 ^ n23904;
  assign n24151 = n24100 ^ n23976;
  assign n23894 = n23827 & n23893;
  assign n23895 = n23894 ^ n23892;
  assign n24150 = n23970 ^ n23895;
  assign n24152 = n24151 ^ n24150;
  assign n20694 = n20376 & n20683;
  assign n20692 = n20683 ^ n20679;
  assign n20693 = n20632 & n20692;
  assign n20695 = n20694 ^ n20693;
  assign n20699 = n20698 ^ n20695;
  assign n20674 = n20618 & n20673;
  assign n20689 = n20688 ^ n20674;
  assign n20691 = n20690 ^ n20689;
  assign n20700 = n20699 ^ n20691;
  assign n18442 = n17020 & n18357;
  assign n18358 = n18357 ^ n18354;
  assign n18362 = n18317 & n18358;
  assign n18443 = n18442 ^ n18362;
  assign n18500 = n18499 ^ n18443;
  assign n18494 = n18306 & n18446;
  assign n18495 = n18494 ^ n18382;
  assign n18496 = n18495 ^ n18447;
  assign n18501 = n18500 ^ n18496;
  assign n18502 = n18501 ^ n14299;
  assign n20701 = n20700 ^ n18502;
  assign n24153 = n24152 ^ n20701;
  assign n26651 = n26650 ^ n24153;
  assign n18503 = n18502 ^ n14300;
  assign n20702 = n20701 ^ n18503;
  assign n24154 = n24153 ^ n20702;
  assign n26652 = n26651 ^ n24154;
  assign n18504 = n18503 ^ n16884;
  assign n22896 = n20702 ^ n18504;
  assign n26122 = n24154 ^ n22896;
  assign n26653 = n26652 ^ n26122;
  assign n18506 = n18505 ^ n18504;
  assign n22897 = n22896 ^ n18506;
  assign n26123 = n26122 ^ n22897;
  assign n26654 = n26653 ^ n26123;
  assign n26597 = n26546 & n26584;
  assign n26638 = n26597 ^ n26593;
  assign n26611 = n26530 & n26589;
  assign n26613 = n26612 ^ n26611;
  assign n26601 = n26547 & n26584;
  assign n26600 = n26539 & n26599;
  assign n26602 = n26601 ^ n26600;
  assign n26604 = n26603 ^ n26602;
  assign n26637 = n26613 ^ n26604;
  assign n26639 = n26638 ^ n26637;
  assign n23898 = n23858 & n23884;
  assign n24068 = n23898 ^ n23892;
  assign n24015 = n23836 & n23879;
  assign n24039 = n24015 ^ n23972;
  assign n23902 = n23856 & n23884;
  assign n23901 = n23860 & n23900;
  assign n23903 = n23902 ^ n23901;
  assign n23905 = n23904 ^ n23903;
  assign n24067 = n24039 ^ n23905;
  assign n24069 = n24068 ^ n24067;
  assign n20786 = n20649 & n20679;
  assign n20953 = n20786 ^ n20688;
  assign n20877 = n20650 & n20679;
  assign n20784 = n20641 & n20692;
  assign n20878 = n20877 ^ n20784;
  assign n20928 = n20878 ^ n20693;
  assign n20788 = n20630 & n20684;
  assign n20789 = n20788 ^ n20743;
  assign n20952 = n20928 ^ n20789;
  assign n20954 = n20953 ^ n20952;
  assign n18379 = n18346 & n18354;
  assign n18383 = n18382 ^ n18379;
  assign n18376 = n18321 & n18373;
  assign n18377 = n18376 ^ n18375;
  assign n18360 = n18344 & n18354;
  assign n18359 = n18303 & n18358;
  assign n18361 = n18360 ^ n18359;
  assign n18363 = n18362 ^ n18361;
  assign n18378 = n18377 ^ n18363;
  assign n18384 = n18383 ^ n18378;
  assign n18385 = n18384 ^ n14213;
  assign n20955 = n20954 ^ n18385;
  assign n24070 = n24069 ^ n20955;
  assign n26640 = n26639 ^ n24070;
  assign n18386 = n18385 ^ n14214;
  assign n20956 = n20955 ^ n18386;
  assign n24071 = n24070 ^ n20956;
  assign n26641 = n26640 ^ n24071;
  assign n18387 = n18386 ^ n16875;
  assign n22893 = n20956 ^ n18387;
  assign n26119 = n24071 ^ n22893;
  assign n26642 = n26641 ^ n26119;
  assign n18389 = n18388 ^ n18387;
  assign n22894 = n22893 ^ n18389;
  assign n26120 = n26119 ^ n22894;
  assign n26643 = n26642 ^ n26120;
  assign n26632 = n26611 ^ n26592;
  assign n26629 = n26521 & n26585;
  assign n24016 = n24015 ^ n23880;
  assign n24012 = n23840 & n23889;
  assign n20865 = n20788 ^ n20687;
  assign n20862 = n20634 & n20680;
  assign n18453 = n18381 ^ n18376;
  assign n18450 = n18316 & n18369;
  assign n18451 = n18450 ^ n14279;
  assign n18441 = n18312 & n18372;
  assign n18444 = n18443 ^ n18441;
  assign n18449 = n18448 ^ n18444;
  assign n18452 = n18451 ^ n18449;
  assign n18454 = n18453 ^ n18452;
  assign n20863 = n20862 ^ n18454;
  assign n20829 = n20624 & n20672;
  assign n20830 = n20829 ^ n20695;
  assign n20861 = n20830 ^ n20742;
  assign n20864 = n20863 ^ n20861;
  assign n20866 = n20865 ^ n20864;
  assign n24013 = n24012 ^ n20866;
  assign n23974 = n23830 & n23878;
  assign n23977 = n23976 ^ n23974;
  assign n24011 = n23977 ^ n23971;
  assign n24014 = n24013 ^ n24011;
  assign n24017 = n24016 ^ n24014;
  assign n26630 = n26629 ^ n24017;
  assign n26621 = n26558 & n26573;
  assign n26624 = n26623 ^ n26621;
  assign n26628 = n26627 ^ n26624;
  assign n26631 = n26630 ^ n26628;
  assign n26633 = n26632 ^ n26631;
  assign n18455 = n18454 ^ n14280;
  assign n20867 = n20866 ^ n18455;
  assign n24018 = n24017 ^ n20867;
  assign n26634 = n26633 ^ n24018;
  assign n18456 = n18455 ^ n16853;
  assign n22884 = n20867 ^ n18456;
  assign n26110 = n24018 ^ n22884;
  assign n26635 = n26634 ^ n26110;
  assign n18458 = n18457 ^ n18456;
  assign n22885 = n22884 ^ n18458;
  assign n26111 = n26110 ^ n22885;
  assign n26636 = n26635 ^ n26111;
  assign n26644 = n26643 ^ n26636;
  assign n26655 = n26654 ^ n26644;
  assign n26719 = n26683 ^ n26655;
  assign n26662 = n26535 & n26588;
  assign n26598 = n26597 ^ n26596;
  assign n26663 = n26662 ^ n26598;
  assign n26660 = n26659 ^ n26624;
  assign n23980 = n23829 & n23874;
  assign n23899 = n23898 ^ n23897;
  assign n23981 = n23980 ^ n23899;
  assign n23978 = n23977 ^ n23973;
  assign n20833 = n20622 & n20683;
  assign n20787 = n20786 ^ n20746;
  assign n20834 = n20833 ^ n20787;
  assign n20831 = n20830 ^ n20744;
  assign n18657 = n18310 & n18357;
  assign n18535 = n18534 ^ n18379;
  assign n18658 = n18657 ^ n18535;
  assign n18655 = n18566 ^ n18444;
  assign n18654 = n18495 ^ n14394;
  assign n18656 = n18655 ^ n18654;
  assign n18659 = n18658 ^ n18656;
  assign n20828 = n20689 ^ n18659;
  assign n20832 = n20831 ^ n20828;
  assign n20835 = n20834 ^ n20832;
  assign n23968 = n23895 ^ n20835;
  assign n23979 = n23978 ^ n23968;
  assign n23982 = n23981 ^ n23979;
  assign n26658 = n26594 ^ n23982;
  assign n26661 = n26660 ^ n26658;
  assign n26664 = n26663 ^ n26661;
  assign n18660 = n18659 ^ n14395;
  assign n20836 = n20835 ^ n18660;
  assign n23983 = n23982 ^ n20836;
  assign n26665 = n26664 ^ n23983;
  assign n18661 = n18660 ^ n16848;
  assign n22881 = n20836 ^ n18661;
  assign n26107 = n23983 ^ n22881;
  assign n26666 = n26665 ^ n26107;
  assign n18663 = n18662 ^ n18661;
  assign n22882 = n22881 ^ n18663;
  assign n26108 = n26107 ^ n22882;
  assign n26667 = n26666 ^ n26108;
  assign n26614 = n26613 ^ n26598;
  assign n26610 = n26600 ^ n26594;
  assign n26615 = n26614 ^ n26610;
  assign n24040 = n24039 ^ n23899;
  assign n24038 = n23901 ^ n23895;
  assign n24041 = n24040 ^ n24038;
  assign n20790 = n20789 ^ n20787;
  assign n20785 = n20784 ^ n20689;
  assign n20791 = n20790 ^ n20785;
  assign n18626 = n18535 ^ n18377;
  assign n18625 = n18495 ^ n18359;
  assign n18627 = n18626 ^ n18625;
  assign n18628 = n18627 ^ n14412;
  assign n20792 = n20791 ^ n18628;
  assign n24042 = n24041 ^ n20792;
  assign n26616 = n26615 ^ n24042;
  assign n18629 = n18628 ^ n14413;
  assign n20793 = n20792 ^ n18629;
  assign n24043 = n24042 ^ n20793;
  assign n26617 = n26616 ^ n24043;
  assign n18630 = n18629 ^ n16860;
  assign n22901 = n20793 ^ n18630;
  assign n26127 = n24043 ^ n22901;
  assign n26618 = n26617 ^ n26127;
  assign n18632 = n18631 ^ n18630;
  assign n22902 = n22901 ^ n18632;
  assign n26128 = n26127 ^ n22902;
  assign n26619 = n26618 ^ n26128;
  assign n26691 = n26667 ^ n26619;
  assign n26720 = n26719 ^ n26691;
  assign n26708 = ~n26655 & n26683;
  assign n26672 = n26646 ^ n26622;
  assign n26670 = n26602 ^ n26598;
  assign n24114 = n24099 ^ n23975;
  assign n24112 = n23903 ^ n23899;
  assign n20881 = n20697 ^ n20694;
  assign n20879 = n20878 ^ n20787;
  assign n18584 = n18498 ^ n18442;
  assign n18582 = n18535 ^ n18361;
  assign n18581 = n18382 ^ n14425;
  assign n18583 = n18582 ^ n18581;
  assign n18585 = n18584 ^ n18583;
  assign n20876 = n20688 ^ n18585;
  assign n20880 = n20879 ^ n20876;
  assign n20882 = n20881 ^ n20880;
  assign n24111 = n23892 ^ n20882;
  assign n24113 = n24112 ^ n24111;
  assign n24115 = n24114 ^ n24113;
  assign n26669 = n26593 ^ n24115;
  assign n26671 = n26670 ^ n26669;
  assign n26673 = n26672 ^ n26671;
  assign n18586 = n18585 ^ n14426;
  assign n20883 = n20882 ^ n18586;
  assign n24116 = n24115 ^ n20883;
  assign n26674 = n26673 ^ n24116;
  assign n18587 = n18586 ^ n16836;
  assign n22887 = n20883 ^ n18587;
  assign n26113 = n24116 ^ n22887;
  assign n26675 = n26674 ^ n26113;
  assign n18589 = n18588 ^ n18587;
  assign n22888 = n22887 ^ n18589;
  assign n26114 = n26113 ^ n22888;
  assign n26676 = n26675 ^ n26114;
  assign n26684 = n26683 ^ n26676;
  assign n26668 = n26667 ^ n26636;
  assign n26685 = n26684 ^ n26668;
  assign n26688 = n26683 ^ n26619;
  assign n26689 = n26685 & ~n26688;
  assign n26709 = n26708 ^ n26689;
  assign n26706 = n26688 ^ n26685;
  assign n26605 = n26604 ^ n26598;
  assign n23906 = n23905 ^ n23899;
  assign n20929 = n20928 ^ n20787;
  assign n18536 = n18535 ^ n18363;
  assign n18533 = n18495 ^ n14464;
  assign n18537 = n18536 ^ n18533;
  assign n20927 = n20689 ^ n18537;
  assign n20930 = n20929 ^ n20927;
  assign n23896 = n23895 ^ n20930;
  assign n23907 = n23906 ^ n23896;
  assign n26595 = n26594 ^ n23907;
  assign n26606 = n26605 ^ n26595;
  assign n18538 = n18537 ^ n14465;
  assign n20931 = n20930 ^ n18538;
  assign n23908 = n23907 ^ n20931;
  assign n26607 = n26606 ^ n23908;
  assign n18539 = n18538 ^ n16868;
  assign n22879 = n20931 ^ n18539;
  assign n26105 = n23908 ^ n22879;
  assign n26608 = n26607 ^ n26105;
  assign n18541 = n18540 ^ n18539;
  assign n22880 = n22879 ^ n18541;
  assign n26106 = n26105 ^ n22880;
  assign n26609 = n26608 ^ n26106;
  assign n26702 = n26667 ^ n26609;
  assign n26620 = n26619 ^ n26609;
  assign n26703 = n26668 ^ n26620;
  assign n26704 = n26702 & ~n26703;
  assign n26695 = n26667 ^ n26643;
  assign n26696 = n26695 ^ n26684;
  assign n26697 = n26620 & n26696;
  assign n26705 = n26704 ^ n26697;
  assign n26707 = n26706 ^ n26705;
  assign n26710 = n26709 ^ n26707;
  assign n26692 = n26684 ^ n26620;
  assign n26724 = n26695 ^ n26692;
  assign n26725 = n26724 ^ n26705;
  assign n26721 = n26692 ^ n26654;
  assign n26722 = n26720 & n26721;
  assign n26713 = n26702 ^ n26688;
  assign n26714 = ~n26692 & ~n26713;
  assign n26723 = n26722 ^ n26714;
  assign n26726 = n26725 ^ n26723;
  assign n26727 = ~n26710 & n26726;
  assign n26686 = n26685 ^ n26655;
  assign n26656 = n26655 ^ n26609;
  assign n26657 = n26656 ^ n26620;
  assign n26700 = n26686 ^ n26657;
  assign n26693 = n26692 ^ n26644;
  assign n26694 = n26691 & ~n26693;
  assign n26698 = n26697 ^ n26694;
  assign n26687 = ~n26657 & ~n26686;
  assign n26690 = n26689 ^ n26687;
  assign n26699 = n26698 ^ n26690;
  assign n26701 = n26700 ^ n26699;
  assign n26711 = n26710 ^ n26701;
  assign n26743 = n26727 ^ n26711;
  assign n26716 = n26693 ^ n26691;
  assign n26712 = ~n26654 & ~n26656;
  assign n26715 = n26714 ^ n26712;
  assign n26717 = n26716 ^ n26715;
  assign n26718 = n26717 ^ n26698;
  assign n26741 = ~n26710 & ~n26718;
  assign n26742 = ~n26701 & n26741;
  assign n26744 = n26743 ^ n26742;
  assign n26759 = n26720 & ~n26744;
  assign n26738 = n26718 & n26726;
  assign n26739 = n26701 & n26738;
  assign n26731 = n26726 ^ n26718;
  assign n26737 = n26731 ^ n26727;
  assign n26740 = n26739 ^ n26737;
  assign n26758 = ~n26655 & ~n26740;
  assign n26760 = n26759 ^ n26758;
  assign n26745 = n26744 ^ n26740;
  assign n26732 = n26727 ^ n26701;
  assign n26733 = ~n26731 & n26732;
  assign n26734 = n26733 ^ n26718;
  assign n26728 = n26727 ^ n26718;
  assign n26729 = ~n26711 & ~n26728;
  assign n26730 = n26729 ^ n26701;
  assign n26735 = n26734 ^ n26730;
  assign n26746 = n26745 ^ n26735;
  assign n26756 = ~n26703 & ~n26746;
  assign n26755 = n26696 & ~n26735;
  assign n26757 = n26756 ^ n26755;
  assign n26761 = n26760 ^ n26757;
  assign n26752 = n26744 ^ n26730;
  assign n26753 = ~n26713 & ~n26752;
  assign n26749 = n26740 ^ n26734;
  assign n26750 = n26685 & n26749;
  assign n26747 = n26702 & ~n26746;
  assign n26736 = n26620 & ~n26735;
  assign n26748 = n26747 ^ n26736;
  assign n26751 = n26750 ^ n26748;
  assign n26754 = n26753 ^ n26751;
  assign n26762 = n26761 ^ n26754;
  assign n26139 = n26120 ^ n26108;
  assign n26117 = n26116 ^ n26114;
  assign n26140 = n26139 ^ n26117;
  assign n26129 = n26128 ^ n26106;
  assign n26136 = n26129 ^ n26117;
  assign n26121 = n26120 ^ n26111;
  assign n26137 = n26136 ^ n26121;
  assign n26135 = n26128 ^ n26108;
  assign n26161 = n26137 ^ n26135;
  assign n26124 = n26123 ^ n26121;
  assign n26126 = n26124 ^ n26106;
  assign n26159 = n26123 & n26126;
  assign n26132 = n26128 ^ n26116;
  assign n26109 = n26108 ^ n26106;
  assign n26146 = n26132 ^ n26109;
  assign n26147 = n26136 & n26146;
  assign n26160 = n26159 ^ n26147;
  assign n26162 = n26161 ^ n26160;
  assign n26141 = n26129 & n26140;
  assign n26138 = n26135 & n26137;
  assign n26142 = n26141 ^ n26138;
  assign n26163 = n26162 ^ n26142;
  assign n26156 = n26139 ^ n26136;
  assign n26112 = n26111 ^ n26108;
  assign n26153 = n26129 ^ n26112;
  assign n26154 = n26109 & n26153;
  assign n26155 = n26154 ^ n26141;
  assign n26157 = n26156 ^ n26155;
  assign n26148 = n26124 ^ n26116;
  assign n26149 = n26148 ^ n26135;
  assign n26150 = n26136 ^ n26123;
  assign n26151 = n26149 & n26150;
  assign n26152 = n26151 ^ n26147;
  assign n26158 = n26157 ^ n26152;
  assign n26172 = n26163 ^ n26158;
  assign n26168 = ~n26116 & n26124;
  assign n26118 = n26117 ^ n26112;
  assign n26133 = n26118 & n26132;
  assign n26169 = n26168 ^ n26133;
  assign n26166 = n26132 ^ n26118;
  assign n26167 = n26166 ^ n26155;
  assign n26170 = n26169 ^ n26167;
  assign n26171 = n26158 & n26170;
  assign n26130 = n26129 ^ n26126;
  assign n26125 = n26124 ^ n26118;
  assign n26144 = n26130 ^ n26125;
  assign n26131 = n26125 & n26130;
  assign n26134 = n26133 ^ n26131;
  assign n26143 = n26142 ^ n26134;
  assign n26145 = n26144 ^ n26143;
  assign n26184 = n26171 ^ n26145;
  assign n26185 = n26172 & n26184;
  assign n26186 = n26185 ^ n26163;
  assign n26177 = n26170 ^ n26145;
  assign n26181 = n26171 ^ n26163;
  assign n26182 = n26177 & n26181;
  assign n26183 = n26182 ^ n26145;
  assign n26187 = n26186 ^ n26183;
  assign n26360 = n26140 & n26187;
  assign n26178 = n26177 ^ n26171;
  assign n26175 = n26163 & n26170;
  assign n26176 = ~n26145 & n26175;
  assign n26179 = n26178 ^ n26176;
  assign n26173 = n26172 ^ n26171;
  assign n26164 = n26158 & ~n26163;
  assign n26165 = n26145 & n26164;
  assign n26174 = n26173 ^ n26165;
  assign n26180 = n26179 ^ n26174;
  assign n26188 = n26187 ^ n26180;
  assign n26199 = n26153 & n26188;
  assign n26361 = n26360 ^ n26199;
  assign n26211 = n26149 & n26179;
  assign n26210 = n26124 & n26174;
  assign n26212 = n26211 ^ n26210;
  assign n26362 = n26361 ^ n26212;
  assign n26202 = n26183 ^ n26179;
  assign n26269 = n26146 & n26202;
  assign n26192 = n26186 ^ n26174;
  assign n26193 = n26118 & n26192;
  assign n26190 = n26129 & n26187;
  assign n26189 = n26109 & n26188;
  assign n26191 = n26190 ^ n26189;
  assign n26194 = n26193 ^ n26191;
  assign n26359 = n26269 ^ n26194;
  assign n26363 = n26362 ^ n26359;
  assign n22913 = n22894 ^ n22882;
  assign n22891 = n22890 ^ n22888;
  assign n22914 = n22913 ^ n22891;
  assign n22903 = n22902 ^ n22880;
  assign n22910 = n22903 ^ n22891;
  assign n22895 = n22894 ^ n22885;
  assign n22911 = n22910 ^ n22895;
  assign n22909 = n22902 ^ n22882;
  assign n22935 = n22911 ^ n22909;
  assign n22898 = n22897 ^ n22895;
  assign n22900 = n22898 ^ n22880;
  assign n22933 = n22897 & n22900;
  assign n22906 = n22902 ^ n22890;
  assign n22883 = n22882 ^ n22880;
  assign n22920 = n22906 ^ n22883;
  assign n22921 = n22910 & n22920;
  assign n22934 = n22933 ^ n22921;
  assign n22936 = n22935 ^ n22934;
  assign n22915 = n22903 & n22914;
  assign n22912 = n22909 & n22911;
  assign n22916 = n22915 ^ n22912;
  assign n22937 = n22936 ^ n22916;
  assign n22930 = n22913 ^ n22910;
  assign n22886 = n22885 ^ n22882;
  assign n22927 = n22903 ^ n22886;
  assign n22928 = n22883 & n22927;
  assign n22929 = n22928 ^ n22915;
  assign n22931 = n22930 ^ n22929;
  assign n22922 = n22910 ^ n22897;
  assign n22923 = n22898 ^ n22890;
  assign n22924 = n22923 ^ n22909;
  assign n22925 = n22922 & n22924;
  assign n22926 = n22925 ^ n22921;
  assign n22932 = n22931 ^ n22926;
  assign n22946 = n22937 ^ n22932;
  assign n22942 = ~n22890 & n22898;
  assign n22892 = n22891 ^ n22886;
  assign n22907 = n22892 & n22906;
  assign n22943 = n22942 ^ n22907;
  assign n22940 = n22906 ^ n22892;
  assign n22941 = n22940 ^ n22929;
  assign n22944 = n22943 ^ n22941;
  assign n22945 = n22932 & n22944;
  assign n22904 = n22903 ^ n22900;
  assign n22899 = n22898 ^ n22892;
  assign n22918 = n22904 ^ n22899;
  assign n22905 = n22899 & n22904;
  assign n22908 = n22907 ^ n22905;
  assign n22917 = n22916 ^ n22908;
  assign n22919 = n22918 ^ n22917;
  assign n22958 = n22945 ^ n22919;
  assign n22959 = n22946 & n22958;
  assign n22960 = n22959 ^ n22937;
  assign n22951 = n22944 ^ n22919;
  assign n22955 = n22945 ^ n22937;
  assign n22956 = n22951 & n22955;
  assign n22957 = n22956 ^ n22919;
  assign n22961 = n22960 ^ n22957;
  assign n23034 = n22914 & n22961;
  assign n22952 = n22951 ^ n22945;
  assign n22949 = n22937 & n22944;
  assign n22950 = ~n22919 & n22949;
  assign n22953 = n22952 ^ n22950;
  assign n22947 = n22946 ^ n22945;
  assign n22938 = n22932 & ~n22937;
  assign n22939 = n22919 & n22938;
  assign n22948 = n22947 ^ n22939;
  assign n22954 = n22953 ^ n22948;
  assign n22962 = n22961 ^ n22954;
  assign n22973 = n22927 & n22962;
  assign n23102 = n23034 ^ n22973;
  assign n22985 = n22924 & n22953;
  assign n22984 = n22898 & n22948;
  assign n22986 = n22985 ^ n22984;
  assign n23103 = n23102 ^ n22986;
  assign n22976 = n22957 ^ n22953;
  assign n23077 = n22920 & n22976;
  assign n22966 = n22960 ^ n22948;
  assign n22967 = n22892 & n22966;
  assign n22964 = n22903 & n22961;
  assign n22963 = n22883 & n22962;
  assign n22965 = n22964 ^ n22963;
  assign n22968 = n22967 ^ n22965;
  assign n23101 = n23077 ^ n22968;
  assign n23104 = n23103 ^ n23101;
  assign n21561 = n18663 ^ n18389;
  assign n21556 = n18589 ^ n18574;
  assign n21562 = n21561 ^ n21556;
  assign n21558 = n18458 ^ n18389;
  assign n21565 = n21558 ^ n18506;
  assign n21599 = ~n18574 & n21565;
  assign n21553 = n18632 ^ n18574;
  assign n21580 = n18663 ^ n18458;
  assign n21588 = n21580 ^ n21556;
  assign n21592 = n21553 & n21588;
  assign n21600 = n21599 ^ n21592;
  assign n21597 = n21588 ^ n21553;
  assign n21568 = n18663 ^ n18541;
  assign n21555 = n18632 ^ n18541;
  assign n21581 = n21580 ^ n21555;
  assign n21582 = n21568 & n21581;
  assign n21563 = n21555 & n21562;
  assign n21583 = n21582 ^ n21563;
  assign n21598 = n21597 ^ n21583;
  assign n21601 = n21600 ^ n21598;
  assign n21566 = n21565 ^ n18541;
  assign n21590 = n21566 ^ n21555;
  assign n21589 = n21588 ^ n21565;
  assign n21595 = n21590 ^ n21589;
  assign n21591 = n21589 & n21590;
  assign n21593 = n21592 ^ n21591;
  assign n21554 = n18663 ^ n18632;
  assign n21557 = n21556 ^ n21555;
  assign n21559 = n21558 ^ n21557;
  assign n21560 = n21554 & n21559;
  assign n21564 = n21563 ^ n21560;
  assign n21594 = n21593 ^ n21564;
  assign n21596 = n21595 ^ n21594;
  assign n21614 = n21601 ^ n21596;
  assign n21584 = n21561 ^ n21557;
  assign n21585 = n21584 ^ n21583;
  assign n21575 = n21565 ^ n18574;
  assign n21576 = n21575 ^ n21554;
  assign n21577 = n21557 ^ n18506;
  assign n21578 = n21576 & n21577;
  assign n21569 = n21568 ^ n21553;
  assign n21570 = n21557 & n21569;
  assign n21579 = n21578 ^ n21570;
  assign n21586 = n21585 ^ n21579;
  assign n21602 = n21586 & n21601;
  assign n21572 = n21559 ^ n21554;
  assign n21567 = n18506 & n21566;
  assign n21571 = n21570 ^ n21567;
  assign n21573 = n21572 ^ n21571;
  assign n21574 = n21573 ^ n21564;
  assign n21620 = n21602 ^ n21574;
  assign n21621 = n21614 & n21620;
  assign n21622 = n21621 ^ n21596;
  assign n21587 = n21586 ^ n21574;
  assign n21603 = n21602 ^ n21596;
  assign n21604 = n21587 & n21603;
  assign n21605 = n21604 ^ n21574;
  assign n21623 = n21622 ^ n21605;
  assign n21779 = n21562 & n21623;
  assign n21615 = n21614 ^ n21602;
  assign n21612 = n21574 & n21601;
  assign n21613 = ~n21596 & n21612;
  assign n21616 = n21615 ^ n21613;
  assign n21608 = n21602 ^ n21587;
  assign n21606 = ~n21574 & n21586;
  assign n21607 = n21596 & n21606;
  assign n21609 = n21608 ^ n21607;
  assign n21617 = n21616 ^ n21609;
  assign n21624 = n21623 ^ n21617;
  assign n21625 = n21581 & n21624;
  assign n21807 = n21779 ^ n21625;
  assign n21695 = n21576 & n21616;
  assign n21634 = n21565 & n21609;
  assign n21696 = n21695 ^ n21634;
  assign n21857 = n21807 ^ n21696;
  assign n21610 = n21609 ^ n21605;
  assign n21716 = n21588 & n21610;
  assign n21632 = n21555 & n21623;
  assign n21631 = n21568 & n21624;
  assign n21633 = n21632 ^ n21631;
  assign n21717 = n21716 ^ n21633;
  assign n21692 = n21622 ^ n21616;
  assign n21693 = n21569 & n21692;
  assign n21856 = n21717 ^ n21693;
  assign n21858 = n21857 ^ n21856;
  assign n21859 = n21858 ^ n19452;
  assign n23105 = n23104 ^ n21859;
  assign n26364 = n26363 ^ n23105;
  assign n26763 = n26762 ^ n26364;
  assign n26431 = n26360 ^ n26190;
  assign n26428 = n26135 & n26180;
  assign n23035 = n23034 ^ n22964;
  assign n23031 = n22909 & n22954;
  assign n21780 = n21779 ^ n21632;
  assign n21776 = n21554 & n21617;
  assign n21777 = n21776 ^ n19302;
  assign n21721 = n21590 & n21605;
  assign n21719 = n21557 & n21692;
  assign n21699 = n18506 & n21622;
  assign n21720 = n21719 ^ n21699;
  assign n21722 = n21721 ^ n21720;
  assign n21618 = n21559 & n21617;
  assign n21611 = n21553 & n21610;
  assign n21619 = n21618 ^ n21611;
  assign n21775 = n21722 ^ n21619;
  assign n21778 = n21777 ^ n21775;
  assign n21781 = n21780 ^ n21778;
  assign n23032 = n23031 ^ n21781;
  assign n22978 = n22897 & n22957;
  assign n22977 = n22910 & n22976;
  assign n22979 = n22978 ^ n22977;
  assign n22975 = n22904 & n22960;
  assign n22980 = n22979 ^ n22975;
  assign n22971 = n22906 & n22966;
  assign n22970 = n22911 & n22954;
  assign n22972 = n22971 ^ n22970;
  assign n23030 = n22980 ^ n22972;
  assign n23033 = n23032 ^ n23030;
  assign n23036 = n23035 ^ n23033;
  assign n26429 = n26428 ^ n23036;
  assign n26204 = n26123 & n26183;
  assign n26203 = n26136 & n26202;
  assign n26205 = n26204 ^ n26203;
  assign n26201 = n26130 & n26186;
  assign n26206 = n26205 ^ n26201;
  assign n26197 = n26132 & n26192;
  assign n26196 = n26137 & n26180;
  assign n26198 = n26197 ^ n26196;
  assign n26427 = n26206 ^ n26198;
  assign n26430 = n26429 ^ n26427;
  assign n26432 = n26431 ^ n26430;
  assign n23741 = n21781 ^ n19303;
  assign n24279 = n23741 ^ n19304;
  assign n25444 = n24279 ^ n21965;
  assign n21725 = n21566 & n21622;
  assign n21726 = n21725 ^ n21696;
  assign n21626 = n21625 ^ n21619;
  assign n21723 = n21722 ^ n21626;
  assign n21718 = n21717 ^ n19379;
  assign n21724 = n21723 ^ n21718;
  assign n21727 = n21726 ^ n21724;
  assign n23727 = n21727 ^ n19380;
  assign n24244 = n23727 ^ n19381;
  assign n25414 = n24244 ^ n21982;
  assign n25668 = n25444 ^ n25414;
  assign n23692 = n21859 ^ n19453;
  assign n24288 = n23692 ^ n19454;
  assign n25452 = n24288 ^ n21988;
  assign n21691 = n21577 & n21616;
  assign n21694 = n21693 ^ n21691;
  assign n21806 = n21719 ^ n21694;
  assign n21847 = n21806 ^ n21696;
  assign n21846 = n21717 ^ n19426;
  assign n21848 = n21847 ^ n21846;
  assign n23698 = n21848 ^ n19427;
  assign n24275 = n23698 ^ n19428;
  assign n25440 = n24275 ^ n21995;
  assign n25664 = n25452 ^ n25440;
  assign n25671 = n25668 ^ n25664;
  assign n21809 = n21695 ^ n21633;
  assign n21808 = n21807 ^ n21806;
  assign n21810 = n21809 ^ n21808;
  assign n21811 = n21810 ^ n19479;
  assign n23732 = n21811 ^ n19480;
  assign n24248 = n23732 ^ n19481;
  assign n25418 = n24248 ^ n21961;
  assign n25679 = n25444 ^ n25418;
  assign n21628 = n21589 & n21605;
  assign n21700 = n21699 ^ n21628;
  assign n21697 = n21696 ^ n21694;
  assign n21690 = n21633 ^ n19561;
  assign n21698 = n21697 ^ n21690;
  assign n21701 = n21700 ^ n21698;
  assign n23712 = n21701 ^ n19562;
  assign n24262 = n23712 ^ n19563;
  assign n25429 = n24262 ^ n21977;
  assign n21635 = n21634 ^ n21633;
  assign n21627 = n21575 & n21609;
  assign n21629 = n21628 ^ n21627;
  assign n21630 = n21629 ^ n21626;
  assign n21636 = n21635 ^ n21630;
  assign n21637 = n21636 ^ n19534;
  assign n23705 = n21637 ^ n19535;
  assign n24255 = n23705 ^ n19536;
  assign n25424 = n24255 ^ n21957;
  assign n25665 = n25429 ^ n25424;
  assign n25666 = n25665 ^ n25664;
  assign n25702 = n25679 ^ n25666;
  assign n25687 = n25452 ^ n25414;
  assign n25712 = n25702 ^ n25687;
  assign n21796 = n21720 ^ n21629;
  assign n21795 = n21717 ^ n21611;
  assign n21797 = n21796 ^ n21795;
  assign n21798 = n21797 ^ n19509;
  assign n23720 = n21798 ^ n19510;
  assign n24269 = n23720 ^ n19511;
  assign n25435 = n24269 ^ n21969;
  assign n25680 = n25679 ^ n25435;
  assign n25698 = n25680 ^ n25440;
  assign n25710 = n25435 & ~n25698;
  assign n25672 = n25440 ^ n25414;
  assign n25667 = n25452 ^ n25424;
  assign n25690 = n25672 ^ n25667;
  assign n25691 = n25666 & ~n25690;
  assign n25711 = n25710 ^ n25691;
  assign n25713 = n25712 ^ n25711;
  assign n25703 = ~n25687 & ~n25702;
  assign n25674 = n25418 ^ n25414;
  assign n25675 = n25674 ^ n25665;
  assign n25676 = n25664 & n25675;
  assign n25704 = n25703 ^ n25676;
  assign n25714 = n25713 ^ n25704;
  assign n25693 = n25674 ^ n25666;
  assign n25673 = ~n25671 & ~n25672;
  assign n25677 = n25676 ^ n25673;
  assign n25694 = n25693 ^ n25677;
  assign n25685 = n25666 ^ n25435;
  assign n25686 = n25680 ^ n25424;
  assign n25688 = n25687 ^ n25686;
  assign n25689 = n25685 & n25688;
  assign n25692 = n25691 ^ n25689;
  assign n25695 = n25694 ^ n25692;
  assign n25725 = n25714 ^ n25695;
  assign n25699 = n25698 ^ n25664;
  assign n25669 = n25668 ^ n25665;
  assign n25697 = n25680 ^ n25669;
  assign n25706 = n25699 ^ n25697;
  assign n25700 = n25697 & ~n25699;
  assign n25682 = n25667 & ~n25669;
  assign n25701 = n25700 ^ n25682;
  assign n25705 = n25704 ^ n25701;
  assign n25707 = n25706 ^ n25705;
  assign n25681 = ~n25424 & ~n25680;
  assign n25683 = n25682 ^ n25681;
  assign n25670 = n25669 ^ n25667;
  assign n25678 = n25677 ^ n25670;
  assign n25684 = n25683 ^ n25678;
  assign n25696 = ~n25684 & n25695;
  assign n25726 = n25707 ^ n25696;
  assign n25727 = n25725 & ~n25726;
  assign n25728 = n25727 ^ n25714;
  assign n25708 = n25707 ^ n25684;
  assign n25718 = n25714 ^ n25696;
  assign n25719 = n25708 & n25718;
  assign n25720 = n25719 ^ n25707;
  assign n25744 = n25728 ^ n25720;
  assign n25733 = n25725 ^ n25696;
  assign n25731 = n25695 & ~n25714;
  assign n25732 = ~n25707 & n25731;
  assign n25734 = n25733 ^ n25732;
  assign n25715 = ~n25684 & n25714;
  assign n25716 = n25707 & n25715;
  assign n25709 = n25708 ^ n25696;
  assign n25717 = n25716 ^ n25709;
  assign n25737 = n25734 ^ n25717;
  assign n25811 = n25744 ^ n25737;
  assign n25812 = ~n25671 & ~n25811;
  assign n25745 = n25675 & ~n25744;
  assign n25898 = n25812 ^ n25745;
  assign n25822 = ~n25680 & n25734;
  assign n25821 = n25688 & n25717;
  assign n25823 = n25822 ^ n25821;
  assign n25899 = n25898 ^ n25823;
  assign n25721 = n25720 ^ n25717;
  assign n25869 = ~n25690 & ~n25721;
  assign n25735 = n25734 ^ n25728;
  assign n25817 = ~n25669 & n25735;
  assign n25815 = ~n25672 & ~n25811;
  assign n25746 = n25664 & ~n25744;
  assign n25816 = n25815 ^ n25746;
  assign n25818 = n25817 ^ n25816;
  assign n25897 = n25869 ^ n25818;
  assign n25900 = n25899 ^ n25897;
  assign n25901 = n25900 ^ n22743;
  assign n25902 = n25901 ^ n22744;
  assign n25903 = n25902 ^ n22745;
  assign n25904 = n25903 ^ n22746;
  assign n3074 = x193 ^ x65;
  assign n3073 = x194 ^ x66;
  assign n3075 = n3074 ^ n3073;
  assign n3072 = x199 ^ x71;
  assign n3076 = n3075 ^ n3072;
  assign n3069 = x197 ^ x69;
  assign n3095 = n3074 ^ n3069;
  assign n3084 = x195 ^ x67;
  assign n3068 = x192 ^ x64;
  assign n3086 = n3084 ^ n3068;
  assign n3079 = x196 ^ x68;
  assign n3071 = x198 ^ x70;
  assign n3080 = n3079 ^ n3071;
  assign n3092 = n3086 ^ n3080;
  assign n3124 = n3095 ^ n3092;
  assign n3103 = n3084 ^ n3069;
  assign n3081 = n3073 ^ n3069;
  assign n3104 = n3086 ^ n3081;
  assign n3105 = n3103 & n3104;
  assign n3096 = n3095 ^ n3080;
  assign n3097 = n3086 & n3096;
  assign n3106 = n3105 ^ n3097;
  assign n3125 = n3124 ^ n3106;
  assign n3077 = n3076 ^ n3071;
  assign n3070 = n3069 ^ n3068;
  assign n3078 = n3077 ^ n3070;
  assign n3121 = n3092 ^ n3072;
  assign n3122 = n3078 & n3121;
  assign n3089 = n3071 ^ n3068;
  assign n3112 = n3103 ^ n3089;
  assign n3113 = n3092 & n3112;
  assign n3123 = n3122 ^ n3113;
  assign n3126 = n3125 ^ n3123;
  assign n3093 = n3092 ^ n3075;
  assign n3115 = n3093 ^ n3070;
  assign n3085 = n3084 ^ n3076;
  assign n3111 = n3072 & n3085;
  assign n3114 = n3113 ^ n3111;
  assign n3116 = n3115 ^ n3114;
  assign n3094 = n3070 & n3093;
  assign n3098 = n3097 ^ n3094;
  assign n3117 = n3116 ^ n3098;
  assign n3133 = n3126 ^ n3117;
  assign n3108 = ~n3071 & n3076;
  assign n3082 = n3081 ^ n3080;
  assign n3090 = n3082 & n3089;
  assign n3109 = n3108 ^ n3090;
  assign n3102 = n3089 ^ n3082;
  assign n3107 = n3106 ^ n3102;
  assign n3110 = n3109 ^ n3107;
  assign n3127 = n3110 & n3126;
  assign n3134 = n3133 ^ n3127;
  assign n3087 = n3086 ^ n3085;
  assign n3083 = n3082 ^ n3076;
  assign n3100 = n3087 ^ n3083;
  assign n3088 = n3083 & n3087;
  assign n3091 = n3090 ^ n3088;
  assign n3099 = n3098 ^ n3091;
  assign n3101 = n3100 ^ n3099;
  assign n3131 = ~n3117 & n3126;
  assign n3132 = n3101 & n3131;
  assign n3135 = n3134 ^ n3132;
  assign n3204 = n3076 & n3135;
  assign n3120 = n3110 ^ n3101;
  assign n3128 = n3127 ^ n3120;
  assign n3118 = n3110 & n3117;
  assign n3119 = ~n3101 & n3118;
  assign n3129 = n3128 ^ n3119;
  assign n3130 = n3078 & n3129;
  assign n3205 = n3204 ^ n3130;
  assign n3140 = n3127 ^ n3117;
  assign n3141 = n3120 & n3140;
  assign n3142 = n3141 ^ n3101;
  assign n3137 = n3127 ^ n3101;
  assign n3138 = n3133 & n3137;
  assign n3139 = n3138 ^ n3117;
  assign n3143 = n3142 ^ n3139;
  assign n3136 = n3135 ^ n3129;
  assign n3144 = n3143 ^ n3136;
  assign n3156 = n3104 & n3144;
  assign n3155 = n3096 & n3143;
  assign n3157 = n3156 ^ n3155;
  assign n3206 = n3205 ^ n3157;
  assign n3191 = n3139 ^ n3135;
  assign n3192 = n3082 & n3191;
  assign n3146 = n3086 & n3143;
  assign n3145 = n3103 & n3144;
  assign n3147 = n3146 ^ n3145;
  assign n3193 = n3192 ^ n3147;
  assign n3150 = n3142 ^ n3129;
  assign n3151 = n3112 & n3150;
  assign n3203 = n3193 ^ n3151;
  assign n3207 = n3206 ^ n3203;
  assign n2997 = x239 ^ x111;
  assign n2986 = x234 ^ x106;
  assign n2985 = x233 ^ x105;
  assign n2987 = n2986 ^ n2985;
  assign n2998 = n2997 ^ n2987;
  assign n2974 = x237 ^ x109;
  assign n2991 = n2985 ^ n2974;
  assign n2978 = x232 ^ x104;
  assign n2975 = x235 ^ x107;
  assign n2983 = n2978 ^ n2975;
  assign n2981 = x236 ^ x108;
  assign n2977 = x238 ^ x110;
  assign n2982 = n2981 ^ n2977;
  assign n2984 = n2983 ^ n2982;
  assign n3028 = n2991 ^ n2984;
  assign n2976 = n2975 ^ n2974;
  assign n2995 = n2986 ^ n2974;
  assign n3008 = n2995 ^ n2983;
  assign n3009 = n2976 & n3008;
  assign n2992 = n2991 ^ n2982;
  assign n2993 = n2983 & n2992;
  assign n3010 = n3009 ^ n2993;
  assign n3029 = n3028 ^ n3010;
  assign n3023 = n2997 ^ n2984;
  assign n3024 = n2998 ^ n2977;
  assign n2989 = n2978 ^ n2974;
  assign n3025 = n3024 ^ n2989;
  assign n3026 = n3023 & n3025;
  assign n2979 = n2978 ^ n2977;
  assign n2980 = n2979 ^ n2976;
  assign n3018 = n2980 & n2984;
  assign n3027 = n3026 ^ n3018;
  assign n3030 = n3029 ^ n3027;
  assign n2988 = n2987 ^ n2984;
  assign n3020 = n2989 ^ n2988;
  assign n3000 = n2998 ^ n2975;
  assign n3017 = n2997 & n3000;
  assign n3019 = n3018 ^ n3017;
  assign n3021 = n3020 ^ n3019;
  assign n2990 = n2988 & n2989;
  assign n2994 = n2993 ^ n2990;
  assign n3022 = n3021 ^ n2994;
  assign n3041 = n3030 ^ n3022;
  assign n3013 = ~n2977 & n2998;
  assign n2996 = n2995 ^ n2982;
  assign n3003 = n2979 & n2996;
  assign n3014 = n3013 ^ n3003;
  assign n3011 = n2996 ^ n2979;
  assign n3012 = n3011 ^ n3010;
  assign n3015 = n3014 ^ n3012;
  assign n3031 = n3015 & n3030;
  assign n3047 = n3041 ^ n3031;
  assign n3001 = n3000 ^ n2983;
  assign n2999 = n2998 ^ n2996;
  assign n3006 = n3001 ^ n2999;
  assign n3002 = n2999 & n3001;
  assign n3004 = n3003 ^ n3002;
  assign n3005 = n3004 ^ n2994;
  assign n3007 = n3006 ^ n3005;
  assign n3045 = ~n3022 & n3030;
  assign n3046 = n3007 & n3045;
  assign n3048 = n3047 ^ n3046;
  assign n3063 = n2998 & n3048;
  assign n3016 = n3015 ^ n3007;
  assign n3037 = n3031 ^ n3016;
  assign n3035 = n3015 & n3022;
  assign n3036 = ~n3007 & n3035;
  assign n3038 = n3037 ^ n3036;
  assign n3062 = n3025 & n3038;
  assign n3064 = n3063 ^ n3062;
  assign n3052 = n3048 ^ n3038;
  assign n3042 = n3031 ^ n3007;
  assign n3043 = n3041 & n3042;
  assign n3044 = n3043 ^ n3022;
  assign n3032 = n3031 ^ n3022;
  assign n3033 = n3016 & n3032;
  assign n3034 = n3033 ^ n3007;
  assign n3051 = n3044 ^ n3034;
  assign n3053 = n3052 ^ n3051;
  assign n3060 = n3008 & n3053;
  assign n3059 = n2992 & n3051;
  assign n3061 = n3060 ^ n3059;
  assign n3065 = n3064 ^ n3061;
  assign n3055 = n2983 & n3051;
  assign n3054 = n2976 & n3053;
  assign n3056 = n3055 ^ n3054;
  assign n3049 = n3048 ^ n3044;
  assign n3050 = n2996 & n3049;
  assign n3057 = n3056 ^ n3050;
  assign n3039 = n3038 ^ n3034;
  assign n3040 = n2980 & n3039;
  assign n3058 = n3057 ^ n3040;
  assign n3066 = n3065 ^ n3058;
  assign n3437 = n3207 ^ n3066;
  assign n2890 = x148 ^ x20;
  assign n2885 = x150 ^ x22;
  assign n2891 = n2890 ^ n2885;
  assign n2884 = x144 ^ x16;
  assign n2882 = x147 ^ x19;
  assign n2889 = n2884 ^ n2882;
  assign n2892 = n2891 ^ n2889;
  assign n2905 = x151 ^ x23;
  assign n2894 = x146 ^ x18;
  assign n2893 = x145 ^ x17;
  assign n2895 = n2894 ^ n2893;
  assign n2906 = n2905 ^ n2895;
  assign n2920 = ~n2885 & n2906;
  assign n2886 = n2885 ^ n2884;
  assign n2881 = x149 ^ x21;
  assign n2902 = n2894 ^ n2881;
  assign n2903 = n2902 ^ n2891;
  assign n2904 = n2886 & n2903;
  assign n2921 = n2920 ^ n2904;
  assign n2918 = n2903 ^ n2886;
  assign n2883 = n2882 ^ n2881;
  assign n2915 = n2902 ^ n2889;
  assign n2916 = n2883 & n2915;
  assign n2898 = n2893 ^ n2881;
  assign n2899 = n2898 ^ n2891;
  assign n2900 = n2889 & n2899;
  assign n2917 = n2916 ^ n2900;
  assign n2919 = n2918 ^ n2917;
  assign n2922 = n2921 ^ n2919;
  assign n2908 = n2906 ^ n2882;
  assign n2909 = n2908 ^ n2889;
  assign n2907 = n2906 ^ n2903;
  assign n2913 = n2909 ^ n2907;
  assign n2910 = n2907 & n2909;
  assign n2911 = n2910 ^ n2904;
  assign n2888 = n2884 ^ n2881;
  assign n2896 = n2895 ^ n2892;
  assign n2897 = n2888 & n2896;
  assign n2901 = n2900 ^ n2897;
  assign n2912 = n2911 ^ n2901;
  assign n2914 = n2913 ^ n2912;
  assign n2940 = n2922 ^ n2914;
  assign n2936 = n2898 ^ n2892;
  assign n2937 = n2936 ^ n2917;
  assign n2931 = n2905 ^ n2892;
  assign n2932 = n2906 ^ n2885;
  assign n2933 = n2932 ^ n2888;
  assign n2934 = n2931 & n2933;
  assign n2887 = n2886 ^ n2883;
  assign n2924 = n2887 & n2892;
  assign n2935 = n2934 ^ n2924;
  assign n2938 = n2937 ^ n2935;
  assign n2939 = n2922 & n2938;
  assign n2926 = n2896 ^ n2888;
  assign n2923 = n2905 & n2908;
  assign n2925 = n2924 ^ n2923;
  assign n2927 = n2926 ^ n2925;
  assign n2928 = n2927 ^ n2901;
  assign n2943 = n2939 ^ n2928;
  assign n2944 = n2940 & n2943;
  assign n2945 = n2944 ^ n2914;
  assign n2941 = n2940 ^ n2939;
  assign n2929 = n2922 & n2928;
  assign n2930 = ~n2914 & n2929;
  assign n2942 = n2941 ^ n2930;
  assign n2946 = n2945 ^ n2942;
  assign n3269 = n2892 & n2946;
  assign n3268 = n2905 & n2945;
  assign n3270 = n3269 ^ n3268;
  assign n2950 = n2938 ^ n2928;
  assign n2951 = n2950 ^ n2939;
  assign n2948 = ~n2928 & n2938;
  assign n2949 = n2914 & n2948;
  assign n2952 = n2951 ^ n2949;
  assign n3172 = n2932 & n2952;
  assign n2954 = n2939 ^ n2914;
  assign n2955 = n2950 & n2954;
  assign n2956 = n2955 ^ n2928;
  assign n3171 = n2907 & n2956;
  assign n3173 = n3172 ^ n3171;
  assign n3434 = n3270 ^ n3173;
  assign n2962 = n2956 ^ n2952;
  assign n3174 = n2886 & n2962;
  assign n2963 = n2903 & n2962;
  assign n2957 = n2956 ^ n2945;
  assign n2960 = n2889 & n2957;
  assign n2953 = n2952 ^ n2942;
  assign n2958 = n2957 ^ n2953;
  assign n2959 = n2883 & n2958;
  assign n2961 = n2960 ^ n2959;
  assign n2964 = n2963 ^ n2961;
  assign n3433 = n3174 ^ n2964;
  assign n3435 = n3434 ^ n3433;
  assign n3210 = n2997 & n3034;
  assign n3162 = n2984 & n3039;
  assign n3211 = n3210 ^ n3162;
  assign n3182 = n3024 & n3048;
  assign n3181 = n2999 & n3044;
  assign n3183 = n3182 ^ n3181;
  assign n3212 = n3211 ^ n3183;
  assign n3184 = n2979 & n3049;
  assign n3209 = n3184 ^ n3057;
  assign n3213 = n3212 ^ n3209;
  assign n3436 = n3435 ^ n3213;
  assign n3438 = n3437 ^ n3436;
  assign n2711 = x191 ^ x63;
  assign n2703 = x190 ^ x62;
  assign n2712 = x185 ^ x57;
  assign n2706 = x186 ^ x58;
  assign n2713 = n2712 ^ n2706;
  assign n2714 = n2713 ^ n2711;
  assign n2738 = ~n2703 & n2714;
  assign n2702 = x184 ^ x56;
  assign n2704 = n2703 ^ n2702;
  assign n2708 = x188 ^ x60;
  assign n2709 = n2708 ^ n2703;
  assign n2699 = x189 ^ x61;
  assign n2707 = n2706 ^ n2699;
  assign n2710 = n2709 ^ n2707;
  assign n2720 = n2704 & n2710;
  assign n2739 = n2738 ^ n2720;
  assign n2700 = x187 ^ x59;
  assign n2701 = n2700 ^ n2699;
  assign n2716 = n2702 ^ n2700;
  assign n2734 = n2716 ^ n2707;
  assign n2735 = n2701 & n2734;
  assign n2726 = n2712 ^ n2699;
  assign n2727 = n2726 ^ n2709;
  assign n2728 = n2716 & n2727;
  assign n2736 = n2735 ^ n2728;
  assign n2733 = n2710 ^ n2704;
  assign n2737 = n2736 ^ n2733;
  assign n2740 = n2739 ^ n2737;
  assign n2717 = n2714 ^ n2700;
  assign n2718 = n2717 ^ n2716;
  assign n2715 = n2714 ^ n2710;
  assign n2731 = n2718 ^ n2715;
  assign n2722 = n2716 ^ n2709;
  assign n2723 = n2722 ^ n2713;
  assign n2724 = n2702 ^ n2699;
  assign n2725 = n2723 & n2724;
  assign n2729 = n2728 ^ n2725;
  assign n2719 = n2715 & n2718;
  assign n2721 = n2720 ^ n2719;
  assign n2730 = n2729 ^ n2721;
  assign n2732 = n2731 ^ n2730;
  assign n2758 = n2740 ^ n2732;
  assign n2754 = n2726 ^ n2722;
  assign n2755 = n2754 ^ n2736;
  assign n2749 = n2722 ^ n2711;
  assign n2750 = n2714 ^ n2703;
  assign n2751 = n2750 ^ n2724;
  assign n2752 = n2749 & n2751;
  assign n2705 = n2704 ^ n2701;
  assign n2742 = n2705 & n2722;
  assign n2753 = n2752 ^ n2742;
  assign n2756 = n2755 ^ n2753;
  assign n2757 = n2740 & n2756;
  assign n2744 = n2724 ^ n2723;
  assign n2741 = n2711 & n2717;
  assign n2743 = n2742 ^ n2741;
  assign n2745 = n2744 ^ n2743;
  assign n2746 = n2745 ^ n2729;
  assign n2761 = n2757 ^ n2746;
  assign n2762 = n2758 & n2761;
  assign n2763 = n2762 ^ n2732;
  assign n3245 = n2711 & n2763;
  assign n2759 = n2758 ^ n2757;
  assign n2747 = n2740 & n2746;
  assign n2748 = ~n2732 & n2747;
  assign n2760 = n2759 ^ n2748;
  assign n2764 = n2763 ^ n2760;
  assign n3244 = n2722 & n2764;
  assign n3246 = n3245 ^ n3244;
  assign n2766 = n2756 ^ n2746;
  assign n2767 = n2757 ^ n2732;
  assign n2768 = n2766 & n2767;
  assign n2769 = n2768 ^ n2746;
  assign n3218 = n2715 & n2769;
  assign n2773 = n2766 ^ n2757;
  assign n2771 = ~n2746 & n2756;
  assign n2772 = n2732 & n2771;
  assign n2774 = n2773 ^ n2772;
  assign n3217 = n2750 & n2774;
  assign n3219 = n3218 ^ n3217;
  assign n3424 = n3246 ^ n3219;
  assign n2780 = n2774 ^ n2769;
  assign n3220 = n2704 & n2780;
  assign n2781 = n2710 & n2780;
  assign n2770 = n2769 ^ n2763;
  assign n2778 = n2716 & n2770;
  assign n2775 = n2774 ^ n2760;
  assign n2776 = n2775 ^ n2770;
  assign n2777 = n2701 & n2776;
  assign n2779 = n2778 ^ n2777;
  assign n2782 = n2781 ^ n2779;
  assign n3423 = n3220 ^ n2782;
  assign n3425 = n3424 ^ n3423;
  assign n3432 = n3431 ^ n3425;
  assign n3439 = n3438 ^ n3432;
  assign n3408 = n3070 & n3136;
  assign n3285 = n3093 & n3136;
  assign n3194 = n3089 & n3191;
  assign n3286 = n3285 ^ n3194;
  assign n3409 = n3408 ^ n3286;
  assign n3406 = n3155 ^ n3146;
  assign n3352 = n3087 & n3139;
  assign n3196 = n3072 & n3142;
  assign n3153 = n3092 & n3150;
  assign n3197 = n3196 ^ n3153;
  assign n3353 = n3352 ^ n3197;
  assign n3407 = n3406 ^ n3353;
  assign n3410 = n3409 ^ n3407;
  assign n3383 = n2989 & n3052;
  assign n3185 = n2988 & n3052;
  assign n3186 = n3185 ^ n3184;
  assign n3384 = n3383 ^ n3186;
  assign n3381 = n3059 ^ n3055;
  assign n3278 = n3001 & n3044;
  assign n3279 = n3278 ^ n3211;
  assign n3382 = n3381 ^ n3279;
  assign n3385 = n3384 ^ n3382;
  assign n3411 = n3410 ^ n3385;
  assign n3309 = n2931 & n2942;
  assign n2947 = n2887 & n2946;
  assign n3310 = n3309 ^ n2947;
  assign n3311 = n3310 ^ n3269;
  assign n2967 = n2915 & n2958;
  assign n2966 = n2899 & n2957;
  assign n2968 = n2967 ^ n2966;
  assign n3403 = n3311 ^ n2968;
  assign n2969 = n2933 & n2942;
  assign n3402 = n2969 ^ n2961;
  assign n3404 = n3403 ^ n3402;
  assign n3165 = n3062 ^ n3056;
  assign n3160 = n3023 & n3038;
  assign n3161 = n3160 ^ n3040;
  assign n3163 = n3162 ^ n3161;
  assign n3164 = n3163 ^ n3061;
  assign n3166 = n3165 ^ n3164;
  assign n3405 = n3404 ^ n3166;
  assign n3412 = n3411 ^ n3405;
  assign n2788 = n2751 & n2760;
  assign n3393 = n2788 ^ n2779;
  assign n3295 = n2749 & n2760;
  assign n2765 = n2705 & n2764;
  assign n3296 = n3295 ^ n2765;
  assign n3297 = n3296 ^ n3244;
  assign n2785 = n2734 & n2776;
  assign n2784 = n2727 & n2770;
  assign n2786 = n2785 ^ n2784;
  assign n3392 = n3297 ^ n2786;
  assign n3394 = n3393 ^ n3392;
  assign n3401 = n3400 ^ n3394;
  assign n3413 = n3412 ^ n3401;
  assign n3149 = n3121 & n3129;
  assign n3152 = n3151 ^ n3149;
  assign n3154 = n3153 ^ n3152;
  assign n3387 = n3205 ^ n3154;
  assign n3388 = n3387 ^ n3193;
  assign n3314 = n3163 ^ n3064;
  assign n3315 = n3314 ^ n3057;
  assign n3389 = n3388 ^ n3315;
  assign n3378 = n2888 & n2953;
  assign n3175 = n2896 & n2953;
  assign n3176 = n3175 ^ n3174;
  assign n3379 = n3378 ^ n3176;
  assign n3376 = n2966 ^ n2960;
  assign n3271 = n2909 & n2956;
  assign n3272 = n3271 ^ n3270;
  assign n3377 = n3376 ^ n3272;
  assign n3380 = n3379 ^ n3377;
  assign n3386 = n3385 ^ n3380;
  assign n3390 = n3389 ^ n3386;
  assign n3364 = n2724 & n2775;
  assign n3221 = n2723 & n2775;
  assign n3222 = n3221 ^ n3220;
  assign n3365 = n3364 ^ n3222;
  assign n3362 = n2784 ^ n2778;
  assign n3247 = n2718 & n2769;
  assign n3248 = n3247 ^ n3246;
  assign n3363 = n3362 ^ n3248;
  assign n3366 = n3365 ^ n3363;
  assign n3375 = n3374 ^ n3366;
  assign n3391 = n3390 ^ n3375;
  assign n3414 = n3413 ^ n3391;
  assign n3440 = n3439 ^ n3414;
  assign n3323 = n3210 ^ n3181;
  assign n3324 = n3323 ^ n3161;
  assign n3322 = n3064 ^ n3056;
  assign n3325 = n3324 ^ n3322;
  assign n3326 = n3325 ^ n3066;
  assign n3199 = n3083 & n3139;
  assign n3318 = n3199 ^ n3196;
  assign n3319 = n3318 ^ n3152;
  assign n3317 = n3205 ^ n3147;
  assign n3320 = n3319 ^ n3317;
  assign n3321 = n3320 ^ n3207;
  assign n3327 = n3326 ^ n3321;
  assign n2970 = n2906 & n2952;
  assign n2971 = n2970 ^ n2969;
  assign n3312 = n3311 ^ n2971;
  assign n3313 = n3312 ^ n2964;
  assign n3316 = n3315 ^ n3313;
  assign n3328 = n3327 ^ n3316;
  assign n2787 = n2714 & n2774;
  assign n2789 = n2788 ^ n2787;
  assign n3298 = n3297 ^ n2789;
  assign n3299 = n3298 ^ n2782;
  assign n3308 = n3307 ^ n3299;
  assign n3329 = n3328 ^ n3308;
  assign n3289 = n3204 ^ n3147;
  assign n3287 = n3286 ^ n3156;
  assign n3198 = n3077 & n3135;
  assign n3200 = n3199 ^ n3198;
  assign n3288 = n3287 ^ n3200;
  assign n3290 = n3289 ^ n3288;
  assign n3187 = n3186 ^ n3060;
  assign n3188 = n3187 ^ n3183;
  assign n3180 = n3063 ^ n3056;
  assign n3189 = n3188 ^ n3180;
  assign n3291 = n3290 ^ n3189;
  assign n3280 = n3000 & n3034;
  assign n3281 = n3280 ^ n3064;
  assign n3282 = n3281 ^ n3279;
  assign n3277 = n3187 ^ n3057;
  assign n3283 = n3282 ^ n3277;
  assign n3273 = n2908 & n2945;
  assign n3274 = n3273 ^ n2971;
  assign n3275 = n3274 ^ n3272;
  assign n3177 = n3176 ^ n2967;
  assign n3267 = n3177 ^ n2964;
  assign n3276 = n3275 ^ n3267;
  assign n3284 = n3283 ^ n3276;
  assign n3292 = n3291 ^ n3284;
  assign n3249 = n2717 & n2763;
  assign n3250 = n3249 ^ n2789;
  assign n3251 = n3250 ^ n3248;
  assign n3223 = n3222 ^ n2785;
  assign n3243 = n3223 ^ n2782;
  assign n3252 = n3251 ^ n3243;
  assign n3266 = n3265 ^ n3252;
  assign n3293 = n3292 ^ n3266;
  assign n3454 = n3329 ^ n3293;
  assign n3421 = n3391 ^ n3293;
  assign n3158 = n3157 ^ n3154;
  assign n3148 = n3147 ^ n3130;
  assign n3159 = n3158 ^ n3148;
  assign n3167 = n3166 ^ n3159;
  assign n2972 = n2971 ^ n2968;
  assign n2965 = n2964 ^ n2947;
  assign n2973 = n2972 ^ n2965;
  assign n3067 = n3066 ^ n2973;
  assign n3168 = n3167 ^ n3067;
  assign n2790 = n2789 ^ n2786;
  assign n2783 = n2782 ^ n2765;
  assign n2791 = n2790 ^ n2783;
  assign n2880 = n2879 ^ n2791;
  assign n3169 = n3168 ^ n2880;
  assign n3330 = n3329 ^ n3169;
  assign n3459 = n3421 ^ n3330;
  assign n3460 = n3454 & n3459;
  assign n3417 = n3413 ^ n3293;
  assign n3357 = n3283 ^ n3066;
  assign n3350 = n3085 & n3142;
  assign n3351 = n3350 ^ n3205;
  assign n3354 = n3353 ^ n3351;
  assign n3349 = n3287 ^ n3193;
  assign n3355 = n3354 ^ n3349;
  assign n3356 = n3355 ^ n3207;
  assign n3358 = n3357 ^ n3356;
  assign n3338 = n3245 ^ n3218;
  assign n3339 = n3338 ^ n3296;
  assign n3337 = n2789 ^ n2779;
  assign n3340 = n3339 ^ n3337;
  assign n3348 = n3347 ^ n3340;
  assign n3359 = n3358 ^ n3348;
  assign n3332 = n3268 ^ n3171;
  assign n3333 = n3332 ^ n3310;
  assign n3331 = n2971 ^ n2961;
  assign n3334 = n3333 ^ n3331;
  assign n3335 = n3334 ^ n3325;
  assign n3225 = n2787 ^ n2779;
  assign n3224 = n3223 ^ n3219;
  assign n3226 = n3225 ^ n3224;
  assign n3240 = n3239 ^ n3226;
  assign n3214 = n3213 ^ n3066;
  assign n3201 = n3200 ^ n3197;
  assign n3195 = n3194 ^ n3193;
  assign n3202 = n3201 ^ n3195;
  assign n3208 = n3207 ^ n3202;
  assign n3215 = n3214 ^ n3208;
  assign n3178 = n3177 ^ n3173;
  assign n3170 = n2970 ^ n2961;
  assign n3179 = n3178 ^ n3170;
  assign n3190 = n3189 ^ n3179;
  assign n3216 = n3215 ^ n3190;
  assign n3241 = n3240 ^ n3216;
  assign n3336 = n3335 ^ n3241;
  assign n3360 = n3359 ^ n3336;
  assign n3418 = n3417 ^ n3360;
  assign n3419 = n3330 & n3418;
  assign n3461 = n3460 ^ n3419;
  assign n3361 = n3360 ^ n3330;
  assign n3458 = n3417 ^ n3361;
  assign n3462 = n3461 ^ n3458;
  assign n3242 = n3241 ^ n3169;
  assign n3455 = n3454 ^ n3242;
  assign n3456 = n3361 & n3455;
  assign n3450 = n3439 ^ n3361;
  assign n3451 = n3440 ^ n3241;
  assign n3294 = n3293 ^ n3169;
  assign n3452 = n3451 ^ n3294;
  assign n3453 = ~n3450 & ~n3452;
  assign n3457 = n3456 ^ n3453;
  assign n3463 = n3462 ^ n3457;
  assign n3474 = ~n3241 & ~n3440;
  assign n3422 = n3421 ^ n3360;
  assign n3445 = n3242 & n3422;
  assign n3475 = n3474 ^ n3445;
  assign n3472 = n3422 ^ n3242;
  assign n3473 = n3472 ^ n3461;
  assign n3476 = n3475 ^ n3473;
  assign n3477 = n3463 & n3476;
  assign n3415 = n3414 ^ n3361;
  assign n3466 = n3415 ^ n3294;
  assign n3442 = n3440 ^ n3329;
  assign n3464 = ~n3439 & ~n3442;
  assign n3465 = n3464 ^ n3456;
  assign n3467 = n3466 ^ n3465;
  assign n3416 = n3294 & n3415;
  assign n3420 = n3419 ^ n3416;
  assign n3468 = n3467 ^ n3420;
  assign n3471 = n3468 ^ n3463;
  assign n3478 = n3477 ^ n3471;
  assign n3443 = n3442 ^ n3330;
  assign n3441 = n3440 ^ n3422;
  assign n3448 = n3443 ^ n3441;
  assign n3444 = ~n3441 & ~n3443;
  assign n3446 = n3445 ^ n3444;
  assign n3447 = n3446 ^ n3420;
  assign n3449 = n3448 ^ n3447;
  assign n3469 = n3463 & ~n3468;
  assign n3470 = n3449 & n3469;
  assign n3479 = n3478 ^ n3470;
  assign n3507 = ~n3440 & n3479;
  assign n3487 = n3476 ^ n3449;
  assign n3493 = n3477 ^ n3468;
  assign n3494 = n3487 & n3493;
  assign n3495 = n3494 ^ n3449;
  assign n3480 = n3477 ^ n3449;
  assign n3481 = n3471 & n3480;
  assign n3482 = n3481 ^ n3468;
  assign n3496 = n3495 ^ n3482;
  assign n3501 = n3330 & n3496;
  assign n3488 = n3487 ^ n3477;
  assign n3485 = n3468 & n3476;
  assign n3486 = ~n3449 & n3485;
  assign n3489 = n3488 ^ n3486;
  assign n3490 = n3489 ^ n3479;
  assign n3497 = n3496 ^ n3490;
  assign n3500 = n3454 & n3497;
  assign n3502 = n3501 ^ n3500;
  assign n3734 = n3507 ^ n3502;
  assign n3731 = ~n3441 & n3482;
  assign n3730 = ~n3451 & n3479;
  assign n3732 = n3731 ^ n3730;
  assign n3498 = n3459 & n3497;
  assign n3491 = n3415 & n3490;
  assign n3483 = n3482 ^ n3479;
  assign n3484 = n3242 & n3483;
  assign n3492 = n3491 ^ n3484;
  assign n3499 = n3498 ^ n3492;
  assign n3733 = n3732 ^ n3499;
  assign n3735 = n3734 ^ n3733;
  assign n1476 = x183 ^ x55;
  assign n1460 = x176 ^ x48;
  assign n1458 = x179 ^ x51;
  assign n1465 = n1460 ^ n1458;
  assign n1463 = x180 ^ x52;
  assign n1462 = x182 ^ x54;
  assign n1464 = n1463 ^ n1462;
  assign n1466 = n1465 ^ n1464;
  assign n1487 = n1476 ^ n1466;
  assign n1468 = x177 ^ x49;
  assign n1467 = x178 ^ x50;
  assign n1469 = n1468 ^ n1467;
  assign n1477 = n1476 ^ n1469;
  assign n1511 = ~n1462 & n1477;
  assign n1480 = n1462 ^ n1460;
  assign n1457 = x181 ^ x53;
  assign n1492 = n1467 ^ n1457;
  assign n1501 = n1492 ^ n1464;
  assign n1504 = n1480 & n1501;
  assign n1512 = n1511 ^ n1504;
  assign n1509 = n1501 ^ n1480;
  assign n1459 = n1458 ^ n1457;
  assign n1493 = n1492 ^ n1465;
  assign n1494 = n1459 & n1493;
  assign n1472 = n1468 ^ n1457;
  assign n1473 = n1472 ^ n1464;
  assign n1474 = n1465 & n1473;
  assign n1495 = n1494 ^ n1474;
  assign n1510 = n1509 ^ n1495;
  assign n1513 = n1512 ^ n1510;
  assign n1502 = n1501 ^ n1477;
  assign n1478 = n1477 ^ n1458;
  assign n1500 = n1478 ^ n1465;
  assign n1507 = n1502 ^ n1500;
  assign n1503 = n1500 & n1502;
  assign n1505 = n1504 ^ n1503;
  assign n1461 = n1460 ^ n1457;
  assign n1470 = n1469 ^ n1466;
  assign n1471 = n1461 & n1470;
  assign n1475 = n1474 ^ n1471;
  assign n1506 = n1505 ^ n1475;
  assign n1508 = n1507 ^ n1506;
  assign n1518 = n1513 ^ n1508;
  assign n1496 = n1472 ^ n1466;
  assign n1497 = n1496 ^ n1495;
  assign n1488 = n1477 ^ n1462;
  assign n1489 = n1488 ^ n1461;
  assign n1490 = n1487 & n1489;
  assign n1481 = n1480 ^ n1459;
  assign n1482 = n1466 & n1481;
  assign n1491 = n1490 ^ n1482;
  assign n1498 = n1497 ^ n1491;
  assign n1514 = n1498 & n1513;
  assign n1525 = n1518 ^ n1514;
  assign n1484 = n1470 ^ n1461;
  assign n1479 = n1476 & n1478;
  assign n1483 = n1482 ^ n1479;
  assign n1485 = n1484 ^ n1483;
  assign n1486 = n1485 ^ n1475;
  assign n1523 = n1486 & n1513;
  assign n1524 = ~n1508 & n1523;
  assign n1526 = n1525 ^ n1524;
  assign n1581 = n1487 & n1526;
  assign n1519 = n1514 ^ n1486;
  assign n1520 = n1518 & n1519;
  assign n1521 = n1520 ^ n1508;
  assign n1553 = n1526 ^ n1521;
  assign n1558 = n1481 & n1553;
  assign n1582 = n1581 ^ n1558;
  assign n1554 = n1466 & n1553;
  assign n1631 = n1582 ^ n1554;
  assign n1499 = n1498 ^ n1486;
  assign n1515 = n1514 ^ n1508;
  assign n1516 = n1499 & n1515;
  assign n1517 = n1516 ^ n1486;
  assign n1522 = n1521 ^ n1517;
  assign n1560 = n1473 & n1522;
  assign n1529 = n1514 ^ n1499;
  assign n1527 = ~n1486 & n1498;
  assign n1528 = n1508 & n1527;
  assign n1530 = n1529 ^ n1528;
  assign n1531 = n1530 ^ n1526;
  assign n1532 = n1531 ^ n1522;
  assign n1542 = n1493 & n1532;
  assign n1561 = n1560 ^ n1542;
  assign n1675 = n1631 ^ n1561;
  assign n1562 = n1489 & n1526;
  assign n1534 = n1465 & n1522;
  assign n1533 = n1459 & n1532;
  assign n1535 = n1534 ^ n1533;
  assign n1674 = n1562 ^ n1535;
  assign n1676 = n1675 ^ n1674;
  assign n1536 = n1477 & n1530;
  assign n1563 = n1562 ^ n1536;
  assign n1564 = n1563 ^ n1561;
  assign n1539 = n1530 ^ n1517;
  assign n1549 = n1501 & n1539;
  assign n1550 = n1549 ^ n1535;
  assign n1559 = n1558 ^ n1550;
  assign n1565 = n1564 ^ n1559;
  assign n1677 = n1676 ^ n1565;
  assign n1373 = x143 ^ x15;
  assign n1363 = x138 ^ x10;
  assign n1362 = x137 ^ x9;
  assign n1364 = n1363 ^ n1362;
  assign n1374 = n1373 ^ n1364;
  assign n1352 = x142 ^ x14;
  assign n1385 = n1374 ^ n1352;
  assign n1355 = x141 ^ x13;
  assign n1353 = x136 ^ x8;
  assign n1356 = n1355 ^ n1353;
  assign n1386 = n1385 ^ n1356;
  assign n1408 = ~n1352 & n1374;
  assign n1354 = n1353 ^ n1352;
  assign n1371 = n1363 ^ n1355;
  assign n1357 = x140 ^ x12;
  assign n1358 = n1357 ^ n1352;
  assign n1372 = n1371 ^ n1358;
  assign n1379 = n1354 & n1372;
  assign n1409 = n1408 ^ n1379;
  assign n1406 = n1372 ^ n1354;
  assign n1359 = x139 ^ x11;
  assign n1388 = n1359 ^ n1355;
  assign n1360 = n1359 ^ n1353;
  assign n1393 = n1371 ^ n1360;
  assign n1394 = n1388 & n1393;
  assign n1367 = n1362 ^ n1355;
  assign n1368 = n1367 ^ n1358;
  assign n1369 = n1360 & n1368;
  assign n1395 = n1394 ^ n1369;
  assign n1407 = n1406 ^ n1395;
  assign n1410 = n1409 ^ n1407;
  assign n1376 = n1374 ^ n1359;
  assign n1377 = n1376 ^ n1360;
  assign n1375 = n1374 ^ n1372;
  assign n1382 = n1377 ^ n1375;
  assign n1378 = n1375 & n1377;
  assign n1380 = n1379 ^ n1378;
  assign n1361 = n1360 ^ n1358;
  assign n1365 = n1364 ^ n1361;
  assign n1366 = n1356 & n1365;
  assign n1370 = n1369 ^ n1366;
  assign n1381 = n1380 ^ n1370;
  assign n1383 = n1382 ^ n1381;
  assign n1422 = n1410 ^ n1383;
  assign n1392 = n1367 ^ n1361;
  assign n1396 = n1395 ^ n1392;
  assign n1389 = n1388 ^ n1354;
  assign n1390 = n1361 & n1389;
  assign n1384 = n1373 ^ n1361;
  assign n1387 = n1384 & n1386;
  assign n1391 = n1390 ^ n1387;
  assign n1397 = n1396 ^ n1391;
  assign n1411 = n1397 & n1410;
  assign n1423 = n1422 ^ n1411;
  assign n1400 = n1365 ^ n1356;
  assign n1398 = n1373 & n1376;
  assign n1399 = n1398 ^ n1390;
  assign n1401 = n1400 ^ n1399;
  assign n1402 = n1401 ^ n1370;
  assign n1420 = n1402 & n1410;
  assign n1421 = ~n1383 & n1420;
  assign n1424 = n1423 ^ n1421;
  assign n1447 = n1386 & n1424;
  assign n1426 = n1411 ^ n1402;
  assign n1427 = n1422 & n1426;
  assign n1428 = n1427 ^ n1383;
  assign n1405 = n1402 ^ n1397;
  assign n1414 = n1411 ^ n1383;
  assign n1415 = n1405 & n1414;
  assign n1416 = n1415 ^ n1402;
  assign n1429 = n1428 ^ n1416;
  assign n1432 = n1360 & n1429;
  assign n1412 = n1411 ^ n1405;
  assign n1403 = n1397 & ~n1402;
  assign n1404 = n1383 & n1403;
  assign n1413 = n1412 ^ n1404;
  assign n1425 = n1424 ^ n1413;
  assign n1430 = n1429 ^ n1425;
  assign n1431 = n1388 & n1430;
  assign n1433 = n1432 ^ n1431;
  assign n1671 = n1447 ^ n1433;
  assign n1619 = n1384 & n1424;
  assign n1439 = n1428 ^ n1424;
  assign n1445 = n1389 & n1439;
  assign n1620 = n1619 ^ n1445;
  assign n1440 = n1361 & n1439;
  assign n1669 = n1620 ^ n1440;
  assign n1451 = n1393 & n1430;
  assign n1450 = n1368 & n1429;
  assign n1452 = n1451 ^ n1450;
  assign n1670 = n1669 ^ n1452;
  assign n1672 = n1671 ^ n1670;
  assign n1268 = x229 ^ x101;
  assign n1262 = x225 ^ x97;
  assign n1285 = n1268 ^ n1262;
  assign n1266 = x228 ^ x100;
  assign n1265 = x230 ^ x102;
  assign n1267 = n1266 ^ n1265;
  assign n1286 = n1285 ^ n1267;
  assign n1274 = x224 ^ x96;
  assign n1272 = x227 ^ x99;
  assign n1275 = n1274 ^ n1272;
  assign n1282 = n1275 ^ n1267;
  assign n1261 = x226 ^ x98;
  assign n1263 = n1262 ^ n1261;
  assign n1283 = n1282 ^ n1263;
  assign n1281 = n1274 ^ n1268;
  assign n1308 = n1283 ^ n1281;
  assign n1260 = x231 ^ x103;
  assign n1264 = n1263 ^ n1260;
  assign n1273 = n1272 ^ n1264;
  assign n1306 = n1260 & n1273;
  assign n1292 = n1272 ^ n1268;
  assign n1278 = n1274 ^ n1265;
  assign n1293 = n1292 ^ n1278;
  assign n1294 = n1282 & n1293;
  assign n1307 = n1306 ^ n1294;
  assign n1309 = n1308 ^ n1307;
  assign n1287 = n1275 & n1286;
  assign n1284 = n1281 & n1283;
  assign n1288 = n1287 ^ n1284;
  assign n1310 = n1309 ^ n1288;
  assign n1303 = n1285 ^ n1282;
  assign n1269 = n1268 ^ n1261;
  assign n1300 = n1275 ^ n1269;
  assign n1301 = n1292 & n1300;
  assign n1302 = n1301 ^ n1287;
  assign n1304 = n1303 ^ n1302;
  assign n1295 = n1282 ^ n1260;
  assign n1296 = n1265 ^ n1264;
  assign n1297 = n1296 ^ n1281;
  assign n1298 = n1295 & n1297;
  assign n1299 = n1298 ^ n1294;
  assign n1305 = n1304 ^ n1299;
  assign n1319 = n1310 ^ n1305;
  assign n1315 = n1264 & ~n1265;
  assign n1270 = n1269 ^ n1267;
  assign n1279 = n1270 & n1278;
  assign n1316 = n1315 ^ n1279;
  assign n1313 = n1278 ^ n1270;
  assign n1314 = n1313 ^ n1302;
  assign n1317 = n1316 ^ n1314;
  assign n1318 = n1305 & n1317;
  assign n1276 = n1275 ^ n1273;
  assign n1271 = n1270 ^ n1264;
  assign n1290 = n1276 ^ n1271;
  assign n1277 = n1271 & n1276;
  assign n1280 = n1279 ^ n1277;
  assign n1289 = n1288 ^ n1280;
  assign n1291 = n1290 ^ n1289;
  assign n1332 = n1318 ^ n1291;
  assign n1333 = n1319 & n1332;
  assign n1334 = n1333 ^ n1310;
  assign n1325 = n1317 ^ n1291;
  assign n1329 = n1318 ^ n1310;
  assign n1330 = n1325 & n1329;
  assign n1331 = n1330 ^ n1291;
  assign n1335 = n1334 ^ n1331;
  assign n1665 = n1286 & n1335;
  assign n1326 = n1325 ^ n1318;
  assign n1323 = n1310 & n1317;
  assign n1324 = ~n1291 & n1323;
  assign n1327 = n1326 ^ n1324;
  assign n1320 = n1319 ^ n1318;
  assign n1311 = n1305 & ~n1310;
  assign n1312 = n1291 & n1311;
  assign n1321 = n1320 ^ n1312;
  assign n1328 = n1327 ^ n1321;
  assign n1336 = n1335 ^ n1328;
  assign n1345 = n1300 & n1336;
  assign n1666 = n1665 ^ n1345;
  assign n1597 = n1297 & n1327;
  assign n1322 = n1264 & n1321;
  assign n1598 = n1597 ^ n1322;
  assign n1667 = n1666 ^ n1598;
  assign n1342 = n1334 ^ n1321;
  assign n1614 = n1270 & n1342;
  assign n1338 = n1275 & n1335;
  assign n1337 = n1292 & n1336;
  assign n1339 = n1338 ^ n1337;
  assign n1615 = n1614 ^ n1339;
  assign n1602 = n1331 ^ n1327;
  assign n1603 = n1293 & n1602;
  assign n1664 = n1615 ^ n1603;
  assign n1668 = n1667 ^ n1664;
  assign n1673 = n1672 ^ n1668;
  assign n1678 = n1677 ^ n1673;
  assign n1057 = x221 ^ x93;
  assign n1052 = x217 ^ x89;
  assign n1077 = n1057 ^ n1052;
  assign n1060 = x222 ^ x94;
  assign n1059 = x220 ^ x92;
  assign n1061 = n1060 ^ n1059;
  assign n1078 = n1077 ^ n1061;
  assign n1066 = x216 ^ x88;
  assign n1064 = x219 ^ x91;
  assign n1067 = n1066 ^ n1064;
  assign n1074 = n1067 ^ n1061;
  assign n1053 = x218 ^ x90;
  assign n1054 = n1053 ^ n1052;
  assign n1075 = n1074 ^ n1054;
  assign n1073 = n1066 ^ n1057;
  assign n1100 = n1075 ^ n1073;
  assign n1055 = x223 ^ x95;
  assign n1056 = n1055 ^ n1054;
  assign n1065 = n1064 ^ n1056;
  assign n1098 = n1055 & n1065;
  assign n1084 = n1064 ^ n1057;
  assign n1070 = n1066 ^ n1060;
  assign n1085 = n1084 ^ n1070;
  assign n1086 = n1074 & n1085;
  assign n1099 = n1098 ^ n1086;
  assign n1101 = n1100 ^ n1099;
  assign n1079 = n1067 & n1078;
  assign n1076 = n1073 & n1075;
  assign n1080 = n1079 ^ n1076;
  assign n1102 = n1101 ^ n1080;
  assign n1095 = n1077 ^ n1074;
  assign n1058 = n1057 ^ n1053;
  assign n1092 = n1067 ^ n1058;
  assign n1093 = n1084 & n1092;
  assign n1094 = n1093 ^ n1079;
  assign n1096 = n1095 ^ n1094;
  assign n1087 = n1074 ^ n1055;
  assign n1088 = n1060 ^ n1056;
  assign n1089 = n1088 ^ n1073;
  assign n1090 = n1087 & n1089;
  assign n1091 = n1090 ^ n1086;
  assign n1097 = n1096 ^ n1091;
  assign n1111 = n1102 ^ n1097;
  assign n1107 = n1056 & ~n1060;
  assign n1062 = n1061 ^ n1058;
  assign n1071 = n1062 & n1070;
  assign n1108 = n1107 ^ n1071;
  assign n1105 = n1070 ^ n1062;
  assign n1106 = n1105 ^ n1094;
  assign n1109 = n1108 ^ n1106;
  assign n1110 = n1097 & n1109;
  assign n1068 = n1067 ^ n1065;
  assign n1063 = n1062 ^ n1056;
  assign n1082 = n1068 ^ n1063;
  assign n1069 = n1063 & n1068;
  assign n1072 = n1071 ^ n1069;
  assign n1081 = n1080 ^ n1072;
  assign n1083 = n1082 ^ n1081;
  assign n1126 = n1110 ^ n1083;
  assign n1127 = n1111 & n1126;
  assign n1128 = n1127 ^ n1102;
  assign n1117 = n1109 ^ n1083;
  assign n1123 = n1110 ^ n1102;
  assign n1124 = n1117 & n1123;
  assign n1125 = n1124 ^ n1083;
  assign n1129 = n1128 ^ n1125;
  assign n1650 = n1078 & n1129;
  assign n1118 = n1117 ^ n1110;
  assign n1115 = n1102 & n1109;
  assign n1116 = ~n1083 & n1115;
  assign n1119 = n1118 ^ n1116;
  assign n1112 = n1111 ^ n1110;
  assign n1103 = n1097 & ~n1102;
  assign n1104 = n1083 & n1103;
  assign n1113 = n1112 ^ n1104;
  assign n1122 = n1119 ^ n1113;
  assign n1130 = n1129 ^ n1122;
  assign n1237 = n1092 & n1130;
  assign n1651 = n1650 ^ n1237;
  assign n1120 = n1089 & n1119;
  assign n1114 = n1056 & n1113;
  assign n1121 = n1120 ^ n1114;
  assign n1652 = n1651 ^ n1121;
  assign n1234 = n1128 ^ n1113;
  assign n1628 = n1062 & n1234;
  assign n1132 = n1067 & n1129;
  assign n1131 = n1084 & n1130;
  assign n1133 = n1132 ^ n1131;
  assign n1629 = n1628 ^ n1133;
  assign n1139 = n1125 ^ n1119;
  assign n1140 = n1085 & n1139;
  assign n1649 = n1629 ^ n1140;
  assign n1653 = n1652 ^ n1649;
  assign n1663 = n1662 ^ n1653;
  assign n1679 = n1678 ^ n1663;
  assign n1632 = n1631 ^ n1563;
  assign n1633 = n1632 ^ n1550;
  assign n1625 = n1074 & n1139;
  assign n1138 = n1087 & n1119;
  assign n1141 = n1140 ^ n1138;
  assign n1626 = n1625 ^ n1141;
  assign n1627 = n1626 ^ n1121;
  assign n1630 = n1629 ^ n1627;
  assign n1634 = n1633 ^ n1630;
  assign n1552 = n1476 & n1521;
  assign n1545 = n1502 & n1517;
  assign n1580 = n1552 ^ n1545;
  assign n1583 = n1582 ^ n1580;
  assign n1579 = n1563 ^ n1535;
  assign n1584 = n1583 ^ n1579;
  assign n1624 = n1584 ^ n1565;
  assign n1635 = n1634 ^ n1624;
  assign n1441 = n1373 & n1428;
  assign n1437 = n1375 & n1416;
  assign n1618 = n1441 ^ n1437;
  assign n1621 = n1620 ^ n1618;
  assign n1448 = n1374 & n1413;
  assign n1449 = n1448 ^ n1447;
  assign n1617 = n1449 ^ n1433;
  assign n1622 = n1621 ^ n1617;
  assign n1453 = n1452 ^ n1449;
  assign n1417 = n1416 ^ n1413;
  assign n1419 = n1372 & n1417;
  assign n1434 = n1433 ^ n1419;
  assign n1446 = n1445 ^ n1434;
  assign n1454 = n1453 ^ n1446;
  assign n1623 = n1622 ^ n1454;
  assign n1636 = n1635 ^ n1623;
  assign n1611 = n1282 & n1602;
  assign n1604 = n1295 & n1327;
  assign n1605 = n1604 ^ n1603;
  assign n1612 = n1611 ^ n1605;
  assign n1613 = n1612 ^ n1598;
  assign n1616 = n1615 ^ n1613;
  assign n1637 = n1636 ^ n1616;
  assign n1648 = n1647 ^ n1637;
  assign n1680 = n1679 ^ n1648;
  assign n1555 = n1554 ^ n1552;
  assign n1544 = n1488 & n1530;
  assign n1546 = n1545 ^ n1544;
  assign n1556 = n1555 ^ n1546;
  assign n1540 = n1480 & n1539;
  assign n1551 = n1550 ^ n1540;
  assign n1557 = n1556 ^ n1551;
  assign n1566 = n1565 ^ n1557;
  assign n1538 = n1470 & n1531;
  assign n1541 = n1540 ^ n1538;
  assign n1543 = n1542 ^ n1541;
  assign n1547 = n1546 ^ n1543;
  assign n1537 = n1536 ^ n1535;
  assign n1548 = n1547 ^ n1537;
  assign n1567 = n1566 ^ n1548;
  assign n1442 = n1441 ^ n1440;
  assign n1436 = n1385 & n1413;
  assign n1438 = n1437 ^ n1436;
  assign n1443 = n1442 ^ n1438;
  assign n1418 = n1354 & n1417;
  assign n1435 = n1434 ^ n1418;
  assign n1444 = n1443 ^ n1435;
  assign n1455 = n1454 ^ n1444;
  assign n1348 = n1271 & n1334;
  assign n1347 = n1296 & n1321;
  assign n1349 = n1348 ^ n1347;
  assign n1343 = n1278 & n1342;
  assign n1341 = n1283 & n1328;
  assign n1344 = n1343 ^ n1341;
  assign n1346 = n1345 ^ n1344;
  assign n1350 = n1349 ^ n1346;
  assign n1340 = n1339 ^ n1322;
  assign n1351 = n1350 ^ n1340;
  assign n1456 = n1455 ^ n1351;
  assign n1568 = n1567 ^ n1456;
  assign n1242 = n1133 ^ n1114;
  assign n1239 = n1088 & n1113;
  assign n1136 = n1063 & n1128;
  assign n1240 = n1239 ^ n1136;
  assign n1235 = n1070 & n1234;
  assign n1233 = n1075 & n1122;
  assign n1236 = n1235 ^ n1233;
  assign n1238 = n1237 ^ n1236;
  assign n1241 = n1240 ^ n1238;
  assign n1243 = n1242 ^ n1241;
  assign n1259 = n1258 ^ n1243;
  assign n1569 = n1568 ^ n1259;
  assign n1600 = n1260 & n1331;
  assign n1686 = n1611 ^ n1600;
  assign n1759 = n1686 ^ n1349;
  assign n1758 = n1615 ^ n1343;
  assign n1760 = n1759 ^ n1758;
  assign n1761 = n1760 ^ n1454;
  assign n1762 = n1761 ^ n1566;
  assign n1135 = n1055 & n1125;
  assign n1694 = n1625 ^ n1135;
  assign n1748 = n1694 ^ n1240;
  assign n1747 = n1629 ^ n1235;
  assign n1749 = n1748 ^ n1747;
  assign n1757 = n1756 ^ n1749;
  assign n1763 = n1762 ^ n1757;
  assign n1732 = n1133 ^ n1120;
  assign n1731 = n1651 ^ n1626;
  assign n1733 = n1732 ^ n1731;
  assign n1734 = n1733 ^ n1676;
  assign n1727 = n1356 & n1425;
  assign n1586 = n1365 & n1425;
  assign n1587 = n1586 ^ n1418;
  assign n1728 = n1727 ^ n1587;
  assign n1725 = n1450 ^ n1432;
  assign n1592 = n1377 & n1416;
  assign n1593 = n1592 ^ n1442;
  assign n1726 = n1725 ^ n1593;
  assign n1729 = n1728 ^ n1726;
  assign n1703 = n1461 & n1531;
  assign n1704 = n1703 ^ n1541;
  assign n1701 = n1560 ^ n1534;
  assign n1574 = n1500 & n1517;
  assign n1575 = n1574 ^ n1555;
  assign n1702 = n1701 ^ n1575;
  assign n1705 = n1704 ^ n1702;
  assign n1730 = n1729 ^ n1705;
  assign n1735 = n1734 ^ n1730;
  assign n1723 = n1597 ^ n1339;
  assign n1722 = n1666 ^ n1612;
  assign n1724 = n1723 ^ n1722;
  assign n1736 = n1735 ^ n1724;
  assign n1744 = n1743 ^ n1736;
  assign n1698 = n1073 & n1122;
  assign n1699 = n1698 ^ n1236;
  assign n1696 = n1650 ^ n1132;
  assign n1693 = n1068 & n1128;
  assign n1695 = n1694 ^ n1693;
  assign n1697 = n1696 ^ n1695;
  assign n1700 = n1699 ^ n1697;
  assign n1706 = n1705 ^ n1700;
  assign n1690 = n1281 & n1328;
  assign n1691 = n1690 ^ n1344;
  assign n1688 = n1665 ^ n1338;
  assign n1685 = n1276 & n1334;
  assign n1687 = n1686 ^ n1685;
  assign n1689 = n1688 ^ n1687;
  assign n1692 = n1691 ^ n1689;
  assign n1707 = n1706 ^ n1692;
  assign n1682 = n1669 ^ n1449;
  assign n1683 = n1682 ^ n1434;
  assign n1684 = n1683 ^ n1633;
  assign n1708 = n1707 ^ n1684;
  assign n1721 = n1720 ^ n1708;
  assign n1745 = n1744 ^ n1721;
  assign n1764 = n1763 ^ n1745;
  assign n1823 = ~n1569 & n1764;
  assign n1778 = n1448 ^ n1433;
  assign n1588 = n1587 ^ n1451;
  assign n1777 = n1588 ^ n1438;
  assign n1779 = n1778 ^ n1777;
  assign n1780 = n1779 ^ n1548;
  assign n1773 = n1065 & n1125;
  assign n1774 = n1773 ^ n1121;
  assign n1775 = n1774 ^ n1695;
  assign n1772 = n1629 ^ n1238;
  assign n1776 = n1775 ^ n1772;
  assign n1781 = n1780 ^ n1776;
  assign n1572 = n1478 & n1521;
  assign n1573 = n1572 ^ n1563;
  assign n1576 = n1575 ^ n1573;
  assign n1571 = n1550 ^ n1543;
  assign n1577 = n1576 ^ n1571;
  assign n1782 = n1781 ^ n1577;
  assign n1768 = n1273 & n1331;
  assign n1769 = n1768 ^ n1598;
  assign n1770 = n1769 ^ n1687;
  assign n1767 = n1615 ^ n1346;
  assign n1771 = n1770 ^ n1767;
  assign n1783 = n1782 ^ n1771;
  assign n1793 = n1792 ^ n1783;
  assign n1794 = n1793 ^ n1721;
  assign n1601 = n1600 ^ n1348;
  assign n1606 = n1605 ^ n1601;
  assign n1599 = n1598 ^ n1339;
  assign n1607 = n1606 ^ n1599;
  assign n1590 = n1376 & n1428;
  assign n1591 = n1590 ^ n1449;
  assign n1594 = n1593 ^ n1591;
  assign n1589 = n1588 ^ n1434;
  assign n1595 = n1594 ^ n1589;
  assign n1596 = n1595 ^ n1454;
  assign n1608 = n1607 ^ n1596;
  assign n1578 = n1577 ^ n1565;
  assign n1585 = n1584 ^ n1578;
  assign n1609 = n1608 ^ n1585;
  assign n1137 = n1136 ^ n1135;
  assign n1142 = n1141 ^ n1137;
  assign n1134 = n1133 ^ n1121;
  assign n1143 = n1142 ^ n1134;
  assign n1232 = n1231 ^ n1143;
  assign n1570 = n1569 ^ n1232;
  assign n1610 = n1609 ^ n1570;
  assign n1795 = n1794 ^ n1610;
  assign n1798 = n1679 ^ n1569;
  assign n1799 = n1795 & n1798;
  assign n1824 = n1823 ^ n1799;
  assign n1810 = n1793 ^ n1648;
  assign n1819 = n1794 ^ n1680;
  assign n1820 = n1810 & n1819;
  assign n1803 = n1793 ^ n1744;
  assign n1804 = n1803 ^ n1610;
  assign n1805 = n1680 & n1804;
  assign n1821 = n1820 ^ n1805;
  assign n1818 = n1798 ^ n1795;
  assign n1822 = n1821 ^ n1818;
  assign n1825 = n1824 ^ n1822;
  assign n1796 = n1795 ^ n1764;
  assign n1765 = n1764 ^ n1648;
  assign n1766 = n1765 ^ n1680;
  assign n1808 = n1796 ^ n1766;
  assign n1681 = n1680 ^ n1610;
  assign n1746 = n1745 ^ n1681;
  assign n1801 = n1793 ^ n1679;
  assign n1802 = n1746 & n1801;
  assign n1806 = n1805 ^ n1802;
  assign n1797 = n1766 & n1796;
  assign n1800 = n1799 ^ n1797;
  assign n1807 = n1806 ^ n1800;
  assign n1809 = n1808 ^ n1807;
  assign n1828 = n1825 ^ n1809;
  assign n1831 = n1764 ^ n1569;
  assign n1832 = n1831 ^ n1801;
  assign n1833 = n1763 ^ n1681;
  assign n1834 = n1832 & n1833;
  assign n1811 = n1810 ^ n1798;
  assign n1812 = n1681 & n1811;
  assign n1835 = n1834 ^ n1812;
  assign n1829 = n1803 ^ n1681;
  assign n1830 = n1829 ^ n1821;
  assign n1836 = n1835 ^ n1830;
  assign n1837 = n1825 & n1836;
  assign n1815 = n1801 ^ n1746;
  assign n1813 = n1763 & n1765;
  assign n1814 = n1813 ^ n1812;
  assign n1816 = n1815 ^ n1814;
  assign n1817 = n1816 ^ n1806;
  assign n1853 = n1837 ^ n1817;
  assign n1854 = n1828 & n1853;
  assign n1855 = n1854 ^ n1809;
  assign n1842 = n1836 ^ n1817;
  assign n1847 = n1837 ^ n1809;
  assign n1848 = n1842 & n1847;
  assign n1849 = n1848 ^ n1817;
  assign n1856 = n1855 ^ n1849;
  assign n1866 = n1680 & n1856;
  assign n1843 = n1842 ^ n1837;
  assign n1840 = ~n1817 & n1836;
  assign n1841 = n1809 & n1840;
  assign n1844 = n1843 ^ n1841;
  assign n1838 = n1837 ^ n1828;
  assign n1826 = n1817 & n1825;
  assign n1827 = ~n1809 & n1826;
  assign n1839 = n1838 ^ n1827;
  assign n1845 = n1844 ^ n1839;
  assign n1857 = n1856 ^ n1845;
  assign n1865 = n1810 & n1857;
  assign n1867 = n1866 ^ n1865;
  assign n1864 = n1764 & n1844;
  assign n1868 = n1867 ^ n1864;
  assign n1861 = n1831 & n1844;
  assign n1860 = n1796 & n1849;
  assign n1862 = n1861 ^ n1860;
  assign n1858 = n1819 & n1857;
  assign n1850 = n1849 ^ n1844;
  assign n1851 = n1798 & n1850;
  assign n1846 = n1746 & n1845;
  assign n1852 = n1851 ^ n1846;
  assign n1859 = n1858 ^ n1852;
  assign n1863 = n1862 ^ n1859;
  assign n1869 = n1868 ^ n1863;
  assign n7607 = n3735 ^ n1869;
  assign n3763 = n1765 & n1855;
  assign n3722 = n1832 & n1839;
  assign n3723 = n3722 ^ n1864;
  assign n3764 = n3763 ^ n3723;
  assign n3667 = n1855 ^ n1839;
  assign n3668 = n1681 & n3667;
  assign n3666 = n1763 & n1855;
  assign n3669 = n3668 ^ n3666;
  assign n3665 = n1766 & n1849;
  assign n3670 = n3669 ^ n3665;
  assign n3765 = n3764 ^ n3670;
  assign n3718 = n1795 & n1850;
  assign n3719 = n3718 ^ n1867;
  assign n3762 = n3719 ^ n1859;
  assign n3766 = n3765 ^ n3762;
  assign n268 = x254 ^ x126;
  assign n267 = x252 ^ x124;
  assign n269 = n268 ^ n267;
  assign n265 = x251 ^ x123;
  assign n262 = x248 ^ x120;
  assign n266 = n265 ^ n262;
  assign n270 = n269 ^ n266;
  assign n259 = x250 ^ x122;
  assign n258 = x249 ^ x121;
  assign n260 = n259 ^ n258;
  assign n257 = x255 ^ x127;
  assign n261 = n260 ^ n257;
  assign n313 = n261 & ~n268;
  assign n263 = x253 ^ x125;
  assign n277 = n263 ^ n259;
  assign n278 = n277 ^ n269;
  assign n283 = n268 ^ n262;
  assign n284 = n278 & n283;
  assign n314 = n313 ^ n284;
  assign n311 = n283 ^ n278;
  assign n293 = n265 ^ n263;
  assign n298 = n277 ^ n266;
  assign n299 = n293 & n298;
  assign n273 = n263 ^ n258;
  assign n274 = n273 ^ n269;
  assign n275 = n266 & n274;
  assign n300 = n299 ^ n275;
  assign n312 = n311 ^ n300;
  assign n315 = n314 ^ n312;
  assign n280 = n265 ^ n261;
  assign n281 = n280 ^ n266;
  assign n279 = n278 ^ n261;
  assign n287 = n281 ^ n279;
  assign n282 = n279 & n281;
  assign n285 = n284 ^ n282;
  assign n264 = n263 ^ n262;
  assign n271 = n270 ^ n260;
  assign n272 = n264 & n271;
  assign n276 = n275 ^ n272;
  assign n286 = n285 ^ n276;
  assign n288 = n287 ^ n286;
  assign n322 = n315 ^ n288;
  assign n297 = n273 ^ n270;
  assign n301 = n300 ^ n297;
  assign n294 = n293 ^ n283;
  assign n295 = n270 & n294;
  assign n289 = n270 ^ n257;
  assign n290 = n268 ^ n261;
  assign n291 = n290 ^ n264;
  assign n292 = n289 & n291;
  assign n296 = n295 ^ n292;
  assign n302 = n301 ^ n296;
  assign n316 = n302 & n315;
  assign n305 = n271 ^ n264;
  assign n303 = n257 & n280;
  assign n304 = n303 ^ n295;
  assign n306 = n305 ^ n304;
  assign n307 = n306 ^ n276;
  assign n327 = n316 ^ n307;
  assign n328 = n322 & n327;
  assign n329 = n328 ^ n288;
  assign n323 = n322 ^ n316;
  assign n320 = n307 & n315;
  assign n321 = ~n288 & n320;
  assign n324 = n323 ^ n321;
  assign n343 = n329 ^ n324;
  assign n552 = n270 & n343;
  assign n345 = n289 & n324;
  assign n344 = n294 & n343;
  assign n346 = n345 ^ n344;
  assign n817 = n552 ^ n346;
  assign n325 = n291 & n324;
  assign n310 = n307 ^ n302;
  assign n317 = n316 ^ n310;
  assign n308 = n302 & ~n307;
  assign n309 = n288 & n308;
  assign n318 = n317 ^ n309;
  assign n319 = n261 & n318;
  assign n326 = n325 ^ n319;
  assign n864 = n817 ^ n326;
  assign n330 = n316 ^ n288;
  assign n331 = n310 & n330;
  assign n332 = n331 ^ n307;
  assign n539 = n332 ^ n318;
  assign n540 = n278 & n539;
  assign n333 = n332 ^ n329;
  assign n337 = n266 & n333;
  assign n334 = n324 ^ n318;
  assign n335 = n334 ^ n333;
  assign n336 = n293 & n335;
  assign n338 = n337 ^ n336;
  assign n541 = n540 ^ n338;
  assign n865 = n864 ^ n541;
  assign n871 = n870 ^ n865;
  assign n572 = x168 ^ x40;
  assign n570 = x171 ^ x43;
  assign n573 = n572 ^ n570;
  assign n566 = x172 ^ x44;
  assign n565 = x174 ^ x46;
  assign n567 = n566 ^ n565;
  assign n580 = n573 ^ n567;
  assign n560 = x169 ^ x41;
  assign n559 = x170 ^ x42;
  assign n561 = n560 ^ n559;
  assign n558 = x175 ^ x47;
  assign n562 = n561 ^ n558;
  assign n614 = n562 & ~n565;
  assign n563 = x173 ^ x45;
  assign n564 = n563 ^ n559;
  assign n568 = n567 ^ n564;
  assign n576 = n572 ^ n565;
  assign n577 = n568 & n576;
  assign n615 = n614 ^ n577;
  assign n612 = n576 ^ n568;
  assign n590 = n570 ^ n563;
  assign n599 = n573 ^ n564;
  assign n600 = n590 & n599;
  assign n583 = n563 ^ n560;
  assign n584 = n583 ^ n567;
  assign n585 = n573 & n584;
  assign n601 = n600 ^ n585;
  assign n613 = n612 ^ n601;
  assign n616 = n615 ^ n613;
  assign n571 = n570 ^ n562;
  assign n574 = n573 ^ n571;
  assign n569 = n568 ^ n562;
  assign n588 = n574 ^ n569;
  assign n579 = n572 ^ n563;
  assign n581 = n580 ^ n561;
  assign n582 = n579 & n581;
  assign n586 = n585 ^ n582;
  assign n575 = n569 & n574;
  assign n578 = n577 ^ n575;
  assign n587 = n586 ^ n578;
  assign n589 = n588 ^ n587;
  assign n623 = n616 ^ n589;
  assign n598 = n583 ^ n580;
  assign n602 = n601 ^ n598;
  assign n593 = n580 ^ n558;
  assign n594 = n565 ^ n562;
  assign n595 = n594 ^ n579;
  assign n596 = n593 & n595;
  assign n591 = n590 ^ n576;
  assign n592 = n580 & n591;
  assign n597 = n596 ^ n592;
  assign n603 = n602 ^ n597;
  assign n617 = n603 & n616;
  assign n606 = n581 ^ n579;
  assign n604 = n558 & n571;
  assign n605 = n604 ^ n592;
  assign n607 = n606 ^ n605;
  assign n608 = n607 ^ n586;
  assign n630 = n617 ^ n608;
  assign n631 = n623 & n630;
  assign n632 = n631 ^ n589;
  assign n624 = n623 ^ n617;
  assign n621 = n608 & n616;
  assign n622 = ~n589 & n621;
  assign n625 = n624 ^ n622;
  assign n790 = n632 ^ n625;
  assign n858 = n580 & n790;
  assign n792 = n593 & n625;
  assign n791 = n591 & n790;
  assign n793 = n792 ^ n791;
  assign n859 = n858 ^ n793;
  assign n785 = n595 & n625;
  assign n611 = n608 ^ n603;
  assign n618 = n617 ^ n611;
  assign n609 = n603 & ~n608;
  assign n610 = n589 & n609;
  assign n619 = n618 ^ n610;
  assign n620 = n562 & n619;
  assign n786 = n785 ^ n620;
  assign n860 = n859 ^ n786;
  assign n627 = n617 ^ n589;
  assign n628 = n611 & n627;
  assign n629 = n628 ^ n608;
  assign n639 = n629 ^ n619;
  assign n821 = n568 & n639;
  assign n633 = n632 ^ n629;
  assign n636 = n573 & n633;
  assign n626 = n625 ^ n619;
  assign n634 = n633 ^ n626;
  assign n635 = n590 & n634;
  assign n637 = n636 ^ n635;
  assign n822 = n821 ^ n637;
  assign n861 = n860 ^ n822;
  assign n664 = x131 ^ x3;
  assign n650 = x128 ^ x0;
  assign n666 = n664 ^ n650;
  assign n656 = x132 ^ x4;
  assign n651 = x134 ^ x6;
  assign n657 = n656 ^ n651;
  assign n672 = n666 ^ n657;
  assign n661 = x135 ^ x7;
  assign n659 = x129 ^ x1;
  assign n653 = x130 ^ x2;
  assign n660 = n659 ^ n653;
  assign n662 = n661 ^ n660;
  assign n705 = ~n651 & n662;
  assign n652 = n651 ^ n650;
  assign n654 = x133 ^ x5;
  assign n655 = n654 ^ n653;
  assign n658 = n657 ^ n655;
  assign n669 = n652 & n658;
  assign n706 = n705 ^ n669;
  assign n703 = n658 ^ n652;
  assign n682 = n664 ^ n654;
  assign n690 = n666 ^ n655;
  assign n691 = n682 & n690;
  assign n675 = n659 ^ n654;
  assign n676 = n675 ^ n657;
  assign n677 = n666 & n676;
  assign n692 = n691 ^ n677;
  assign n704 = n703 ^ n692;
  assign n707 = n706 ^ n704;
  assign n665 = n664 ^ n662;
  assign n667 = n666 ^ n665;
  assign n663 = n662 ^ n658;
  assign n680 = n667 ^ n663;
  assign n671 = n654 ^ n650;
  assign n673 = n672 ^ n660;
  assign n674 = n671 & n673;
  assign n678 = n677 ^ n674;
  assign n668 = n663 & n667;
  assign n670 = n669 ^ n668;
  assign n679 = n678 ^ n670;
  assign n681 = n680 ^ n679;
  assign n719 = n707 ^ n681;
  assign n693 = n675 ^ n672;
  assign n694 = n693 ^ n692;
  assign n685 = n672 ^ n661;
  assign n686 = n662 ^ n651;
  assign n687 = n686 ^ n671;
  assign n688 = n685 & n687;
  assign n683 = n682 ^ n652;
  assign n684 = n672 & n683;
  assign n689 = n688 ^ n684;
  assign n695 = n694 ^ n689;
  assign n708 = n695 & n707;
  assign n698 = n673 ^ n671;
  assign n696 = n661 & n665;
  assign n697 = n696 ^ n684;
  assign n699 = n698 ^ n697;
  assign n700 = n699 ^ n678;
  assign n725 = n708 ^ n700;
  assign n726 = n719 & n725;
  assign n727 = n726 ^ n681;
  assign n720 = n719 ^ n708;
  assign n717 = n700 & n707;
  assign n718 = ~n681 & n717;
  assign n721 = n720 ^ n718;
  assign n801 = n727 ^ n721;
  assign n854 = n672 & n801;
  assign n803 = n685 & n721;
  assign n802 = n683 & n801;
  assign n804 = n803 ^ n802;
  assign n855 = n854 ^ n804;
  assign n796 = n687 & n721;
  assign n709 = n700 ^ n695;
  assign n710 = n709 ^ n708;
  assign n701 = n695 & ~n700;
  assign n702 = n681 & n701;
  assign n711 = n710 ^ n702;
  assign n736 = n662 & n711;
  assign n797 = n796 ^ n736;
  assign n856 = n855 ^ n797;
  assign n712 = n708 ^ n681;
  assign n713 = n709 & n712;
  assign n714 = n713 ^ n700;
  assign n715 = n714 ^ n711;
  assign n828 = n658 & n715;
  assign n728 = n727 ^ n714;
  assign n738 = n666 & n728;
  assign n722 = n721 ^ n711;
  assign n729 = n728 ^ n722;
  assign n737 = n682 & n729;
  assign n739 = n738 ^ n737;
  assign n829 = n828 ^ n739;
  assign n857 = n856 ^ n829;
  assign n862 = n861 ^ n857;
  assign n544 = n274 & n333;
  assign n543 = n298 & n335;
  assign n545 = n544 ^ n543;
  assign n546 = n545 ^ n326;
  assign n542 = n541 ^ n344;
  assign n547 = n546 ^ n542;
  assign n341 = n257 & n329;
  assign n340 = n279 & n332;
  assign n342 = n341 ^ n340;
  assign n347 = n346 ^ n342;
  assign n339 = n338 ^ n326;
  assign n348 = n347 ^ n339;
  assign n852 = n547 ^ n348;
  assign n442 = x215 ^ x87;
  assign n449 = x208 ^ x80;
  assign n443 = x211 ^ x83;
  assign n450 = n449 ^ n443;
  assign n444 = x209 ^ x81;
  assign n435 = x210 ^ x82;
  assign n445 = n444 ^ n435;
  assign n446 = n445 ^ n442;
  assign n447 = n446 ^ n443;
  assign n487 = n450 ^ n447;
  assign n439 = x214 ^ x86;
  assign n438 = x212 ^ x84;
  assign n440 = n439 ^ n438;
  assign n436 = x213 ^ x85;
  assign n437 = n436 ^ n435;
  assign n441 = n440 ^ n437;
  assign n486 = n446 ^ n441;
  assign n491 = n487 ^ n486;
  assign n488 = n486 & n487;
  assign n453 = n449 ^ n439;
  assign n481 = n441 & n453;
  assign n489 = n488 ^ n481;
  assign n462 = n444 ^ n436;
  assign n463 = n462 ^ n440;
  assign n464 = n450 & n463;
  assign n451 = n450 ^ n440;
  assign n457 = n451 ^ n445;
  assign n458 = n449 ^ n436;
  assign n461 = n457 & n458;
  assign n465 = n464 ^ n461;
  assign n490 = n489 ^ n465;
  assign n492 = n491 ^ n490;
  assign n482 = ~n439 & n446;
  assign n483 = n482 ^ n481;
  assign n479 = n453 ^ n441;
  assign n452 = n443 ^ n436;
  assign n473 = n450 ^ n437;
  assign n474 = n452 & n473;
  assign n475 = n474 ^ n464;
  assign n480 = n479 ^ n475;
  assign n484 = n483 ^ n480;
  assign n502 = n492 ^ n484;
  assign n472 = n462 ^ n451;
  assign n476 = n475 ^ n472;
  assign n467 = n451 ^ n442;
  assign n468 = n446 ^ n439;
  assign n469 = n468 ^ n458;
  assign n470 = n467 & n469;
  assign n454 = n453 ^ n452;
  assign n455 = n451 & n454;
  assign n471 = n470 ^ n455;
  assign n477 = n476 ^ n471;
  assign n485 = n477 & n484;
  assign n459 = n458 ^ n457;
  assign n448 = n442 & n447;
  assign n456 = n455 ^ n448;
  assign n460 = n459 ^ n456;
  assign n466 = n465 ^ n460;
  assign n503 = n485 ^ n466;
  assign n504 = n502 & n503;
  assign n505 = n504 ^ n492;
  assign n522 = n442 & n505;
  assign n478 = n477 ^ n466;
  assign n493 = n492 ^ n485;
  assign n494 = n478 & n493;
  assign n495 = n494 ^ n466;
  assign n519 = n486 & n495;
  assign n848 = n522 ^ n519;
  assign n509 = n502 ^ n485;
  assign n507 = n466 & n484;
  assign n508 = ~n492 & n507;
  assign n510 = n509 ^ n508;
  assign n811 = n467 & n510;
  assign n523 = n510 ^ n505;
  assign n528 = n454 & n523;
  assign n812 = n811 ^ n528;
  assign n849 = n848 ^ n812;
  assign n534 = n469 & n510;
  assign n498 = n485 ^ n478;
  assign n496 = ~n466 & n477;
  assign n497 = n492 & n496;
  assign n499 = n498 ^ n497;
  assign n533 = n446 & n499;
  assign n535 = n534 ^ n533;
  assign n506 = n505 ^ n495;
  assign n514 = n450 & n506;
  assign n511 = n510 ^ n499;
  assign n512 = n511 ^ n506;
  assign n513 = n452 & n512;
  assign n515 = n514 ^ n513;
  assign n847 = n535 ^ n515;
  assign n850 = n849 ^ n847;
  assign n531 = n463 & n506;
  assign n530 = n473 & n512;
  assign n532 = n531 ^ n530;
  assign n536 = n535 ^ n532;
  assign n500 = n499 ^ n495;
  assign n501 = n441 & n500;
  assign n516 = n515 ^ n501;
  assign n529 = n528 ^ n516;
  assign n537 = n536 ^ n529;
  assign n851 = n850 ^ n537;
  assign n853 = n852 ^ n851;
  assign n863 = n862 ^ n853;
  assign n872 = n871 ^ n863;
  assign n845 = n844 ^ n547;
  assign n831 = n676 & n728;
  assign n730 = n690 & n729;
  assign n832 = n831 ^ n730;
  assign n833 = n832 ^ n797;
  assign n830 = n829 ^ n802;
  assign n834 = n833 ^ n830;
  assign n824 = n584 & n633;
  assign n643 = n599 & n634;
  assign n825 = n824 ^ n643;
  assign n826 = n825 ^ n786;
  assign n823 = n822 ^ n791;
  assign n827 = n826 ^ n823;
  assign n835 = n834 ^ n827;
  assign n818 = n817 ^ n545;
  assign n816 = n338 ^ n325;
  assign n819 = n818 ^ n816;
  assign n524 = n451 & n523;
  assign n813 = n812 ^ n524;
  assign n814 = n813 ^ n532;
  assign n810 = n534 ^ n515;
  assign n815 = n814 ^ n810;
  assign n820 = n819 ^ n815;
  assign n836 = n835 ^ n820;
  assign n846 = n845 ^ n836;
  assign n873 = n872 ^ n846;
  assign n799 = n661 & n727;
  assign n733 = n663 & n714;
  assign n800 = n799 ^ n733;
  assign n805 = n804 ^ n800;
  assign n798 = n797 ^ n739;
  assign n806 = n805 ^ n798;
  assign n788 = n558 & n632;
  assign n645 = n569 & n629;
  assign n789 = n788 ^ n645;
  assign n794 = n793 ^ n789;
  assign n787 = n786 ^ n637;
  assign n795 = n794 ^ n787;
  assign n807 = n806 ^ n795;
  assign n779 = n281 & n332;
  assign n553 = n552 ^ n341;
  assign n780 = n779 ^ n553;
  assign n777 = n280 & n329;
  assign n778 = n777 ^ n326;
  assign n781 = n780 ^ n778;
  assign n744 = n271 & n334;
  assign n548 = n283 & n539;
  assign n745 = n744 ^ n548;
  assign n746 = n745 ^ n543;
  assign n776 = n746 ^ n541;
  assign n782 = n781 ^ n776;
  assign n783 = n782 ^ n547;
  assign n771 = n487 & n495;
  assign n525 = n524 ^ n522;
  assign n772 = n771 ^ n525;
  assign n769 = n447 & n505;
  assign n770 = n769 ^ n535;
  assign n773 = n772 ^ n770;
  assign n765 = n457 & n511;
  assign n517 = n453 & n500;
  assign n766 = n765 ^ n517;
  assign n767 = n766 ^ n530;
  assign n768 = n767 ^ n516;
  assign n774 = n773 ^ n768;
  assign n775 = n774 ^ n537;
  assign n784 = n783 ^ n775;
  assign n808 = n807 ^ n784;
  assign n748 = n338 ^ n319;
  assign n550 = n290 & n318;
  assign n551 = n550 ^ n340;
  assign n747 = n746 ^ n551;
  assign n749 = n748 ^ n747;
  assign n762 = n761 ^ n749;
  assign n740 = n739 ^ n736;
  assign n732 = n686 & n711;
  assign n734 = n733 ^ n732;
  assign n723 = n673 & n722;
  assign n716 = n652 & n715;
  assign n724 = n723 ^ n716;
  assign n731 = n730 ^ n724;
  assign n735 = n734 ^ n731;
  assign n741 = n740 ^ n735;
  assign n646 = n594 & n619;
  assign n647 = n646 ^ n645;
  assign n641 = n581 & n626;
  assign n640 = n576 & n639;
  assign n642 = n641 ^ n640;
  assign n644 = n643 ^ n642;
  assign n648 = n647 ^ n644;
  assign n638 = n637 ^ n620;
  assign n649 = n648 ^ n638;
  assign n742 = n741 ^ n649;
  assign n554 = n553 ^ n551;
  assign n549 = n548 ^ n541;
  assign n555 = n554 ^ n549;
  assign n556 = n555 ^ n547;
  assign n520 = n468 & n499;
  assign n521 = n520 ^ n519;
  assign n526 = n525 ^ n521;
  assign n518 = n517 ^ n516;
  assign n527 = n526 ^ n518;
  assign n538 = n537 ^ n527;
  assign n557 = n556 ^ n538;
  assign n743 = n742 ^ n557;
  assign n763 = n762 ^ n743;
  assign n434 = n433 ^ n348;
  assign n764 = n763 ^ n434;
  assign n809 = n808 ^ n764;
  assign n874 = n873 ^ n809;
  assign n947 = n946 ^ n555;
  assign n878 = n854 ^ n799;
  assign n939 = n878 ^ n734;
  assign n938 = n829 ^ n716;
  assign n940 = n939 ^ n938;
  assign n886 = n858 ^ n788;
  assign n936 = n886 ^ n647;
  assign n935 = n822 ^ n640;
  assign n937 = n936 ^ n935;
  assign n941 = n940 ^ n937;
  assign n934 = n547 ^ n537;
  assign n942 = n941 ^ n934;
  assign n948 = n947 ^ n942;
  assign n927 = n855 ^ n832;
  assign n926 = n796 ^ n739;
  assign n928 = n927 ^ n926;
  assign n924 = n859 ^ n825;
  assign n923 = n785 ^ n637;
  assign n925 = n924 ^ n923;
  assign n929 = n928 ^ n925;
  assign n919 = n458 & n511;
  assign n920 = n919 ^ n766;
  assign n917 = n531 ^ n514;
  assign n918 = n917 ^ n772;
  assign n921 = n920 ^ n918;
  assign n898 = n264 & n334;
  assign n899 = n898 ^ n745;
  assign n896 = n544 ^ n337;
  assign n897 = n896 ^ n780;
  assign n900 = n899 ^ n897;
  assign n922 = n921 ^ n900;
  assign n930 = n929 ^ n922;
  assign n916 = n915 ^ n819;
  assign n931 = n930 ^ n916;
  assign n910 = n909 ^ n900;
  assign n891 = n579 & n626;
  assign n892 = n891 ^ n642;
  assign n889 = n824 ^ n636;
  assign n887 = n574 & n629;
  assign n888 = n887 ^ n886;
  assign n890 = n889 ^ n888;
  assign n893 = n892 ^ n890;
  assign n883 = n671 & n722;
  assign n884 = n883 ^ n724;
  assign n881 = n831 ^ n738;
  assign n879 = n667 & n714;
  assign n880 = n879 ^ n878;
  assign n882 = n881 ^ n880;
  assign n885 = n884 ^ n882;
  assign n894 = n893 ^ n885;
  assign n875 = n813 ^ n535;
  assign n876 = n875 ^ n516;
  assign n877 = n876 ^ n865;
  assign n895 = n894 ^ n877;
  assign n911 = n910 ^ n895;
  assign n932 = n931 ^ n911;
  assign n949 = n948 ^ n932;
  assign n1005 = ~n763 & n949;
  assign n974 = n973 ^ n782;
  assign n964 = n767 ^ n521;
  assign n963 = n533 ^ n515;
  assign n965 = n964 ^ n963;
  assign n966 = n965 ^ n749;
  assign n958 = n571 & n632;
  assign n959 = n958 ^ n786;
  assign n960 = n959 ^ n888;
  assign n957 = n822 ^ n644;
  assign n961 = n960 ^ n957;
  assign n953 = n665 & n727;
  assign n954 = n953 ^ n797;
  assign n955 = n954 ^ n880;
  assign n952 = n829 ^ n731;
  assign n956 = n955 ^ n952;
  assign n962 = n961 ^ n956;
  assign n967 = n966 ^ n962;
  assign n975 = n974 ^ n967;
  assign n976 = n975 ^ n911;
  assign n977 = n976 ^ n809;
  assign n980 = n846 ^ n763;
  assign n981 = n977 & n980;
  assign n1006 = n1005 ^ n981;
  assign n993 = n975 ^ n872;
  assign n1001 = n976 ^ n873;
  assign n1002 = n993 & n1001;
  assign n985 = n975 ^ n931;
  assign n986 = n985 ^ n809;
  assign n987 = n873 & n986;
  assign n1003 = n1002 ^ n987;
  assign n1000 = n980 ^ n977;
  assign n1004 = n1003 ^ n1000;
  assign n1007 = n1006 ^ n1004;
  assign n978 = n977 ^ n949;
  assign n950 = n949 ^ n872;
  assign n951 = n950 ^ n873;
  assign n990 = n978 ^ n951;
  assign n933 = n932 ^ n874;
  assign n983 = n975 ^ n846;
  assign n984 = n933 & n983;
  assign n988 = n987 ^ n984;
  assign n979 = n951 & n978;
  assign n982 = n981 ^ n979;
  assign n989 = n988 ^ n982;
  assign n991 = n990 ^ n989;
  assign n1010 = n1007 ^ n991;
  assign n1016 = n985 ^ n874;
  assign n1017 = n1016 ^ n1003;
  assign n1011 = n949 ^ n763;
  assign n1012 = n1011 ^ n983;
  assign n1013 = n948 ^ n874;
  assign n1014 = n1012 & n1013;
  assign n994 = n993 ^ n980;
  assign n995 = n874 & n994;
  assign n1015 = n1014 ^ n995;
  assign n1018 = n1017 ^ n1015;
  assign n1019 = n1007 & n1018;
  assign n997 = n983 ^ n933;
  assign n992 = n948 & n950;
  assign n996 = n995 ^ n992;
  assign n998 = n997 ^ n996;
  assign n999 = n998 ^ n988;
  assign n1035 = n1019 ^ n999;
  assign n1036 = n1010 & n1035;
  assign n1037 = n1036 ^ n991;
  assign n1020 = n1019 ^ n1010;
  assign n1008 = n999 & n1007;
  assign n1009 = ~n991 & n1008;
  assign n1021 = n1020 ^ n1009;
  assign n2692 = n1037 ^ n1021;
  assign n2693 = n874 & n2692;
  assign n2691 = n948 & n1037;
  assign n2694 = n2693 ^ n2691;
  assign n1024 = n1018 ^ n999;
  assign n1029 = n1019 ^ n991;
  assign n1030 = n1024 & n1029;
  assign n1031 = n1030 ^ n999;
  assign n2690 = n951 & n1031;
  assign n2695 = n2694 ^ n2690;
  assign n2687 = n1012 & n1021;
  assign n1025 = n1024 ^ n1019;
  assign n1022 = ~n999 & n1018;
  assign n1023 = n991 & n1022;
  assign n1026 = n1025 ^ n1023;
  assign n1046 = n949 & n1026;
  assign n2688 = n2687 ^ n1046;
  assign n2686 = n950 & n1037;
  assign n2689 = n2688 ^ n2686;
  assign n2696 = n2695 ^ n2689;
  assign n1032 = n1031 ^ n1026;
  assign n2683 = n977 & n1032;
  assign n1038 = n1037 ^ n1031;
  assign n1048 = n873 & n1038;
  assign n1027 = n1026 ^ n1021;
  assign n1039 = n1038 ^ n1027;
  assign n1047 = n993 & n1039;
  assign n1049 = n1048 ^ n1047;
  assign n2684 = n2683 ^ n1049;
  assign n1040 = n1001 & n1039;
  assign n1033 = n980 & n1032;
  assign n1028 = n933 & n1027;
  assign n1034 = n1033 ^ n1028;
  assign n1041 = n1040 ^ n1034;
  assign n2685 = n2684 ^ n1041;
  assign n2697 = n2696 ^ n2685;
  assign n7606 = n3766 ^ n2697;
  assign n7608 = n7607 ^ n7606;
  assign n1885 = x157 ^ x29;
  assign n1875 = x154 ^ x26;
  assign n1907 = n1885 ^ n1875;
  assign n1872 = x152 ^ x24;
  assign n1871 = x155 ^ x27;
  assign n1873 = n1872 ^ n1871;
  assign n1908 = n1907 ^ n1873;
  assign n1886 = n1885 ^ n1871;
  assign n1909 = n1886 & n1908;
  assign n1876 = x153 ^ x25;
  assign n1896 = n1885 ^ n1876;
  assign n1882 = x158 ^ x30;
  assign n1881 = x156 ^ x28;
  assign n1883 = n1882 ^ n1881;
  assign n1897 = n1896 ^ n1883;
  assign n1898 = n1873 & n1897;
  assign n1910 = n1909 ^ n1898;
  assign n1884 = n1883 ^ n1873;
  assign n1906 = n1896 ^ n1884;
  assign n1911 = n1910 ^ n1906;
  assign n1874 = x159 ^ x31;
  assign n1901 = n1884 ^ n1874;
  assign n1877 = n1876 ^ n1875;
  assign n1878 = n1877 ^ n1874;
  assign n1902 = n1882 ^ n1878;
  assign n1892 = n1885 ^ n1872;
  assign n1903 = n1902 ^ n1892;
  assign n1904 = n1901 & n1903;
  assign n1887 = n1882 ^ n1872;
  assign n1888 = n1887 ^ n1886;
  assign n1889 = n1884 & n1888;
  assign n1905 = n1904 ^ n1889;
  assign n1912 = n1911 ^ n1905;
  assign n1918 = n1878 & ~n1882;
  assign n1914 = n1907 ^ n1883;
  assign n1917 = n1887 & n1914;
  assign n1919 = n1918 ^ n1917;
  assign n1915 = n1914 ^ n1887;
  assign n1916 = n1915 ^ n1910;
  assign n1920 = n1919 ^ n1916;
  assign n1921 = n1912 & n1920;
  assign n1891 = n1884 ^ n1877;
  assign n1895 = n1891 & n1892;
  assign n1899 = n1898 ^ n1895;
  assign n1893 = n1892 ^ n1891;
  assign n1879 = n1878 ^ n1871;
  assign n1880 = n1874 & n1879;
  assign n1890 = n1889 ^ n1880;
  assign n1894 = n1893 ^ n1890;
  assign n1900 = n1899 ^ n1894;
  assign n1913 = n1912 ^ n1900;
  assign n1953 = n1921 ^ n1913;
  assign n1923 = n1879 ^ n1873;
  assign n1922 = n1914 ^ n1878;
  assign n1927 = n1923 ^ n1922;
  assign n1924 = n1922 & n1923;
  assign n1925 = n1924 ^ n1917;
  assign n1926 = n1925 ^ n1899;
  assign n1928 = n1927 ^ n1926;
  assign n1951 = ~n1900 & n1912;
  assign n1952 = n1928 & n1951;
  assign n1954 = n1953 ^ n1952;
  assign n1932 = n1928 ^ n1920;
  assign n1943 = n1932 ^ n1921;
  assign n1941 = n1900 & n1920;
  assign n1942 = ~n1928 & n1941;
  assign n1944 = n1943 ^ n1942;
  assign n1955 = n1954 ^ n1944;
  assign n1933 = n1921 ^ n1900;
  assign n1934 = n1932 & n1933;
  assign n1935 = n1934 ^ n1928;
  assign n1929 = n1928 ^ n1921;
  assign n1930 = n1913 & n1929;
  assign n1931 = n1930 ^ n1900;
  assign n1936 = n1935 ^ n1931;
  assign n2387 = n1955 ^ n1936;
  assign n2461 = n1908 & n2387;
  assign n1938 = n1897 & n1936;
  assign n2462 = n2461 ^ n1938;
  assign n2382 = n1901 & n1944;
  assign n1945 = n1944 ^ n1935;
  assign n2381 = n1888 & n1945;
  assign n2383 = n2382 ^ n2381;
  assign n1946 = n1884 & n1945;
  assign n2384 = n2383 ^ n1946;
  assign n2542 = n2462 ^ n2384;
  assign n2388 = n1886 & n2387;
  assign n1937 = n1873 & n1936;
  assign n2389 = n2388 ^ n1937;
  assign n2379 = n1903 & n1944;
  assign n2541 = n2389 ^ n2379;
  assign n2543 = n2542 ^ n2541;
  assign n2549 = n2548 ^ n2543;
  assign n2061 = x161 ^ x33;
  assign n2053 = x162 ^ x34;
  assign n2062 = n2061 ^ n2053;
  assign n2060 = x167 ^ x39;
  assign n2063 = n2062 ^ n2060;
  assign n2054 = x165 ^ x37;
  assign n2051 = x160 ^ x32;
  assign n2073 = n2054 ^ n2051;
  assign n2057 = x166 ^ x38;
  assign n2056 = x164 ^ x36;
  assign n2058 = n2057 ^ n2056;
  assign n2050 = x163 ^ x35;
  assign n2052 = n2051 ^ n2050;
  assign n2071 = n2058 ^ n2052;
  assign n2072 = n2071 ^ n2062;
  assign n2105 = n2073 ^ n2072;
  assign n2065 = n2063 ^ n2050;
  assign n2103 = n2060 & n2065;
  assign n2083 = n2054 ^ n2050;
  assign n2068 = n2057 ^ n2051;
  assign n2096 = n2083 ^ n2068;
  assign n2097 = n2071 & n2096;
  assign n2104 = n2103 ^ n2097;
  assign n2106 = n2105 ^ n2104;
  assign n2075 = n2061 ^ n2054;
  assign n2076 = n2075 ^ n2058;
  assign n2077 = n2052 & n2076;
  assign n2074 = n2072 & n2073;
  assign n2078 = n2077 ^ n2074;
  assign n2107 = n2106 ^ n2078;
  assign n2099 = n2075 ^ n2071;
  assign n2055 = n2054 ^ n2053;
  assign n2084 = n2055 ^ n2052;
  assign n2085 = n2083 & n2084;
  assign n2086 = n2085 ^ n2077;
  assign n2100 = n2099 ^ n2086;
  assign n2092 = n2071 ^ n2060;
  assign n2093 = n2063 ^ n2057;
  assign n2094 = n2093 ^ n2073;
  assign n2095 = n2092 & n2094;
  assign n2098 = n2097 ^ n2095;
  assign n2101 = n2100 ^ n2098;
  assign n2111 = n2107 ^ n2101;
  assign n2088 = ~n2057 & n2063;
  assign n2059 = n2058 ^ n2055;
  assign n2069 = n2059 & n2068;
  assign n2089 = n2088 ^ n2069;
  assign n2082 = n2068 ^ n2059;
  assign n2087 = n2086 ^ n2082;
  assign n2090 = n2089 ^ n2087;
  assign n2102 = n2090 & n2101;
  assign n2132 = n2111 ^ n2102;
  assign n2066 = n2065 ^ n2052;
  assign n2064 = n2063 ^ n2059;
  assign n2080 = n2066 ^ n2064;
  assign n2067 = n2064 & n2066;
  assign n2070 = n2069 ^ n2067;
  assign n2079 = n2078 ^ n2070;
  assign n2081 = n2080 ^ n2079;
  assign n2130 = n2101 & ~n2107;
  assign n2131 = n2081 & n2130;
  assign n2133 = n2132 ^ n2131;
  assign n2343 = n2063 & n2133;
  assign n2091 = n2090 ^ n2081;
  assign n2122 = n2102 ^ n2091;
  assign n2120 = n2090 & n2107;
  assign n2121 = ~n2081 & n2120;
  assign n2123 = n2122 ^ n2121;
  assign n2145 = n2094 & n2123;
  assign n2344 = n2343 ^ n2145;
  assign n2134 = n2133 ^ n2123;
  assign n2112 = n2102 ^ n2081;
  assign n2113 = n2111 & n2112;
  assign n2114 = n2113 ^ n2107;
  assign n2108 = n2107 ^ n2102;
  assign n2109 = n2091 & n2108;
  assign n2110 = n2109 ^ n2081;
  assign n2115 = n2114 ^ n2110;
  assign n2142 = n2134 ^ n2115;
  assign n2151 = n2084 & n2142;
  assign n2117 = n2076 & n2115;
  assign n2152 = n2151 ^ n2117;
  assign n2436 = n2344 ^ n2152;
  assign n2136 = n2133 ^ n2114;
  assign n2346 = n2059 & n2136;
  assign n2143 = n2083 & n2142;
  assign n2116 = n2052 & n2115;
  assign n2144 = n2143 ^ n2116;
  assign n2347 = n2346 ^ n2144;
  assign n2124 = n2123 ^ n2110;
  assign n2148 = n2096 & n2124;
  assign n2435 = n2347 ^ n2148;
  assign n2437 = n2436 ^ n2435;
  assign n2147 = n2092 & n2123;
  assign n2149 = n2148 ^ n2147;
  assign n2125 = n2071 & n2124;
  assign n2150 = n2149 ^ n2125;
  assign n2153 = n2152 ^ n2150;
  assign n2146 = n2145 ^ n2144;
  assign n2154 = n2153 ^ n2146;
  assign n2539 = n2437 ^ n2154;
  assign n2169 = x201 ^ x73;
  assign n2165 = x202 ^ x74;
  assign n2170 = n2169 ^ n2165;
  assign n2163 = x207 ^ x79;
  assign n2171 = n2170 ^ n2163;
  assign n2166 = x205 ^ x77;
  assign n2182 = n2169 ^ n2166;
  assign n2160 = x206 ^ x78;
  assign n2159 = x204 ^ x76;
  assign n2161 = n2160 ^ n2159;
  assign n2157 = x200 ^ x72;
  assign n2156 = x203 ^ x75;
  assign n2158 = n2157 ^ n2156;
  assign n2162 = n2161 ^ n2158;
  assign n2211 = n2182 ^ n2162;
  assign n2167 = n2166 ^ n2165;
  assign n2189 = n2167 ^ n2158;
  assign n2190 = n2166 ^ n2156;
  assign n2191 = n2189 & n2190;
  assign n2183 = n2182 ^ n2161;
  assign n2184 = n2158 & n2183;
  assign n2192 = n2191 ^ n2184;
  assign n2212 = n2211 ^ n2192;
  assign n2164 = n2163 ^ n2162;
  assign n2207 = n2171 ^ n2160;
  assign n2179 = n2166 ^ n2157;
  assign n2208 = n2207 ^ n2179;
  assign n2209 = n2164 & n2208;
  assign n2176 = n2160 ^ n2157;
  assign n2199 = n2190 ^ n2176;
  assign n2200 = n2162 & n2199;
  assign n2210 = n2209 ^ n2200;
  assign n2213 = n2212 ^ n2210;
  assign n2180 = n2170 ^ n2162;
  assign n2202 = n2180 ^ n2179;
  assign n2173 = n2171 ^ n2156;
  assign n2198 = n2163 & n2173;
  assign n2201 = n2200 ^ n2198;
  assign n2203 = n2202 ^ n2201;
  assign n2181 = n2179 & n2180;
  assign n2185 = n2184 ^ n2181;
  assign n2204 = n2203 ^ n2185;
  assign n2229 = n2213 ^ n2204;
  assign n2195 = ~n2160 & n2171;
  assign n2168 = n2167 ^ n2161;
  assign n2177 = n2168 & n2176;
  assign n2196 = n2195 ^ n2177;
  assign n2193 = n2176 ^ n2168;
  assign n2194 = n2193 ^ n2192;
  assign n2197 = n2196 ^ n2194;
  assign n2214 = n2197 & n2213;
  assign n2230 = n2229 ^ n2214;
  assign n2174 = n2173 ^ n2158;
  assign n2172 = n2171 ^ n2168;
  assign n2187 = n2174 ^ n2172;
  assign n2175 = n2172 & n2174;
  assign n2178 = n2177 ^ n2175;
  assign n2186 = n2185 ^ n2178;
  assign n2188 = n2187 ^ n2186;
  assign n2227 = ~n2204 & n2213;
  assign n2228 = n2188 & n2227;
  assign n2231 = n2230 ^ n2228;
  assign n2410 = n2171 & n2231;
  assign n2215 = n2197 ^ n2188;
  assign n2216 = n2215 ^ n2214;
  assign n2205 = n2197 & n2204;
  assign n2206 = ~n2188 & n2205;
  assign n2217 = n2216 ^ n2206;
  assign n2245 = n2208 & n2217;
  assign n2411 = n2410 ^ n2245;
  assign n2233 = n2214 ^ n2188;
  assign n2234 = n2229 & n2233;
  assign n2235 = n2234 ^ n2204;
  assign n2219 = n2214 ^ n2204;
  assign n2220 = n2215 & n2219;
  assign n2221 = n2220 ^ n2188;
  assign n2236 = n2235 ^ n2221;
  assign n2239 = n2183 & n2236;
  assign n2232 = n2231 ^ n2217;
  assign n2237 = n2236 ^ n2232;
  assign n2238 = n2189 & n2237;
  assign n2240 = n2239 ^ n2238;
  assign n2536 = n2411 ^ n2240;
  assign n2357 = n2235 ^ n2231;
  assign n2514 = n2168 & n2357;
  assign n2243 = n2158 & n2236;
  assign n2242 = n2190 & n2237;
  assign n2244 = n2243 ^ n2242;
  assign n2515 = n2514 ^ n2244;
  assign n2222 = n2221 ^ n2217;
  assign n2223 = n2199 & n2222;
  assign n2535 = n2515 ^ n2223;
  assign n2537 = n2536 ^ n2535;
  assign n2259 = x247 ^ x119;
  assign n2257 = x241 ^ x113;
  assign n2254 = x242 ^ x114;
  assign n2258 = n2257 ^ n2254;
  assign n2260 = n2259 ^ n2258;
  assign n2249 = x245 ^ x117;
  assign n2248 = x243 ^ x115;
  assign n2250 = n2249 ^ n2248;
  assign n2263 = x240 ^ x112;
  assign n2264 = n2263 ^ n2248;
  assign n2255 = n2254 ^ n2249;
  assign n2289 = n2264 ^ n2255;
  assign n2290 = n2250 & n2289;
  assign n2274 = n2257 ^ n2249;
  assign n2252 = x246 ^ x118;
  assign n2251 = x244 ^ x116;
  assign n2253 = n2252 ^ n2251;
  assign n2275 = n2274 ^ n2253;
  assign n2276 = n2264 & n2275;
  assign n2291 = n2290 ^ n2276;
  assign n2271 = n2264 ^ n2253;
  assign n2288 = n2274 ^ n2271;
  assign n2292 = n2291 ^ n2288;
  assign n2283 = n2260 ^ n2252;
  assign n2270 = n2263 ^ n2249;
  assign n2284 = n2283 ^ n2270;
  assign n2285 = n2271 ^ n2259;
  assign n2286 = n2284 & n2285;
  assign n2267 = n2263 ^ n2252;
  assign n2281 = n2267 ^ n2250;
  assign n2282 = n2271 & n2281;
  assign n2287 = n2286 ^ n2282;
  assign n2293 = n2292 ^ n2287;
  assign n2304 = ~n2252 & n2260;
  assign n2256 = n2255 ^ n2253;
  assign n2268 = n2256 & n2267;
  assign n2305 = n2304 ^ n2268;
  assign n2302 = n2267 ^ n2256;
  assign n2303 = n2302 ^ n2291;
  assign n2306 = n2305 ^ n2303;
  assign n2307 = n2293 & n2306;
  assign n2272 = n2271 ^ n2258;
  assign n2296 = n2272 ^ n2270;
  assign n2262 = n2260 ^ n2248;
  assign n2294 = n2259 & n2262;
  assign n2295 = n2294 ^ n2282;
  assign n2297 = n2296 ^ n2295;
  assign n2273 = n2270 & n2272;
  assign n2277 = n2276 ^ n2273;
  assign n2298 = n2297 ^ n2277;
  assign n2301 = n2298 ^ n2293;
  assign n2308 = n2307 ^ n2301;
  assign n2265 = n2264 ^ n2262;
  assign n2261 = n2260 ^ n2256;
  assign n2279 = n2265 ^ n2261;
  assign n2266 = n2261 & n2265;
  assign n2269 = n2268 ^ n2266;
  assign n2278 = n2277 ^ n2269;
  assign n2280 = n2279 ^ n2278;
  assign n2299 = n2293 & ~n2298;
  assign n2300 = n2280 & n2299;
  assign n2309 = n2308 ^ n2300;
  assign n2417 = n2260 & n2309;
  assign n2312 = n2306 ^ n2280;
  assign n2313 = n2312 ^ n2307;
  assign n2310 = n2298 & n2306;
  assign n2311 = ~n2280 & n2310;
  assign n2314 = n2313 ^ n2311;
  assign n2327 = n2284 & n2314;
  assign n2418 = n2417 ^ n2327;
  assign n2319 = n2307 ^ n2280;
  assign n2320 = n2301 & n2319;
  assign n2321 = n2320 ^ n2298;
  assign n2316 = n2307 ^ n2298;
  assign n2317 = n2312 & n2316;
  assign n2318 = n2317 ^ n2280;
  assign n2322 = n2321 ^ n2318;
  assign n2336 = n2275 & n2322;
  assign n2315 = n2314 ^ n2309;
  assign n2323 = n2322 ^ n2315;
  assign n2335 = n2289 & n2323;
  assign n2337 = n2336 ^ n2335;
  assign n2533 = n2418 ^ n2337;
  assign n2370 = n2321 ^ n2309;
  assign n2510 = n2256 & n2370;
  assign n2325 = n2264 & n2322;
  assign n2324 = n2250 & n2323;
  assign n2326 = n2325 ^ n2324;
  assign n2511 = n2510 ^ n2326;
  assign n2329 = n2318 ^ n2314;
  assign n2332 = n2281 & n2329;
  assign n2532 = n2511 ^ n2332;
  assign n2534 = n2533 ^ n2532;
  assign n2538 = n2537 ^ n2534;
  assign n2540 = n2539 ^ n2538;
  assign n2550 = n2549 ^ n2540;
  assign n2456 = n1922 & n1931;
  assign n1940 = n1874 & n1935;
  assign n2520 = n2456 ^ n1940;
  assign n2521 = n2520 ^ n2383;
  assign n2378 = n1878 & n1954;
  assign n2380 = n2379 ^ n2378;
  assign n2519 = n2389 ^ n2380;
  assign n2522 = n2521 ^ n2519;
  assign n2463 = n2462 ^ n2380;
  assign n1957 = n1954 ^ n1931;
  assign n2386 = n1914 & n1957;
  assign n2390 = n2389 ^ n2386;
  assign n2460 = n2390 ^ n2381;
  assign n2464 = n2463 ^ n2460;
  assign n2523 = n2522 ^ n2464;
  assign n2530 = n2529 ^ n2523;
  assign n2225 = n2162 & n2222;
  assign n2218 = n2164 & n2217;
  assign n2224 = n2223 ^ n2218;
  assign n2226 = n2225 ^ n2224;
  assign n2513 = n2411 ^ n2226;
  assign n2516 = n2515 ^ n2513;
  assign n2331 = n2285 & n2314;
  assign n2333 = n2332 ^ n2331;
  assign n2330 = n2271 & n2329;
  assign n2334 = n2333 ^ n2330;
  assign n2509 = n2418 ^ n2334;
  assign n2512 = n2511 ^ n2509;
  assign n2517 = n2516 ^ n2512;
  assign n2427 = n2064 & n2114;
  assign n2119 = n2060 & n2110;
  assign n2501 = n2427 ^ n2119;
  assign n2502 = n2501 ^ n2149;
  assign n2500 = n2344 ^ n2144;
  assign n2503 = n2502 ^ n2500;
  assign n2507 = n2503 ^ n2437;
  assign n2345 = n2344 ^ n2150;
  assign n2348 = n2347 ^ n2345;
  assign n2508 = n2507 ^ n2348;
  assign n2518 = n2517 ^ n2508;
  assign n2531 = n2530 ^ n2518;
  assign n2551 = n2550 ^ n2531;
  assign n2495 = n2065 & n2110;
  assign n2496 = n2495 ^ n2344;
  assign n2127 = n2066 & n2114;
  assign n2126 = n2125 ^ n2119;
  assign n2128 = n2127 ^ n2126;
  assign n2497 = n2496 ^ n2128;
  assign n2138 = n2072 & n2134;
  assign n2137 = n2068 & n2136;
  assign n2139 = n2138 ^ n2137;
  assign n2429 = n2151 ^ n2139;
  assign n2494 = n2429 ^ n2347;
  assign n2498 = n2497 ^ n2494;
  assign n2499 = n2498 ^ n2437;
  assign n2504 = n2503 ^ n2499;
  assign n2481 = n1879 & n1935;
  assign n2482 = n2481 ^ n2380;
  assign n1948 = n1923 & n1931;
  assign n1947 = n1946 ^ n1940;
  assign n1949 = n1948 ^ n1947;
  assign n2483 = n2482 ^ n1949;
  assign n1959 = n1891 & n1955;
  assign n1958 = n1887 & n1957;
  assign n1960 = n1959 ^ n1958;
  assign n2479 = n2461 ^ n1960;
  assign n2480 = n2479 ^ n2390;
  assign n2484 = n2483 ^ n2480;
  assign n2485 = n2484 ^ n2464;
  assign n2493 = n2492 ^ n2485;
  assign n2505 = n2504 ^ n2493;
  assign n2455 = n1902 & n1954;
  assign n2457 = n2456 ^ n2455;
  assign n2458 = n2457 ^ n1947;
  assign n2454 = n2390 ^ n1958;
  assign n2459 = n2458 ^ n2454;
  assign n2465 = n2464 ^ n2459;
  assign n2476 = n2475 ^ n2465;
  assign n2450 = n2417 ^ n2326;
  assign n2372 = n2272 & n2315;
  assign n2371 = n2267 & n2370;
  assign n2373 = n2372 ^ n2371;
  assign n2448 = n2373 ^ n2335;
  assign n2446 = n2283 & n2309;
  assign n2420 = n2261 & n2321;
  assign n2447 = n2446 ^ n2420;
  assign n2449 = n2448 ^ n2447;
  assign n2451 = n2450 ^ n2449;
  assign n2444 = n2410 ^ n2244;
  assign n2441 = n2207 & n2231;
  assign n2413 = n2172 & n2235;
  assign n2442 = n2441 ^ n2413;
  assign n2359 = n2180 & n2232;
  assign n2358 = n2176 & n2357;
  assign n2360 = n2359 ^ n2358;
  assign n2440 = n2360 ^ n2238;
  assign n2443 = n2442 ^ n2440;
  assign n2445 = n2444 ^ n2443;
  assign n2452 = n2451 ^ n2445;
  assign n2426 = n2093 & n2133;
  assign n2428 = n2427 ^ n2426;
  assign n2433 = n2428 ^ n2126;
  assign n2432 = n2347 ^ n2137;
  assign n2434 = n2433 ^ n2432;
  assign n2438 = n2437 ^ n2434;
  assign n2430 = n2429 ^ n2428;
  assign n2425 = n2343 ^ n2144;
  assign n2431 = n2430 ^ n2425;
  assign n2439 = n2438 ^ n2431;
  assign n2453 = n2452 ^ n2439;
  assign n2477 = n2476 ^ n2453;
  assign n2363 = n2259 & n2318;
  assign n2421 = n2420 ^ n2363;
  assign n2422 = n2421 ^ n2333;
  assign n2419 = n2418 ^ n2326;
  assign n2423 = n2422 ^ n2419;
  assign n2350 = n2163 & n2221;
  assign n2414 = n2413 ^ n2350;
  assign n2415 = n2414 ^ n2224;
  assign n2412 = n2411 ^ n2244;
  assign n2416 = n2415 ^ n2412;
  assign n2424 = n2423 ^ n2416;
  assign n2478 = n2477 ^ n2424;
  assign n2506 = n2505 ^ n2478;
  assign n2552 = n2551 ^ n2506;
  assign n2351 = n2350 ^ n2225;
  assign n2564 = n2442 ^ n2351;
  assign n2563 = n2515 ^ n2358;
  assign n2565 = n2564 ^ n2563;
  assign n2364 = n2363 ^ n2330;
  assign n2561 = n2447 ^ n2364;
  assign n2560 = n2511 ^ n2371;
  assign n2562 = n2561 ^ n2560;
  assign n2566 = n2565 ^ n2562;
  assign n2567 = n2566 ^ n2438;
  assign n2559 = n2558 ^ n2464;
  assign n2568 = n2567 ^ n2559;
  assign n2385 = n2384 ^ n2380;
  assign n2391 = n2390 ^ n2385;
  assign n2407 = n2406 ^ n2391;
  assign n2369 = n2270 & n2315;
  assign n2374 = n2373 ^ n2369;
  assign n2367 = n2336 ^ n2325;
  assign n2365 = n2265 & n2321;
  assign n2366 = n2365 ^ n2364;
  assign n2368 = n2367 ^ n2366;
  assign n2375 = n2374 ^ n2368;
  assign n2356 = n2179 & n2232;
  assign n2361 = n2360 ^ n2356;
  assign n2354 = n2243 ^ n2239;
  assign n2352 = n2174 & n2235;
  assign n2353 = n2352 ^ n2351;
  assign n2355 = n2354 ^ n2353;
  assign n2362 = n2361 ^ n2355;
  assign n2376 = n2375 ^ n2362;
  assign n2135 = n2073 & n2134;
  assign n2140 = n2139 ^ n2135;
  assign n2118 = n2117 ^ n2116;
  assign n2129 = n2128 ^ n2118;
  assign n2141 = n2140 ^ n2129;
  assign n2349 = n2348 ^ n2141;
  assign n2377 = n2376 ^ n2349;
  assign n2408 = n2407 ^ n2377;
  assign n2338 = n2337 ^ n2334;
  assign n2328 = n2327 ^ n2326;
  assign n2339 = n2338 ^ n2328;
  assign n2246 = n2245 ^ n2244;
  assign n2241 = n2240 ^ n2226;
  assign n2247 = n2246 ^ n2241;
  assign n2340 = n2339 ^ n2247;
  assign n2155 = n2154 ^ n2141;
  assign n2341 = n2340 ^ n2155;
  assign n1956 = n1892 & n1955;
  assign n1961 = n1960 ^ n1956;
  assign n1939 = n1938 ^ n1937;
  assign n1950 = n1949 ^ n1939;
  assign n1962 = n1961 ^ n1950;
  assign n2049 = n2048 ^ n1962;
  assign n2342 = n2341 ^ n2049;
  assign n2409 = n2408 ^ n2342;
  assign n2569 = n2568 ^ n2409;
  assign n2637 = ~n2477 & n2569;
  assign n2594 = n2498 ^ n2431;
  assign n2589 = n2173 & n2221;
  assign n2590 = n2589 ^ n2411;
  assign n2591 = n2590 ^ n2353;
  assign n2588 = n2515 ^ n2440;
  assign n2592 = n2591 ^ n2588;
  assign n2584 = n2262 & n2318;
  assign n2585 = n2584 ^ n2418;
  assign n2586 = n2585 ^ n2366;
  assign n2583 = n2511 ^ n2448;
  assign n2587 = n2586 ^ n2583;
  assign n2593 = n2592 ^ n2587;
  assign n2595 = n2594 ^ n2593;
  assign n2573 = n2389 ^ n2378;
  assign n2572 = n2479 ^ n2457;
  assign n2574 = n2573 ^ n2572;
  assign n2582 = n2581 ^ n2574;
  assign n2596 = n2595 ^ n2582;
  assign n2597 = n2596 ^ n2408;
  assign n2598 = n2597 ^ n2506;
  assign n2601 = n2550 ^ n2477;
  assign n2602 = n2598 & n2601;
  assign n2638 = n2637 ^ n2602;
  assign n2635 = n2601 ^ n2598;
  assign n2614 = n2596 ^ n2531;
  assign n2615 = n2597 ^ n2551;
  assign n2616 = n2614 & n2615;
  assign n2606 = n2596 ^ n2342;
  assign n2607 = n2606 ^ n2506;
  assign n2608 = n2551 & n2607;
  assign n2617 = n2616 ^ n2608;
  assign n2636 = n2635 ^ n2617;
  assign n2639 = n2638 ^ n2636;
  assign n2599 = n2598 ^ n2569;
  assign n2570 = n2569 ^ n2531;
  assign n2571 = n2570 ^ n2551;
  assign n2611 = n2599 ^ n2571;
  assign n2553 = n2552 ^ n2409;
  assign n2604 = n2596 ^ n2550;
  assign n2605 = n2553 & n2604;
  assign n2609 = n2608 ^ n2605;
  assign n2600 = n2571 & n2599;
  assign n2603 = n2602 ^ n2600;
  assign n2610 = n2609 ^ n2603;
  assign n2612 = n2611 ^ n2610;
  assign n2645 = n2639 ^ n2612;
  assign n2621 = n2569 ^ n2477;
  assign n2622 = n2621 ^ n2604;
  assign n2623 = n2568 ^ n2552;
  assign n2624 = n2622 & n2623;
  assign n2619 = n2614 ^ n2601;
  assign n2620 = n2552 & n2619;
  assign n2625 = n2624 ^ n2620;
  assign n2613 = n2606 ^ n2552;
  assign n2618 = n2617 ^ n2613;
  assign n2626 = n2625 ^ n2618;
  assign n2640 = n2626 & n2639;
  assign n2629 = n2604 ^ n2553;
  assign n2627 = n2568 & n2570;
  assign n2628 = n2627 ^ n2620;
  assign n2630 = n2629 ^ n2628;
  assign n2631 = n2630 ^ n2609;
  assign n2656 = n2640 ^ n2631;
  assign n2657 = n2645 & n2656;
  assign n2658 = n2657 ^ n2612;
  assign n2646 = n2645 ^ n2640;
  assign n2643 = n2631 & n2639;
  assign n2644 = ~n2612 & n2643;
  assign n2647 = n2646 ^ n2644;
  assign n2676 = n2658 ^ n2647;
  assign n2677 = n2552 & n2676;
  assign n2675 = n2568 & n2658;
  assign n2678 = n2677 ^ n2675;
  assign n2634 = n2631 ^ n2626;
  assign n2650 = n2640 ^ n2612;
  assign n2651 = n2634 & n2650;
  assign n2652 = n2651 ^ n2631;
  assign n2674 = n2571 & n2652;
  assign n2679 = n2678 ^ n2674;
  assign n2671 = n2622 & n2647;
  assign n2641 = n2640 ^ n2634;
  assign n2632 = n2626 & ~n2631;
  assign n2633 = n2612 & n2632;
  assign n2642 = n2641 ^ n2633;
  assign n2670 = n2569 & n2642;
  assign n2672 = n2671 ^ n2670;
  assign n2669 = n2570 & n2658;
  assign n2673 = n2672 ^ n2669;
  assign n2680 = n2679 ^ n2673;
  assign n2653 = n2652 ^ n2642;
  assign n2666 = n2598 & n2653;
  assign n2659 = n2658 ^ n2652;
  assign n2664 = n2551 & n2659;
  assign n2648 = n2647 ^ n2642;
  assign n2660 = n2659 ^ n2648;
  assign n2663 = n2614 & n2660;
  assign n2665 = n2664 ^ n2663;
  assign n2667 = n2666 ^ n2665;
  assign n2661 = n2615 & n2660;
  assign n2654 = n2601 & n2653;
  assign n2649 = n2553 & n2648;
  assign n2655 = n2654 ^ n2649;
  assign n2662 = n2661 ^ n2655;
  assign n2668 = n2667 ^ n2662;
  assign n2681 = n2680 ^ n2668;
  assign n7605 = n7604 ^ n2681;
  assign n7609 = n7608 ^ n7605;
  assign n3643 = n2623 & n2647;
  assign n3642 = n2619 & n2676;
  assign n3644 = n3643 ^ n3642;
  assign n3645 = n3644 ^ n2677;
  assign n3801 = n3645 ^ n2672;
  assign n3802 = n3801 ^ n2667;
  assign n7580 = n7579 ^ n3802;
  assign n3683 = n3418 & n3496;
  assign n3684 = n3683 ^ n3498;
  assign n3508 = ~n3452 & n3489;
  assign n3509 = n3508 ^ n3507;
  assign n3867 = n3684 ^ n3509;
  assign n3512 = n3495 ^ n3489;
  assign n3680 = n3455 & n3512;
  assign n3503 = n3422 & n3483;
  assign n3504 = n3503 ^ n3502;
  assign n3866 = n3680 ^ n3504;
  assign n3868 = n3867 ^ n3866;
  assign n3511 = ~n3439 & n3495;
  assign n3769 = n3731 ^ n3511;
  assign n3679 = ~n3450 & n3489;
  assign n3681 = n3680 ^ n3679;
  assign n3770 = n3769 ^ n3681;
  assign n3768 = n3509 ^ n3502;
  assign n3771 = n3770 ^ n3768;
  assign n7576 = n3868 ^ n3771;
  assign n3807 = n1833 & n1839;
  assign n3717 = n1811 & n3667;
  assign n3808 = n3807 ^ n3717;
  assign n3806 = n3666 ^ n1860;
  assign n3809 = n3808 ^ n3806;
  assign n3805 = n3723 ^ n1867;
  assign n3810 = n3809 ^ n3805;
  assign n3671 = n1804 & n1856;
  assign n3721 = n3671 ^ n1858;
  assign n3724 = n3723 ^ n3721;
  assign n3720 = n3719 ^ n3717;
  assign n3725 = n3724 ^ n3720;
  assign n3811 = n3810 ^ n3725;
  assign n7577 = n7576 ^ n3811;
  assign n3834 = n3808 ^ n3668;
  assign n3835 = n3834 ^ n3723;
  assign n3836 = n3835 ^ n3719;
  assign n3654 = n1013 & n1021;
  assign n3653 = n994 & n2692;
  assign n3655 = n3654 ^ n3653;
  assign n3656 = n3655 ^ n2693;
  assign n3799 = n3656 ^ n2688;
  assign n3800 = n3799 ^ n2684;
  assign n3837 = n3836 ^ n3800;
  assign n7578 = n7577 ^ n3837;
  assign n7581 = n7580 ^ n7578;
  assign n7615 = n7609 ^ n7581;
  assign n3830 = n3294 & n3490;
  assign n3831 = n3830 ^ n3492;
  assign n3828 = n3683 ^ n3501;
  assign n3515 = ~n3443 & n3482;
  assign n3513 = n3361 & n3512;
  assign n3514 = n3513 ^ n3511;
  assign n3516 = n3515 ^ n3514;
  assign n3829 = n3828 ^ n3516;
  assign n3832 = n3831 ^ n3829;
  assign n3674 = n1801 & n1845;
  assign n3675 = n3674 ^ n1852;
  assign n3672 = n3671 ^ n1866;
  assign n3673 = n3672 ^ n3670;
  assign n3676 = n3675 ^ n3673;
  assign n7598 = n3832 ^ n3676;
  assign n3863 = n3834 ^ n3721;
  assign n3862 = n3722 ^ n1867;
  assign n3864 = n3863 ^ n3862;
  assign n3651 = n986 & n1038;
  assign n3652 = n3651 ^ n1040;
  assign n3657 = n3656 ^ n3652;
  assign n3650 = n2687 ^ n1049;
  assign n3658 = n3657 ^ n3650;
  assign n3865 = n3864 ^ n3658;
  assign n7599 = n7598 ^ n3865;
  assign n3646 = n2607 & n2659;
  assign n3647 = n3646 ^ n2661;
  assign n3648 = n3647 ^ n3645;
  assign n3641 = n2671 ^ n2665;
  assign n3649 = n3648 ^ n3641;
  assign n7597 = n7596 ^ n3649;
  assign n7600 = n7599 ^ n7597;
  assign n3682 = n3681 ^ n3513;
  assign n3813 = n3682 ^ n3509;
  assign n3814 = n3813 ^ n3504;
  assign n7593 = n3836 ^ n3814;
  assign n3662 = n983 & n1027;
  assign n3663 = n3662 ^ n1034;
  assign n3660 = n3651 ^ n1048;
  assign n3661 = n3660 ^ n2695;
  assign n3664 = n3663 ^ n3661;
  assign n3677 = n3676 ^ n3664;
  assign n7594 = n7593 ^ n3677;
  assign n3824 = n2604 & n2648;
  assign n3825 = n3824 ^ n2655;
  assign n3822 = n3646 ^ n2664;
  assign n3823 = n3822 ^ n2679;
  assign n3826 = n3825 ^ n3823;
  assign n7592 = n7591 ^ n3826;
  assign n7595 = n7594 ^ n7592;
  assign n7601 = n7600 ^ n7595;
  assign n3686 = n3508 ^ n3502;
  assign n3685 = n3684 ^ n3682;
  assign n3687 = n3686 ^ n3685;
  assign n7573 = n3864 ^ n3687;
  assign n3738 = n3652 ^ n2688;
  assign n3737 = n3653 ^ n2684;
  assign n3739 = n3738 ^ n3737;
  assign n7572 = n3739 ^ n3725;
  assign n7574 = n7573 ^ n7572;
  assign n3853 = n3647 ^ n2672;
  assign n3852 = n3642 ^ n2667;
  assign n3854 = n3853 ^ n3852;
  assign n7571 = n7570 ^ n3854;
  assign n7575 = n7574 ^ n7571;
  assign n7582 = n7581 ^ n7575;
  assign n3506 = ~n3442 & n3495;
  assign n3510 = n3509 ^ n3506;
  assign n3517 = n3516 ^ n3510;
  assign n3505 = n3504 ^ n3499;
  assign n3518 = n3517 ^ n3505;
  assign n7566 = n3868 ^ n3518;
  assign n3767 = n3766 ^ n3725;
  assign n7567 = n7566 ^ n3767;
  assign n3704 = n2599 & n2652;
  assign n3705 = n3704 ^ n2675;
  assign n3706 = n3705 ^ n3644;
  assign n3703 = n2672 ^ n2665;
  assign n3707 = n3706 ^ n3703;
  assign n7565 = n7564 ^ n3707;
  assign n7568 = n7567 ^ n7565;
  assign n1042 = n978 & n1031;
  assign n3775 = n2691 ^ n1042;
  assign n3776 = n3775 ^ n3655;
  assign n3774 = n2688 ^ n1049;
  assign n3777 = n3776 ^ n3774;
  assign n7562 = n3810 ^ n3777;
  assign n3749 = n2670 ^ n2665;
  assign n3746 = n2621 & n2642;
  assign n3747 = n3746 ^ n3704;
  assign n3748 = n3747 ^ n2662;
  assign n3750 = n3749 ^ n3748;
  assign n7560 = n7559 ^ n3750;
  assign n3793 = n3732 ^ n3514;
  assign n3792 = n3504 ^ n3484;
  assign n3794 = n3793 ^ n3792;
  assign n7556 = n3868 ^ n3794;
  assign n3727 = n3669 ^ n1862;
  assign n3726 = n3719 ^ n1851;
  assign n3728 = n3727 ^ n3726;
  assign n3729 = n3728 ^ n3725;
  assign n7557 = n7556 ^ n3729;
  assign n1050 = n1049 ^ n1046;
  assign n1043 = n1011 & n1026;
  assign n1044 = n1043 ^ n1042;
  assign n1045 = n1044 ^ n1041;
  assign n1051 = n1050 ^ n1045;
  assign n1870 = n1869 ^ n1051;
  assign n7558 = n7557 ^ n1870;
  assign n7561 = n7560 ^ n7558;
  assign n7563 = n7562 ^ n7561;
  assign n7569 = n7568 ^ n7563;
  assign n7583 = n7582 ^ n7569;
  assign n7641 = n7601 ^ n7583;
  assign n7628 = n7609 ^ n7575;
  assign n7651 = n7641 ^ n7628;
  assign n3741 = n2694 ^ n1044;
  assign n3740 = n2684 ^ n1033;
  assign n3742 = n3741 ^ n3740;
  assign n7587 = n3742 ^ n3728;
  assign n7586 = n3868 ^ n3725;
  assign n7588 = n7587 ^ n7586;
  assign n3783 = n3747 ^ n2678;
  assign n3782 = n2667 ^ n2654;
  assign n3784 = n3783 ^ n3782;
  assign n7585 = n7584 ^ n3784;
  assign n7589 = n7588 ^ n7585;
  assign n7602 = n7601 ^ n7589;
  assign n7636 = n7602 ^ n7581;
  assign n7649 = n7589 & n7636;
  assign n7612 = n7575 ^ n7561;
  assign n7631 = n7615 ^ n7612;
  assign n7632 = n7583 & n7631;
  assign n7650 = n7649 ^ n7632;
  assign n7652 = n7651 ^ n7650;
  assign n7642 = n7628 & n7641;
  assign n7618 = n7609 ^ n7600;
  assign n7619 = n7618 ^ n7569;
  assign n7620 = n7582 & ~n7619;
  assign n7643 = n7642 ^ n7620;
  assign n7653 = n7652 ^ n7643;
  assign n7590 = n7589 ^ n7583;
  assign n7627 = n7602 ^ n7561;
  assign n7629 = n7628 ^ n7627;
  assign n7630 = n7590 & n7629;
  assign n7633 = n7632 ^ n7630;
  assign n7625 = n7618 ^ n7583;
  assign n7610 = n7609 ^ n7595;
  assign n7616 = n7610 ^ n7582;
  assign n7617 = n7615 & ~n7616;
  assign n7621 = n7620 ^ n7617;
  assign n7626 = n7625 ^ n7621;
  assign n7634 = n7633 ^ n7626;
  assign n7669 = n7653 ^ n7634;
  assign n7611 = n7610 ^ n7569;
  assign n7622 = n7612 ^ n7611;
  assign n7623 = n7622 ^ n7621;
  assign n7613 = ~n7611 & n7612;
  assign n7603 = ~n7561 & n7602;
  assign n7614 = n7613 ^ n7603;
  assign n7624 = n7623 ^ n7614;
  assign n7635 = ~n7624 & ~n7634;
  assign n7670 = n7669 ^ n7635;
  assign n7638 = n7611 ^ n7602;
  assign n7637 = n7636 ^ n7582;
  assign n7645 = n7638 ^ n7637;
  assign n7639 = n7637 & ~n7638;
  assign n7640 = n7639 ^ n7613;
  assign n7644 = n7643 ^ n7640;
  assign n7646 = n7645 ^ n7644;
  assign n7667 = ~n7634 & ~n7653;
  assign n7668 = ~n7646 & n7667;
  assign n7671 = n7670 ^ n7668;
  assign n7654 = ~n7624 & n7653;
  assign n7655 = n7646 & n7654;
  assign n7647 = n7646 ^ n7624;
  assign n7648 = n7647 ^ n7635;
  assign n7656 = n7655 ^ n7648;
  assign n7680 = n7671 ^ n7656;
  assign n7675 = n7646 ^ n7635;
  assign n7676 = ~n7669 & ~n7675;
  assign n7677 = n7676 ^ n7653;
  assign n7658 = n7653 ^ n7635;
  assign n7659 = n7647 & n7658;
  assign n7660 = n7659 ^ n7646;
  assign n7678 = n7677 ^ n7660;
  assign n7681 = n7680 ^ n7678;
  assign n7682 = n7615 & n7681;
  assign n7679 = n7582 & ~n7678;
  assign n7683 = n7682 ^ n7679;
  assign n7672 = n7602 & ~n7671;
  assign n7945 = n7683 ^ n7672;
  assign n7942 = n7627 & ~n7671;
  assign n7941 = ~n7638 & n7677;
  assign n7943 = n7942 ^ n7941;
  assign n7684 = n7677 ^ n7671;
  assign n7839 = n7612 & ~n7684;
  assign n7838 = n7641 & ~n7680;
  assign n7840 = n7839 ^ n7838;
  assign n7789 = ~n7616 & n7681;
  assign n7899 = n7840 ^ n7789;
  assign n7944 = n7943 ^ n7899;
  assign n7946 = n7945 ^ n7944;
  assign n7901 = n7636 & ~n7660;
  assign n7666 = n7629 & n7656;
  assign n7673 = n7672 ^ n7666;
  assign n7902 = n7901 ^ n7673;
  assign n7844 = n7589 & ~n7660;
  assign n7661 = n7660 ^ n7656;
  assign n7664 = n7583 & ~n7661;
  assign n7845 = n7844 ^ n7664;
  assign n7843 = n7637 & n7677;
  assign n7846 = n7845 ^ n7843;
  assign n7903 = n7902 ^ n7846;
  assign n7685 = ~n7611 & ~n7684;
  assign n7686 = n7685 ^ n7683;
  assign n7900 = n7899 ^ n7686;
  assign n7904 = n7903 ^ n7900;
  assign n12664 = n7946 ^ n7904;
  assign n4336 = n1753 ^ n555;
  assign n4334 = n940 ^ n827;
  assign n4335 = n4334 ^ n538;
  assign n4337 = n4336 ^ n4335;
  assign n4331 = n1740 ^ n819;
  assign n4328 = n921 ^ n893;
  assign n4329 = n4328 ^ n928;
  assign n4330 = n4329 ^ n815;
  assign n4332 = n4331 ^ n4330;
  assign n4325 = n876 ^ n861;
  assign n4324 = n922 ^ n885;
  assign n4326 = n4325 ^ n4324;
  assign n4327 = n4326 ^ n1717;
  assign n4333 = n4332 ^ n4327;
  assign n4338 = n4337 ^ n4333;
  assign n4360 = n1255 ^ n749;
  assign n4357 = n937 ^ n827;
  assign n4358 = n4357 ^ n741;
  assign n4356 = n965 ^ n538;
  assign n4359 = n4358 ^ n4356;
  assign n4361 = n4360 ^ n4359;
  assign n4411 = n4338 & ~n4361;
  assign n4343 = n965 ^ n649;
  assign n4344 = n4343 ^ n782;
  assign n4345 = n4344 ^ n774;
  assign n4346 = n4345 ^ n956;
  assign n4347 = n4346 ^ n1789;
  assign n4377 = n4347 ^ n4327;
  assign n4365 = n850 ^ n775;
  assign n4363 = n961 ^ n827;
  assign n4364 = n4363 ^ n806;
  assign n4366 = n4365 ^ n4364;
  assign n4355 = n1228 ^ n348;
  assign n4362 = n4361 ^ n4355;
  assign n4367 = n4366 ^ n4362;
  assign n4378 = n4377 ^ n4367;
  assign n4339 = n925 ^ n815;
  assign n4340 = n4339 ^ n834;
  assign n4341 = n4340 ^ n934;
  assign n4342 = n4341 ^ n1659;
  assign n4381 = n4361 ^ n4342;
  assign n4382 = n4378 & n4381;
  assign n4412 = n4411 ^ n4382;
  assign n4409 = n4381 ^ n4378;
  assign n4350 = n827 ^ n795;
  assign n4349 = n877 ^ n851;
  assign n4351 = n4350 ^ n4349;
  assign n4352 = n4351 ^ n857;
  assign n4353 = n4352 ^ n1644;
  assign n4387 = n4353 ^ n4347;
  assign n4354 = n4353 ^ n4342;
  assign n4396 = n4377 ^ n4354;
  assign n4397 = n4387 & n4396;
  assign n4371 = n4347 ^ n4332;
  assign n4372 = n4371 ^ n4367;
  assign n4373 = n4354 & n4372;
  assign n4398 = n4397 ^ n4373;
  assign n4410 = n4409 ^ n4398;
  assign n4413 = n4412 ^ n4410;
  assign n4379 = n4378 ^ n4338;
  assign n4375 = n4353 ^ n4338;
  assign n4376 = n4375 ^ n4354;
  assign n4385 = n4379 ^ n4376;
  assign n4380 = n4376 & n4379;
  assign n4383 = n4382 ^ n4380;
  assign n4348 = n4347 ^ n4342;
  assign n4368 = n4367 ^ n4354;
  assign n4369 = n4368 ^ n4333;
  assign n4370 = n4348 & n4369;
  assign n4374 = n4373 ^ n4370;
  assign n4384 = n4383 ^ n4374;
  assign n4386 = n4385 ^ n4384;
  assign n4420 = n4413 ^ n4386;
  assign n4395 = n4371 ^ n4368;
  assign n4399 = n4398 ^ n4395;
  assign n4390 = n4361 ^ n4338;
  assign n4391 = n4390 ^ n4348;
  assign n4392 = n4368 ^ n4337;
  assign n4393 = n4391 & n4392;
  assign n4388 = n4387 ^ n4381;
  assign n4389 = n4368 & n4388;
  assign n4394 = n4393 ^ n4389;
  assign n4400 = n4399 ^ n4394;
  assign n4414 = n4400 & n4413;
  assign n4403 = n4369 ^ n4348;
  assign n4401 = n4337 & n4375;
  assign n4402 = n4401 ^ n4389;
  assign n4404 = n4403 ^ n4402;
  assign n4405 = n4404 ^ n4374;
  assign n4425 = n4414 ^ n4405;
  assign n4426 = n4420 & n4425;
  assign n4427 = n4426 ^ n4386;
  assign n4718 = n4337 & n4427;
  assign n4408 = n4405 ^ n4400;
  assign n4435 = n4414 ^ n4386;
  assign n4436 = n4408 & n4435;
  assign n4437 = n4436 ^ n4405;
  assign n4669 = n4379 & n4437;
  assign n4719 = n4718 ^ n4669;
  assign n4421 = n4420 ^ n4414;
  assign n4418 = n4405 & n4413;
  assign n4419 = ~n4386 & n4418;
  assign n4422 = n4421 ^ n4419;
  assign n4430 = n4392 & n4422;
  assign n4428 = n4427 ^ n4422;
  assign n4429 = n4388 & n4428;
  assign n4431 = n4430 ^ n4429;
  assign n4720 = n4719 ^ n4431;
  assign n4441 = n4437 ^ n4427;
  assign n4444 = n4354 & n4441;
  assign n4415 = n4414 ^ n4408;
  assign n4406 = n4400 & ~n4405;
  assign n4407 = n4386 & n4406;
  assign n4416 = n4415 ^ n4407;
  assign n4440 = n4422 ^ n4416;
  assign n4442 = n4441 ^ n4440;
  assign n4443 = n4387 & n4442;
  assign n4445 = n4444 ^ n4443;
  assign n4423 = n4391 & n4422;
  assign n4417 = n4338 & n4416;
  assign n4424 = n4423 ^ n4417;
  assign n4717 = n4445 ^ n4424;
  assign n4721 = n4720 ^ n4717;
  assign n4597 = n4372 & n4441;
  assign n4596 = n4396 & n4442;
  assign n4598 = n4597 ^ n4596;
  assign n4599 = n4598 ^ n4424;
  assign n4438 = n4437 ^ n4416;
  assign n4439 = n4378 & n4438;
  assign n4446 = n4445 ^ n4439;
  assign n4595 = n4446 ^ n4429;
  assign n4600 = n4599 ^ n4595;
  assign n7440 = n4721 ^ n4600;
  assign n4231 = n2503 ^ n2416;
  assign n4229 = n2587 ^ n2534;
  assign n4230 = n4229 ^ n2485;
  assign n4232 = n4231 ^ n4230;
  assign n4226 = n3523 ^ n2574;
  assign n4223 = n2562 ^ n2534;
  assign n4224 = n4223 ^ n2465;
  assign n4222 = n2445 ^ n2431;
  assign n4225 = n4224 ^ n4222;
  assign n4227 = n4226 ^ n4225;
  assign n4221 = n3520 ^ n2522;
  assign n4228 = n4227 ^ n4221;
  assign n4233 = n4232 ^ n4228;
  assign n4218 = n3543 ^ n2391;
  assign n4215 = n2534 ^ n2423;
  assign n4216 = n4215 ^ n2523;
  assign n4214 = n2516 ^ n2348;
  assign n4217 = n4216 ^ n4214;
  assign n4219 = n4218 ^ n4217;
  assign n4210 = n2543 ^ n2339;
  assign n4209 = n2537 ^ n2437;
  assign n4211 = n4210 ^ n4209;
  assign n4208 = n3548 ^ n2464;
  assign n4212 = n4211 ^ n4208;
  assign n4220 = n4219 ^ n4212;
  assign n4234 = n4233 ^ n4220;
  assign n4198 = n2375 ^ n1962;
  assign n4197 = n2247 ^ n2154;
  assign n4199 = n4198 ^ n4197;
  assign n4196 = n3538 ^ n2543;
  assign n4200 = n4199 ^ n4196;
  assign n4193 = n2512 ^ n2391;
  assign n4192 = n2362 ^ n2141;
  assign n4194 = n4193 ^ n4192;
  assign n4191 = n3527 ^ n1962;
  assign n4195 = n4194 ^ n4191;
  assign n4201 = n4200 ^ n4195;
  assign n4187 = n2534 ^ n2465;
  assign n4188 = n4187 ^ n2565;
  assign n4189 = n4188 ^ n2434;
  assign n4190 = n4189 ^ n3535;
  assign n4202 = n4201 ^ n4190;
  assign n4277 = n4202 & ~n4227;
  assign n4205 = n2574 ^ n2451;
  assign n4204 = n2592 ^ n2498;
  assign n4206 = n4205 ^ n4204;
  assign n4203 = n3530 ^ n2484;
  assign n4207 = n4206 ^ n4203;
  assign n4243 = n4207 ^ n4195;
  assign n4244 = n4243 ^ n4233;
  assign n4247 = n4227 ^ n4212;
  assign n4248 = n4244 & n4247;
  assign n4278 = n4277 ^ n4248;
  assign n4275 = n4247 ^ n4244;
  assign n4254 = n4219 ^ n4207;
  assign n4255 = n4243 ^ n4220;
  assign n4256 = n4254 & n4255;
  assign n4237 = n4207 ^ n4200;
  assign n4238 = n4237 ^ n4233;
  assign n4239 = n4220 & n4238;
  assign n4257 = n4256 ^ n4239;
  assign n4276 = n4275 ^ n4257;
  assign n4279 = n4278 ^ n4276;
  assign n4245 = n4244 ^ n4202;
  assign n4241 = n4219 ^ n4202;
  assign n4242 = n4241 ^ n4220;
  assign n4251 = n4245 ^ n4242;
  assign n4246 = n4242 & n4245;
  assign n4249 = n4248 ^ n4246;
  assign n4213 = n4212 ^ n4207;
  assign n4235 = n4234 ^ n4201;
  assign n4236 = n4213 & n4235;
  assign n4240 = n4239 ^ n4236;
  assign n4250 = n4249 ^ n4240;
  assign n4252 = n4251 ^ n4250;
  assign n4286 = n4279 ^ n4252;
  assign n4261 = n4227 ^ n4202;
  assign n4262 = n4261 ^ n4213;
  assign n4263 = n4234 ^ n4190;
  assign n4264 = n4262 & n4263;
  assign n4259 = n4254 ^ n4247;
  assign n4260 = n4234 & n4259;
  assign n4265 = n4264 ^ n4260;
  assign n4253 = n4237 ^ n4234;
  assign n4258 = n4257 ^ n4253;
  assign n4266 = n4265 ^ n4258;
  assign n4280 = n4266 & n4279;
  assign n4269 = n4235 ^ n4213;
  assign n4267 = n4190 & n4241;
  assign n4268 = n4267 ^ n4260;
  assign n4270 = n4269 ^ n4268;
  assign n4271 = n4270 ^ n4240;
  assign n4295 = n4280 ^ n4271;
  assign n4296 = n4286 & n4295;
  assign n4297 = n4296 ^ n4252;
  assign n4287 = n4286 ^ n4280;
  assign n4284 = n4271 & n4279;
  assign n4285 = ~n4252 & n4284;
  assign n4288 = n4287 ^ n4285;
  assign n4307 = n4297 ^ n4288;
  assign n4611 = n4234 & n4307;
  assign n4309 = n4263 & n4288;
  assign n4308 = n4259 & n4307;
  assign n4310 = n4309 ^ n4308;
  assign n4612 = n4611 ^ n4310;
  assign n4289 = n4262 & n4288;
  assign n4274 = n4271 ^ n4266;
  assign n4281 = n4280 ^ n4274;
  assign n4272 = n4266 & ~n4271;
  assign n4273 = n4252 & n4272;
  assign n4282 = n4281 ^ n4273;
  assign n4283 = n4202 & n4282;
  assign n4290 = n4289 ^ n4283;
  assign n4789 = n4612 ^ n4290;
  assign n4292 = n4280 ^ n4252;
  assign n4293 = n4274 & n4292;
  assign n4294 = n4293 ^ n4271;
  assign n4313 = n4294 ^ n4282;
  assign n4314 = n4244 & n4313;
  assign n4298 = n4297 ^ n4294;
  assign n4301 = n4220 & n4298;
  assign n4291 = n4288 ^ n4282;
  assign n4299 = n4298 ^ n4291;
  assign n4300 = n4254 & n4299;
  assign n4302 = n4301 ^ n4300;
  assign n4315 = n4314 ^ n4302;
  assign n4790 = n4789 ^ n4315;
  assign n3988 = n3410 ^ n3388;
  assign n3989 = n3988 ^ n3386;
  assign n3987 = n3986 ^ n3299;
  assign n3990 = n3989 ^ n3987;
  assign n3982 = n3355 ^ n3290;
  assign n3983 = n3982 ^ n3284;
  assign n3981 = n3980 ^ n3226;
  assign n3984 = n3983 ^ n3981;
  assign n4003 = n3990 ^ n3984;
  assign n3969 = n3252 ^ n2791;
  assign n3971 = n3970 ^ n3969;
  assign n3968 = n3356 ^ n3320;
  assign n3972 = n3971 ^ n3968;
  assign n3963 = n3425 ^ n2791;
  assign n3965 = n3964 ^ n3963;
  assign n3961 = n3290 ^ n3208;
  assign n3962 = n3961 ^ n3190;
  assign n3966 = n3965 ^ n3962;
  assign n3967 = n3966 ^ n3335;
  assign n3973 = n3972 ^ n3967;
  assign n4004 = n4003 ^ n3973;
  assign n3993 = n3410 ^ n3159;
  assign n3994 = n3993 ^ n3405;
  assign n3992 = n3991 ^ n3366;
  assign n3995 = n3994 ^ n3992;
  assign n3999 = n3995 ^ n3984;
  assign n3957 = n3207 ^ n3159;
  assign n3958 = n3957 ^ n3067;
  assign n3956 = n3955 ^ n3394;
  assign n3959 = n3958 ^ n3956;
  assign n3951 = n3340 ^ n2791;
  assign n3953 = n3952 ^ n3951;
  assign n3949 = n3388 ^ n3321;
  assign n3950 = n3949 ^ n3316;
  assign n3954 = n3953 ^ n3950;
  assign n3960 = n3959 ^ n3954;
  assign n3974 = n3973 ^ n3960;
  assign n4038 = n3999 ^ n3974;
  assign n4016 = n3984 ^ n3954;
  assign n4017 = n4003 ^ n3960;
  assign n4018 = n4016 & n4017;
  assign n4000 = n3999 ^ n3973;
  assign n4001 = n3960 & n4000;
  assign n4019 = n4018 ^ n4001;
  assign n4039 = n4038 ^ n4019;
  assign n3977 = n3436 ^ n3208;
  assign n3976 = n3975 ^ n2791;
  assign n3978 = n3977 ^ n3976;
  assign n3979 = n3978 ^ n3974;
  assign n3996 = n3995 ^ n3990;
  assign n4005 = n3996 ^ n3978;
  assign n4034 = n4005 ^ n3966;
  assign n3985 = n3984 ^ n3959;
  assign n4035 = n4034 ^ n3985;
  assign n4036 = n3979 & n4035;
  assign n4010 = n3966 ^ n3959;
  assign n4026 = n4016 ^ n4010;
  assign n4027 = n3974 & n4026;
  assign n4037 = n4036 ^ n4027;
  assign n4040 = n4039 ^ n4037;
  assign n3997 = n3996 ^ n3974;
  assign n4029 = n3997 ^ n3985;
  assign n4007 = n4005 ^ n3954;
  assign n4025 = n3978 & n4007;
  assign n4028 = n4027 ^ n4025;
  assign n4030 = n4029 ^ n4028;
  assign n3998 = n3985 & n3997;
  assign n4002 = n4001 ^ n3998;
  assign n4031 = n4030 ^ n4002;
  assign n4056 = n4040 ^ n4031;
  assign n4022 = ~n3966 & n4005;
  assign n4011 = n4004 & n4010;
  assign n4023 = n4022 ^ n4011;
  assign n4020 = n4010 ^ n4004;
  assign n4021 = n4020 ^ n4019;
  assign n4024 = n4023 ^ n4021;
  assign n4041 = n4024 & n4040;
  assign n4008 = n4007 ^ n3960;
  assign n4006 = n4005 ^ n4004;
  assign n4014 = n4008 ^ n4006;
  assign n4009 = n4006 & n4008;
  assign n4012 = n4011 ^ n4009;
  assign n4013 = n4012 ^ n4002;
  assign n4015 = n4014 ^ n4013;
  assign n4064 = n4041 ^ n4015;
  assign n4065 = n4056 & n4064;
  assign n4066 = n4065 ^ n4031;
  assign n4057 = n4056 ^ n4041;
  assign n4054 = ~n4031 & n4040;
  assign n4055 = n4015 & n4054;
  assign n4058 = n4057 ^ n4055;
  assign n4072 = n4066 ^ n4058;
  assign n4073 = n4004 & n4072;
  assign n4042 = n4024 ^ n4015;
  assign n4046 = n4041 ^ n4031;
  assign n4047 = n4042 & n4046;
  assign n4048 = n4047 ^ n4015;
  assign n4067 = n4066 ^ n4048;
  assign n4070 = n3960 & n4067;
  assign n4043 = n4042 ^ n4041;
  assign n4032 = n4024 & n4031;
  assign n4033 = ~n4015 & n4032;
  assign n4044 = n4043 ^ n4033;
  assign n4063 = n4058 ^ n4044;
  assign n4068 = n4067 ^ n4063;
  assign n4069 = n4016 & n4068;
  assign n4071 = n4070 ^ n4069;
  assign n4074 = n4073 ^ n4071;
  assign n4060 = n4035 & n4044;
  assign n4059 = n4005 & n4058;
  assign n4061 = n4060 ^ n4059;
  assign n4049 = n4048 ^ n4044;
  assign n4052 = n3974 & n4049;
  assign n4050 = n4026 & n4049;
  assign n4045 = n3979 & n4044;
  assign n4051 = n4050 ^ n4045;
  assign n4053 = n4052 ^ n4051;
  assign n4062 = n4061 ^ n4053;
  assign n4075 = n4074 ^ n4062;
  assign n4791 = n4790 ^ n4075;
  assign n4318 = n4238 & n4298;
  assign n4317 = n4255 & n4299;
  assign n4319 = n4318 ^ n4317;
  assign n4320 = n4319 ^ n4290;
  assign n4316 = n4315 ^ n4308;
  assign n4321 = n4320 ^ n4316;
  assign n4305 = n4190 & n4297;
  assign n4304 = n4245 & n4294;
  assign n4306 = n4305 ^ n4304;
  assign n4311 = n4310 ^ n4306;
  assign n4303 = n4302 ^ n4290;
  assign n4312 = n4311 ^ n4303;
  assign n4322 = n4321 ^ n4312;
  assign n7439 = n4791 ^ n4322;
  assign n7441 = n7440 ^ n7439;
  assign n4501 = n1595 ^ n1577;
  assign n4500 = n1779 ^ n1351;
  assign n4502 = n4501 ^ n4500;
  assign n4499 = n4498 ^ n1776;
  assign n4503 = n4502 ^ n4499;
  assign n4485 = n1683 ^ n1616;
  assign n4486 = n4485 ^ n1730;
  assign n4484 = n4483 ^ n1700;
  assign n4487 = n4486 ^ n4484;
  assign n4504 = n4503 ^ n4487;
  assign n4477 = n1771 ^ n1668;
  assign n4478 = n4477 ^ n1596;
  assign n4476 = n4475 ^ n1143;
  assign n4479 = n4478 ^ n4476;
  assign n4473 = n1622 ^ n1584;
  assign n4469 = n1760 ^ n1668;
  assign n4470 = n4469 ^ n1455;
  assign n4471 = n4470 ^ n1780;
  assign n4468 = n4467 ^ n1243;
  assign n4472 = n4471 ^ n4468;
  assign n4474 = n4473 ^ n4472;
  assign n4480 = n4479 ^ n4474;
  assign n4505 = n4504 ^ n4480;
  assign n4491 = n1676 ^ n1672;
  assign n4490 = n1729 ^ n1692;
  assign n4492 = n4491 ^ n4490;
  assign n4489 = n4488 ^ n1733;
  assign n4493 = n4492 ^ n4489;
  assign n4514 = n4503 ^ n4493;
  assign n4463 = n1565 ^ n1454;
  assign n4462 = n1724 ^ n1672;
  assign n4464 = n4463 ^ n4462;
  assign n4461 = n4460 ^ n1653;
  assign n4465 = n4464 ^ n4461;
  assign n4456 = n1668 ^ n1607;
  assign n4457 = n4456 ^ n1623;
  assign n4458 = n4457 ^ n1684;
  assign n4455 = n4454 ^ n1630;
  assign n4459 = n4458 ^ n4455;
  assign n4466 = n4465 ^ n4459;
  assign n4481 = n4480 ^ n4466;
  assign n4544 = n4514 ^ n4481;
  assign n4521 = n4503 ^ n4459;
  assign n4530 = n4504 ^ n4466;
  assign n4531 = n4521 & n4530;
  assign n4515 = n4514 ^ n4480;
  assign n4516 = n4466 & n4515;
  assign n4532 = n4531 ^ n4516;
  assign n4545 = n4544 ^ n4532;
  assign n4451 = n1557 ^ n1444;
  assign n4450 = n1668 ^ n1454;
  assign n4452 = n4451 ^ n4450;
  assign n4449 = n4448 ^ n1749;
  assign n4453 = n4452 ^ n4449;
  assign n4482 = n4481 ^ n4453;
  assign n4494 = n4493 ^ n4487;
  assign n4495 = n4494 ^ n4453;
  assign n4540 = n4495 ^ n4472;
  assign n4512 = n4503 ^ n4465;
  assign n4541 = n4540 ^ n4512;
  assign n4542 = ~n4482 & ~n4541;
  assign n4508 = n4472 ^ n4465;
  assign n4522 = n4521 ^ n4508;
  assign n4523 = n4481 & n4522;
  assign n4543 = n4542 ^ n4523;
  assign n4546 = n4545 ^ n4543;
  assign n4511 = n4494 ^ n4481;
  assign n4526 = n4512 ^ n4511;
  assign n4496 = n4495 ^ n4459;
  assign n4524 = ~n4453 & ~n4496;
  assign n4525 = n4524 ^ n4523;
  assign n4527 = n4526 ^ n4525;
  assign n4513 = n4511 & n4512;
  assign n4517 = n4516 ^ n4513;
  assign n4528 = n4527 ^ n4517;
  assign n4561 = n4546 ^ n4528;
  assign n4534 = ~n4472 & ~n4495;
  assign n4509 = n4505 & n4508;
  assign n4535 = n4534 ^ n4509;
  assign n4529 = n4508 ^ n4505;
  assign n4533 = n4532 ^ n4529;
  assign n4536 = n4535 ^ n4533;
  assign n4547 = n4536 & n4546;
  assign n4506 = n4505 ^ n4495;
  assign n4497 = n4496 ^ n4466;
  assign n4519 = n4506 ^ n4497;
  assign n4507 = ~n4497 & ~n4506;
  assign n4510 = n4509 ^ n4507;
  assign n4518 = n4517 ^ n4510;
  assign n4520 = n4519 ^ n4518;
  assign n4569 = n4547 ^ n4520;
  assign n4570 = n4561 & n4569;
  assign n4571 = n4570 ^ n4528;
  assign n4562 = n4561 ^ n4547;
  assign n4559 = ~n4528 & n4546;
  assign n4560 = n4520 & n4559;
  assign n4563 = n4562 ^ n4560;
  assign n4577 = n4571 ^ n4563;
  assign n4578 = n4505 & n4577;
  assign n4539 = n4536 ^ n4520;
  assign n4551 = n4547 ^ n4528;
  assign n4552 = n4539 & n4551;
  assign n4553 = n4552 ^ n4520;
  assign n4572 = n4571 ^ n4553;
  assign n4575 = n4466 & n4572;
  assign n4548 = n4547 ^ n4539;
  assign n4537 = n4528 & n4536;
  assign n4538 = ~n4520 & n4537;
  assign n4549 = n4548 ^ n4538;
  assign n4568 = n4563 ^ n4549;
  assign n4573 = n4572 ^ n4568;
  assign n4574 = n4521 & n4573;
  assign n4576 = n4575 ^ n4574;
  assign n4579 = n4578 ^ n4576;
  assign n4565 = ~n4541 & n4549;
  assign n4564 = ~n4495 & n4563;
  assign n4566 = n4565 ^ n4564;
  assign n4554 = n4553 ^ n4549;
  assign n4557 = n4481 & n4554;
  assign n4555 = n4522 & n4554;
  assign n4550 = ~n4482 & n4549;
  assign n4556 = n4555 ^ n4550;
  assign n4558 = n4557 ^ n4556;
  assign n4567 = n4566 ^ n4558;
  assign n4580 = n4579 ^ n4567;
  assign n7442 = n7441 ^ n4580;
  assign n7443 = n7442 ^ n6727;
  assign n4806 = n4445 ^ n4423;
  assign n4432 = n4368 & n4428;
  assign n4433 = n4432 ^ n4431;
  assign n4805 = n4598 ^ n4433;
  assign n4807 = n4806 ^ n4805;
  assign n4614 = n4302 ^ n4289;
  assign n4613 = n4612 ^ n4319;
  assign n4615 = n4614 ^ n4613;
  assign n7428 = n4807 ^ n4615;
  assign n7429 = n7428 ^ n6726;
  assign n7430 = n7429 ^ n4321;
  assign n4603 = n4515 & n4572;
  assign n4602 = n4530 & n4573;
  assign n4604 = n4603 ^ n4602;
  assign n4605 = n4604 ^ n4566;
  assign n4601 = n4579 ^ n4555;
  assign n4606 = n4605 ^ n4601;
  assign n7431 = n7430 ^ n4606;
  assign n4182 = n4000 & n4067;
  assign n4181 = n4017 & n4068;
  assign n4183 = n4182 ^ n4181;
  assign n4184 = n4183 ^ n4061;
  assign n4180 = n4074 ^ n4050;
  assign n4185 = n4184 ^ n4180;
  assign n7432 = n7431 ^ n4185;
  assign n7461 = n7443 ^ n7432;
  assign n4811 = n4213 & n4291;
  assign n4700 = n4235 & n4291;
  assign n4659 = n4247 & n4313;
  assign n4701 = n4700 ^ n4659;
  assign n4812 = n4811 ^ n4701;
  assign n4809 = n4318 ^ n4301;
  assign n4706 = n4242 & n4294;
  assign n4663 = n4611 ^ n4305;
  assign n4707 = n4706 ^ n4663;
  assign n4810 = n4809 ^ n4707;
  assign n4813 = n4812 ^ n4810;
  assign n4785 = n4348 & n4440;
  assign n4672 = n4369 & n4440;
  assign n4671 = n4381 & n4438;
  assign n4673 = n4672 ^ n4671;
  assign n4786 = n4785 ^ n4673;
  assign n4783 = n4597 ^ n4444;
  assign n4751 = n4376 & n4437;
  assign n4750 = n4718 ^ n4432;
  assign n4752 = n4751 ^ n4750;
  assign n4784 = n4783 ^ n4752;
  assign n4787 = n4786 ^ n4784;
  assign n7454 = n4813 ^ n4787;
  assign n4609 = n4183 ^ n4053;
  assign n4608 = n4071 ^ n4060;
  assign n4610 = n4609 ^ n4608;
  assign n4616 = n4615 ^ n4610;
  assign n7455 = n7454 ^ n4616;
  assign n4803 = n4576 ^ n4565;
  assign n4802 = n4604 ^ n4558;
  assign n4804 = n4803 ^ n4802;
  assign n7456 = n7455 ^ n4804;
  assign n7457 = n7456 ^ n6734;
  assign n4434 = n4433 ^ n4424;
  assign n4447 = n4446 ^ n4434;
  assign n7451 = n4790 ^ n4447;
  assign n4765 = n3985 & n4063;
  assign n4632 = n3997 & n4063;
  assign n4631 = n4010 & n4072;
  assign n4633 = n4632 ^ n4631;
  assign n4766 = n4765 ^ n4633;
  assign n4763 = n4182 ^ n4070;
  assign n4695 = n4008 & n4066;
  assign n4176 = n3978 & n4048;
  assign n4655 = n4176 ^ n4052;
  assign n4696 = n4695 ^ n4655;
  assign n4764 = n4763 ^ n4696;
  assign n4767 = n4766 ^ n4764;
  assign n4814 = n4813 ^ n4767;
  assign n4780 = n4512 & n4568;
  assign n4680 = n4511 & n4568;
  assign n4679 = n4508 & n4577;
  assign n4681 = n4680 ^ n4679;
  assign n4781 = n4780 ^ n4681;
  assign n4778 = n4603 ^ n4575;
  assign n4743 = ~n4497 & n4571;
  assign n4713 = ~n4453 & n4553;
  assign n4742 = n4713 ^ n4557;
  assign n4744 = n4743 ^ n4742;
  assign n4779 = n4778 ^ n4744;
  assign n4782 = n4781 ^ n4779;
  assign n7450 = n4814 ^ n4782;
  assign n7452 = n7451 ^ n7450;
  assign n7453 = n7452 ^ n6733;
  assign n7458 = n7457 ^ n7453;
  assign n4684 = ~n4506 & n4571;
  assign n4683 = ~n4540 & n4563;
  assign n4685 = n4684 ^ n4683;
  assign n4832 = n4742 ^ n4685;
  assign n4831 = n4679 ^ n4579;
  assign n4833 = n4832 ^ n4831;
  assign n7447 = n4833 ^ n4600;
  assign n4661 = n4261 & n4282;
  assign n4662 = n4661 ^ n4304;
  assign n4664 = n4663 ^ n4662;
  assign n4660 = n4659 ^ n4315;
  assign n4665 = n4664 ^ n4660;
  assign n4666 = n4665 ^ n4321;
  assign n7448 = n7447 ^ n4666;
  assign n4635 = n4034 & n4058;
  assign n4175 = n4006 & n4066;
  assign n4636 = n4635 ^ n4175;
  assign n4656 = n4655 ^ n4636;
  assign n4654 = n4631 ^ n4074;
  assign n4657 = n4656 ^ n4654;
  assign n7446 = n6737 ^ n4657;
  assign n7449 = n7448 ^ n7446;
  assign n7459 = n7458 ^ n7449;
  assign n7460 = n7459 ^ n7443;
  assign n7462 = n7461 ^ n7460;
  assign n4668 = n4390 & n4416;
  assign n4670 = n4669 ^ n4668;
  assign n4828 = n4750 ^ n4670;
  assign n4827 = n4671 ^ n4446;
  assign n4829 = n4828 ^ n4827;
  assign n7424 = n4829 ^ n4600;
  assign n4682 = n4681 ^ n4602;
  assign n4686 = n4685 ^ n4682;
  assign n4678 = n4576 ^ n4564;
  assign n4687 = n4686 ^ n4678;
  assign n7425 = n7424 ^ n4687;
  assign n4702 = n4701 ^ n4317;
  assign n4757 = n4702 ^ n4662;
  assign n4756 = n4302 ^ n4283;
  assign n4758 = n4757 ^ n4756;
  assign n7423 = n4758 ^ n4666;
  assign n7426 = n7425 ^ n7423;
  assign n4638 = n4071 ^ n4059;
  assign n4634 = n4633 ^ n4181;
  assign n4637 = n4636 ^ n4634;
  assign n4639 = n4638 ^ n4637;
  assign n7422 = n6729 ^ n4639;
  assign n7427 = n7426 ^ n7422;
  assign n7506 = n7459 ^ n7427;
  assign n4676 = n4445 ^ n4417;
  assign n4674 = n4673 ^ n4596;
  assign n4675 = n4674 ^ n4670;
  assign n4677 = n4676 ^ n4675;
  assign n7434 = n4758 ^ n4677;
  assign n4693 = n4007 & n4048;
  assign n4694 = n4693 ^ n4061;
  assign n4697 = n4696 ^ n4694;
  assign n4692 = n4634 ^ n4074;
  assign n4698 = n4697 ^ n4692;
  assign n7435 = n7434 ^ n4698;
  assign n4704 = n4241 & n4297;
  assign n4705 = n4704 ^ n4290;
  assign n4708 = n4707 ^ n4705;
  assign n4703 = n4702 ^ n4315;
  assign n4709 = n4708 ^ n4703;
  assign n7436 = n7435 ^ n4709;
  assign n4740 = ~n4496 & n4553;
  assign n4741 = n4740 ^ n4566;
  assign n4745 = n4744 ^ n4741;
  assign n4739 = n4682 ^ n4579;
  assign n4746 = n4745 ^ n4739;
  assign n7437 = n7436 ^ n4746;
  assign n7438 = n7437 ^ n6741;
  assign n7478 = n7438 ^ n7432;
  assign n7507 = n7506 ^ n7478;
  assign n4710 = n4709 ^ n4321;
  assign n7468 = n4710 ^ n4312;
  assign n4748 = n4375 & n4427;
  assign n4749 = n4748 ^ n4424;
  assign n4753 = n4752 ^ n4749;
  assign n4747 = n4674 ^ n4446;
  assign n4754 = n4753 ^ n4747;
  assign n7466 = n4754 ^ n4600;
  assign n4714 = n4713 ^ n4684;
  assign n4715 = n4714 ^ n4556;
  assign n4712 = n4576 ^ n4566;
  assign n4716 = n4715 ^ n4712;
  assign n7467 = n7466 ^ n4716;
  assign n7469 = n7468 ^ n7467;
  assign n4177 = n4176 ^ n4175;
  assign n4178 = n4177 ^ n4051;
  assign n4174 = n4071 ^ n4061;
  assign n4179 = n4178 ^ n4174;
  assign n7464 = n6730 ^ n4179;
  assign n7465 = n7464 ^ n7427;
  assign n7470 = n7469 ^ n7465;
  assign n7476 = n7470 ^ n7461;
  assign n7508 = n7476 ^ n7449;
  assign n7509 = n7507 & n7508;
  assign n7444 = n7443 ^ n7438;
  assign n7433 = n7432 ^ n7427;
  assign n7445 = n7444 ^ n7433;
  assign n7487 = n7445 & n7476;
  assign n7510 = n7509 ^ n7487;
  assign n7480 = n7457 ^ n7438;
  assign n7504 = n7480 ^ n7476;
  assign n7463 = n7453 ^ n7438;
  assign n7494 = n7463 ^ n7461;
  assign n7495 = n7444 & n7494;
  assign n7481 = n7480 ^ n7470;
  assign n7482 = n7461 & n7481;
  assign n7496 = n7495 ^ n7482;
  assign n7505 = n7504 ^ n7496;
  assign n7511 = n7510 ^ n7505;
  assign n7477 = n7476 ^ n7458;
  assign n7490 = n7478 ^ n7477;
  assign n7488 = n7449 & n7460;
  assign n7489 = n7488 ^ n7487;
  assign n7491 = n7490 ^ n7489;
  assign n7479 = n7477 & n7478;
  assign n7483 = n7482 ^ n7479;
  assign n7492 = n7491 ^ n7483;
  assign n7520 = n7511 ^ n7492;
  assign n7498 = ~n7427 & n7459;
  assign n7471 = n7470 ^ n7463;
  assign n7474 = n7433 & n7471;
  assign n7499 = n7498 ^ n7474;
  assign n7493 = n7471 ^ n7433;
  assign n7497 = n7496 ^ n7493;
  assign n7500 = n7499 ^ n7497;
  assign n7512 = n7500 & n7511;
  assign n7472 = n7471 ^ n7459;
  assign n7485 = n7472 ^ n7462;
  assign n7473 = n7462 & n7472;
  assign n7475 = n7474 ^ n7473;
  assign n7484 = n7483 ^ n7475;
  assign n7486 = n7485 ^ n7484;
  assign n7521 = n7512 ^ n7486;
  assign n7522 = n7520 & n7521;
  assign n7523 = n7522 ^ n7492;
  assign n7970 = n7462 & n7523;
  assign n7503 = n7500 ^ n7486;
  assign n7515 = n7512 ^ n7492;
  assign n7516 = n7503 & n7515;
  assign n7517 = n7516 ^ n7486;
  assign n7513 = n7512 ^ n7503;
  assign n7501 = n7492 & n7500;
  assign n7502 = ~n7486 & n7501;
  assign n7514 = n7513 ^ n7502;
  assign n7518 = n7517 ^ n7514;
  assign n7782 = n7476 & n7518;
  assign n7548 = n7449 & n7517;
  assign n7937 = n7782 ^ n7548;
  assign n7971 = n7970 ^ n7937;
  assign n7968 = n7460 & n7517;
  assign n7542 = n7507 & n7514;
  assign n7527 = n7520 ^ n7512;
  assign n7525 = ~n7492 & n7511;
  assign n7526 = n7486 & n7525;
  assign n7528 = n7527 ^ n7526;
  assign n7541 = n7459 & n7528;
  assign n7543 = n7542 ^ n7541;
  assign n7969 = n7968 ^ n7543;
  assign n7972 = n7971 ^ n7969;
  assign n7529 = n7528 ^ n7514;
  assign n7879 = n7477 & n7529;
  assign n7534 = n7528 ^ n7523;
  assign n7878 = n7433 & n7534;
  assign n7880 = n7879 ^ n7878;
  assign n7524 = n7523 ^ n7517;
  assign n7530 = n7529 ^ n7524;
  assign n7539 = n7494 & n7530;
  assign n7881 = n7880 ^ n7539;
  assign n7535 = n7471 & n7534;
  assign n7532 = n7461 & n7524;
  assign n7531 = n7444 & n7530;
  assign n7533 = n7532 ^ n7531;
  assign n7536 = n7535 ^ n7533;
  assign n7967 = n7881 ^ n7536;
  assign n7973 = n7972 ^ n7967;
  assign n5877 = n1724 ^ n1692;
  assign n5878 = n5877 ^ n4491;
  assign n5876 = n4086 ^ n1700;
  assign n5879 = n5878 ^ n5876;
  assign n5848 = n1771 ^ n1351;
  assign n5849 = n5848 ^ n4501;
  assign n5847 = n4080 ^ n1243;
  assign n5850 = n5849 ^ n5847;
  assign n5889 = n5879 ^ n5850;
  assign n5869 = n4477 ^ n1607;
  assign n5406 = n1776 ^ n1653;
  assign n5868 = n5406 ^ n4083;
  assign n5870 = n5869 ^ n5868;
  assign n5400 = n1749 ^ n1653;
  assign n5858 = n5400 ^ n4082;
  assign n5856 = n4469 ^ n1351;
  assign n5857 = n5856 ^ n1780;
  assign n5859 = n5858 ^ n5857;
  assign n5867 = n5859 ^ n4473;
  assign n5871 = n5870 ^ n5867;
  assign n5890 = n5889 ^ n5871;
  assign n5853 = n1724 ^ n1668;
  assign n5854 = n5853 ^ n4463;
  assign n5852 = n4077 ^ n1733;
  assign n5855 = n5854 ^ n5852;
  assign n5844 = n4456 ^ n1616;
  assign n5845 = n5844 ^ n1684;
  assign n5394 = n1653 ^ n1143;
  assign n5843 = n5394 ^ n4076;
  assign n5846 = n5845 ^ n5843;
  assign n5884 = n5855 ^ n5846;
  assign n5893 = n5884 ^ n5871;
  assign n5922 = n5893 ^ n5889;
  assign n5851 = n5850 ^ n5846;
  assign n5863 = n1692 ^ n1616;
  assign n5864 = n5863 ^ n1730;
  assign n5862 = n4079 ^ n1630;
  assign n5865 = n5864 ^ n5862;
  assign n5866 = n5865 ^ n5850;
  assign n5907 = n5884 ^ n5866;
  assign n5908 = n5851 & n5907;
  assign n5891 = n5884 & n5890;
  assign n5909 = n5908 ^ n5891;
  assign n5923 = n5922 ^ n5909;
  assign n5874 = n4469 ^ n4451;
  assign n5873 = n4088 ^ n1653;
  assign n5875 = n5874 ^ n5873;
  assign n5917 = n5893 ^ n5875;
  assign n5880 = n5879 ^ n5865;
  assign n5881 = n5880 ^ n5875;
  assign n5918 = n5881 ^ n5859;
  assign n5892 = n5855 ^ n5850;
  assign n5919 = n5918 ^ n5892;
  assign n5920 = n5917 & n5919;
  assign n5860 = n5859 ^ n5855;
  assign n5861 = n5860 ^ n5851;
  assign n5900 = n5861 & n5893;
  assign n5921 = n5920 ^ n5900;
  assign n5924 = n5923 ^ n5921;
  assign n5894 = n5893 ^ n5880;
  assign n5903 = n5894 ^ n5892;
  assign n5883 = n5881 ^ n5846;
  assign n5901 = n5875 & n5883;
  assign n5902 = n5901 ^ n5900;
  assign n5904 = n5903 ^ n5902;
  assign n5895 = n5892 & n5894;
  assign n5896 = n5895 ^ n5891;
  assign n5905 = n5904 ^ n5896;
  assign n5935 = n5924 ^ n5905;
  assign n5911 = ~n5859 & n5881;
  assign n5872 = n5871 ^ n5866;
  assign n5887 = n5860 & n5872;
  assign n5912 = n5911 ^ n5887;
  assign n5906 = n5872 ^ n5860;
  assign n5910 = n5909 ^ n5906;
  assign n5913 = n5912 ^ n5910;
  assign n5925 = n5913 & n5924;
  assign n5885 = n5884 ^ n5883;
  assign n5882 = n5881 ^ n5872;
  assign n5898 = n5885 ^ n5882;
  assign n5886 = n5882 & n5885;
  assign n5888 = n5887 ^ n5886;
  assign n5897 = n5896 ^ n5888;
  assign n5899 = n5898 ^ n5897;
  assign n5939 = n5925 ^ n5899;
  assign n5940 = n5935 & n5939;
  assign n5941 = n5940 ^ n5905;
  assign n5916 = n5913 ^ n5899;
  assign n5928 = n5925 ^ n5905;
  assign n5929 = n5916 & n5928;
  assign n5930 = n5929 ^ n5899;
  assign n5942 = n5941 ^ n5930;
  assign n5955 = n5890 & n5942;
  assign n5936 = n5935 ^ n5925;
  assign n5933 = ~n5905 & n5924;
  assign n5934 = n5899 & n5933;
  assign n5937 = n5936 ^ n5934;
  assign n5926 = n5925 ^ n5916;
  assign n5914 = n5905 & n5913;
  assign n5915 = ~n5899 & n5914;
  assign n5927 = n5926 ^ n5915;
  assign n5938 = n5937 ^ n5927;
  assign n5943 = n5942 ^ n5938;
  assign n5954 = n5907 & n5943;
  assign n5956 = n5955 ^ n5954;
  assign n5952 = n5919 & n5927;
  assign n5951 = n5881 & n5937;
  assign n5953 = n5952 ^ n5951;
  assign n5957 = n5956 ^ n5953;
  assign n5947 = n5941 ^ n5937;
  assign n5948 = n5872 & n5947;
  assign n5945 = n5884 & n5942;
  assign n5944 = n5851 & n5943;
  assign n5946 = n5945 ^ n5944;
  assign n5949 = n5948 ^ n5946;
  assign n5931 = n5930 ^ n5927;
  assign n5932 = n5861 & n5931;
  assign n5950 = n5949 ^ n5932;
  assign n5958 = n5957 ^ n5950;
  assign n7300 = n5958 ^ n4590;
  assign n6066 = n4210 ^ n2376;
  assign n6067 = n6066 ^ n2154;
  assign n6068 = n6067 ^ n1741;
  assign n6062 = n2484 ^ n2452;
  assign n6063 = n6062 ^ n2587;
  assign n6064 = n6063 ^ n2498;
  assign n6065 = n6064 ^ n1790;
  assign n6069 = n6068 ^ n6065;
  assign n5273 = n2592 ^ n2537;
  assign n6059 = n5273 ^ n2503;
  assign n6058 = n4229 ^ n2423;
  assign n6060 = n6059 ^ n6058;
  assign n6056 = n2522 ^ n1229;
  assign n6053 = n2574 ^ n1256;
  assign n6051 = n4223 ^ n2451;
  assign n5267 = n2565 ^ n2537;
  assign n6050 = n5267 ^ n2431;
  assign n6052 = n6051 ^ n6050;
  assign n6054 = n6053 ^ n6052;
  assign n6057 = n6056 ^ n6054;
  assign n6061 = n6060 ^ n6057;
  assign n6070 = n6069 ^ n6061;
  assign n6091 = n2459 ^ n1754;
  assign n6089 = n2537 ^ n2434;
  assign n6090 = n6089 ^ n4223;
  assign n6092 = n6091 ^ n6090;
  assign n6078 = n4198 ^ n2141;
  assign n6079 = n6078 ^ n2517;
  assign n6080 = n6079 ^ n1718;
  assign n6081 = n6080 ^ n6068;
  assign n6093 = n6092 ^ n6081;
  assign n6126 = ~n6054 & n6093;
  assign n6047 = n2437 ^ n2340;
  assign n6048 = n6047 ^ n2534;
  assign n6046 = n2464 ^ n1660;
  assign n6049 = n6048 ^ n6046;
  assign n6055 = n6054 ^ n6049;
  assign n6086 = n6080 ^ n6065;
  assign n6087 = n6086 ^ n6061;
  assign n6088 = n6055 & n6087;
  assign n6127 = n6126 ^ n6088;
  assign n6124 = n6087 ^ n6055;
  assign n6071 = n4215 ^ n4193;
  assign n5287 = n2537 ^ n2416;
  assign n6072 = n6071 ^ n5287;
  assign n6073 = n6072 ^ n2348;
  assign n6074 = n6073 ^ n1645;
  assign n6102 = n6074 ^ n6065;
  assign n6075 = n6074 ^ n6049;
  assign n6111 = n6086 ^ n6075;
  assign n6112 = n6102 & n6111;
  assign n6076 = n6070 & n6075;
  assign n6113 = n6112 ^ n6076;
  assign n6125 = n6124 ^ n6113;
  assign n6128 = n6127 ^ n6125;
  assign n6095 = n6093 ^ n6074;
  assign n6096 = n6095 ^ n6075;
  assign n6094 = n6093 ^ n6087;
  assign n6100 = n6096 ^ n6094;
  assign n6097 = n6094 & n6096;
  assign n6098 = n6097 ^ n6088;
  assign n6077 = n6075 ^ n6061;
  assign n6082 = n6081 ^ n6077;
  assign n6083 = n6065 ^ n6049;
  assign n6084 = n6082 & n6083;
  assign n6085 = n6084 ^ n6076;
  assign n6099 = n6098 ^ n6085;
  assign n6101 = n6100 ^ n6099;
  assign n6139 = n6128 ^ n6101;
  assign n6110 = n6077 ^ n6069;
  assign n6114 = n6113 ^ n6110;
  assign n6105 = n6092 ^ n6077;
  assign n6106 = n6093 ^ n6054;
  assign n6107 = n6106 ^ n6083;
  assign n6108 = n6105 & n6107;
  assign n6103 = n6102 ^ n6055;
  assign n6104 = n6077 & n6103;
  assign n6109 = n6108 ^ n6104;
  assign n6115 = n6114 ^ n6109;
  assign n6129 = n6115 & n6128;
  assign n6118 = n6083 ^ n6082;
  assign n6116 = n6092 & n6095;
  assign n6117 = n6116 ^ n6104;
  assign n6119 = n6118 ^ n6117;
  assign n6120 = n6119 ^ n6085;
  assign n6143 = n6129 ^ n6120;
  assign n6144 = n6139 & n6143;
  assign n6145 = n6144 ^ n6101;
  assign n6123 = n6120 ^ n6115;
  assign n6132 = n6129 ^ n6101;
  assign n6133 = n6123 & n6132;
  assign n6134 = n6133 ^ n6120;
  assign n6146 = n6145 ^ n6134;
  assign n6469 = n6070 & n6146;
  assign n6140 = n6139 ^ n6129;
  assign n6137 = n6120 & n6128;
  assign n6138 = ~n6101 & n6137;
  assign n6141 = n6140 ^ n6138;
  assign n6130 = n6129 ^ n6123;
  assign n6121 = n6115 & ~n6120;
  assign n6122 = n6101 & n6121;
  assign n6131 = n6130 ^ n6122;
  assign n6142 = n6141 ^ n6131;
  assign n6147 = n6146 ^ n6142;
  assign n6468 = n6111 & n6147;
  assign n6470 = n6469 ^ n6468;
  assign n6450 = n6107 & n6141;
  assign n6449 = n6093 & n6131;
  assign n6451 = n6450 ^ n6449;
  assign n6471 = n6470 ^ n6451;
  assign n6155 = n6145 ^ n6141;
  assign n6446 = n6103 & n6155;
  assign n6135 = n6134 ^ n6131;
  assign n6151 = n6087 & n6135;
  assign n6149 = n6075 & n6146;
  assign n6148 = n6102 & n6147;
  assign n6150 = n6149 ^ n6148;
  assign n6152 = n6151 ^ n6150;
  assign n6467 = n6446 ^ n6152;
  assign n6472 = n6471 ^ n6467;
  assign n6297 = n3398 ^ n819;
  assign n6296 = n4339 ^ n894;
  assign n6298 = n6297 ^ n6296;
  assign n6294 = n3263 ^ n782;
  assign n4930 = n961 ^ n774;
  assign n6293 = n4930 ^ n742;
  assign n6295 = n6294 ^ n6293;
  assign n6299 = n6298 ^ n6295;
  assign n6290 = n3345 ^ n348;
  assign n4971 = n956 ^ n834;
  assign n6289 = n4971 ^ n4363;
  assign n6291 = n6290 ^ n6289;
  assign n6285 = n3237 ^ n749;
  assign n4958 = n940 ^ n834;
  assign n6283 = n4958 ^ n4357;
  assign n6284 = n6283 ^ n4343;
  assign n6286 = n6285 ^ n6284;
  assign n4968 = n850 ^ n795;
  assign n6288 = n6286 ^ n4968;
  assign n6292 = n6291 ^ n6288;
  assign n6300 = n6299 ^ n6292;
  assign n6320 = n3429 ^ n555;
  assign n4957 = n937 ^ n527;
  assign n6319 = n4957 ^ n835;
  assign n6321 = n6320 ^ n6319;
  assign n6309 = n3372 ^ n900;
  assign n6308 = n4328 ^ n862;
  assign n6310 = n6309 ^ n6308;
  assign n6311 = n6310 ^ n6298;
  assign n6322 = n6321 ^ n6311;
  assign n6355 = ~n6286 & ~n6322;
  assign n6281 = n2877 ^ n547;
  assign n4945 = n827 ^ n537;
  assign n6280 = n4945 ^ n929;
  assign n6282 = n6281 ^ n6280;
  assign n6287 = n6286 ^ n6282;
  assign n6316 = n6310 ^ n6295;
  assign n6317 = n6316 ^ n6292;
  assign n6318 = n6287 & n6317;
  assign n6356 = n6355 ^ n6318;
  assign n6353 = n6317 ^ n6287;
  assign n6303 = n3305 ^ n865;
  assign n4939 = n834 ^ n806;
  assign n6301 = n4939 ^ n4350;
  assign n6302 = n6301 ^ n4325;
  assign n6304 = n6303 ^ n6302;
  assign n6331 = n6304 ^ n6295;
  assign n6305 = n6304 ^ n6282;
  assign n6340 = n6316 ^ n6305;
  assign n6341 = n6331 & n6340;
  assign n6306 = n6300 & n6305;
  assign n6342 = n6341 ^ n6306;
  assign n6354 = n6353 ^ n6342;
  assign n6357 = n6356 ^ n6354;
  assign n6325 = n6322 ^ n6317;
  assign n6323 = n6322 ^ n6304;
  assign n6324 = n6323 ^ n6305;
  assign n6329 = n6325 ^ n6324;
  assign n6326 = ~n6324 & ~n6325;
  assign n6327 = n6326 ^ n6318;
  assign n6307 = n6305 ^ n6292;
  assign n6312 = n6311 ^ n6307;
  assign n6313 = n6295 ^ n6282;
  assign n6314 = n6312 & n6313;
  assign n6315 = n6314 ^ n6306;
  assign n6328 = n6327 ^ n6315;
  assign n6330 = n6329 ^ n6328;
  assign n6368 = n6357 ^ n6330;
  assign n6339 = n6307 ^ n6299;
  assign n6343 = n6342 ^ n6339;
  assign n6334 = n6322 ^ n6286;
  assign n6335 = n6334 ^ n6313;
  assign n6336 = n6321 ^ n6307;
  assign n6337 = ~n6335 & ~n6336;
  assign n6332 = n6331 ^ n6287;
  assign n6333 = n6307 & n6332;
  assign n6338 = n6337 ^ n6333;
  assign n6344 = n6343 ^ n6338;
  assign n6358 = n6344 & n6357;
  assign n6347 = n6313 ^ n6312;
  assign n6345 = ~n6321 & ~n6323;
  assign n6346 = n6345 ^ n6333;
  assign n6348 = n6347 ^ n6346;
  assign n6349 = n6348 ^ n6315;
  assign n6372 = n6358 ^ n6349;
  assign n6373 = n6368 & n6372;
  assign n6374 = n6373 ^ n6330;
  assign n6352 = n6349 ^ n6344;
  assign n6361 = n6358 ^ n6330;
  assign n6362 = n6352 & n6361;
  assign n6363 = n6362 ^ n6349;
  assign n6375 = n6374 ^ n6363;
  assign n6398 = n6300 & n6375;
  assign n6369 = n6368 ^ n6358;
  assign n6366 = n6349 & n6357;
  assign n6367 = ~n6330 & n6366;
  assign n6370 = n6369 ^ n6367;
  assign n6359 = n6358 ^ n6352;
  assign n6350 = n6344 & ~n6349;
  assign n6351 = n6330 & n6350;
  assign n6360 = n6359 ^ n6351;
  assign n6371 = n6370 ^ n6360;
  assign n6376 = n6375 ^ n6371;
  assign n6397 = n6340 & n6376;
  assign n6399 = n6398 ^ n6397;
  assign n6395 = ~n6335 & n6370;
  assign n6394 = ~n6322 & n6360;
  assign n6396 = n6395 ^ n6394;
  assign n6400 = n6399 ^ n6396;
  assign n6384 = n6374 ^ n6370;
  assign n6392 = n6332 & n6384;
  assign n6364 = n6363 ^ n6360;
  assign n6380 = n6317 & n6364;
  assign n6378 = n6305 & n6375;
  assign n6377 = n6331 & n6376;
  assign n6379 = n6378 ^ n6377;
  assign n6381 = n6380 ^ n6379;
  assign n6393 = n6392 ^ n6381;
  assign n6401 = n6400 ^ n6393;
  assign n7298 = n6472 ^ n6401;
  assign n6193 = n3226 ^ n3179;
  assign n6192 = n3355 ^ n3283;
  assign n6194 = n6193 ^ n6192;
  assign n6191 = n3531 ^ n3252;
  assign n6195 = n6194 ^ n6191;
  assign n5153 = n3380 ^ n3366;
  assign n6175 = n5153 ^ n3167;
  assign n6174 = n3539 ^ n3394;
  assign n6176 = n6175 ^ n6174;
  assign n6198 = n6195 ^ n6176;
  assign n6181 = n3325 ^ n3320;
  assign n5167 = n3276 ^ n2973;
  assign n6180 = n5167 ^ n3969;
  assign n6182 = n6181 ^ n6180;
  assign n6178 = n3521 ^ n3340;
  assign n6165 = n3524 ^ n3226;
  assign n5158 = n3435 ^ n2973;
  assign n6163 = n5158 ^ n3963;
  assign n6164 = n6163 ^ n3291;
  assign n6166 = n6165 ^ n6164;
  assign n6179 = n6178 ^ n6166;
  assign n6183 = n6182 ^ n6179;
  assign n6199 = n6198 ^ n6183;
  assign n6204 = n3963 ^ n2973;
  assign n6205 = n6204 ^ n3213;
  assign n6206 = n6205 ^ n3202;
  assign n6207 = n6206 ^ n3536;
  assign n5142 = n3313 ^ n3299;
  assign n6172 = n5142 ^ n3411;
  assign n6171 = n3528 ^ n3366;
  assign n6173 = n6172 ^ n6171;
  assign n6177 = n6176 ^ n6173;
  assign n6208 = n6207 ^ n6177;
  assign n6242 = ~n6166 & n6208;
  assign n5176 = n3404 ^ n3394;
  assign n6168 = n5176 ^ n3437;
  assign n6167 = n3549 ^ n2791;
  assign n6169 = n6168 ^ n6167;
  assign n6170 = n6169 ^ n6166;
  assign n6202 = n6195 ^ n6173;
  assign n6203 = n6202 ^ n6183;
  assign n6213 = n6170 & n6203;
  assign n6243 = n6242 ^ n6213;
  assign n6240 = n6203 ^ n6170;
  assign n6186 = n3544 ^ n3299;
  assign n5143 = n3334 ^ n2973;
  assign n6184 = n5143 ^ n3951;
  assign n6185 = n6184 ^ n3389;
  assign n6187 = n6186 ^ n6185;
  assign n6218 = n6195 ^ n6187;
  assign n6188 = n6187 ^ n6169;
  assign n6227 = n6202 ^ n6188;
  assign n6228 = n6218 & n6227;
  assign n6200 = n6188 & n6199;
  assign n6229 = n6228 ^ n6200;
  assign n6241 = n6240 ^ n6229;
  assign n6244 = n6243 ^ n6241;
  assign n6210 = n6208 ^ n6187;
  assign n6211 = n6210 ^ n6188;
  assign n6209 = n6208 ^ n6203;
  assign n6216 = n6211 ^ n6209;
  assign n6212 = n6209 & n6211;
  assign n6214 = n6213 ^ n6212;
  assign n6189 = n6188 ^ n6183;
  assign n6190 = n6189 ^ n6177;
  assign n6196 = n6195 ^ n6169;
  assign n6197 = n6190 & n6196;
  assign n6201 = n6200 ^ n6197;
  assign n6215 = n6214 ^ n6201;
  assign n6217 = n6216 ^ n6215;
  assign n6256 = n6244 ^ n6217;
  assign n6226 = n6198 ^ n6189;
  assign n6230 = n6229 ^ n6226;
  assign n6221 = n6207 ^ n6189;
  assign n6222 = n6208 ^ n6166;
  assign n6223 = n6222 ^ n6196;
  assign n6224 = n6221 & n6223;
  assign n6219 = n6218 ^ n6170;
  assign n6220 = n6189 & n6219;
  assign n6225 = n6224 ^ n6220;
  assign n6231 = n6230 ^ n6225;
  assign n6245 = n6231 & n6244;
  assign n6234 = n6196 ^ n6190;
  assign n6232 = n6207 & n6210;
  assign n6233 = n6232 ^ n6220;
  assign n6235 = n6234 ^ n6233;
  assign n6236 = n6235 ^ n6201;
  assign n6260 = n6245 ^ n6236;
  assign n6261 = n6256 & n6260;
  assign n6262 = n6261 ^ n6217;
  assign n6239 = n6236 ^ n6231;
  assign n6248 = n6245 ^ n6217;
  assign n6249 = n6239 & n6248;
  assign n6250 = n6249 ^ n6236;
  assign n6263 = n6262 ^ n6250;
  assign n6463 = n6199 & n6263;
  assign n6257 = n6256 ^ n6245;
  assign n6254 = n6236 & n6244;
  assign n6255 = ~n6217 & n6254;
  assign n6258 = n6257 ^ n6255;
  assign n6246 = n6245 ^ n6239;
  assign n6237 = n6231 & ~n6236;
  assign n6238 = n6217 & n6237;
  assign n6247 = n6246 ^ n6238;
  assign n6259 = n6258 ^ n6247;
  assign n6264 = n6263 ^ n6259;
  assign n6462 = n6227 & n6264;
  assign n6464 = n6463 ^ n6462;
  assign n6440 = n6221 & n6258;
  assign n6274 = n6262 ^ n6258;
  assign n6439 = n6219 & n6274;
  assign n6441 = n6440 ^ n6439;
  assign n6275 = n6189 & n6274;
  assign n6442 = n6441 ^ n6275;
  assign n6616 = n6464 ^ n6442;
  assign n6437 = n6223 & n6258;
  assign n6266 = n6188 & n6263;
  assign n6265 = n6218 & n6264;
  assign n6267 = n6266 ^ n6265;
  assign n6615 = n6437 ^ n6267;
  assign n6617 = n6616 ^ n6615;
  assign n6476 = n5893 & n5931;
  assign n6409 = n5917 & n5927;
  assign n6410 = n6409 ^ n5932;
  assign n6477 = n6476 ^ n6410;
  assign n6478 = n6477 ^ n5956;
  assign n6475 = n5952 ^ n5946;
  assign n6479 = n6478 ^ n6475;
  assign n7297 = n6617 ^ n6479;
  assign n7299 = n7298 ^ n7297;
  assign n7301 = n7300 ^ n7299;
  assign n6567 = n6477 ^ n5953;
  assign n6568 = n6567 ^ n5949;
  assign n7288 = n6568 ^ n4169;
  assign n6445 = n6105 & n6141;
  assign n6447 = n6446 ^ n6445;
  assign n6156 = n6077 & n6155;
  assign n6448 = n6447 ^ n6156;
  assign n6452 = n6451 ^ n6448;
  assign n6453 = n6452 ^ n6152;
  assign n6427 = ~n6336 & n6370;
  assign n6428 = n6427 ^ n6392;
  assign n6385 = n6307 & n6384;
  assign n6432 = n6428 ^ n6385;
  assign n6433 = n6432 ^ n6396;
  assign n6434 = n6433 ^ n6381;
  assign n7286 = n6453 ^ n6434;
  assign n6273 = n6207 & n6262;
  assign n6271 = n6209 & n6250;
  assign n6533 = n6273 ^ n6271;
  assign n6534 = n6533 ^ n6441;
  assign n6436 = n6208 & n6247;
  assign n6438 = n6437 ^ n6436;
  assign n6532 = n6438 ^ n6267;
  assign n6535 = n6534 ^ n6532;
  assign n6465 = n6464 ^ n6438;
  assign n6251 = n6250 ^ n6247;
  assign n6253 = n6203 & n6251;
  assign n6268 = n6267 ^ n6253;
  assign n6461 = n6439 ^ n6268;
  assign n6466 = n6465 ^ n6461;
  assign n7284 = n6535 ^ n6466;
  assign n6407 = n5875 & n5930;
  assign n6406 = n5882 & n5941;
  assign n6408 = n6407 ^ n6406;
  assign n6411 = n6410 ^ n6408;
  assign n6405 = n5953 ^ n5946;
  assign n6412 = n6411 ^ n6405;
  assign n6413 = n6412 ^ n5958;
  assign n7285 = n7284 ^ n6413;
  assign n7287 = n7286 ^ n7285;
  assign n7289 = n7288 ^ n7287;
  assign n7319 = n7301 ^ n7289;
  assign n6159 = n6094 & n6134;
  assign n6154 = n6092 & n6145;
  assign n6529 = n6159 ^ n6154;
  assign n6530 = n6529 ^ n6447;
  assign n6528 = n6451 ^ n6150;
  assign n6531 = n6530 ^ n6528;
  assign n6388 = ~n6325 & n6363;
  assign n6383 = ~n6321 & n6374;
  assign n6426 = n6388 ^ n6383;
  assign n6429 = n6428 ^ n6426;
  assign n6425 = n6396 ^ n6379;
  assign n6430 = n6429 ^ n6425;
  assign n7314 = n6531 ^ n6430;
  assign n6630 = n6210 & n6262;
  assign n6631 = n6630 ^ n6438;
  assign n6585 = n6211 & n6250;
  assign n6276 = n6275 ^ n6273;
  assign n6586 = n6585 ^ n6276;
  assign n6632 = n6631 ^ n6586;
  assign n6513 = n6190 & n6259;
  assign n6252 = n6170 & n6251;
  assign n6514 = n6513 ^ n6252;
  assign n6515 = n6514 ^ n6462;
  assign n6629 = n6515 ^ n6268;
  assign n6633 = n6632 ^ n6629;
  assign n7312 = n6633 ^ n6466;
  assign n6544 = n5883 & n5930;
  assign n6545 = n6544 ^ n5953;
  assign n6542 = n5885 & n5941;
  assign n6494 = n6476 ^ n6407;
  assign n6543 = n6542 ^ n6494;
  assign n6546 = n6545 ^ n6543;
  assign n6538 = n5894 & n5938;
  assign n6490 = n5860 & n5947;
  assign n6539 = n6538 ^ n6490;
  assign n6540 = n6539 ^ n5954;
  assign n6541 = n6540 ^ n5949;
  assign n6547 = n6546 ^ n6541;
  assign n6548 = n6547 ^ n5958;
  assign n7313 = n7312 ^ n6548;
  assign n7315 = n7314 ^ n7313;
  assign n7310 = n6412 ^ n4626;
  assign n6492 = n5918 & n5937;
  assign n6493 = n6492 ^ n6406;
  assign n6637 = n6540 ^ n6493;
  assign n6636 = n5951 ^ n5946;
  assign n6638 = n6637 ^ n6636;
  assign n7295 = n6638 ^ n4649;
  assign n6523 = n6449 ^ n6150;
  assign n6519 = n6082 & n6142;
  assign n6136 = n6055 & n6135;
  assign n6520 = n6519 ^ n6136;
  assign n6521 = n6520 ^ n6468;
  assign n6158 = n6106 & n6131;
  assign n6160 = n6159 ^ n6158;
  assign n6522 = n6521 ^ n6160;
  assign n6524 = n6523 ^ n6522;
  assign n6507 = n6312 & n6371;
  assign n6365 = n6287 & n6364;
  assign n6508 = n6507 ^ n6365;
  assign n6509 = n6508 ^ n6397;
  assign n6387 = ~n6334 & n6360;
  assign n6389 = n6388 ^ n6387;
  assign n6510 = n6509 ^ n6389;
  assign n6506 = n6394 ^ n6379;
  assign n6511 = n6510 ^ n6506;
  assign n7293 = n6524 ^ n6511;
  assign n6270 = n6222 & n6247;
  assign n6272 = n6271 ^ n6270;
  assign n6277 = n6276 ^ n6272;
  assign n6269 = n6268 ^ n6252;
  assign n6278 = n6277 ^ n6269;
  assign n7291 = n6466 ^ n6278;
  assign n6495 = n6494 ^ n6493;
  assign n6491 = n6490 ^ n5949;
  assign n6496 = n6495 ^ n6491;
  assign n6497 = n6496 ^ n5958;
  assign n7292 = n7291 ^ n6497;
  assign n7294 = n7293 ^ n7292;
  assign n7296 = n7295 ^ n7294;
  assign n7311 = n7310 ^ n7296;
  assign n7316 = n7315 ^ n7311;
  assign n7348 = n7319 ^ n7316;
  assign n7325 = n6479 ^ n4797;
  assign n6613 = n6470 ^ n6448;
  assign n6612 = n6450 ^ n6150;
  assign n6614 = n6613 ^ n6612;
  assign n6458 = n6432 ^ n6399;
  assign n6457 = n6395 ^ n6379;
  assign n6459 = n6458 ^ n6457;
  assign n7323 = n6614 ^ n6459;
  assign n6603 = n5892 & n5938;
  assign n6604 = n6603 ^ n6539;
  assign n6601 = n5955 ^ n5945;
  assign n6602 = n6601 ^ n6543;
  assign n6605 = n6604 ^ n6602;
  assign n6588 = n6196 & n6259;
  assign n6589 = n6588 ^ n6514;
  assign n6584 = n6463 ^ n6266;
  assign n6587 = n6586 ^ n6584;
  assign n6590 = n6589 ^ n6587;
  assign n7322 = n6605 ^ n6590;
  assign n7324 = n7323 ^ n7322;
  assign n7326 = n7325 ^ n7324;
  assign n7307 = n6605 ^ n4773;
  assign n6595 = n6083 & n6142;
  assign n6596 = n6595 ^ n6520;
  assign n6593 = n6469 ^ n6149;
  assign n6591 = n6096 & n6134;
  assign n6157 = n6156 ^ n6154;
  assign n6592 = n6591 ^ n6157;
  assign n6594 = n6593 ^ n6592;
  assign n6597 = n6596 ^ n6594;
  assign n6580 = n6313 & n6371;
  assign n6581 = n6580 ^ n6508;
  assign n6578 = n6398 ^ n6378;
  assign n6558 = ~n6324 & n6363;
  assign n6386 = n6385 ^ n6383;
  assign n6559 = n6558 ^ n6386;
  assign n6579 = n6578 ^ n6559;
  assign n6582 = n6581 ^ n6579;
  assign n7305 = n6597 ^ n6582;
  assign n6443 = n6442 ^ n6438;
  assign n6444 = n6443 ^ n6268;
  assign n7304 = n6568 ^ n6444;
  assign n7306 = n7305 ^ n7304;
  assign n7308 = n7307 ^ n7306;
  assign n7337 = n7326 ^ n7308;
  assign n7349 = n7348 ^ n7337;
  assign n7335 = n6496 ^ n4838;
  assign n6390 = n6389 ^ n6386;
  assign n6382 = n6381 ^ n6365;
  assign n6391 = n6390 ^ n6382;
  assign n6161 = n6160 ^ n6157;
  assign n6153 = n6152 ^ n6136;
  assign n6162 = n6161 ^ n6153;
  assign n7333 = n6391 ^ n6162;
  assign n7332 = n6466 ^ n5958;
  assign n7334 = n7333 ^ n7332;
  assign n7336 = n7335 ^ n7334;
  assign n7338 = n7337 ^ n7336;
  assign n6625 = n6095 & n6145;
  assign n6626 = n6625 ^ n6451;
  assign n6627 = n6626 ^ n6592;
  assign n6624 = n6521 ^ n6152;
  assign n6628 = n6627 ^ n6624;
  assign n6556 = ~n6323 & n6374;
  assign n6557 = n6556 ^ n6396;
  assign n6560 = n6559 ^ n6557;
  assign n6555 = n6509 ^ n6381;
  assign n6561 = n6560 ^ n6555;
  assign n7281 = n6628 ^ n6561;
  assign n6517 = n6436 ^ n6267;
  assign n6516 = n6515 ^ n6272;
  assign n6518 = n6517 ^ n6516;
  assign n7280 = n6638 ^ n6518;
  assign n7282 = n7281 ^ n7280;
  assign n7279 = n6547 ^ n4734;
  assign n7283 = n7282 ^ n7279;
  assign n7309 = n7308 ^ n7283;
  assign n7317 = n7316 ^ n7309;
  assign n7345 = n7338 ^ n7317;
  assign n7343 = n7338 ^ n7289;
  assign n7344 = n7343 ^ n7319;
  assign n7354 = n7345 ^ n7344;
  assign n7350 = n7301 ^ n7283;
  assign n7351 = ~n7349 & n7350;
  assign n7327 = n7326 ^ n7283;
  assign n7328 = n7327 ^ n7316;
  assign n7329 = n7319 & n7328;
  assign n7352 = n7351 ^ n7329;
  assign n7346 = ~n7344 & ~n7345;
  assign n7302 = n7301 ^ n7296;
  assign n7340 = ~n7302 & n7317;
  assign n7347 = n7346 ^ n7340;
  assign n7353 = n7352 ^ n7347;
  assign n7355 = n7354 ^ n7353;
  assign n7363 = n7348 ^ n7327;
  assign n7290 = n7289 ^ n7283;
  assign n7320 = n7319 ^ n7309;
  assign n7321 = n7290 & ~n7320;
  assign n7330 = n7329 ^ n7321;
  assign n7364 = n7363 ^ n7330;
  assign n7303 = n7302 ^ n7290;
  assign n7361 = ~n7303 & ~n7348;
  assign n7357 = n7338 ^ n7296;
  assign n7358 = n7357 ^ n7350;
  assign n7359 = n7348 ^ n7336;
  assign n7360 = n7358 & n7359;
  assign n7362 = n7361 ^ n7360;
  assign n7365 = n7364 ^ n7362;
  assign n7369 = n7350 ^ n7349;
  assign n7367 = ~n7336 & ~n7343;
  assign n7368 = n7367 ^ n7361;
  assign n7370 = n7369 ^ n7368;
  assign n7371 = n7370 ^ n7352;
  assign n7387 = n7365 & n7371;
  assign n7388 = n7355 & n7387;
  assign n7385 = n7371 ^ n7365;
  assign n7339 = n7296 & ~n7338;
  assign n7341 = n7340 ^ n7339;
  assign n7318 = n7317 ^ n7302;
  assign n7331 = n7330 ^ n7318;
  assign n7342 = n7341 ^ n7331;
  assign n7366 = ~n7342 & n7365;
  assign n7386 = n7385 ^ n7366;
  assign n7389 = n7388 ^ n7386;
  assign n7356 = n7355 ^ n7342;
  assign n7377 = n7366 ^ n7356;
  assign n7375 = ~n7342 & ~n7371;
  assign n7376 = ~n7355 & n7375;
  assign n7378 = n7377 ^ n7376;
  assign n7399 = n7389 ^ n7378;
  assign n7832 = ~n7349 & n7399;
  assign n7394 = n7366 ^ n7355;
  assign n7395 = ~n7385 & n7394;
  assign n7396 = n7395 ^ n7371;
  assign n7403 = n7396 ^ n7389;
  assign n7831 = ~n7302 & n7403;
  assign n7833 = n7832 ^ n7831;
  assign n7372 = n7371 ^ n7366;
  assign n7373 = ~n7356 & ~n7372;
  assign n7374 = n7373 ^ n7355;
  assign n7397 = n7396 ^ n7374;
  assign n7400 = n7399 ^ n7397;
  assign n7410 = ~n7320 & ~n7400;
  assign n7872 = n7833 ^ n7410;
  assign n7404 = n7317 & n7403;
  assign n7401 = n7290 & ~n7400;
  assign n7398 = n7319 & ~n7397;
  assign n7402 = n7401 ^ n7398;
  assign n7405 = n7404 ^ n7402;
  assign n7896 = n7872 ^ n7405;
  assign n7893 = ~n7343 & n7374;
  assign n7391 = n7358 & ~n7378;
  assign n7390 = ~n7338 & ~n7389;
  assign n7392 = n7391 ^ n7390;
  assign n7894 = n7893 ^ n7392;
  assign n7827 = ~n7344 & ~n7396;
  assign n7415 = ~n7336 & n7374;
  assign n7379 = n7378 ^ n7374;
  assign n7383 = ~n7348 & ~n7379;
  assign n7826 = n7415 ^ n7383;
  assign n7828 = n7827 ^ n7826;
  assign n7895 = n7894 ^ n7828;
  assign n7897 = n7896 ^ n7895;
  assign n11690 = n7973 ^ n7897;
  assign n12665 = n12664 ^ n11690;
  assign n4959 = n4958 ^ n4957;
  assign n4956 = n2557 ^ n547;
  assign n4960 = n4959 ^ n4956;
  assign n4953 = n2047 ^ n900;
  assign n4951 = n928 ^ n885;
  assign n4952 = n4951 ^ n4339;
  assign n4954 = n4953 ^ n4952;
  assign n4936 = n2405 ^ n865;
  assign n4934 = n885 ^ n857;
  assign n4935 = n4934 ^ n4328;
  assign n4937 = n4936 ^ n4935;
  assign n4955 = n4954 ^ n4937;
  assign n4961 = n4960 ^ n4955;
  assign n4965 = n4958 ^ n741;
  assign n4966 = n4965 ^ n4343;
  assign n4964 = n2474 ^ n556;
  assign n4967 = n4966 ^ n4964;
  assign n5012 = n4967 ^ n4961;
  assign n4947 = n2547 ^ n819;
  assign n4944 = n928 ^ n834;
  assign n4946 = n4945 ^ n4944;
  assign n4948 = n4947 ^ n4946;
  assign n4932 = n2580 ^ n749;
  assign n4929 = n956 ^ n741;
  assign n4931 = n4930 ^ n4929;
  assign n4933 = n4932 ^ n4931;
  assign n4981 = n4948 ^ n4933;
  assign n5013 = n5012 ^ n4981;
  assign n4972 = n4971 ^ n806;
  assign n4970 = n2491 ^ n783;
  assign n4973 = n4972 ^ n4970;
  assign n4969 = n4968 ^ n4967;
  assign n4974 = n4973 ^ n4969;
  assign n4942 = n2528 ^ n852;
  assign n4940 = n4939 ^ n857;
  assign n4941 = n4940 ^ n4325;
  assign n4943 = n4942 ^ n4941;
  assign n4949 = n4948 ^ n4943;
  assign n4982 = n4974 ^ n4949;
  assign n5014 = n4982 ^ n4960;
  assign n5015 = n5013 & n5014;
  assign n4993 = n4943 ^ n4933;
  assign n4978 = n4967 ^ n4948;
  assign n4994 = n4993 ^ n4978;
  assign n4995 = n4982 & n4994;
  assign n5016 = n5015 ^ n4995;
  assign n4985 = n4954 ^ n4933;
  assign n5010 = n4985 ^ n4982;
  assign n4938 = n4937 ^ n4933;
  assign n4950 = n4949 ^ n4938;
  assign n5001 = n4950 & n4993;
  assign n4986 = n4985 ^ n4974;
  assign n4987 = n4949 & n4986;
  assign n5002 = n5001 ^ n4987;
  assign n5011 = n5010 ^ n5002;
  assign n5017 = n5016 ^ n5011;
  assign n4983 = n4982 ^ n4955;
  assign n4997 = n4983 ^ n4981;
  assign n4962 = n4961 ^ n4943;
  assign n4992 = n4960 & n4962;
  assign n4996 = n4995 ^ n4992;
  assign n4998 = n4997 ^ n4996;
  assign n4984 = n4981 & n4983;
  assign n4988 = n4987 ^ n4984;
  assign n4999 = n4998 ^ n4988;
  assign n5023 = n5017 ^ n4999;
  assign n5004 = n4961 & ~n4967;
  assign n4975 = n4974 ^ n4938;
  assign n4979 = n4975 & n4978;
  assign n5005 = n5004 ^ n4979;
  assign n5000 = n4978 ^ n4975;
  assign n5003 = n5002 ^ n5000;
  assign n5006 = n5005 ^ n5003;
  assign n5018 = n5006 & n5017;
  assign n5024 = n5023 ^ n5018;
  assign n4976 = n4975 ^ n4961;
  assign n4963 = n4962 ^ n4949;
  assign n4990 = n4976 ^ n4963;
  assign n4977 = n4963 & n4976;
  assign n4980 = n4979 ^ n4977;
  assign n4989 = n4988 ^ n4980;
  assign n4991 = n4990 ^ n4989;
  assign n5021 = ~n4999 & n5017;
  assign n5022 = n4991 & n5021;
  assign n5025 = n5024 ^ n5022;
  assign n5625 = n4961 & n5025;
  assign n5009 = n5006 ^ n4991;
  assign n5019 = n5018 ^ n5009;
  assign n5007 = n4999 & n5006;
  assign n5008 = ~n4991 & n5007;
  assign n5020 = n5019 ^ n5008;
  assign n5048 = n5013 & n5020;
  assign n5626 = n5625 ^ n5048;
  assign n5041 = n5014 & n5020;
  assign n5030 = n5018 ^ n4999;
  assign n5031 = n5009 & n5030;
  assign n5032 = n5031 ^ n4991;
  assign n5038 = n5032 ^ n5020;
  assign n5040 = n4994 & n5038;
  assign n5042 = n5041 ^ n5040;
  assign n5039 = n4982 & n5038;
  assign n5043 = n5042 ^ n5039;
  assign n5704 = n5626 ^ n5043;
  assign n5027 = n5018 ^ n4991;
  assign n5028 = n5023 & n5027;
  assign n5029 = n5028 ^ n4999;
  assign n5516 = n5029 ^ n5025;
  assign n5576 = n4975 & n5516;
  assign n5033 = n5032 ^ n5029;
  assign n5046 = n4949 & n5033;
  assign n5026 = n5025 ^ n5020;
  assign n5034 = n5033 ^ n5026;
  assign n5045 = n4993 & n5034;
  assign n5047 = n5046 ^ n5045;
  assign n5577 = n5576 ^ n5047;
  assign n5705 = n5704 ^ n5577;
  assign n7190 = n7189 ^ n5705;
  assign n5290 = n3306 ^ n2391;
  assign n5288 = n5287 ^ n2507;
  assign n5289 = n5288 ^ n2517;
  assign n5291 = n5290 ^ n5289;
  assign n5264 = n4222 ^ n2593;
  assign n5263 = n3264 ^ n2484;
  assign n5265 = n5264 ^ n5263;
  assign n5300 = n5291 ^ n5265;
  assign n5283 = n3373 ^ n1962;
  assign n5282 = n4214 ^ n2376;
  assign n5284 = n5283 ^ n5282;
  assign n5318 = n5284 ^ n5265;
  assign n5295 = n4197 ^ n2538;
  assign n5294 = n2878 ^ n2464;
  assign n5296 = n5295 ^ n5294;
  assign n5297 = n5296 ^ n5291;
  assign n5319 = n5318 ^ n5297;
  assign n5320 = n5300 & n5319;
  assign n5275 = n3346 ^ n2522;
  assign n5274 = n5273 ^ n2499;
  assign n5276 = n5275 ^ n5274;
  assign n5270 = n3238 ^ n2574;
  assign n5268 = n5267 ^ n2438;
  assign n5269 = n5268 ^ n2452;
  assign n5271 = n5270 ^ n5269;
  assign n5272 = n5271 ^ n2424;
  assign n5277 = n5276 ^ n5272;
  assign n5261 = n4192 ^ n2340;
  assign n5260 = n3399 ^ n2543;
  assign n5262 = n5261 ^ n5260;
  assign n5266 = n5265 ^ n5262;
  assign n5278 = n5277 ^ n5266;
  assign n5309 = n5278 & n5297;
  assign n5321 = n5320 ^ n5309;
  assign n5298 = n5297 ^ n5277;
  assign n5317 = n5298 ^ n5266;
  assign n5322 = n5321 ^ n5317;
  assign n5285 = n5284 ^ n5262;
  assign n5280 = n3430 ^ n2459;
  assign n5279 = n4209 ^ n2566;
  assign n5281 = n5280 ^ n5279;
  assign n5286 = n5285 ^ n5281;
  assign n5312 = n5286 ^ n5271;
  assign n5305 = n5296 ^ n5265;
  assign n5313 = n5312 ^ n5305;
  assign n5314 = n5298 ^ n5281;
  assign n5315 = ~n5313 & ~n5314;
  assign n5299 = n5296 ^ n5271;
  assign n5301 = n5300 ^ n5299;
  assign n5302 = n5298 & n5301;
  assign n5316 = n5315 ^ n5302;
  assign n5323 = n5322 ^ n5316;
  assign n5336 = ~n5271 & ~n5286;
  assign n5326 = n5318 ^ n5277;
  assign n5329 = n5299 & n5326;
  assign n5337 = n5336 ^ n5329;
  assign n5334 = n5326 ^ n5299;
  assign n5335 = n5334 ^ n5321;
  assign n5338 = n5337 ^ n5335;
  assign n5339 = n5323 & n5338;
  assign n5304 = n5298 ^ n5285;
  assign n5308 = n5304 & n5305;
  assign n5310 = n5309 ^ n5308;
  assign n5306 = n5305 ^ n5304;
  assign n5292 = n5291 ^ n5286;
  assign n5293 = ~n5281 & ~n5292;
  assign n5303 = n5302 ^ n5293;
  assign n5307 = n5306 ^ n5303;
  assign n5311 = n5310 ^ n5307;
  assign n5324 = n5323 ^ n5311;
  assign n5364 = n5339 ^ n5324;
  assign n5327 = n5326 ^ n5286;
  assign n5325 = n5297 ^ n5292;
  assign n5332 = n5327 ^ n5325;
  assign n5328 = ~n5325 & ~n5327;
  assign n5330 = n5329 ^ n5328;
  assign n5331 = n5330 ^ n5310;
  assign n5333 = n5332 ^ n5331;
  assign n5362 = ~n5311 & n5323;
  assign n5363 = n5333 & n5362;
  assign n5365 = n5364 ^ n5363;
  assign n5343 = n5338 ^ n5333;
  assign n5354 = n5343 ^ n5339;
  assign n5352 = n5311 & n5338;
  assign n5353 = ~n5333 & n5352;
  assign n5355 = n5354 ^ n5353;
  assign n5366 = n5365 ^ n5355;
  assign n5344 = n5339 ^ n5311;
  assign n5345 = n5343 & n5344;
  assign n5346 = n5345 ^ n5333;
  assign n5340 = n5339 ^ n5333;
  assign n5341 = n5324 & n5340;
  assign n5342 = n5341 ^ n5311;
  assign n5347 = n5346 ^ n5342;
  assign n5553 = n5366 ^ n5347;
  assign n5554 = n5300 & n5553;
  assign n5349 = n5297 & n5347;
  assign n5555 = n5554 ^ n5349;
  assign n5368 = n5365 ^ n5342;
  assign n5552 = n5326 & n5368;
  assign n5556 = n5555 ^ n5552;
  assign n5548 = ~n5314 & n5355;
  assign n5356 = n5355 ^ n5346;
  assign n5547 = n5301 & n5356;
  assign n5549 = n5548 ^ n5547;
  assign n5357 = n5298 & n5356;
  assign n5550 = n5549 ^ n5357;
  assign n5545 = ~n5313 & n5355;
  assign n5544 = ~n5286 & n5365;
  assign n5546 = n5545 ^ n5544;
  assign n5551 = n5550 ^ n5546;
  assign n5557 = n5556 ^ n5551;
  assign n5370 = n5304 & n5366;
  assign n5369 = n5299 & n5368;
  assign n5371 = n5370 ^ n5369;
  assign n5367 = n5305 & n5366;
  assign n5372 = n5371 ^ n5367;
  assign n5359 = ~n5325 & n5342;
  assign n5351 = ~n5281 & n5346;
  assign n5358 = n5357 ^ n5351;
  assign n5360 = n5359 ^ n5358;
  assign n5348 = n5278 & n5347;
  assign n5350 = n5349 ^ n5348;
  assign n5361 = n5360 ^ n5350;
  assign n5373 = n5372 ^ n5361;
  assign n7187 = n5557 ^ n5373;
  assign n5420 = n4490 ^ n1634;
  assign n5419 = n3529 ^ n1700;
  assign n5421 = n5420 ^ n5419;
  assign n5417 = n4462 ^ n1706;
  assign n5416 = n3540 ^ n1733;
  assign n5418 = n5417 ^ n5416;
  assign n5422 = n5421 ^ n5418;
  assign n5412 = n4450 ^ n1734;
  assign n5411 = n3550 ^ n1653;
  assign n5413 = n5412 ^ n5411;
  assign n5395 = n5394 ^ n1624;
  assign n5396 = n5395 ^ n4485;
  assign n5393 = n3545 ^ n1630;
  assign n5397 = n5396 ^ n5393;
  assign n5414 = n5413 ^ n5397;
  assign n5408 = n1622 ^ n1607;
  assign n5407 = n5406 ^ n1578;
  assign n5409 = n5408 ^ n5407;
  assign n5404 = n3522 ^ n1143;
  assign n5401 = n5400 ^ n1566;
  assign n5402 = n5401 ^ n4500;
  assign n5399 = n3525 ^ n1243;
  assign n5403 = n5402 ^ n5399;
  assign n5405 = n5404 ^ n5403;
  assign n5410 = n5409 ^ n5405;
  assign n5415 = n5414 ^ n5410;
  assign n5423 = n5422 ^ n5415;
  assign n5432 = n5400 ^ n1565;
  assign n5433 = n5432 ^ n1444;
  assign n5434 = n5433 ^ n1760;
  assign n5435 = n5434 ^ n3537;
  assign n5436 = n5435 ^ n5422;
  assign n5452 = ~n5403 & n5436;
  assign n5390 = n1548 ^ n1243;
  assign n5389 = n1771 ^ n1595;
  assign n5391 = n5390 ^ n5389;
  assign n5388 = n3532 ^ n1776;
  assign n5392 = n5391 ^ n5388;
  assign n5430 = n5421 ^ n5392;
  assign n5431 = n5430 ^ n5410;
  assign n5441 = n5413 ^ n5403;
  assign n5442 = n5431 & n5441;
  assign n5453 = n5452 ^ n5442;
  assign n5450 = n5441 ^ n5431;
  assign n5398 = n5397 ^ n5392;
  assign n5447 = n5430 ^ n5414;
  assign n5448 = n5398 & n5447;
  assign n5426 = n5418 ^ n5392;
  assign n5427 = n5426 ^ n5410;
  assign n5428 = n5414 & n5427;
  assign n5449 = n5448 ^ n5428;
  assign n5451 = n5450 ^ n5449;
  assign n5454 = n5453 ^ n5451;
  assign n5468 = n5426 ^ n5415;
  assign n5469 = n5468 ^ n5449;
  assign n5463 = n5435 ^ n5415;
  assign n5464 = n5436 ^ n5403;
  assign n5424 = n5413 ^ n5392;
  assign n5465 = n5464 ^ n5424;
  assign n5466 = n5463 & n5465;
  assign n5457 = n5441 ^ n5398;
  assign n5458 = n5415 & n5457;
  assign n5467 = n5466 ^ n5458;
  assign n5470 = n5469 ^ n5467;
  assign n5471 = n5454 & n5470;
  assign n5438 = n5436 ^ n5397;
  assign n5439 = n5438 ^ n5414;
  assign n5437 = n5436 ^ n5431;
  assign n5445 = n5439 ^ n5437;
  assign n5440 = n5437 & n5439;
  assign n5443 = n5442 ^ n5440;
  assign n5425 = n5423 & n5424;
  assign n5429 = n5428 ^ n5425;
  assign n5444 = n5443 ^ n5429;
  assign n5446 = n5445 ^ n5444;
  assign n5455 = n5454 ^ n5446;
  assign n5486 = n5471 ^ n5455;
  assign n5460 = n5424 ^ n5423;
  assign n5456 = n5435 & n5438;
  assign n5459 = n5458 ^ n5456;
  assign n5461 = n5460 ^ n5459;
  assign n5462 = n5461 ^ n5429;
  assign n5484 = n5454 & n5462;
  assign n5485 = ~n5446 & n5484;
  assign n5487 = n5486 ^ n5485;
  assign n5475 = n5470 ^ n5462;
  assign n5482 = n5475 ^ n5471;
  assign n5480 = ~n5462 & n5470;
  assign n5481 = n5446 & n5480;
  assign n5483 = n5482 ^ n5481;
  assign n5488 = n5487 ^ n5483;
  assign n5568 = n5423 & n5488;
  assign n5476 = n5471 ^ n5446;
  assign n5477 = n5475 & n5476;
  assign n5478 = n5477 ^ n5462;
  assign n5566 = n5483 ^ n5478;
  assign n5567 = n5441 & n5566;
  assign n5569 = n5568 ^ n5567;
  assign n5565 = n5424 & n5488;
  assign n5570 = n5569 ^ n5565;
  assign n5562 = n5439 & n5478;
  assign n5472 = n5471 ^ n5462;
  assign n5473 = n5455 & n5472;
  assign n5474 = n5473 ^ n5446;
  assign n5560 = n5435 & n5474;
  assign n5496 = n5487 ^ n5474;
  assign n5499 = n5415 & n5496;
  assign n5561 = n5560 ^ n5499;
  assign n5563 = n5562 ^ n5561;
  assign n5479 = n5478 ^ n5474;
  assign n5502 = n5427 & n5479;
  assign n5491 = n5414 & n5479;
  assign n5559 = n5502 ^ n5491;
  assign n5564 = n5563 ^ n5559;
  assign n5571 = n5570 ^ n5564;
  assign n5168 = n5167 ^ n3334;
  assign n5166 = n3357 ^ n3320;
  assign n5169 = n5168 ^ n5166;
  assign n5164 = n3340 ^ n1230;
  assign n5162 = n3226 ^ n1257;
  assign n5160 = n3290 ^ n3214;
  assign n5159 = n5158 ^ n3179;
  assign n5161 = n5160 ^ n5159;
  assign n5163 = n5162 ^ n5161;
  assign n5165 = n5164 ^ n5163;
  assign n5170 = n5169 ^ n5165;
  assign n5144 = n5143 ^ n5142;
  assign n5145 = n5144 ^ n3326;
  assign n5146 = n5145 ^ n3388;
  assign n5147 = n5146 ^ n1646;
  assign n5138 = n3405 ^ n1661;
  assign n5139 = n5138 ^ n2973;
  assign n5140 = n5139 ^ n3207;
  assign n5141 = n5140 ^ n2791;
  assign n5148 = n5147 ^ n5141;
  assign n5189 = n5170 ^ n5148;
  assign n5177 = n5176 ^ n3386;
  assign n5178 = n5177 ^ n3159;
  assign n5179 = n5178 ^ n1742;
  assign n5154 = n5153 ^ n3410;
  assign n5155 = n5154 ^ n3316;
  assign n5156 = n5155 ^ n1719;
  assign n5180 = n5179 ^ n5156;
  assign n5190 = n5189 ^ n5180;
  assign n5173 = n3202 ^ n3066;
  assign n5174 = n5173 ^ n5158;
  assign n5172 = n3425 ^ n1755;
  assign n5175 = n5174 ^ n5172;
  assign n5181 = n5180 ^ n5175;
  assign n5219 = n5181 ^ n5163;
  assign n5149 = n3252 ^ n3190;
  assign n5150 = n5149 ^ n3276;
  assign n5151 = n5150 ^ n3355;
  assign n5152 = n5151 ^ n1791;
  assign n5191 = n5152 ^ n5141;
  assign n5220 = n5219 ^ n5191;
  assign n5221 = n5189 ^ n5175;
  assign n5222 = n5220 & n5221;
  assign n5201 = n5152 ^ n5147;
  assign n5186 = n5163 ^ n5141;
  assign n5211 = n5201 ^ n5186;
  assign n5212 = n5189 & n5211;
  assign n5223 = n5222 ^ n5212;
  assign n5193 = n5179 ^ n5152;
  assign n5217 = n5193 ^ n5189;
  assign n5157 = n5156 ^ n5152;
  assign n5202 = n5157 ^ n5148;
  assign n5203 = n5201 & n5202;
  assign n5194 = n5193 ^ n5170;
  assign n5195 = n5148 & n5194;
  assign n5204 = n5203 ^ n5195;
  assign n5218 = n5217 ^ n5204;
  assign n5224 = n5223 ^ n5218;
  assign n5214 = n5191 ^ n5190;
  assign n5183 = n5181 ^ n5147;
  assign n5210 = n5175 & n5183;
  assign n5213 = n5212 ^ n5210;
  assign n5215 = n5214 ^ n5213;
  assign n5192 = n5190 & n5191;
  assign n5196 = n5195 ^ n5192;
  assign n5216 = n5215 ^ n5196;
  assign n5229 = n5224 ^ n5216;
  assign n5206 = ~n5163 & n5181;
  assign n5171 = n5170 ^ n5157;
  assign n5187 = n5171 & n5186;
  assign n5207 = n5206 ^ n5187;
  assign n5200 = n5186 ^ n5171;
  assign n5205 = n5204 ^ n5200;
  assign n5208 = n5207 ^ n5205;
  assign n5225 = n5208 & n5224;
  assign n5250 = n5229 ^ n5225;
  assign n5184 = n5183 ^ n5148;
  assign n5182 = n5181 ^ n5171;
  assign n5198 = n5184 ^ n5182;
  assign n5185 = n5182 & n5184;
  assign n5188 = n5187 ^ n5185;
  assign n5197 = n5196 ^ n5188;
  assign n5199 = n5198 ^ n5197;
  assign n5248 = ~n5216 & n5224;
  assign n5249 = n5199 & n5248;
  assign n5251 = n5250 ^ n5249;
  assign n5209 = n5208 ^ n5199;
  assign n5239 = n5225 ^ n5209;
  assign n5237 = n5208 & n5216;
  assign n5238 = ~n5199 & n5237;
  assign n5240 = n5239 ^ n5238;
  assign n5252 = n5251 ^ n5240;
  assign n5256 = n5190 & n5252;
  assign n5230 = n5225 ^ n5199;
  assign n5231 = n5229 & n5230;
  assign n5232 = n5231 ^ n5216;
  assign n5254 = n5251 ^ n5232;
  assign n5255 = n5186 & n5254;
  assign n5257 = n5256 ^ n5255;
  assign n5253 = n5191 & n5252;
  assign n5258 = n5257 ^ n5253;
  assign n5245 = n5184 & n5232;
  assign n5226 = n5225 ^ n5216;
  assign n5227 = n5209 & n5226;
  assign n5228 = n5227 ^ n5199;
  assign n5243 = n5175 & n5228;
  assign n5241 = n5240 ^ n5228;
  assign n5242 = n5189 & n5241;
  assign n5244 = n5243 ^ n5242;
  assign n5246 = n5245 ^ n5244;
  assign n5233 = n5232 ^ n5228;
  assign n5235 = n5194 & n5233;
  assign n5234 = n5148 & n5233;
  assign n5236 = n5235 ^ n5234;
  assign n5247 = n5246 ^ n5236;
  assign n5259 = n5258 ^ n5247;
  assign n5572 = n5571 ^ n5259;
  assign n7188 = n7187 ^ n5572;
  assign n7191 = n7190 ^ n7188;
  assign n5518 = n4983 & n5026;
  assign n5517 = n4978 & n5516;
  assign n5519 = n5518 ^ n5517;
  assign n5515 = n4981 & n5026;
  assign n5520 = n5519 ^ n5515;
  assign n5036 = n4986 & n5033;
  assign n5513 = n5046 ^ n5036;
  assign n5510 = n4960 & n5032;
  assign n5511 = n5510 ^ n5039;
  assign n5509 = n4963 & n5029;
  assign n5512 = n5511 ^ n5509;
  assign n5514 = n5513 ^ n5512;
  assign n5521 = n5520 ^ n5514;
  assign n7185 = n7184 ^ n5521;
  assign n5679 = n5555 ^ n5545;
  assign n5599 = n5319 & n5553;
  assign n5600 = n5599 ^ n5348;
  assign n5678 = n5600 ^ n5550;
  assign n5680 = n5679 ^ n5678;
  assign n7182 = n5680 ^ n5373;
  assign n5489 = n5488 ^ n5479;
  assign n5501 = n5447 & n5489;
  assign n5503 = n5502 ^ n5501;
  assign n5497 = n5457 & n5496;
  assign n5495 = n5463 & n5487;
  assign n5498 = n5497 ^ n5495;
  assign n5500 = n5499 ^ n5498;
  assign n5504 = n5503 ^ n5500;
  assign n5493 = n5465 & n5487;
  assign n5490 = n5398 & n5489;
  assign n5492 = n5491 ^ n5490;
  assign n5494 = n5493 ^ n5492;
  assign n5505 = n5504 ^ n5494;
  assign n5375 = n5252 ^ n5233;
  assign n5384 = n5202 & n5375;
  assign n5385 = n5384 ^ n5235;
  assign n5381 = n5211 & n5241;
  assign n5380 = n5221 & n5240;
  assign n5382 = n5381 ^ n5380;
  assign n5383 = n5382 ^ n5242;
  assign n5386 = n5385 ^ n5383;
  assign n5378 = n5220 & n5240;
  assign n5376 = n5201 & n5375;
  assign n5377 = n5376 ^ n5234;
  assign n5379 = n5378 ^ n5377;
  assign n5387 = n5386 ^ n5379;
  assign n5506 = n5505 ^ n5387;
  assign n7183 = n7182 ^ n5506;
  assign n7186 = n7185 ^ n7183;
  assign n7192 = n7191 ^ n7186;
  assign n5035 = n4950 & n5034;
  assign n5037 = n5036 ^ n5035;
  assign n5670 = n5626 ^ n5037;
  assign n5669 = n5577 ^ n5040;
  assign n5671 = n5670 ^ n5669;
  assign n7180 = n7179 ^ n5671;
  assign n5647 = ~n5327 & n5342;
  assign n5646 = ~n5312 & n5365;
  assign n5648 = n5647 ^ n5646;
  assign n5715 = n5648 ^ n5358;
  assign n5714 = n5556 ^ n5369;
  assign n5716 = n5715 ^ n5714;
  assign n5601 = n5600 ^ n5546;
  assign n5598 = n5556 ^ n5547;
  assign n5602 = n5601 ^ n5598;
  assign n5717 = n5716 ^ n5602;
  assign n5614 = n5437 & n5478;
  assign n5613 = n5464 & n5483;
  assign n5615 = n5614 ^ n5613;
  assign n5616 = n5615 ^ n5561;
  assign n5610 = n5431 & n5566;
  assign n5611 = n5610 ^ n5492;
  assign n5612 = n5611 ^ n5567;
  assign n5617 = n5616 ^ n5612;
  assign n5606 = n5182 & n5232;
  assign n5605 = n5219 & n5251;
  assign n5607 = n5606 ^ n5605;
  assign n5608 = n5607 ^ n5244;
  assign n5541 = n5171 & n5254;
  assign n5542 = n5541 ^ n5377;
  assign n5604 = n5542 ^ n5255;
  assign n5609 = n5608 ^ n5604;
  assign n5618 = n5617 ^ n5609;
  assign n7178 = n5717 ^ n5618;
  assign n7181 = n7180 ^ n7178;
  assign n7193 = n7192 ^ n7181;
  assign n5580 = n4976 & n5029;
  assign n5579 = n5012 & n5025;
  assign n5581 = n5580 ^ n5579;
  assign n5582 = n5581 ^ n5511;
  assign n5578 = n5577 ^ n5517;
  assign n5583 = n5582 ^ n5578;
  assign n7166 = n5671 ^ n5583;
  assign n7168 = n7167 ^ n7166;
  assign n5650 = n5555 ^ n5544;
  assign n5645 = n5599 ^ n5371;
  assign n5649 = n5648 ^ n5645;
  assign n5651 = n5650 ^ n5649;
  assign n7164 = n5717 ^ n5651;
  assign n5653 = n5569 ^ n5501;
  assign n5720 = n5653 ^ n5615;
  assign n5656 = n5436 & n5483;
  assign n5719 = n5656 ^ n5492;
  assign n5721 = n5720 ^ n5719;
  assign n5538 = n5181 & n5251;
  assign n5643 = n5538 ^ n5377;
  assign n5641 = n5384 ^ n5257;
  assign n5642 = n5641 ^ n5607;
  assign n5644 = n5643 ^ n5642;
  assign n5722 = n5721 ^ n5644;
  assign n7165 = n7164 ^ n5722;
  assign n7169 = n7168 ^ n7165;
  assign n7231 = n7193 ^ n7169;
  assign n5753 = ~n5292 & n5346;
  assign n5754 = n5753 ^ n5546;
  assign n5755 = n5754 ^ n5360;
  assign n5752 = n5645 ^ n5556;
  assign n5756 = n5755 ^ n5752;
  assign n5757 = n5756 ^ n5602;
  assign n5695 = n5647 ^ n5351;
  assign n5696 = n5695 ^ n5549;
  assign n5694 = n5555 ^ n5546;
  assign n5697 = n5696 ^ n5694;
  assign n7174 = n5757 ^ n5697;
  assign n5624 = n4962 & n5032;
  assign n5627 = n5626 ^ n5624;
  assign n5628 = n5627 ^ n5512;
  assign n5622 = n5519 ^ n5035;
  assign n5623 = n5622 ^ n5577;
  assign n5629 = n5628 ^ n5623;
  assign n7171 = n5671 ^ n5629;
  assign n7173 = n7172 ^ n7171;
  assign n7175 = n7174 ^ n7173;
  assign n5735 = n5614 ^ n5560;
  assign n5736 = n5735 ^ n5498;
  assign n5657 = n5656 ^ n5493;
  assign n5734 = n5657 ^ n5492;
  assign n5737 = n5736 ^ n5734;
  assign n5690 = n5606 ^ n5243;
  assign n5691 = n5690 ^ n5382;
  assign n5539 = n5538 ^ n5378;
  assign n5689 = n5539 ^ n5377;
  assign n5692 = n5691 ^ n5689;
  assign n5738 = n5737 ^ n5692;
  assign n7170 = n7169 ^ n5738;
  assign n7176 = n7175 ^ n7170;
  assign n5049 = n5048 ^ n5047;
  assign n5044 = n5043 ^ n5037;
  assign n5050 = n5049 ^ n5044;
  assign n7161 = n7160 ^ n5050;
  assign n7158 = n5680 ^ n5602;
  assign n5683 = n5657 ^ n5503;
  assign n5682 = n5611 ^ n5497;
  assign n5684 = n5683 ^ n5682;
  assign n5596 = n5539 ^ n5385;
  assign n5595 = n5542 ^ n5381;
  assign n5597 = n5596 ^ n5595;
  assign n5685 = n5684 ^ n5597;
  assign n7159 = n7158 ^ n5685;
  assign n7162 = n7161 ^ n7159;
  assign n5741 = n5580 ^ n5510;
  assign n5742 = n5741 ^ n5042;
  assign n5740 = n5626 ^ n5047;
  assign n5743 = n5742 ^ n5740;
  assign n7154 = n5743 ^ n5671;
  assign n7156 = n7155 ^ n7154;
  assign n5698 = n5697 ^ n5602;
  assign n7152 = n5698 ^ n5557;
  assign n5700 = n5657 ^ n5500;
  assign n5701 = n5700 ^ n5611;
  assign n5540 = n5539 ^ n5383;
  assign n5543 = n5542 ^ n5540;
  assign n5702 = n5701 ^ n5543;
  assign n7153 = n7152 ^ n5702;
  assign n7157 = n7156 ^ n7153;
  assign n7163 = n7162 ^ n7157;
  assign n7177 = n7176 ^ n7163;
  assign n7209 = n7192 ^ n7177;
  assign n5725 = n5622 ^ n5581;
  assign n5724 = n5625 ^ n5047;
  assign n5726 = n5725 ^ n5724;
  assign n7199 = n7198 ^ n5726;
  assign n7196 = n5756 ^ n5651;
  assign n5662 = n5183 & n5228;
  assign n5663 = n5662 ^ n5539;
  assign n5664 = n5663 ^ n5246;
  assign n5661 = n5641 ^ n5542;
  assign n5665 = n5664 ^ n5661;
  assign n5655 = n5438 & n5474;
  assign n5658 = n5657 ^ n5655;
  assign n5659 = n5658 ^ n5563;
  assign n5654 = n5653 ^ n5611;
  assign n5660 = n5659 ^ n5654;
  assign n5666 = n5665 ^ n5660;
  assign n7197 = n7196 ^ n5666;
  assign n7200 = n7199 ^ n7197;
  assign n7208 = n7200 ^ n7162;
  assign n7241 = n7209 ^ n7208;
  assign n7194 = n7193 ^ n7157;
  assign n7239 = n7181 & n7194;
  assign n7219 = n7200 ^ n7157;
  assign n7205 = n7169 ^ n7162;
  assign n7228 = n7219 ^ n7205;
  assign n7229 = n7177 & n7228;
  assign n7240 = n7239 ^ n7229;
  assign n7242 = n7241 ^ n7240;
  assign n7211 = n7200 ^ n7186;
  assign n7212 = n7211 ^ n7176;
  assign n7213 = n7163 & n7212;
  assign n7210 = n7208 & n7209;
  assign n7214 = n7213 ^ n7210;
  assign n7243 = n7242 ^ n7214;
  assign n7235 = n7211 ^ n7177;
  assign n7201 = n7200 ^ n7191;
  assign n7220 = n7201 ^ n7163;
  assign n7221 = n7219 & n7220;
  assign n7222 = n7221 ^ n7213;
  assign n7236 = n7235 ^ n7222;
  assign n7230 = n7181 ^ n7177;
  assign n7232 = n7231 ^ n7208;
  assign n7233 = n7230 & n7232;
  assign n7234 = n7233 ^ n7229;
  assign n7237 = n7236 ^ n7234;
  assign n7260 = n7243 ^ n7237;
  assign n7224 = ~n7169 & n7193;
  assign n7202 = n7201 ^ n7176;
  assign n7206 = n7202 & n7205;
  assign n7225 = n7224 ^ n7206;
  assign n7218 = n7205 ^ n7202;
  assign n7223 = n7222 ^ n7218;
  assign n7226 = n7225 ^ n7223;
  assign n7238 = n7226 & n7237;
  assign n7261 = n7260 ^ n7238;
  assign n7203 = n7202 ^ n7193;
  assign n7195 = n7194 ^ n7163;
  assign n7216 = n7203 ^ n7195;
  assign n7204 = n7195 & n7203;
  assign n7207 = n7206 ^ n7204;
  assign n7215 = n7214 ^ n7207;
  assign n7217 = n7216 ^ n7215;
  assign n7258 = n7237 & ~n7243;
  assign n7259 = n7217 & n7258;
  assign n7262 = n7261 ^ n7259;
  assign n7950 = n7231 & n7262;
  assign n7266 = n7238 ^ n7217;
  assign n7267 = n7260 & n7266;
  assign n7268 = n7267 ^ n7243;
  assign n7918 = n7203 & n7268;
  assign n7951 = n7950 ^ n7918;
  assign n7227 = n7226 ^ n7217;
  assign n7249 = n7238 ^ n7227;
  assign n7247 = n7226 & n7243;
  assign n7248 = ~n7217 & n7247;
  assign n7250 = n7249 ^ n7248;
  assign n7272 = n7262 ^ n7250;
  assign n7821 = n7209 & n7272;
  assign n7269 = n7268 ^ n7262;
  assign n7820 = n7205 & n7269;
  assign n7822 = n7821 ^ n7820;
  assign n7244 = n7243 ^ n7238;
  assign n7245 = n7227 & n7244;
  assign n7246 = n7245 ^ n7217;
  assign n7271 = n7268 ^ n7246;
  assign n7273 = n7272 ^ n7271;
  assign n7797 = n7220 & n7273;
  assign n7886 = n7822 ^ n7797;
  assign n7952 = n7951 ^ n7886;
  assign n7275 = n7163 & n7271;
  assign n7274 = n7219 & n7273;
  assign n7276 = n7275 ^ n7274;
  assign n7263 = n7193 & n7262;
  assign n7949 = n7276 ^ n7263;
  assign n7953 = n7952 ^ n7949;
  assign n12663 = n10817 ^ n7953;
  assign n12666 = n12665 ^ n12663;
  assign n7976 = n7941 ^ n7844;
  assign n7662 = n7631 & ~n7661;
  assign n7657 = n7590 & n7656;
  assign n7663 = n7662 ^ n7657;
  assign n7977 = n7976 ^ n7663;
  assign n7975 = n7683 ^ n7673;
  assign n7978 = n7977 ^ n7975;
  assign n7788 = ~n7619 & ~n7678;
  assign n7790 = n7789 ^ n7788;
  assign n7791 = n7790 ^ n7673;
  assign n7787 = n7686 ^ n7662;
  assign n7792 = n7791 ^ n7787;
  assign n11661 = n7978 ^ n7792;
  assign n7665 = n7664 ^ n7663;
  assign n7674 = n7673 ^ n7665;
  assign n7687 = n7686 ^ n7674;
  assign n12642 = n11661 ^ n7687;
  assign n7550 = n7508 & n7514;
  assign n7519 = n7445 & n7518;
  assign n7551 = n7550 ^ n7519;
  assign n7783 = n7782 ^ n7551;
  assign n7850 = n7783 ^ n7543;
  assign n7851 = n7850 ^ n7536;
  assign n7381 = n7359 & ~n7378;
  assign n7380 = ~n7303 & ~n7379;
  assign n7382 = n7381 ^ n7380;
  assign n7384 = n7383 ^ n7382;
  assign n7393 = n7392 ^ n7384;
  assign n7406 = n7405 ^ n7393;
  assign n7852 = n7851 ^ n7406;
  assign n12643 = n12642 ^ n7852;
  assign n7814 = n7181 & n7246;
  assign n7919 = n7918 ^ n7814;
  assign n7251 = n7250 ^ n7246;
  assign n7254 = n7228 & n7251;
  assign n7253 = n7230 & n7250;
  assign n7255 = n7254 ^ n7253;
  assign n7920 = n7919 ^ n7255;
  assign n7257 = n7232 & n7250;
  assign n7264 = n7263 ^ n7257;
  assign n7917 = n7276 ^ n7264;
  assign n7921 = n7920 ^ n7917;
  assign n7796 = n7212 & n7271;
  assign n7798 = n7797 ^ n7796;
  assign n7799 = n7798 ^ n7264;
  assign n7270 = n7202 & n7269;
  assign n7277 = n7276 ^ n7270;
  assign n7795 = n7277 ^ n7254;
  assign n7800 = n7799 ^ n7795;
  assign n10625 = n7921 ^ n7800;
  assign n12641 = n10797 ^ n10625;
  assign n12644 = n12643 ^ n12641;
  assign n12667 = n12666 ^ n12644;
  assign n8011 = n7683 ^ n7666;
  assign n8010 = n7790 ^ n7665;
  assign n8012 = n8011 ^ n8010;
  assign n12648 = n8012 ^ n7792;
  assign n7538 = n7481 & n7524;
  assign n7540 = n7539 ^ n7538;
  assign n7544 = n7543 ^ n7540;
  assign n7537 = n7536 ^ n7519;
  assign n7545 = n7544 ^ n7537;
  assign n7409 = n7328 & ~n7397;
  assign n7411 = n7410 ^ n7409;
  assign n7412 = n7411 ^ n7392;
  assign n7408 = n7405 ^ n7380;
  assign n7413 = n7412 ^ n7408;
  assign n11669 = n7545 ^ n7413;
  assign n12649 = n12648 ^ n11669;
  assign n8000 = n7276 ^ n7257;
  assign n7252 = n7177 & n7251;
  assign n7256 = n7255 ^ n7252;
  assign n7999 = n7798 ^ n7256;
  assign n8001 = n8000 ^ n7999;
  assign n12647 = n10806 ^ n8001;
  assign n12650 = n12649 ^ n12647;
  assign n12651 = n12650 ^ n12644;
  assign n7984 = n7943 ^ n7845;
  assign n7983 = n7839 ^ n7686;
  assign n7985 = n7984 ^ n7983;
  assign n11675 = n7985 ^ n7792;
  assign n7876 = n7506 & n7528;
  assign n7547 = n7472 & n7523;
  assign n7877 = n7876 ^ n7547;
  assign n7938 = n7937 ^ n7877;
  assign n7936 = n7878 ^ n7536;
  assign n7939 = n7938 ^ n7936;
  assign n7870 = n7357 & ~n7389;
  assign n7414 = ~n7345 & ~n7396;
  assign n7871 = n7870 ^ n7414;
  assign n7932 = n7871 ^ n7826;
  assign n7931 = n7831 ^ n7405;
  assign n7933 = n7932 ^ n7931;
  assign n11645 = n7939 ^ n7933;
  assign n12638 = n11675 ^ n11645;
  assign n12637 = n10835 ^ n7800;
  assign n12639 = n12638 ^ n12637;
  assign n7265 = n7264 ^ n7256;
  assign n7278 = n7277 ^ n7265;
  assign n12634 = n10769 ^ n7278;
  assign n7842 = n7788 ^ n7679;
  assign n7847 = n7846 ^ n7842;
  assign n7837 = n7628 & ~n7680;
  assign n7841 = n7840 ^ n7837;
  assign n7848 = n7847 ^ n7841;
  assign n12632 = n7848 ^ n7687;
  assign n8005 = n7478 & n7529;
  assign n8006 = n8005 ^ n7880;
  assign n8003 = n7538 ^ n7532;
  assign n8004 = n8003 ^ n7971;
  assign n8007 = n8006 ^ n8004;
  assign n7830 = n7350 & n7399;
  assign n7834 = n7833 ^ n7830;
  assign n7825 = n7409 ^ n7398;
  assign n7829 = n7828 ^ n7825;
  assign n7835 = n7834 ^ n7829;
  assign n8008 = n8007 ^ n7835;
  assign n12633 = n12632 ^ n8008;
  assign n12635 = n12634 ^ n12633;
  assign n12629 = n8012 ^ n7848;
  assign n7785 = n7542 ^ n7533;
  assign n7784 = n7783 ^ n7540;
  assign n7786 = n7785 ^ n7784;
  assign n7779 = n7402 ^ n7391;
  assign n7778 = n7411 ^ n7384;
  assign n7780 = n7779 ^ n7778;
  assign n11654 = n7786 ^ n7780;
  assign n12630 = n12629 ^ n11654;
  assign n7819 = n7208 & n7272;
  assign n7823 = n7822 ^ n7819;
  assign n7816 = n7195 & n7268;
  assign n7815 = n7814 ^ n7252;
  assign n7817 = n7816 ^ n7815;
  assign n7813 = n7796 ^ n7275;
  assign n7818 = n7817 ^ n7813;
  assign n7824 = n7823 ^ n7818;
  assign n12628 = n10761 ^ n7824;
  assign n12631 = n12630 ^ n12628;
  assign n12636 = n12635 ^ n12631;
  assign n12640 = n12639 ^ n12636;
  assign n12645 = n12644 ^ n12640;
  assign n12704 = n12651 ^ n12645;
  assign n12687 = n12666 ^ n12635;
  assign n11683 = n7904 ^ n7792;
  assign n12658 = n11683 ^ n7978;
  assign n7888 = n7194 & n7246;
  assign n7889 = n7888 ^ n7264;
  assign n7890 = n7889 ^ n7817;
  assign n7887 = n7886 ^ n7277;
  assign n7891 = n7890 ^ n7887;
  assign n10639 = n7891 ^ n7800;
  assign n12657 = n10789 ^ n10639;
  assign n12659 = n12658 ^ n12657;
  assign n12653 = n11675 ^ n7946;
  assign n7883 = n7541 ^ n7533;
  assign n7882 = n7881 ^ n7877;
  assign n7884 = n7883 ^ n7882;
  assign n7874 = n7402 ^ n7390;
  assign n7873 = n7872 ^ n7871;
  assign n7875 = n7874 ^ n7873;
  assign n7885 = n7884 ^ n7875;
  assign n12654 = n12653 ^ n7885;
  assign n7989 = n7951 ^ n7815;
  assign n7988 = n7820 ^ n7277;
  assign n7990 = n7989 ^ n7988;
  assign n10632 = n7990 ^ n7800;
  assign n12652 = n10778 ^ n10632;
  assign n12655 = n12654 ^ n12652;
  assign n7549 = n7548 ^ n7547;
  assign n7552 = n7551 ^ n7549;
  assign n7546 = n7543 ^ n7533;
  assign n7553 = n7552 ^ n7546;
  assign n7418 = n7402 ^ n7392;
  assign n7416 = n7415 ^ n7414;
  assign n7417 = n7416 ^ n7382;
  assign n7419 = n7418 ^ n7417;
  assign n11681 = n7553 ^ n7419;
  assign n12656 = n12655 ^ n11681;
  assign n12660 = n12659 ^ n12656;
  assign n12694 = n12687 ^ n12660;
  assign n12703 = n12694 ^ n12640;
  assign n12708 = n12704 ^ n12703;
  assign n12705 = ~n12703 & ~n12704;
  assign n12662 = n12655 ^ n12650;
  assign n12698 = ~n12662 & n12694;
  assign n12706 = n12705 ^ n12698;
  assign n12676 = n12666 ^ n12631;
  assign n12677 = n12676 ^ n12660;
  assign n12678 = n12651 & n12677;
  assign n12671 = n12666 ^ n12650;
  assign n12661 = n12660 ^ n12651;
  assign n12672 = n12661 ^ n12636;
  assign n12675 = n12671 & ~n12672;
  assign n12679 = n12678 ^ n12675;
  assign n12707 = n12706 ^ n12679;
  assign n12709 = n12708 ^ n12707;
  assign n12697 = ~n12640 & n12655;
  assign n12699 = n12698 ^ n12697;
  assign n12695 = n12694 ^ n12662;
  assign n12688 = n12687 ^ n12651;
  assign n12689 = n12667 & ~n12688;
  assign n12690 = n12689 ^ n12678;
  assign n12696 = n12695 ^ n12690;
  assign n12700 = n12699 ^ n12696;
  assign n12716 = n12709 ^ n12700;
  assign n12686 = n12676 ^ n12661;
  assign n12691 = n12690 ^ n12686;
  assign n12681 = n12655 ^ n12640;
  assign n12682 = n12681 ^ n12671;
  assign n12683 = n12661 ^ n12639;
  assign n12684 = n12682 & n12683;
  assign n12668 = n12667 ^ n12662;
  assign n12669 = ~n12661 & ~n12668;
  assign n12685 = n12684 ^ n12669;
  assign n12692 = n12691 ^ n12685;
  assign n12701 = n12692 & ~n12700;
  assign n12717 = n12716 ^ n12701;
  assign n12673 = n12672 ^ n12671;
  assign n12646 = ~n12639 & ~n12645;
  assign n12670 = n12669 ^ n12646;
  assign n12674 = n12673 ^ n12670;
  assign n12680 = n12679 ^ n12674;
  assign n12714 = ~n12680 & ~n12700;
  assign n12715 = ~n12709 & n12714;
  assign n12718 = n12717 ^ n12715;
  assign n12710 = n12680 & n12692;
  assign n12711 = n12709 & n12710;
  assign n12693 = n12692 ^ n12680;
  assign n12702 = n12701 ^ n12693;
  assign n12712 = n12711 ^ n12702;
  assign n12729 = n12718 ^ n12712;
  assign n12724 = n12709 ^ n12701;
  assign n12725 = ~n12693 & n12724;
  assign n12726 = n12725 ^ n12680;
  assign n12721 = n12701 ^ n12680;
  assign n12722 = ~n12716 & ~n12721;
  assign n12723 = n12722 ^ n12709;
  assign n12727 = n12726 ^ n12723;
  assign n12730 = n12729 ^ n12727;
  assign n12731 = n12667 & ~n12730;
  assign n12728 = n12651 & ~n12727;
  assign n12732 = n12731 ^ n12728;
  assign n12719 = n12682 & ~n12718;
  assign n12977 = n12732 ^ n12719;
  assign n12737 = n12723 ^ n12718;
  assign n12942 = ~n12661 & ~n12737;
  assign n12739 = n12683 & ~n12718;
  assign n12738 = ~n12668 & ~n12737;
  assign n12740 = n12739 ^ n12738;
  assign n12975 = n12942 ^ n12740;
  assign n12748 = n12677 & ~n12727;
  assign n12747 = ~n12688 & ~n12730;
  assign n12749 = n12748 ^ n12747;
  assign n12976 = n12975 ^ n12749;
  assign n12978 = n12977 ^ n12976;
  assign n12988 = n12987 ^ n12978;
  assign n9189 = n3735 ^ n3518;
  assign n9190 = n9189 ^ n7606;
  assign n9188 = n8117 ^ n3750;
  assign n9191 = n9190 ^ n9188;
  assign n9178 = n3832 ^ n3687;
  assign n9179 = n9178 ^ n3865;
  assign n9177 = n8111 ^ n3826;
  assign n9180 = n9179 ^ n9177;
  assign n9212 = n9191 ^ n9180;
  assign n9199 = n7566 ^ n3771;
  assign n8610 = n3854 ^ n2681;
  assign n9198 = n8610 ^ n8134;
  assign n9200 = n9199 ^ n9198;
  assign n9194 = n7556 ^ n3735;
  assign n9195 = n9194 ^ n1870;
  assign n8603 = n3854 ^ n3784;
  assign n9193 = n8603 ^ n8125;
  assign n9196 = n9195 ^ n9193;
  assign n9197 = n9196 ^ n7562;
  assign n9201 = n9200 ^ n9197;
  assign n9213 = n9212 ^ n9201;
  assign n9169 = n3868 ^ n3687;
  assign n9170 = n9169 ^ n7572;
  assign n9168 = n8165 ^ n3649;
  assign n9171 = n9170 ^ n9168;
  assign n9165 = n7576 ^ n3814;
  assign n9166 = n9165 ^ n3837;
  assign n8594 = n3854 ^ n3707;
  assign n9164 = n8594 ^ n8156;
  assign n9167 = n9166 ^ n9164;
  assign n9172 = n9171 ^ n9167;
  assign n9209 = n9201 ^ n9172;
  assign n9174 = n3832 ^ n3814;
  assign n9175 = n9174 ^ n3677;
  assign n9173 = n8148 ^ n3802;
  assign n9176 = n9175 ^ n9173;
  assign n9181 = n9180 ^ n9176;
  assign n9210 = n9209 ^ n9181;
  assign n9208 = n9191 ^ n9171;
  assign n9242 = n9210 ^ n9208;
  assign n9183 = n7587 ^ n7556;
  assign n9182 = n8142 ^ n3854;
  assign n9184 = n9183 ^ n9182;
  assign n9185 = n9184 ^ n9181;
  assign n9186 = n9185 ^ n9167;
  assign n9240 = ~n9184 & ~n9186;
  assign n9220 = n9191 ^ n9167;
  assign n9205 = n9196 ^ n9171;
  assign n9229 = n9220 ^ n9205;
  assign n9230 = ~n9209 & ~n9229;
  assign n9241 = n9240 ^ n9230;
  assign n9243 = n9242 ^ n9241;
  assign n9214 = n9172 & n9213;
  assign n9211 = n9208 & ~n9210;
  assign n9215 = n9214 ^ n9211;
  assign n9244 = n9243 ^ n9215;
  assign n9236 = n9212 ^ n9209;
  assign n9192 = n9191 ^ n9176;
  assign n9221 = n9192 ^ n9172;
  assign n9222 = n9220 & ~n9221;
  assign n9223 = n9222 ^ n9214;
  assign n9237 = n9236 ^ n9223;
  assign n9231 = n9196 ^ n9185;
  assign n9232 = n9231 ^ n9208;
  assign n9233 = n9209 ^ n9184;
  assign n9234 = n9232 & n9233;
  assign n9235 = n9234 ^ n9230;
  assign n9238 = n9237 ^ n9235;
  assign n9248 = n9244 ^ n9238;
  assign n9225 = ~n9185 & n9196;
  assign n9202 = n9201 ^ n9192;
  assign n9206 = n9202 & ~n9205;
  assign n9226 = n9225 ^ n9206;
  assign n9219 = n9205 ^ n9202;
  assign n9224 = n9223 ^ n9219;
  assign n9227 = n9226 ^ n9224;
  assign n9239 = ~n9227 & n9238;
  assign n9203 = n9202 ^ n9185;
  assign n9187 = n9186 ^ n9172;
  assign n9217 = n9203 ^ n9187;
  assign n9204 = ~n9187 & ~n9203;
  assign n9207 = n9206 ^ n9204;
  assign n9216 = n9215 ^ n9207;
  assign n9218 = n9217 ^ n9216;
  assign n9249 = n9239 ^ n9218;
  assign n9250 = ~n9248 & n9249;
  assign n9251 = n9250 ^ n9244;
  assign n9228 = n9227 ^ n9218;
  assign n9245 = n9244 ^ n9239;
  assign n9246 = ~n9228 & ~n9245;
  assign n9247 = n9246 ^ n9218;
  assign n9252 = n9251 ^ n9247;
  assign n9284 = n9213 & ~n9252;
  assign n9260 = n9239 ^ n9228;
  assign n9258 = ~n9227 & ~n9244;
  assign n9259 = ~n9218 & n9258;
  assign n9261 = n9260 ^ n9259;
  assign n9255 = n9238 & n9244;
  assign n9256 = n9218 & n9255;
  assign n9254 = n9248 ^ n9239;
  assign n9257 = n9256 ^ n9254;
  assign n9262 = n9261 ^ n9257;
  assign n9263 = n9262 ^ n9252;
  assign n9283 = ~n9221 & ~n9263;
  assign n9285 = n9284 ^ n9283;
  assign n9267 = n9232 & ~n9261;
  assign n9266 = ~n9185 & ~n9257;
  assign n9268 = n9267 ^ n9266;
  assign n9286 = n9285 ^ n9268;
  assign n9279 = n9257 ^ n9251;
  assign n9280 = n9202 & n9279;
  assign n9264 = n9220 & ~n9263;
  assign n9253 = n9172 & ~n9252;
  assign n9265 = n9264 ^ n9253;
  assign n9281 = n9280 ^ n9265;
  assign n9274 = n9261 ^ n9247;
  assign n9275 = ~n9229 & ~n9274;
  assign n9282 = n9281 ^ n9275;
  assign n9287 = n9286 ^ n9282;
  assign n12515 = n12514 ^ n9287;
  assign n6525 = n6524 ^ n6518;
  assign n9431 = n6547 ^ n6525;
  assign n9432 = n9431 ^ n6633;
  assign n9433 = n9432 ^ n6561;
  assign n9434 = n9433 ^ n3637;
  assign n9427 = n6479 ^ n3698;
  assign n6598 = n6597 ^ n6590;
  assign n9425 = n6598 ^ n6459;
  assign n9426 = n9425 ^ n6617;
  assign n9428 = n9427 ^ n9426;
  assign n9437 = n9434 ^ n9428;
  assign n8363 = n6628 ^ n6472;
  assign n9418 = n8363 ^ n6430;
  assign n9417 = n7312 ^ n6535;
  assign n9419 = n9418 ^ n9417;
  assign n9415 = n6412 ^ n3713;
  assign n9413 = n6638 ^ n3756;
  assign n8356 = n6472 ^ n6162;
  assign n9411 = n8356 ^ n6511;
  assign n9410 = n7291 ^ n6518;
  assign n9412 = n9411 ^ n9410;
  assign n9414 = n9413 ^ n9412;
  assign n9416 = n9415 ^ n9414;
  assign n9420 = n9419 ^ n9416;
  assign n9438 = n9437 ^ n9420;
  assign n9446 = n6472 ^ n6391;
  assign n9447 = n9446 ^ n7291;
  assign n9445 = n6496 ^ n3788;
  assign n9448 = n9447 ^ n9445;
  assign n9422 = n7322 ^ n6582;
  assign n6454 = n6453 ^ n6444;
  assign n9423 = n9422 ^ n6454;
  assign n9424 = n9423 ^ n3844;
  assign n9429 = n9428 ^ n9424;
  assign n9449 = n9448 ^ n9429;
  assign n9478 = n9449 ^ n9414;
  assign n6618 = n6617 ^ n6614;
  assign n9402 = n6618 ^ n6401;
  assign n9403 = n9402 ^ n7332;
  assign n9404 = n9403 ^ n3858;
  assign n9435 = n9434 ^ n9404;
  assign n9479 = n9478 ^ n9435;
  assign n9405 = n7304 ^ n7284;
  assign n8350 = n6531 ^ n6472;
  assign n9406 = n9405 ^ n8350;
  assign n9407 = n9406 ^ n6434;
  assign n9408 = n9407 ^ n3818;
  assign n9409 = n9408 ^ n9404;
  assign n9421 = n9420 ^ n9409;
  assign n9480 = n9448 ^ n9421;
  assign n9481 = n9479 & n9480;
  assign n9458 = n9434 ^ n9408;
  assign n9443 = n9414 ^ n9404;
  assign n9468 = n9458 ^ n9443;
  assign n9469 = ~n9421 & ~n9468;
  assign n9482 = n9481 ^ n9469;
  assign n9476 = n9437 ^ n9421;
  assign n9441 = n9434 ^ n9424;
  assign n9459 = n9441 ^ n9409;
  assign n9460 = n9458 & ~n9459;
  assign n9439 = n9409 & n9438;
  assign n9461 = n9460 ^ n9439;
  assign n9477 = n9476 ^ n9461;
  assign n9483 = n9482 ^ n9477;
  assign n9430 = n9429 ^ n9421;
  assign n9471 = n9435 ^ n9430;
  assign n9450 = n9449 ^ n9408;
  assign n9467 = ~n9448 & ~n9450;
  assign n9470 = n9469 ^ n9467;
  assign n9472 = n9471 ^ n9470;
  assign n9436 = ~n9430 & n9435;
  assign n9440 = n9439 ^ n9436;
  assign n9473 = n9472 ^ n9440;
  assign n9498 = n9483 ^ n9473;
  assign n9464 = n9414 & ~n9449;
  assign n9442 = n9441 ^ n9420;
  assign n9444 = n9442 & ~n9443;
  assign n9465 = n9464 ^ n9444;
  assign n9462 = n9443 ^ n9442;
  assign n9463 = n9462 ^ n9461;
  assign n9466 = n9465 ^ n9463;
  assign n9484 = ~n9466 & n9483;
  assign n9452 = n9449 ^ n9442;
  assign n9451 = n9450 ^ n9409;
  assign n9456 = n9452 ^ n9451;
  assign n9453 = ~n9451 & ~n9452;
  assign n9454 = n9453 ^ n9444;
  assign n9455 = n9454 ^ n9440;
  assign n9457 = n9456 ^ n9455;
  assign n9506 = n9484 ^ n9457;
  assign n9507 = ~n9498 & n9506;
  assign n9508 = n9507 ^ n9473;
  assign n9485 = n9466 ^ n9457;
  assign n9488 = n9484 ^ n9473;
  assign n9489 = ~n9485 & ~n9488;
  assign n9490 = n9489 ^ n9457;
  assign n9509 = n9508 ^ n9490;
  assign n9633 = n9438 & ~n9509;
  assign n9500 = n9473 & n9483;
  assign n9501 = n9457 & n9500;
  assign n9499 = n9498 ^ n9484;
  assign n9502 = n9501 ^ n9499;
  assign n9486 = n9485 ^ n9484;
  assign n9474 = ~n9466 & ~n9473;
  assign n9475 = ~n9457 & n9474;
  assign n9487 = n9486 ^ n9475;
  assign n9511 = n9502 ^ n9487;
  assign n9512 = n9511 ^ n9509;
  assign n9632 = ~n9459 & ~n9512;
  assign n9634 = n9633 ^ n9632;
  assign n9503 = ~n9449 & ~n9502;
  assign n9497 = n9479 & ~n9487;
  assign n9504 = n9503 ^ n9497;
  assign n9635 = n9634 ^ n9504;
  assign n9515 = n9508 ^ n9502;
  assign n9516 = n9442 & n9515;
  assign n9513 = n9458 & ~n9512;
  assign n9510 = n9409 & ~n9509;
  assign n9514 = n9513 ^ n9510;
  assign n9517 = n9516 ^ n9514;
  assign n9491 = n9490 ^ n9487;
  assign n9494 = ~n9468 & ~n9491;
  assign n9631 = n9517 ^ n9494;
  assign n9636 = n9635 ^ n9631;
  assign n9057 = n5050 ^ n4798;
  assign n8503 = n5571 ^ n5521;
  assign n5681 = n5680 ^ n5387;
  assign n9056 = n8503 ^ n5681;
  assign n9058 = n9057 ^ n9056;
  assign n9045 = n5756 ^ n5665;
  assign n9044 = n5726 ^ n5721;
  assign n9046 = n9045 ^ n9044;
  assign n9043 = n5629 ^ n4735;
  assign n9047 = n9046 ^ n9043;
  assign n9088 = n9058 ^ n9047;
  assign n9075 = n5697 ^ n5692;
  assign n8497 = n5684 ^ n5660;
  assign n9074 = n8497 ^ n7171;
  assign n9076 = n9075 ^ n9074;
  assign n9071 = n5726 ^ n4650;
  assign n8489 = n5684 ^ n5617;
  assign n9069 = n8489 ^ n7166;
  assign n5652 = n5651 ^ n5644;
  assign n9070 = n9069 ^ n5652;
  assign n9072 = n9071 ^ n9070;
  assign n9068 = n5743 ^ n4627;
  assign n9073 = n9072 ^ n9068;
  assign n9077 = n9076 ^ n9073;
  assign n9089 = n9088 ^ n9077;
  assign n9041 = n5705 ^ n4170;
  assign n8471 = n5737 ^ n5684;
  assign n9039 = n8471 ^ n7154;
  assign n5558 = n5557 ^ n5543;
  assign n9040 = n9039 ^ n5558;
  assign n9042 = n9041 ^ n9040;
  assign n9048 = n9047 ^ n9042;
  assign n9054 = n5521 ^ n4774;
  assign n8472 = n5705 ^ n5701;
  assign n5374 = n5373 ^ n5259;
  assign n9053 = n8472 ^ n5374;
  assign n9055 = n9054 ^ n9053;
  assign n9067 = n9055 ^ n9047;
  assign n8507 = n5505 ^ n5050;
  assign n5603 = n5602 ^ n5597;
  assign n9063 = n8507 ^ n5603;
  assign n9062 = n5671 ^ n4591;
  assign n9064 = n9063 ^ n9062;
  assign n9065 = n9064 ^ n9042;
  assign n9108 = n9067 ^ n9065;
  assign n9109 = n9048 & n9108;
  assign n9090 = n9065 & n9089;
  assign n9110 = n9109 ^ n9090;
  assign n9084 = n9077 ^ n9065;
  assign n9107 = n9088 ^ n9084;
  assign n9111 = n9110 ^ n9107;
  assign n9059 = n9058 ^ n9055;
  assign n9049 = n7166 ^ n5684;
  assign n9050 = n9049 ^ n5609;
  assign n9051 = n9050 ^ n5716;
  assign n9052 = n9051 ^ n4839;
  assign n9060 = n9059 ^ n9052;
  assign n9102 = n9072 ^ n9060;
  assign n9086 = n9064 ^ n9047;
  assign n9103 = n9102 ^ n9086;
  assign n9104 = n9084 ^ n9052;
  assign n9105 = n9103 & n9104;
  assign n9081 = n9072 ^ n9064;
  assign n9095 = n9081 ^ n9048;
  assign n9096 = n9084 & n9095;
  assign n9106 = n9105 ^ n9096;
  assign n9112 = n9111 ^ n9106;
  assign n9085 = n9084 ^ n9059;
  assign n9099 = n9086 ^ n9085;
  assign n9061 = n9060 ^ n9042;
  assign n9097 = n9052 & n9061;
  assign n9098 = n9097 ^ n9096;
  assign n9100 = n9099 ^ n9098;
  assign n9087 = n9085 & n9086;
  assign n9091 = n9090 ^ n9087;
  assign n9101 = n9100 ^ n9091;
  assign n9121 = n9112 ^ n9101;
  assign n9117 = n9060 & ~n9072;
  assign n9078 = n9077 ^ n9067;
  assign n9082 = n9078 & n9081;
  assign n9118 = n9117 ^ n9082;
  assign n9115 = n9081 ^ n9078;
  assign n9116 = n9115 ^ n9110;
  assign n9119 = n9118 ^ n9116;
  assign n9120 = n9112 & n9119;
  assign n9079 = n9078 ^ n9060;
  assign n9066 = n9065 ^ n9061;
  assign n9093 = n9079 ^ n9066;
  assign n9080 = n9066 & n9079;
  assign n9083 = n9082 ^ n9080;
  assign n9092 = n9091 ^ n9083;
  assign n9094 = n9093 ^ n9092;
  assign n9133 = n9120 ^ n9094;
  assign n9134 = n9121 & n9133;
  assign n9135 = n9134 ^ n9101;
  assign n9126 = n9119 ^ n9094;
  assign n9130 = n9120 ^ n9101;
  assign n9131 = n9126 & n9130;
  assign n9132 = n9131 ^ n9094;
  assign n9136 = n9135 ^ n9132;
  assign n9159 = n9089 & n9136;
  assign n9127 = n9126 ^ n9120;
  assign n9124 = n9101 & n9119;
  assign n9125 = ~n9094 & n9124;
  assign n9128 = n9127 ^ n9125;
  assign n9122 = n9121 ^ n9120;
  assign n9113 = ~n9101 & n9112;
  assign n9114 = n9094 & n9113;
  assign n9123 = n9122 ^ n9114;
  assign n9129 = n9128 ^ n9123;
  assign n9137 = n9136 ^ n9129;
  assign n9158 = n9108 & n9137;
  assign n9160 = n9159 ^ n9158;
  assign n9142 = n9103 & n9128;
  assign n9141 = n9060 & n9123;
  assign n9143 = n9142 ^ n9141;
  assign n9161 = n9160 ^ n9143;
  assign n9154 = n9135 ^ n9123;
  assign n9155 = n9078 & n9154;
  assign n9139 = n9065 & n9136;
  assign n9138 = n9048 & n9137;
  assign n9140 = n9139 ^ n9138;
  assign n9156 = n9155 ^ n9140;
  assign n9149 = n9132 ^ n9128;
  assign n9150 = n9095 & n9149;
  assign n9157 = n9156 ^ n9150;
  assign n9162 = n9161 ^ n9157;
  assign n10810 = n9636 ^ n9162;
  assign n8159 = n4716 ^ n4606;
  assign n9309 = n8159 ^ n7440;
  assign n9310 = n9309 ^ n7451;
  assign n9308 = n8249 ^ n4075;
  assign n9311 = n9310 ^ n9308;
  assign n8169 = n4600 ^ n4321;
  assign n4808 = n4807 ^ n4804;
  assign n9305 = n8169 ^ n4808;
  assign n9304 = n8250 ^ n4185;
  assign n9306 = n9305 ^ n9304;
  assign n9312 = n9311 ^ n9306;
  assign n8137 = n4746 ^ n4606;
  assign n9319 = n8137 ^ n7466;
  assign n9318 = n8252 ^ n4179;
  assign n9320 = n9319 ^ n9318;
  assign n8128 = n4833 ^ n4606;
  assign n9314 = n8128 ^ n7424;
  assign n9315 = n9314 ^ n7434;
  assign n9313 = n8253 ^ n4639;
  assign n9316 = n9315 ^ n9313;
  assign n8132 = n4721 ^ n4312;
  assign n9317 = n9316 ^ n8132;
  assign n9321 = n9320 ^ n9317;
  assign n9322 = n9321 ^ n9312;
  assign n4788 = n4787 ^ n4782;
  assign n9294 = n7428 ^ n4788;
  assign n9293 = n8262 ^ n4610;
  assign n9295 = n9294 ^ n9293;
  assign n4581 = n4580 ^ n4447;
  assign n9291 = n7454 ^ n4581;
  assign n9290 = n8258 ^ n4767;
  assign n9292 = n9291 ^ n9290;
  assign n9296 = n9295 ^ n9292;
  assign n9323 = n9322 ^ n9296;
  assign n8121 = n4754 ^ n4709;
  assign n4688 = n4687 ^ n4677;
  assign n9302 = n8121 ^ n4688;
  assign n9301 = n8256 ^ n4698;
  assign n9303 = n9302 ^ n9301;
  assign n9307 = n9306 ^ n9303;
  assign n9357 = n9323 ^ n9307;
  assign n8145 = n4829 ^ n4665;
  assign n4607 = n4606 ^ n4600;
  assign n9298 = n8145 ^ n4607;
  assign n9297 = n8271 ^ n4657;
  assign n9299 = n9298 ^ n9297;
  assign n9300 = n9299 ^ n9296;
  assign n9332 = n9311 ^ n9300;
  assign n9355 = n9299 & n9332;
  assign n9342 = n9311 ^ n9303;
  assign n9335 = n9316 ^ n9306;
  assign n9351 = n9342 ^ n9335;
  assign n9352 = ~n9322 & ~n9351;
  assign n9356 = n9355 ^ n9352;
  assign n9358 = n9357 ^ n9356;
  assign n9325 = n9303 ^ n9295;
  assign n9326 = n9325 ^ n9321;
  assign n9327 = n9312 & ~n9326;
  assign n9324 = n9307 & ~n9323;
  assign n9328 = n9327 ^ n9324;
  assign n9359 = n9358 ^ n9328;
  assign n9347 = n9316 ^ n9300;
  assign n9348 = n9347 ^ n9307;
  assign n9349 = n9322 ^ n9299;
  assign n9350 = ~n9348 & ~n9349;
  assign n9353 = n9352 ^ n9350;
  assign n9329 = n9303 ^ n9292;
  assign n9343 = n9329 ^ n9312;
  assign n9344 = n9342 & n9343;
  assign n9345 = n9344 ^ n9327;
  assign n9341 = n9325 ^ n9322;
  assign n9346 = n9345 ^ n9341;
  assign n9354 = n9353 ^ n9346;
  assign n9362 = n9359 ^ n9354;
  assign n9365 = n9300 & n9316;
  assign n9330 = n9329 ^ n9321;
  assign n9336 = ~n9330 & ~n9335;
  assign n9366 = n9365 ^ n9336;
  assign n9363 = n9335 ^ n9330;
  assign n9364 = n9363 ^ n9345;
  assign n9367 = n9366 ^ n9364;
  assign n9368 = ~n9354 & n9367;
  assign n9333 = n9332 ^ n9312;
  assign n9331 = n9330 ^ n9300;
  assign n9339 = n9333 ^ n9331;
  assign n9334 = ~n9331 & n9333;
  assign n9337 = n9336 ^ n9334;
  assign n9338 = n9337 ^ n9328;
  assign n9340 = n9339 ^ n9338;
  assign n9389 = n9368 ^ n9340;
  assign n9390 = n9362 & ~n9389;
  assign n9391 = n9390 ^ n9359;
  assign n9374 = n9367 ^ n9340;
  assign n9379 = n9368 ^ n9359;
  assign n9380 = ~n9374 & ~n9379;
  assign n9381 = n9380 ^ n9340;
  assign n9395 = n9391 ^ n9381;
  assign n9398 = n9312 & n9395;
  assign n9375 = n9374 ^ n9368;
  assign n9372 = ~n9359 & n9367;
  assign n9373 = n9340 & n9372;
  assign n9376 = n9375 ^ n9373;
  assign n9369 = n9368 ^ n9362;
  assign n9360 = ~n9354 & n9359;
  assign n9361 = ~n9340 & n9360;
  assign n9370 = n9369 ^ n9361;
  assign n9394 = n9376 ^ n9370;
  assign n9396 = n9395 ^ n9394;
  assign n9397 = n9342 & ~n9396;
  assign n9399 = n9398 ^ n9397;
  assign n9377 = ~n9348 & ~n9376;
  assign n9854 = n9399 ^ n9377;
  assign n9627 = ~n9326 & n9395;
  assign n9626 = n9343 & ~n9396;
  assign n9628 = n9627 ^ n9626;
  assign n9385 = ~n9349 & ~n9376;
  assign n9382 = n9381 ^ n9376;
  assign n9384 = ~n9351 & n9382;
  assign n9386 = n9385 ^ n9384;
  assign n9383 = ~n9322 & n9382;
  assign n9387 = n9386 ^ n9383;
  assign n9853 = n9628 ^ n9387;
  assign n9855 = n9854 ^ n9853;
  assign n9851 = n9514 ^ n9497;
  assign n9493 = n9480 & ~n9487;
  assign n9495 = n9494 ^ n9493;
  assign n9492 = ~n9421 & ~n9491;
  assign n9496 = n9495 ^ n9492;
  assign n9850 = n9634 ^ n9496;
  assign n9852 = n9851 ^ n9850;
  assign n9856 = n9855 ^ n9852;
  assign n12513 = n10810 ^ n9856;
  assign n12516 = n12515 ^ n12513;
  assign n9521 = ~n9209 & ~n9274;
  assign n9273 = n9233 & ~n9261;
  assign n9276 = n9275 ^ n9273;
  assign n9522 = n9521 ^ n9276;
  assign n9523 = n9522 ^ n9268;
  assign n9524 = n9523 ^ n9281;
  assign n12510 = n12509 ^ n9524;
  assign n9725 = ~n9448 & n9490;
  assign n9681 = ~n9452 & ~n9508;
  assign n9726 = n9725 ^ n9681;
  assign n9727 = n9726 ^ n9495;
  assign n9724 = n9514 ^ n9504;
  assign n9728 = n9727 ^ n9724;
  assign n11543 = n9728 ^ n9636;
  assign n9730 = n9299 & ~n9381;
  assign n9675 = ~n9331 & ~n9391;
  assign n9731 = n9730 ^ n9675;
  assign n9732 = n9731 ^ n9386;
  assign n9371 = n9300 & n9370;
  assign n9378 = n9377 ^ n9371;
  assign n9729 = n9399 ^ n9378;
  assign n9733 = n9732 ^ n9729;
  assign n9629 = n9628 ^ n9378;
  assign n9392 = n9391 ^ n9370;
  assign n9393 = ~n9330 & ~n9392;
  assign n9400 = n9399 ^ n9393;
  assign n9625 = n9400 ^ n9384;
  assign n9630 = n9629 ^ n9625;
  assign n10800 = n9733 ^ n9630;
  assign n12507 = n11543 ^ n10800;
  assign n9616 = n9084 & n9149;
  assign n9148 = n9104 & n9128;
  assign n9151 = n9150 ^ n9148;
  assign n9617 = n9616 ^ n9151;
  assign n9813 = n9617 ^ n9143;
  assign n9814 = n9813 ^ n9156;
  assign n9505 = n9504 ^ n9496;
  assign n9518 = n9517 ^ n9505;
  assign n10802 = n9814 ^ n9518;
  assign n12508 = n12507 ^ n10802;
  assign n12511 = n12510 ^ n12508;
  assign n12517 = n12516 ^ n12511;
  assign n9271 = ~n9184 & n9247;
  assign n9270 = ~n9203 & ~n9251;
  assign n9272 = n9271 ^ n9270;
  assign n9277 = n9276 ^ n9272;
  assign n9269 = n9268 ^ n9265;
  assign n9278 = n9277 ^ n9269;
  assign n12527 = n12526 ^ n9278;
  assign n9789 = ~n9450 & n9490;
  assign n9790 = n9789 ^ n9504;
  assign n9787 = ~n9451 & ~n9508;
  assign n9760 = n9725 ^ n9492;
  assign n9788 = n9787 ^ n9760;
  assign n9791 = n9790 ^ n9788;
  assign n9684 = ~n9430 & n9511;
  assign n9683 = ~n9443 & n9515;
  assign n9685 = n9684 ^ n9683;
  assign n9686 = n9685 ^ n9632;
  assign n9786 = n9686 ^ n9517;
  assign n9792 = n9791 ^ n9786;
  assign n11550 = n9792 ^ n9636;
  assign n9782 = n9333 & ~n9391;
  assign n9765 = n9730 ^ n9383;
  assign n9783 = n9782 ^ n9765;
  assign n9780 = n9332 & ~n9381;
  assign n9781 = n9780 ^ n9378;
  assign n9784 = n9783 ^ n9781;
  assign n9671 = ~n9323 & ~n9394;
  assign n9670 = ~n9335 & ~n9392;
  assign n9672 = n9671 ^ n9670;
  assign n9673 = n9672 ^ n9626;
  assign n9779 = n9673 ^ n9400;
  assign n9785 = n9784 ^ n9779;
  assign n10792 = n9785 ^ n9630;
  assign n12525 = n11550 ^ n10792;
  assign n12528 = n12527 ^ n12525;
  assign n9692 = ~n9210 & n9262;
  assign n9660 = ~n9205 & n9279;
  assign n9693 = n9692 ^ n9660;
  assign n9694 = n9693 ^ n9283;
  assign n9662 = n9231 & ~n9257;
  assign n9663 = n9662 ^ n9270;
  assign n9695 = n9694 ^ n9663;
  assign n9691 = n9266 ^ n9265;
  assign n9696 = n9695 ^ n9691;
  assign n12522 = n12521 ^ n9696;
  assign n9680 = n9478 & ~n9502;
  assign n9682 = n9681 ^ n9680;
  assign n9761 = n9760 ^ n9682;
  assign n9759 = n9683 ^ n9517;
  assign n9762 = n9761 ^ n9759;
  assign n11530 = n9762 ^ n9636;
  assign n9674 = ~n9347 & n9370;
  assign n9676 = n9675 ^ n9674;
  assign n9766 = n9765 ^ n9676;
  assign n9764 = n9670 ^ n9400;
  assign n9767 = n9766 ^ n9764;
  assign n10781 = n9767 ^ n9630;
  assign n12519 = n11530 ^ n10781;
  assign n9735 = n9085 & n9129;
  assign n9652 = n9081 & n9154;
  assign n9736 = n9735 ^ n9652;
  assign n9737 = n9736 ^ n9158;
  assign n9654 = n9102 & n9123;
  assign n9145 = n9079 & n9135;
  assign n9655 = n9654 ^ n9145;
  assign n9795 = n9737 ^ n9655;
  assign n9794 = n9141 ^ n9140;
  assign n9796 = n9795 ^ n9794;
  assign n9687 = n9686 ^ n9682;
  assign n9679 = n9514 ^ n9503;
  assign n9688 = n9687 ^ n9679;
  assign n10783 = n9796 ^ n9688;
  assign n12520 = n12519 ^ n10783;
  assign n12523 = n12522 ^ n12520;
  assign n9146 = n9052 & n9132;
  assign n9147 = n9146 ^ n9145;
  assign n9152 = n9151 ^ n9147;
  assign n9144 = n9143 ^ n9140;
  assign n9153 = n9152 ^ n9144;
  assign n10786 = n9728 ^ n9153;
  assign n12524 = n12523 ^ n10786;
  assign n12529 = n12528 ^ n12524;
  assign n12542 = n12529 ^ n12517;
  assign n9830 = n9208 & n9262;
  assign n9831 = n9830 ^ n9693;
  assign n9828 = n9284 ^ n9253;
  assign n9747 = ~n9187 & ~n9251;
  assign n9664 = n9521 ^ n9271;
  assign n9748 = n9747 ^ n9664;
  assign n9829 = n9828 ^ n9748;
  assign n9832 = n9831 ^ n9829;
  assign n12503 = n12502 ^ n9832;
  assign n9846 = n9086 & n9129;
  assign n9847 = n9846 ^ n9736;
  assign n9844 = n9159 ^ n9139;
  assign n9739 = n9066 & n9135;
  assign n9656 = n9616 ^ n9146;
  assign n9740 = n9739 ^ n9656;
  assign n9845 = n9844 ^ n9740;
  assign n9848 = n9847 ^ n9845;
  assign n9823 = n9435 & n9511;
  assign n9824 = n9823 ^ n9685;
  assign n9821 = n9633 ^ n9510;
  assign n9822 = n9821 ^ n9788;
  assign n9825 = n9824 ^ n9822;
  assign n10773 = n9848 ^ n9825;
  assign n9388 = n9387 ^ n9378;
  assign n9401 = n9400 ^ n9388;
  assign n9519 = n9518 ^ n9401;
  assign n12501 = n10773 ^ n9519;
  assign n12504 = n12503 ^ n12501;
  assign n9622 = n9267 ^ n9265;
  assign n9621 = n9522 ^ n9285;
  assign n9623 = n9622 ^ n9621;
  assign n12499 = n12498 ^ n9623;
  assign n9619 = n9142 ^ n9140;
  assign n9618 = n9617 ^ n9160;
  assign n9620 = n9619 ^ n9618;
  assign n10765 = n9852 ^ n9620;
  assign n9818 = n9307 & ~n9394;
  assign n9819 = n9818 ^ n9672;
  assign n9816 = n9627 ^ n9398;
  assign n9817 = n9816 ^ n9783;
  assign n9820 = n9819 ^ n9817;
  assign n9826 = n9825 ^ n9820;
  assign n12497 = n10765 ^ n9826;
  assign n12500 = n12499 ^ n12497;
  assign n12505 = n12504 ^ n12500;
  assign n12543 = n12542 ^ n12505;
  assign n9749 = ~n9186 & n9247;
  assign n9750 = n9749 ^ n9268;
  assign n9751 = n9750 ^ n9748;
  assign n9746 = n9694 ^ n9281;
  assign n9752 = n9751 ^ n9746;
  assign n12532 = n12531 ^ n9752;
  assign n9741 = n9061 & n9132;
  assign n9742 = n9741 ^ n9143;
  assign n9743 = n9742 ^ n9740;
  assign n9738 = n9737 ^ n9156;
  assign n9744 = n9743 ^ n9738;
  assign n10821 = n9792 ^ n9744;
  assign n9677 = n9676 ^ n9673;
  assign n9669 = n9399 ^ n9371;
  assign n9678 = n9677 ^ n9669;
  assign n9689 = n9688 ^ n9678;
  assign n12530 = n10821 ^ n9689;
  assign n12533 = n12532 ^ n12530;
  assign n12541 = n12533 ^ n12516;
  assign n12568 = n12543 ^ n12541;
  assign n9665 = n9664 ^ n9663;
  assign n9661 = n9660 ^ n9281;
  assign n9666 = n9665 ^ n9661;
  assign n12495 = n12494 ^ n9666;
  assign n9657 = n9656 ^ n9655;
  assign n9653 = n9652 ^ n9156;
  assign n9658 = n9657 ^ n9653;
  assign n10838 = n9762 ^ n9658;
  assign n9637 = n9636 ^ n9630;
  assign n12493 = n10838 ^ n9637;
  assign n12496 = n12495 ^ n12493;
  assign n12506 = n12505 ^ n12496;
  assign n12512 = n12511 ^ n12506;
  assign n12566 = n12496 & n12512;
  assign n12552 = n12533 ^ n12511;
  assign n12538 = n12523 ^ n12516;
  assign n12553 = n12552 ^ n12538;
  assign n12554 = n12542 & ~n12553;
  assign n12567 = n12566 ^ n12554;
  assign n12569 = n12568 ^ n12567;
  assign n12545 = n12533 ^ n12500;
  assign n12546 = n12545 ^ n12529;
  assign n12547 = n12517 & ~n12546;
  assign n12544 = ~n12541 & n12543;
  assign n12548 = n12547 ^ n12544;
  assign n12570 = n12569 ^ n12548;
  assign n12534 = n12533 ^ n12504;
  assign n12561 = n12534 ^ n12517;
  assign n12562 = ~n12552 & ~n12561;
  assign n12563 = n12562 ^ n12547;
  assign n12560 = n12545 ^ n12542;
  assign n12564 = n12563 ^ n12560;
  assign n12555 = n12523 ^ n12506;
  assign n12556 = n12555 ^ n12541;
  assign n12557 = n12542 ^ n12496;
  assign n12558 = ~n12556 & n12557;
  assign n12559 = n12558 ^ n12554;
  assign n12565 = n12564 ^ n12559;
  assign n12579 = n12570 ^ n12565;
  assign n12575 = n12506 & ~n12523;
  assign n12535 = n12534 ^ n12529;
  assign n12539 = ~n12535 & n12538;
  assign n12576 = n12575 ^ n12539;
  assign n12573 = n12538 ^ n12535;
  assign n12574 = n12573 ^ n12563;
  assign n12577 = n12576 ^ n12574;
  assign n12578 = ~n12565 & ~n12577;
  assign n12536 = n12535 ^ n12506;
  assign n12518 = n12517 ^ n12512;
  assign n12550 = n12536 ^ n12518;
  assign n12537 = n12518 & ~n12536;
  assign n12540 = n12539 ^ n12537;
  assign n12549 = n12548 ^ n12540;
  assign n12551 = n12550 ^ n12549;
  assign n12594 = n12578 ^ n12551;
  assign n12595 = n12579 & ~n12594;
  assign n12596 = n12595 ^ n12570;
  assign n12583 = n12577 ^ n12551;
  assign n12591 = n12578 ^ n12570;
  assign n12592 = n12583 & ~n12591;
  assign n12593 = n12592 ^ n12551;
  assign n12597 = n12596 ^ n12593;
  assign n12600 = n12517 & n12597;
  assign n12585 = ~n12570 & ~n12577;
  assign n12586 = n12551 & n12585;
  assign n12584 = n12583 ^ n12578;
  assign n12587 = n12586 ^ n12584;
  assign n12580 = n12579 ^ n12578;
  assign n12571 = ~n12565 & n12570;
  assign n12572 = ~n12551 & n12571;
  assign n12581 = n12580 ^ n12572;
  assign n12590 = n12587 ^ n12581;
  assign n12598 = n12597 ^ n12590;
  assign n12599 = ~n12552 & n12598;
  assign n12601 = n12600 ^ n12599;
  assign n12588 = ~n12556 & n12587;
  assign n12971 = n12601 ^ n12588;
  assign n12606 = n12593 ^ n12587;
  assign n12622 = n12542 & ~n12606;
  assign n12608 = n12557 & n12587;
  assign n12607 = ~n12553 & ~n12606;
  assign n12609 = n12608 ^ n12607;
  assign n12623 = n12622 ^ n12609;
  assign n12617 = ~n12546 & n12597;
  assign n12616 = ~n12561 & n12598;
  assign n12618 = n12617 ^ n12616;
  assign n12970 = n12623 ^ n12618;
  assign n12972 = n12971 ^ n12970;
  assign n12582 = n12506 & n12581;
  assign n12589 = n12588 ^ n12582;
  assign n12619 = n12618 ^ n12589;
  assign n12612 = n12596 ^ n12581;
  assign n12613 = ~n12535 & ~n12612;
  assign n12614 = n12613 ^ n12601;
  assign n12615 = n12614 ^ n12607;
  assign n12620 = n12619 ^ n12615;
  assign n12973 = n12972 ^ n12620;
  assign n8160 = n8159 ^ n4580;
  assign n8161 = n8160 ^ n7451;
  assign n4186 = n4185 ^ n4179;
  assign n8158 = n8157 ^ n4186;
  assign n8162 = n8161 ^ n8158;
  assign n8120 = n4746 ^ n4687;
  assign n8122 = n8121 ^ n8120;
  assign n8119 = n8118 ^ n4639;
  assign n8123 = n8122 ^ n8119;
  assign n8174 = n8162 ^ n8123;
  assign n8151 = n4782 ^ n4580;
  assign n8152 = n8151 ^ n7454;
  assign n8150 = n8149 ^ n4075;
  assign n8153 = n8152 ^ n8150;
  assign n8193 = n8153 ^ n8123;
  assign n8168 = n4804 ^ n4606;
  assign n8170 = n8169 ^ n8168;
  assign n8167 = n8166 ^ n4610;
  assign n8171 = n8170 ^ n8167;
  assign n8172 = n8171 ^ n8162;
  assign n8194 = n8193 ^ n8172;
  assign n8195 = n8174 & n8194;
  assign n8138 = n8137 ^ n4716;
  assign n4699 = n4698 ^ n4185;
  assign n8136 = n8135 ^ n4699;
  assign n8139 = n8138 ^ n8136;
  assign n8129 = n8128 ^ n4687;
  assign n8130 = n8129 ^ n7434;
  assign n4658 = n4657 ^ n4185;
  assign n8127 = n8126 ^ n4658;
  assign n8131 = n8130 ^ n8127;
  assign n8133 = n8132 ^ n8131;
  assign n8140 = n8139 ^ n8133;
  assign n8114 = n4804 ^ n4782;
  assign n8115 = n8114 ^ n7428;
  assign n8113 = n8112 ^ n4767;
  assign n8116 = n8115 ^ n8113;
  assign n8124 = n8123 ^ n8116;
  assign n8141 = n8140 ^ n8124;
  assign n8184 = n8141 & n8172;
  assign n8196 = n8195 ^ n8184;
  assign n8173 = n8172 ^ n8140;
  assign n8192 = n8173 ^ n8124;
  assign n8197 = n8196 ^ n8192;
  assign n8154 = n8153 ^ n8116;
  assign n8146 = n8145 ^ n8128;
  assign n8144 = n8143 ^ n4185;
  assign n8147 = n8146 ^ n8144;
  assign n8155 = n8154 ^ n8147;
  assign n8187 = n8155 ^ n8131;
  assign n8180 = n8171 ^ n8123;
  assign n8188 = n8187 ^ n8180;
  assign n8189 = n8173 ^ n8147;
  assign n8190 = n8188 & n8189;
  assign n8175 = n8171 ^ n8131;
  assign n8176 = n8175 ^ n8174;
  assign n8177 = n8173 & n8176;
  assign n8191 = n8190 ^ n8177;
  assign n8198 = n8197 ^ n8191;
  assign n8204 = ~n8131 & n8155;
  assign n8200 = n8193 ^ n8140;
  assign n8203 = n8175 & n8200;
  assign n8205 = n8204 ^ n8203;
  assign n8201 = n8200 ^ n8175;
  assign n8202 = n8201 ^ n8196;
  assign n8206 = n8205 ^ n8202;
  assign n8207 = n8198 & n8206;
  assign n8179 = n8173 ^ n8154;
  assign n8183 = n8179 & n8180;
  assign n8185 = n8184 ^ n8183;
  assign n8181 = n8180 ^ n8179;
  assign n8163 = n8162 ^ n8155;
  assign n8164 = n8147 & n8163;
  assign n8178 = n8177 ^ n8164;
  assign n8182 = n8181 ^ n8178;
  assign n8186 = n8185 ^ n8182;
  assign n8199 = n8198 ^ n8186;
  assign n8239 = n8207 ^ n8199;
  assign n8209 = n8172 ^ n8163;
  assign n8208 = n8200 ^ n8155;
  assign n8213 = n8209 ^ n8208;
  assign n8210 = n8208 & n8209;
  assign n8211 = n8210 ^ n8203;
  assign n8212 = n8211 ^ n8185;
  assign n8214 = n8213 ^ n8212;
  assign n8237 = ~n8186 & n8198;
  assign n8238 = n8214 & n8237;
  assign n8240 = n8239 ^ n8238;
  assign n8218 = n8214 ^ n8206;
  assign n8228 = n8218 ^ n8207;
  assign n8226 = n8186 & n8206;
  assign n8227 = ~n8214 & n8226;
  assign n8229 = n8228 ^ n8227;
  assign n8241 = n8240 ^ n8229;
  assign n8219 = n8207 ^ n8186;
  assign n8220 = n8218 & n8219;
  assign n8221 = n8220 ^ n8214;
  assign n8215 = n8214 ^ n8207;
  assign n8216 = n8199 & n8215;
  assign n8217 = n8216 ^ n8186;
  assign n8222 = n8221 ^ n8217;
  assign n8724 = n8241 ^ n8222;
  assign n8725 = n8174 & n8724;
  assign n8224 = n8172 & n8222;
  assign n8726 = n8725 ^ n8224;
  assign n8719 = n8188 & n8229;
  assign n8873 = n8726 ^ n8719;
  assign n8782 = n8194 & n8724;
  assign n8223 = n8141 & n8222;
  assign n8783 = n8782 ^ n8223;
  assign n8230 = n8229 ^ n8221;
  assign n8716 = n8176 & n8230;
  assign n8715 = n8189 & n8229;
  assign n8717 = n8716 ^ n8715;
  assign n8231 = n8173 & n8230;
  assign n8718 = n8717 ^ n8231;
  assign n8872 = n8783 ^ n8718;
  assign n8874 = n8873 ^ n8872;
  assign n12410 = n8874 ^ n8017;
  assign n3827 = n3826 ^ n3664;
  assign n8625 = n7573 ^ n3827;
  assign n8624 = n4799 ^ n3649;
  assign n8626 = n8625 ^ n8624;
  assign n8622 = n4775 ^ n3826;
  assign n3803 = n3802 ^ n3800;
  assign n8621 = n7598 ^ n3803;
  assign n8623 = n8622 ^ n8621;
  assign n8627 = n8626 ^ n8623;
  assign n8612 = n3810 ^ n3771;
  assign n3773 = n3739 ^ n2697;
  assign n8611 = n8610 ^ n3773;
  assign n8613 = n8612 ^ n8611;
  assign n8608 = n4628 ^ n3707;
  assign n8606 = n4651 ^ n3750;
  assign n3743 = n3742 ^ n3739;
  assign n8604 = n8603 ^ n3743;
  assign n8605 = n8604 ^ n7607;
  assign n8607 = n8606 ^ n8605;
  assign n8609 = n8608 ^ n8607;
  assign n8614 = n8613 ^ n8609;
  assign n3659 = n3658 ^ n3649;
  assign n8600 = n7586 ^ n3659;
  assign n8599 = n4592 ^ n3854;
  assign n8601 = n8600 ^ n8599;
  assign n8597 = n4171 ^ n3802;
  assign n3798 = n3777 ^ n3739;
  assign n8595 = n8594 ^ n3798;
  assign n8596 = n8595 ^ n7593;
  assign n8598 = n8597 ^ n8596;
  assign n8602 = n8601 ^ n8598;
  assign n8615 = n8614 ^ n8602;
  assign n8628 = n8627 ^ n8615;
  assign n8631 = n3750 ^ n1051;
  assign n8630 = n3766 ^ n3518;
  assign n8632 = n8631 ^ n8630;
  assign n8629 = n4736 ^ n2681;
  assign n8633 = n8632 ^ n8629;
  assign n8643 = n8633 ^ n8623;
  assign n8644 = n8643 ^ n8614;
  assign n8616 = n8603 ^ n3739;
  assign n8617 = n8616 ^ n3728;
  assign n8618 = n8617 ^ n3794;
  assign n8619 = n8618 ^ n4840;
  assign n8640 = n8627 ^ n8619;
  assign n8645 = n8644 ^ n8640;
  assign n8641 = n8640 ^ n8598;
  assign n8642 = n8641 ^ n8602;
  assign n8651 = n8645 ^ n8642;
  assign n8647 = n8607 ^ n8601;
  assign n8648 = n8644 & ~n8647;
  assign n8646 = ~n8642 & ~n8645;
  assign n8649 = n8648 ^ n8646;
  assign n8636 = n8633 ^ n8626;
  assign n8637 = n8636 ^ n8614;
  assign n8638 = n8602 & n8637;
  assign n8634 = n8633 ^ n8601;
  assign n8635 = ~n8628 & n8634;
  assign n8639 = n8638 ^ n8635;
  assign n8650 = n8649 ^ n8639;
  assign n8652 = n8651 ^ n8650;
  assign n8666 = n8634 ^ n8628;
  assign n8653 = n8633 ^ n8598;
  assign n8663 = n8653 ^ n8647;
  assign n8664 = ~n8615 & ~n8663;
  assign n8662 = ~n8619 & ~n8641;
  assign n8665 = n8664 ^ n8662;
  assign n8667 = n8666 ^ n8665;
  assign n8668 = n8667 ^ n8639;
  assign n8675 = n8636 ^ n8615;
  assign n8654 = n8643 ^ n8602;
  assign n8655 = n8653 & ~n8654;
  assign n8656 = n8655 ^ n8638;
  assign n8676 = n8675 ^ n8656;
  assign n8620 = n8619 ^ n8615;
  assign n8671 = n8640 ^ n8607;
  assign n8672 = n8671 ^ n8634;
  assign n8673 = n8620 & n8672;
  assign n8674 = n8673 ^ n8664;
  assign n8677 = n8676 ^ n8674;
  assign n8693 = n8668 & n8677;
  assign n8694 = n8652 & n8693;
  assign n8691 = n8677 ^ n8668;
  assign n8659 = n8607 & ~n8640;
  assign n8660 = n8659 ^ n8648;
  assign n8657 = n8647 ^ n8644;
  assign n8658 = n8657 ^ n8656;
  assign n8661 = n8660 ^ n8658;
  assign n8678 = ~n8661 & n8677;
  assign n8692 = n8691 ^ n8678;
  assign n8695 = n8694 ^ n8692;
  assign n8679 = n8661 ^ n8652;
  assign n8680 = n8679 ^ n8678;
  assign n8669 = ~n8661 & ~n8668;
  assign n8670 = ~n8652 & n8669;
  assign n8681 = n8680 ^ n8670;
  assign n8696 = n8695 ^ n8681;
  assign n8773 = ~n8628 & n8696;
  assign n8697 = n8678 ^ n8652;
  assign n8698 = ~n8691 & n8697;
  assign n8699 = n8698 ^ n8668;
  assign n8771 = n8699 ^ n8695;
  assign n8772 = ~n8647 & n8771;
  assign n8774 = n8773 ^ n8772;
  assign n8770 = n8634 & n8696;
  assign n8775 = n8774 ^ n8770;
  assign n8767 = ~n8642 & ~n8699;
  assign n8683 = n8678 ^ n8668;
  assign n8684 = ~n8679 & ~n8683;
  assign n8685 = n8684 ^ n8652;
  assign n8765 = ~n8619 & n8685;
  assign n8686 = n8685 ^ n8681;
  assign n8689 = ~n8615 & ~n8686;
  assign n8766 = n8765 ^ n8689;
  assign n8768 = n8767 ^ n8766;
  assign n8700 = n8699 ^ n8685;
  assign n8706 = n8602 & ~n8700;
  assign n8703 = n8637 & ~n8700;
  assign n8764 = n8706 ^ n8703;
  assign n8769 = n8768 ^ n8764;
  assign n8776 = n8775 ^ n8769;
  assign n8508 = n8507 ^ n5572;
  assign n8509 = n8508 ^ n5680;
  assign n8510 = n8509 ^ n3699;
  assign n8504 = n8503 ^ n5373;
  assign n8505 = n8504 ^ n5702;
  assign n8506 = n8505 ^ n3845;
  assign n8511 = n8510 ^ n8506;
  assign n5751 = n5665 ^ n5597;
  assign n8499 = n5751 ^ n5697;
  assign n8498 = n8497 ^ n5737;
  assign n8500 = n8499 ^ n8498;
  assign n8495 = n5743 ^ n3714;
  assign n8493 = n5726 ^ n3757;
  assign n5713 = n5609 ^ n5597;
  assign n8491 = n5713 ^ n5651;
  assign n8490 = n8489 ^ n5721;
  assign n8492 = n8491 ^ n8490;
  assign n8494 = n8493 ^ n8492;
  assign n8496 = n8495 ^ n8494;
  assign n8501 = n8500 ^ n8496;
  assign n8485 = n5671 ^ n3859;
  assign n8483 = n5602 ^ n5387;
  assign n8482 = n5684 ^ n5505;
  assign n8484 = n8483 ^ n8482;
  assign n8486 = n8485 ^ n8484;
  assign n8473 = n8472 ^ n8471;
  assign n5693 = n5692 ^ n5597;
  assign n8474 = n8473 ^ n5693;
  assign n8475 = n8474 ^ n5557;
  assign n8476 = n8475 ^ n3819;
  assign n8488 = n8486 ^ n8476;
  assign n8502 = n8501 ^ n8488;
  assign n8512 = n8511 ^ n8502;
  assign n8520 = n5583 ^ n3789;
  assign n8518 = n5716 ^ n5597;
  assign n8519 = n8518 ^ n8489;
  assign n8521 = n8520 ^ n8519;
  assign n8522 = n8521 ^ n8511;
  assign n8558 = ~n8494 & n8522;
  assign n8477 = n5722 ^ n5629;
  assign n8478 = n8477 ^ n5660;
  assign n8479 = n8478 ^ n5756;
  assign n8480 = n8479 ^ n3638;
  assign n8525 = n8506 ^ n8480;
  assign n8526 = n8525 ^ n8501;
  assign n8529 = n8494 ^ n8486;
  assign n8530 = n8526 & n8529;
  assign n8559 = n8558 ^ n8530;
  assign n8556 = n8529 ^ n8526;
  assign n8481 = n8480 ^ n8476;
  assign n8536 = n8525 ^ n8488;
  assign n8537 = n8481 & n8536;
  assign n8514 = n8510 ^ n8480;
  assign n8515 = n8514 ^ n8501;
  assign n8516 = n8488 & n8515;
  assign n8538 = n8537 ^ n8516;
  assign n8557 = n8556 ^ n8538;
  assign n8560 = n8559 ^ n8557;
  assign n8527 = n8526 ^ n8522;
  assign n8523 = n8522 ^ n8476;
  assign n8524 = n8523 ^ n8488;
  assign n8533 = n8527 ^ n8524;
  assign n8528 = n8524 & n8527;
  assign n8531 = n8530 ^ n8528;
  assign n8487 = n8486 ^ n8480;
  assign n8513 = n8487 & n8512;
  assign n8517 = n8516 ^ n8513;
  assign n8532 = n8531 ^ n8517;
  assign n8534 = n8533 ^ n8532;
  assign n8566 = n8560 ^ n8534;
  assign n8544 = n8529 ^ n8481;
  assign n8545 = n8502 & n8544;
  assign n8540 = n8521 ^ n8502;
  assign n8541 = n8522 ^ n8494;
  assign n8542 = n8541 ^ n8487;
  assign n8543 = n8540 & n8542;
  assign n8546 = n8545 ^ n8543;
  assign n8535 = n8514 ^ n8502;
  assign n8539 = n8538 ^ n8535;
  assign n8547 = n8546 ^ n8539;
  assign n8561 = n8547 & n8560;
  assign n8567 = n8566 ^ n8561;
  assign n8550 = n8512 ^ n8487;
  assign n8548 = n8521 & n8523;
  assign n8549 = n8548 ^ n8545;
  assign n8551 = n8550 ^ n8549;
  assign n8552 = n8551 ^ n8517;
  assign n8564 = n8552 & n8560;
  assign n8565 = ~n8534 & n8564;
  assign n8568 = n8567 ^ n8565;
  assign n8555 = n8552 ^ n8547;
  assign n8562 = n8561 ^ n8555;
  assign n8553 = n8547 & ~n8552;
  assign n8554 = n8534 & n8553;
  assign n8563 = n8562 ^ n8554;
  assign n8569 = n8568 ^ n8563;
  assign n8760 = n8512 & n8569;
  assign n8570 = n8561 ^ n8534;
  assign n8571 = n8555 & n8570;
  assign n8572 = n8571 ^ n8552;
  assign n8758 = n8572 ^ n8563;
  assign n8759 = n8529 & n8758;
  assign n8761 = n8760 ^ n8759;
  assign n8757 = n8487 & n8569;
  assign n8762 = n8761 ^ n8757;
  assign n8573 = n8561 ^ n8552;
  assign n8574 = n8566 & n8573;
  assign n8575 = n8574 ^ n8534;
  assign n8753 = n8521 & n8575;
  assign n8584 = n8575 ^ n8568;
  assign n8587 = n8502 & n8584;
  assign n8754 = n8753 ^ n8587;
  assign n8752 = n8524 & n8572;
  assign n8755 = n8754 ^ n8752;
  assign n8576 = n8575 ^ n8572;
  assign n8590 = n8515 & n8576;
  assign n8579 = n8488 & n8576;
  assign n8751 = n8590 ^ n8579;
  assign n8756 = n8755 ^ n8751;
  assign n8763 = n8762 ^ n8756;
  assign n8777 = n8776 ^ n8763;
  assign n8353 = n6568 ^ n5708;
  assign n6431 = n6430 ^ n6401;
  assign n8351 = n8350 ^ n6431;
  assign n8352 = n8351 ^ n6454;
  assign n8354 = n8353 ^ n8352;
  assign n6634 = n6633 ^ n6628;
  assign n8344 = n7293 ^ n6634;
  assign n8343 = n6547 ^ n5638;
  assign n8345 = n8344 ^ n8343;
  assign n8397 = n8354 ^ n8345;
  assign n8359 = n6638 ^ n5730;
  assign n6402 = n6401 ^ n6391;
  assign n8357 = n8356 ^ n6402;
  assign n8358 = n8357 ^ n6525;
  assign n8360 = n8359 ^ n8358;
  assign n6473 = n6472 ^ n6466;
  assign n8347 = n7323 ^ n6473;
  assign n8346 = n5958 ^ n5675;
  assign n8348 = n8347 ^ n8346;
  assign n8391 = n8360 ^ n8348;
  assign n8398 = n8397 ^ n8391;
  assign n6279 = n6278 ^ n6162;
  assign n8382 = n7298 ^ n6279;
  assign n8381 = n6496 ^ n5592;
  assign n8383 = n8382 ^ n8381;
  assign n8372 = n6605 ^ n5535;
  assign n8371 = n7286 ^ n6598;
  assign n8373 = n8372 ^ n8371;
  assign n8369 = n7305 ^ n6618;
  assign n8368 = n6479 ^ n5135;
  assign n8370 = n8369 ^ n8368;
  assign n8374 = n8373 ^ n8370;
  assign n8384 = n8383 ^ n8374;
  assign n8421 = ~n8360 & n8384;
  assign n8387 = n8373 ^ n8345;
  assign n6562 = n6561 ^ n6401;
  assign n8364 = n8363 ^ n6562;
  assign n8362 = n6412 ^ n5748;
  assign n8365 = n8364 ^ n8362;
  assign n6536 = n6535 ^ n6531;
  assign n8361 = n8360 ^ n6536;
  assign n8366 = n8365 ^ n8361;
  assign n8388 = n8387 ^ n8366;
  assign n8392 = ~n8388 & n8391;
  assign n8422 = n8421 ^ n8392;
  assign n8419 = n8391 ^ n8388;
  assign n8355 = n8354 ^ n8348;
  assign n8406 = n8387 ^ n8355;
  assign n8407 = n8397 & ~n8406;
  assign n8377 = n8370 ^ n8345;
  assign n8378 = n8377 ^ n8366;
  assign n8379 = n8355 & ~n8378;
  assign n8408 = n8407 ^ n8379;
  assign n8420 = n8419 ^ n8408;
  assign n8423 = n8422 ^ n8420;
  assign n8389 = n8388 ^ n8384;
  assign n8385 = n8384 ^ n8354;
  assign n8386 = n8385 ^ n8355;
  assign n8395 = n8389 ^ n8386;
  assign n8390 = n8386 & ~n8389;
  assign n8393 = n8392 ^ n8390;
  assign n8349 = n8348 ^ n8345;
  assign n8367 = n8366 ^ n8355;
  assign n8375 = n8374 ^ n8367;
  assign n8376 = n8349 & n8375;
  assign n8380 = n8379 ^ n8376;
  assign n8394 = n8393 ^ n8380;
  assign n8396 = n8395 ^ n8394;
  assign n8427 = n8423 ^ n8396;
  assign n8405 = n8377 ^ n8367;
  assign n8409 = n8408 ^ n8405;
  assign n8400 = n8384 ^ n8360;
  assign n8401 = n8400 ^ n8349;
  assign n8402 = n8383 ^ n8367;
  assign n8403 = n8401 & n8402;
  assign n8399 = n8367 & n8398;
  assign n8404 = n8403 ^ n8399;
  assign n8410 = n8409 ^ n8404;
  assign n8424 = ~n8410 & ~n8423;
  assign n8413 = n8375 ^ n8349;
  assign n8411 = n8383 & n8385;
  assign n8412 = n8411 ^ n8399;
  assign n8414 = n8413 ^ n8412;
  assign n8415 = n8414 ^ n8380;
  assign n8442 = n8424 ^ n8415;
  assign n8443 = n8427 & n8442;
  assign n8444 = n8443 ^ n8396;
  assign n8429 = n8415 & ~n8423;
  assign n8430 = n8396 & n8429;
  assign n8428 = n8427 ^ n8424;
  assign n8431 = n8430 ^ n8428;
  assign n8449 = n8444 ^ n8431;
  assign n8465 = n8398 & ~n8449;
  assign n8464 = n8402 & n8431;
  assign n8466 = n8465 ^ n8464;
  assign n8450 = n8367 & ~n8449;
  assign n8467 = n8466 ^ n8450;
  assign n8418 = n8415 ^ n8410;
  assign n8434 = n8424 ^ n8396;
  assign n8435 = ~n8418 & ~n8434;
  assign n8436 = n8435 ^ n8415;
  assign n8445 = n8444 ^ n8436;
  assign n8425 = n8424 ^ n8418;
  assign n8416 = ~n8410 & ~n8415;
  assign n8417 = ~n8396 & n8416;
  assign n8426 = n8425 ^ n8417;
  assign n8432 = n8431 ^ n8426;
  assign n8457 = n8445 ^ n8432;
  assign n8462 = ~n8406 & n8457;
  assign n8446 = ~n8378 & ~n8445;
  assign n8463 = n8462 ^ n8446;
  assign n8468 = n8467 ^ n8463;
  assign n8460 = n8401 & n8431;
  assign n8458 = n8397 & n8457;
  assign n8447 = n8355 & ~n8445;
  assign n8459 = n8458 ^ n8447;
  assign n8461 = n8460 ^ n8459;
  assign n8469 = n8468 ^ n8461;
  assign n12408 = n8777 ^ n8469;
  assign n8709 = n8672 & ~n8681;
  assign n8701 = n8700 ^ n8696;
  assign n8707 = n8653 & ~n8701;
  assign n8708 = n8707 ^ n8706;
  assign n8710 = n8709 ^ n8708;
  assign n8702 = ~n8654 & ~n8701;
  assign n8704 = n8703 ^ n8702;
  assign n8687 = ~n8663 & ~n8686;
  assign n8682 = n8620 & ~n8681;
  assign n8688 = n8687 ^ n8682;
  assign n8690 = n8689 ^ n8688;
  assign n8705 = n8704 ^ n8690;
  assign n8711 = n8710 ^ n8705;
  assign n12409 = n12408 ^ n8711;
  assign n12411 = n12410 ^ n12409;
  assign n8944 = n8163 & n8221;
  assign n8720 = n8155 & n8240;
  assign n8721 = n8720 ^ n8719;
  assign n8945 = n8944 ^ n8721;
  assign n8234 = n8209 & n8217;
  assign n8232 = n8147 & n8221;
  assign n8233 = n8232 ^ n8231;
  assign n8235 = n8234 ^ n8233;
  assign n8946 = n8945 ^ n8235;
  assign n8245 = n8179 & n8241;
  assign n8243 = n8240 ^ n8217;
  assign n8244 = n8175 & n8243;
  assign n8246 = n8245 ^ n8244;
  assign n8830 = n8782 ^ n8246;
  assign n8723 = n8200 & n8243;
  assign n8727 = n8726 ^ n8723;
  assign n8943 = n8830 ^ n8727;
  assign n8947 = n8946 ^ n8943;
  assign n8853 = n8774 ^ n8702;
  assign n8800 = ~n8645 & ~n8699;
  assign n8799 = n8671 & ~n8695;
  assign n8801 = n8800 ^ n8799;
  assign n8919 = n8853 ^ n8801;
  assign n8856 = ~n8640 & ~n8695;
  assign n8918 = n8856 ^ n8708;
  assign n8920 = n8919 ^ n8918;
  assign n8577 = n8576 ^ n8569;
  assign n8589 = n8536 & n8577;
  assign n8861 = n8761 ^ n8589;
  assign n8808 = n8527 & n8572;
  assign n8807 = n8541 & n8563;
  assign n8809 = n8808 ^ n8807;
  assign n8916 = n8861 ^ n8809;
  assign n8864 = n8522 & n8563;
  assign n8578 = n8481 & n8577;
  assign n8580 = n8579 ^ n8578;
  assign n8915 = n8864 ^ n8580;
  assign n8917 = n8916 ^ n8915;
  assign n8921 = n8920 ^ n8917;
  assign n12400 = n8947 ^ n8921;
  assign n8857 = n8856 ^ n8709;
  assign n8855 = ~n8641 & n8685;
  assign n8858 = n8857 ^ n8855;
  assign n8859 = n8858 ^ n8768;
  assign n8796 = n8644 & n8771;
  assign n8797 = n8796 ^ n8708;
  assign n8854 = n8853 ^ n8797;
  assign n8860 = n8859 ^ n8854;
  assign n12401 = n12400 ^ n8860;
  assign n8845 = n8385 & ~n8444;
  assign n8744 = n8384 & ~n8426;
  assign n8745 = n8744 ^ n8460;
  assign n8846 = n8845 ^ n8745;
  assign n8453 = n8386 & n8436;
  assign n8451 = n8383 & ~n8444;
  assign n8452 = n8451 ^ n8450;
  assign n8454 = n8453 ^ n8452;
  assign n8847 = n8846 ^ n8454;
  assign n8439 = n8375 & ~n8432;
  assign n8437 = n8436 ^ n8426;
  assign n8438 = n8391 & ~n8437;
  assign n8440 = n8439 ^ n8438;
  assign n8843 = n8462 ^ n8440;
  assign n8747 = ~n8388 & ~n8437;
  assign n8748 = n8747 ^ n8459;
  assign n8844 = n8843 ^ n8748;
  assign n8848 = n8847 ^ n8844;
  assign n12402 = n12401 ^ n8848;
  assign n12403 = n12402 ^ n7912;
  assign n12415 = n12411 ^ n12403;
  assign n8581 = n8542 & n8568;
  assign n8865 = n8864 ^ n8581;
  assign n8591 = n8590 ^ n8589;
  assign n8885 = n8865 ^ n8591;
  assign n8804 = n8526 & n8758;
  assign n8805 = n8804 ^ n8580;
  assign n8585 = n8544 & n8584;
  assign n8884 = n8805 ^ n8585;
  assign n8886 = n8885 ^ n8884;
  assign n8863 = n8523 & n8575;
  assign n8866 = n8865 ^ n8863;
  assign n8867 = n8866 ^ n8755;
  assign n8862 = n8861 ^ n8805;
  assign n8868 = n8867 ^ n8862;
  assign n10406 = n8886 ^ n8868;
  assign n8818 = ~n8389 & n8436;
  assign n8892 = n8818 ^ n8451;
  assign n8893 = n8892 ^ n8466;
  assign n8891 = n8745 ^ n8459;
  assign n8894 = n8893 ^ n8891;
  assign n12391 = n10406 ^ n8894;
  assign n8882 = n8857 ^ n8704;
  assign n8881 = n8797 ^ n8687;
  assign n8883 = n8882 ^ n8881;
  assign n11797 = n8883 ^ n8860;
  assign n8938 = n8800 ^ n8765;
  assign n8939 = n8938 ^ n8688;
  assign n8937 = n8857 ^ n8708;
  assign n8940 = n8939 ^ n8937;
  assign n12390 = n11797 ^ n8940;
  assign n12392 = n12391 ^ n12390;
  assign n8828 = n8208 & n8217;
  assign n8827 = n8187 & n8240;
  assign n8829 = n8828 ^ n8827;
  assign n8831 = n8830 ^ n8829;
  assign n8826 = n8726 ^ n8720;
  assign n8832 = n8831 ^ n8826;
  assign n12387 = n8832 ^ n7959;
  assign n8810 = n8809 ^ n8754;
  assign n8806 = n8805 ^ n8759;
  assign n8811 = n8810 ^ n8806;
  assign n10372 = n8886 ^ n8811;
  assign n8817 = n8400 & ~n8426;
  assign n8819 = n8818 ^ n8817;
  assign n8850 = n8843 ^ n8819;
  assign n8849 = n8744 ^ n8459;
  assign n8851 = n8850 ^ n8849;
  assign n12385 = n10372 ^ n8851;
  assign n8802 = n8801 ^ n8766;
  assign n8798 = n8797 ^ n8772;
  assign n8803 = n8802 ^ n8798;
  assign n11791 = n8883 ^ n8803;
  assign n12384 = n11791 ^ n8920;
  assign n12386 = n12385 ^ n12384;
  assign n12388 = n12387 ^ n12386;
  assign n8904 = n8828 ^ n8232;
  assign n8905 = n8904 ^ n8717;
  assign n8903 = n8726 ^ n8721;
  assign n8906 = n8905 ^ n8903;
  assign n12383 = n8906 ^ n7927;
  assign n12389 = n12388 ^ n12383;
  assign n12393 = n12392 ^ n12389;
  assign n12416 = n12415 ^ n12393;
  assign n8814 = n8745 ^ n8463;
  assign n8813 = n8748 ^ n8465;
  assign n8815 = n8814 ^ n8813;
  assign n8583 = n8540 & n8568;
  assign n8586 = n8585 ^ n8583;
  assign n8588 = n8587 ^ n8586;
  assign n8592 = n8591 ^ n8588;
  assign n8582 = n8581 ^ n8580;
  assign n8593 = n8592 ^ n8582;
  assign n8712 = n8711 ^ n8593;
  assign n12379 = n8815 ^ n8712;
  assign n8784 = n8783 ^ n8721;
  assign n8781 = n8727 ^ n8716;
  assign n8785 = n8784 ^ n8781;
  assign n11819 = n8883 ^ n8785;
  assign n12380 = n12379 ^ n11819;
  assign n12381 = n12380 ^ n7807;
  assign n8899 = n8857 ^ n8690;
  assign n8900 = n8899 ^ n8797;
  assign n8722 = n8721 ^ n8718;
  assign n8728 = n8727 ^ n8722;
  assign n11803 = n8900 ^ n8728;
  assign n11773 = n8940 ^ n8883;
  assign n12375 = n11803 ^ n11773;
  assign n8934 = n8808 ^ n8753;
  assign n8935 = n8934 ^ n8586;
  assign n8933 = n8865 ^ n8580;
  assign n8936 = n8935 ^ n8933;
  assign n10378 = n8936 ^ n8886;
  assign n12376 = n12375 ^ n10378;
  assign n8746 = n8745 ^ n8467;
  assign n8749 = n8748 ^ n8746;
  assign n12377 = n12376 ^ n8749;
  assign n12378 = n12377 ^ n7774;
  assign n12382 = n12381 ^ n12378;
  assign n12394 = n12393 ^ n12382;
  assign n12454 = n12415 ^ n12394;
  assign n12432 = n12403 ^ n12378;
  assign n8242 = n8180 & n8241;
  assign n8247 = n8246 ^ n8242;
  assign n8225 = n8224 ^ n8223;
  assign n8236 = n8235 ^ n8225;
  assign n8248 = n8247 ^ n8236;
  assign n11807 = n8776 ^ n8248;
  assign n8448 = n8447 ^ n8446;
  assign n8455 = n8454 ^ n8448;
  assign n8433 = n8349 & ~n8432;
  assign n8441 = n8440 ^ n8433;
  assign n8456 = n8455 ^ n8441;
  assign n12405 = n11807 ^ n8456;
  assign n8897 = n8865 ^ n8588;
  assign n8898 = n8897 ^ n8805;
  assign n8901 = n8900 ^ n8898;
  assign n12406 = n12405 ^ n8901;
  assign n12407 = n12406 ^ n7866;
  assign n12422 = n12407 ^ n12403;
  assign n12433 = n12422 ^ n12382;
  assign n12434 = n12432 & n12433;
  assign n12417 = n12382 & n12416;
  assign n12435 = n12434 ^ n12417;
  assign n12455 = n12454 ^ n12435;
  assign n8924 = n8829 ^ n8233;
  assign n8923 = n8727 ^ n8244;
  assign n8925 = n8924 ^ n8923;
  assign n12397 = n8925 ^ n7994;
  assign n8820 = n8819 ^ n8452;
  assign n8816 = n8748 ^ n8438;
  assign n8821 = n8820 ^ n8816;
  assign n12395 = n8886 ^ n8821;
  assign n12396 = n12395 ^ n11791;
  assign n12398 = n12397 ^ n12396;
  assign n12399 = n12398 ^ n12394;
  assign n12412 = n12411 ^ n12407;
  assign n12419 = n12412 ^ n12398;
  assign n12450 = n12419 ^ n12388;
  assign n12404 = n12403 ^ n12381;
  assign n12451 = n12450 ^ n12404;
  assign n12452 = n12399 & n12451;
  assign n12426 = n12388 ^ n12381;
  assign n12442 = n12432 ^ n12426;
  assign n12443 = n12394 & n12442;
  assign n12453 = n12452 ^ n12443;
  assign n12456 = n12455 ^ n12453;
  assign n12413 = n12412 ^ n12394;
  assign n12445 = n12413 ^ n12404;
  assign n12420 = n12419 ^ n12378;
  assign n12441 = n12398 & n12420;
  assign n12444 = n12443 ^ n12441;
  assign n12446 = n12445 ^ n12444;
  assign n12414 = n12404 & n12413;
  assign n12418 = n12417 ^ n12414;
  assign n12447 = n12446 ^ n12418;
  assign n12472 = n12456 ^ n12447;
  assign n12438 = ~n12388 & n12419;
  assign n12423 = n12422 ^ n12393;
  assign n12427 = n12423 & n12426;
  assign n12439 = n12438 ^ n12427;
  assign n12436 = n12426 ^ n12423;
  assign n12437 = n12436 ^ n12435;
  assign n12440 = n12439 ^ n12437;
  assign n12457 = n12440 & n12456;
  assign n12424 = n12423 ^ n12419;
  assign n12421 = n12420 ^ n12382;
  assign n12430 = n12424 ^ n12421;
  assign n12425 = n12421 & n12424;
  assign n12428 = n12427 ^ n12425;
  assign n12429 = n12428 ^ n12418;
  assign n12431 = n12430 ^ n12429;
  assign n12480 = n12457 ^ n12431;
  assign n12481 = n12472 & n12480;
  assign n12482 = n12481 ^ n12447;
  assign n12458 = n12440 ^ n12431;
  assign n12462 = n12457 ^ n12447;
  assign n12463 = n12458 & n12462;
  assign n12464 = n12463 ^ n12431;
  assign n12483 = n12482 ^ n12464;
  assign n12965 = n12416 & n12483;
  assign n12473 = n12472 ^ n12457;
  assign n12470 = ~n12447 & n12456;
  assign n12471 = n12431 & n12470;
  assign n12474 = n12473 ^ n12471;
  assign n12459 = n12458 ^ n12457;
  assign n12448 = n12440 & n12447;
  assign n12449 = ~n12431 & n12448;
  assign n12460 = n12459 ^ n12449;
  assign n12479 = n12474 ^ n12460;
  assign n12484 = n12483 ^ n12479;
  assign n12861 = n12433 & n12484;
  assign n12966 = n12965 ^ n12861;
  assign n12476 = n12451 & n12460;
  assign n12475 = n12419 & n12474;
  assign n12477 = n12476 ^ n12475;
  assign n12967 = n12966 ^ n12477;
  assign n12488 = n12482 ^ n12474;
  assign n12489 = n12423 & n12488;
  assign n12486 = n12382 & n12483;
  assign n12485 = n12432 & n12484;
  assign n12487 = n12486 ^ n12485;
  assign n12490 = n12489 ^ n12487;
  assign n12465 = n12464 ^ n12460;
  assign n12466 = n12442 & n12465;
  assign n12964 = n12490 ^ n12466;
  assign n12968 = n12967 ^ n12964;
  assign n6645 = n6644 ^ n6638;
  assign n6623 = n6561 ^ n6511;
  assign n6635 = n6634 ^ n6623;
  assign n6646 = n6645 ^ n6635;
  assign n6583 = n6582 ^ n6434;
  assign n6599 = n6598 ^ n6583;
  assign n6577 = n6576 ^ n6568;
  assign n6600 = n6599 ^ n6577;
  assign n6656 = n6646 ^ n6600;
  assign n6487 = n6486 ^ n6479;
  assign n6460 = n6459 ^ n6401;
  assign n6474 = n6473 ^ n6460;
  assign n6488 = n6487 ^ n6474;
  assign n6435 = n6434 ^ n6431;
  assign n6455 = n6454 ^ n6435;
  assign n6424 = n6423 ^ n6413;
  assign n6456 = n6455 ^ n6424;
  assign n6489 = n6488 ^ n6456;
  assign n6667 = n6656 ^ n6489;
  assign n6563 = n6562 ^ n6430;
  assign n6554 = n6553 ^ n6548;
  assign n6564 = n6563 ^ n6554;
  assign n6512 = n6511 ^ n6402;
  assign n6526 = n6525 ^ n6512;
  assign n6505 = n6504 ^ n6497;
  assign n6527 = n6526 ^ n6505;
  assign n6537 = n6536 ^ n6527;
  assign n6565 = n6564 ^ n6537;
  assign n6657 = n6656 ^ n6565;
  assign n6611 = n6582 ^ n6459;
  assign n6619 = n6618 ^ n6611;
  assign n6610 = n6609 ^ n6605;
  assign n6620 = n6619 ^ n6610;
  assign n6621 = n6620 ^ n6600;
  assign n6403 = n6402 ^ n6279;
  assign n6045 = n6044 ^ n5958;
  assign n6404 = n6403 ^ n6045;
  assign n6653 = n6621 ^ n6404;
  assign n6658 = n6657 ^ n6653;
  assign n6654 = n6653 ^ n6456;
  assign n6655 = n6654 ^ n6489;
  assign n6664 = n6658 ^ n6655;
  assign n6660 = n6527 ^ n6488;
  assign n6661 = n6657 & ~n6660;
  assign n6659 = ~n6655 & ~n6658;
  assign n6662 = n6661 ^ n6659;
  assign n6649 = n6646 ^ n6620;
  assign n6650 = n6649 ^ n6565;
  assign n6651 = n6489 & n6650;
  assign n6566 = n6565 ^ n6489;
  assign n6622 = n6621 ^ n6566;
  assign n6647 = n6646 ^ n6488;
  assign n6648 = ~n6622 & n6647;
  assign n6652 = n6651 ^ n6648;
  assign n6663 = n6662 ^ n6652;
  assign n6665 = n6664 ^ n6663;
  assign n6680 = n6647 ^ n6622;
  assign n6666 = n6646 ^ n6456;
  assign n6677 = n6666 ^ n6660;
  assign n6678 = ~n6566 & ~n6677;
  assign n6676 = ~n6404 & ~n6654;
  assign n6679 = n6678 ^ n6676;
  assign n6681 = n6680 ^ n6679;
  assign n6682 = n6681 ^ n6652;
  assign n6685 = n6653 ^ n6527;
  assign n6686 = n6685 ^ n6647;
  assign n6687 = n6566 ^ n6404;
  assign n6688 = n6686 & n6687;
  assign n6689 = n6688 ^ n6678;
  assign n6683 = n6649 ^ n6566;
  assign n6668 = n6666 & ~n6667;
  assign n6669 = n6668 ^ n6651;
  assign n6684 = n6683 ^ n6669;
  assign n6690 = n6689 ^ n6684;
  assign n6715 = n6682 & n6690;
  assign n6716 = n6665 & n6715;
  assign n6703 = n6690 ^ n6682;
  assign n6672 = n6527 & ~n6653;
  assign n6673 = n6672 ^ n6661;
  assign n6670 = n6660 ^ n6657;
  assign n6671 = n6670 ^ n6669;
  assign n6674 = n6673 ^ n6671;
  assign n6691 = ~n6674 & n6690;
  assign n6714 = n6703 ^ n6691;
  assign n6717 = n6716 ^ n6714;
  assign n6675 = n6674 ^ n6665;
  assign n6698 = n6691 ^ n6675;
  assign n6696 = ~n6674 & ~n6682;
  assign n6697 = ~n6665 & n6696;
  assign n6699 = n6698 ^ n6697;
  assign n6718 = n6717 ^ n6699;
  assign n6704 = n6691 ^ n6665;
  assign n6705 = ~n6703 & n6704;
  assign n6706 = n6705 ^ n6682;
  assign n6692 = n6691 ^ n6682;
  assign n6693 = ~n6675 & ~n6692;
  assign n6694 = n6693 ^ n6665;
  assign n6709 = n6706 ^ n6694;
  assign n6856 = n6718 ^ n6709;
  assign n6865 = ~n6667 & ~n6856;
  assign n6711 = n6650 & ~n6709;
  assign n6866 = n6865 ^ n6711;
  assign n6862 = n6687 & ~n6699;
  assign n6700 = n6699 ^ n6694;
  assign n6861 = ~n6677 & ~n6700;
  assign n6863 = n6862 ^ n6861;
  assign n6701 = ~n6566 & ~n6700;
  assign n6864 = n6863 ^ n6701;
  assign n6867 = n6866 ^ n6864;
  assign n6859 = n6686 & ~n6699;
  assign n6857 = n6666 & ~n6856;
  assign n6710 = n6489 & ~n6709;
  assign n6858 = n6857 ^ n6710;
  assign n6860 = n6859 ^ n6858;
  assign n6868 = n6867 ^ n6860;
  assign n12293 = n9862 ^ n6868;
  assign n6723 = n6647 & n6718;
  assign n6720 = n6717 ^ n6706;
  assign n6721 = ~n6660 & n6720;
  assign n6719 = ~n6622 & n6718;
  assign n6722 = n6721 ^ n6719;
  assign n6724 = n6723 ^ n6722;
  assign n6712 = n6711 ^ n6710;
  assign n6707 = ~n6655 & ~n6706;
  assign n6695 = ~n6404 & n6694;
  assign n6702 = n6701 ^ n6695;
  assign n6708 = n6707 ^ n6702;
  assign n6713 = n6712 ^ n6708;
  assign n6725 = n6724 ^ n6713;
  assign n4759 = n4758 ^ n4639;
  assign n4755 = n4754 ^ n4746;
  assign n4760 = n4759 ^ n4755;
  assign n4738 = n4737 ^ n4698;
  assign n4761 = n4760 ^ n4738;
  assign n4617 = n4616 ^ n4607;
  assign n4594 = n4593 ^ n4185;
  assign n4618 = n4617 ^ n4594;
  assign n4762 = n4761 ^ n4618;
  assign n4815 = n4814 ^ n4808;
  assign n4801 = n4800 ^ n4610;
  assign n4816 = n4815 ^ n4801;
  assign n4820 = n4816 ^ n4761;
  assign n4722 = n4721 ^ n4716;
  assign n4711 = n4710 ^ n4699;
  assign n4723 = n4722 ^ n4711;
  assign n4667 = n4666 ^ n4658;
  assign n4689 = n4688 ^ n4667;
  assign n4653 = n4652 ^ n4639;
  assign n4690 = n4689 ^ n4653;
  assign n4630 = n4629 ^ n4179;
  assign n4691 = n4690 ^ n4630;
  assign n4724 = n4723 ^ n4691;
  assign n4323 = n4322 ^ n4186;
  assign n4582 = n4581 ^ n4323;
  assign n4173 = n4172 ^ n4075;
  assign n4583 = n4582 ^ n4173;
  assign n4619 = n4618 ^ n4583;
  assign n4725 = n4724 ^ n4619;
  assign n4876 = n4820 ^ n4725;
  assign n4854 = n4761 ^ n4583;
  assign n4792 = n4791 ^ n4788;
  assign n4777 = n4776 ^ n4767;
  assign n4793 = n4792 ^ n4777;
  assign n4824 = n4793 ^ n4761;
  assign n4855 = n4824 ^ n4619;
  assign n4856 = n4854 & n4855;
  assign n4821 = n4820 ^ n4724;
  assign n4822 = n4619 & n4821;
  assign n4857 = n4856 ^ n4822;
  assign n4877 = n4876 ^ n4857;
  assign n4826 = n4658 ^ n4321;
  assign n4830 = n4829 ^ n4826;
  assign n4834 = n4833 ^ n4830;
  assign n4842 = n4841 ^ n4834;
  assign n4871 = n4842 ^ n4725;
  assign n4817 = n4816 ^ n4793;
  assign n4843 = n4842 ^ n4817;
  assign n4872 = n4843 ^ n4690;
  assign n4873 = n4872 ^ n4762;
  assign n4874 = n4871 & n4873;
  assign n4848 = n4690 ^ n4618;
  assign n4865 = n4854 ^ n4848;
  assign n4866 = n4725 & n4865;
  assign n4875 = n4874 ^ n4866;
  assign n4878 = n4877 ^ n4875;
  assign n4818 = n4817 ^ n4725;
  assign n4868 = n4818 ^ n4762;
  assign n4845 = n4843 ^ n4583;
  assign n4864 = n4842 & n4845;
  assign n4867 = n4866 ^ n4864;
  assign n4869 = n4868 ^ n4867;
  assign n4819 = n4762 & n4818;
  assign n4823 = n4822 ^ n4819;
  assign n4870 = n4869 ^ n4823;
  assign n4891 = n4878 ^ n4870;
  assign n4860 = ~n4690 & n4843;
  assign n4825 = n4824 ^ n4724;
  assign n4849 = n4825 & n4848;
  assign n4861 = n4860 ^ n4849;
  assign n4858 = n4848 ^ n4825;
  assign n4859 = n4858 ^ n4857;
  assign n4862 = n4861 ^ n4859;
  assign n4879 = n4862 & n4878;
  assign n4904 = n4891 ^ n4879;
  assign n4846 = n4845 ^ n4619;
  assign n4844 = n4843 ^ n4825;
  assign n4852 = n4846 ^ n4844;
  assign n4847 = n4844 & n4846;
  assign n4850 = n4849 ^ n4847;
  assign n4851 = n4850 ^ n4823;
  assign n4853 = n4852 ^ n4851;
  assign n4902 = ~n4870 & n4878;
  assign n4903 = n4853 & n4902;
  assign n4905 = n4904 ^ n4903;
  assign n4863 = n4862 ^ n4853;
  assign n4885 = n4879 ^ n4863;
  assign n4883 = n4862 & n4870;
  assign n4884 = ~n4853 & n4883;
  assign n4886 = n4885 ^ n4884;
  assign n4908 = n4905 ^ n4886;
  assign n4911 = n4762 & n4908;
  assign n4909 = n4818 & n4908;
  assign n4892 = n4879 ^ n4853;
  assign n4893 = n4891 & n4892;
  assign n4894 = n4893 ^ n4870;
  assign n4906 = n4905 ^ n4894;
  assign n4907 = n4848 & n4906;
  assign n4910 = n4909 ^ n4907;
  assign n4912 = n4911 ^ n4910;
  assign n4880 = n4879 ^ n4870;
  assign n4881 = n4863 & n4880;
  assign n4882 = n4881 ^ n4853;
  assign n4897 = n4894 ^ n4882;
  assign n4899 = n4821 & n4897;
  assign n4898 = n4619 & n4897;
  assign n4900 = n4899 ^ n4898;
  assign n4895 = n4846 & n4894;
  assign n4889 = n4842 & n4882;
  assign n4887 = n4886 ^ n4882;
  assign n4888 = n4725 & n4887;
  assign n4890 = n4889 ^ n4888;
  assign n4896 = n4895 ^ n4890;
  assign n4901 = n4900 ^ n4896;
  assign n4913 = n4912 ^ n4901;
  assign n10487 = n6725 ^ n4913;
  assign n5710 = n5709 ^ n5705;
  assign n5699 = n5698 ^ n5693;
  assign n5703 = n5702 ^ n5699;
  assign n5711 = n5710 ^ n5703;
  assign n5686 = n5685 ^ n5681;
  assign n5677 = n5676 ^ n5671;
  assign n5687 = n5686 ^ n5677;
  assign n5712 = n5711 ^ n5687;
  assign n5758 = n5757 ^ n5751;
  assign n5750 = n5749 ^ n5743;
  assign n5759 = n5758 ^ n5750;
  assign n5732 = n5731 ^ n5726;
  assign n5718 = n5717 ^ n5713;
  assign n5723 = n5722 ^ n5718;
  assign n5733 = n5732 ^ n5723;
  assign n5739 = n5738 ^ n5733;
  assign n5760 = n5759 ^ n5739;
  assign n5761 = n5760 ^ n5712;
  assign n5573 = n5572 ^ n5558;
  assign n5537 = n5536 ^ n5521;
  assign n5574 = n5573 ^ n5537;
  assign n5507 = n5506 ^ n5374;
  assign n5137 = n5136 ^ n5050;
  assign n5508 = n5507 ^ n5137;
  assign n5575 = n5574 ^ n5508;
  assign n5762 = n5761 ^ n5575;
  assign n5667 = n5666 ^ n5652;
  assign n5640 = n5639 ^ n5629;
  assign n5668 = n5667 ^ n5640;
  assign n5688 = n5687 ^ n5668;
  assign n5796 = n5762 ^ n5688;
  assign n5619 = n5618 ^ n5603;
  assign n5594 = n5593 ^ n5583;
  assign n5620 = n5619 ^ n5594;
  assign n5621 = n5620 ^ n5575;
  assign n5768 = n5711 ^ n5621;
  assign n5794 = n5620 & n5768;
  assign n5784 = n5711 ^ n5668;
  assign n5774 = n5733 ^ n5687;
  assign n5785 = n5784 ^ n5774;
  assign n5786 = ~n5761 & ~n5785;
  assign n5795 = n5794 ^ n5786;
  assign n5797 = n5796 ^ n5795;
  assign n5764 = n5668 ^ n5508;
  assign n5765 = n5764 ^ n5760;
  assign n5766 = n5712 & ~n5765;
  assign n5763 = n5688 & ~n5762;
  assign n5767 = n5766 ^ n5763;
  assign n5798 = n5797 ^ n5767;
  assign n5770 = n5668 ^ n5574;
  assign n5789 = n5770 ^ n5712;
  assign n5790 = n5784 & n5789;
  assign n5791 = n5790 ^ n5766;
  assign n5788 = n5764 ^ n5761;
  assign n5792 = n5791 ^ n5788;
  assign n5780 = n5733 ^ n5621;
  assign n5781 = n5780 ^ n5688;
  assign n5782 = n5761 ^ n5620;
  assign n5783 = ~n5781 & ~n5782;
  assign n5787 = n5786 ^ n5783;
  assign n5793 = n5792 ^ n5787;
  assign n5801 = n5798 ^ n5793;
  assign n5771 = n5770 ^ n5760;
  assign n5804 = n5774 ^ n5771;
  assign n5805 = n5804 ^ n5791;
  assign n5802 = n5621 & n5733;
  assign n5775 = ~n5771 & ~n5774;
  assign n5803 = n5802 ^ n5775;
  assign n5806 = n5805 ^ n5803;
  assign n5807 = ~n5793 & n5806;
  assign n5772 = n5771 ^ n5621;
  assign n5769 = n5768 ^ n5712;
  assign n5778 = n5772 ^ n5769;
  assign n5773 = n5769 & ~n5772;
  assign n5776 = n5775 ^ n5773;
  assign n5777 = n5776 ^ n5767;
  assign n5779 = n5778 ^ n5777;
  assign n5828 = n5807 ^ n5779;
  assign n5829 = n5801 & ~n5828;
  assign n5830 = n5829 ^ n5798;
  assign n5813 = n5806 ^ n5779;
  assign n5818 = n5807 ^ n5798;
  assign n5819 = ~n5813 & ~n5818;
  assign n5820 = n5819 ^ n5779;
  assign n5834 = n5830 ^ n5820;
  assign n5837 = n5712 & n5834;
  assign n5814 = n5813 ^ n5807;
  assign n5811 = ~n5798 & n5806;
  assign n5812 = n5779 & n5811;
  assign n5815 = n5814 ^ n5812;
  assign n5808 = n5807 ^ n5801;
  assign n5799 = ~n5793 & n5798;
  assign n5800 = ~n5779 & n5799;
  assign n5809 = n5808 ^ n5800;
  assign n5833 = n5815 ^ n5809;
  assign n5835 = n5834 ^ n5833;
  assign n5836 = n5784 & ~n5835;
  assign n5838 = n5837 ^ n5836;
  assign n5816 = ~n5781 & ~n5815;
  assign n6940 = n5838 ^ n5816;
  assign n6903 = n5789 & ~n5835;
  assign n6841 = ~n5765 & n5834;
  assign n6904 = n6903 ^ n6841;
  assign n5821 = n5820 ^ n5815;
  assign n5825 = ~n5761 & n5821;
  assign n5823 = ~n5782 & ~n5815;
  assign n5822 = ~n5785 & n5821;
  assign n5824 = n5823 ^ n5822;
  assign n5826 = n5825 ^ n5824;
  assign n6939 = n6904 ^ n5826;
  assign n6941 = n6940 ^ n6939;
  assign n3804 = n3803 ^ n3798;
  assign n3812 = n3811 ^ n3804;
  assign n3815 = n3814 ^ n3812;
  assign n3821 = n3820 ^ n3815;
  assign n2682 = n2681 ^ n1870;
  assign n2698 = n2697 ^ n2682;
  assign n3519 = n3518 ^ n2698;
  assign n3640 = n3639 ^ n3519;
  assign n3874 = n3821 ^ n3640;
  assign n3833 = n3832 ^ n3827;
  assign n3838 = n3837 ^ n3833;
  assign n3847 = n3846 ^ n3838;
  assign n3893 = n3847 ^ n3640;
  assign n3778 = n3777 ^ n3773;
  assign n3772 = n3771 ^ n3767;
  assign n3779 = n3778 ^ n3772;
  assign n3759 = n3758 ^ n3750;
  assign n3744 = n3743 ^ n1051;
  assign n3736 = n3735 ^ n3729;
  assign n3745 = n3744 ^ n3736;
  assign n3760 = n3759 ^ n3745;
  assign n3716 = n3715 ^ n3707;
  assign n3761 = n3760 ^ n3716;
  assign n3780 = n3779 ^ n3761;
  assign n3900 = n3893 ^ n3780;
  assign n3678 = n3677 ^ n3659;
  assign n3688 = n3687 ^ n3678;
  assign n3701 = n3700 ^ n3688;
  assign n3848 = n3847 ^ n3701;
  assign n3795 = n3794 ^ n3725;
  assign n3796 = n3795 ^ n3743;
  assign n3791 = n3790 ^ n3784;
  assign n3797 = n3796 ^ n3791;
  assign n3849 = n3848 ^ n3797;
  assign n3909 = n3900 ^ n3849;
  assign n3869 = n3868 ^ n3865;
  assign n3870 = n3869 ^ n3739;
  assign n3861 = n3860 ^ n3854;
  assign n3871 = n3870 ^ n3861;
  assign n3872 = n3871 ^ n3821;
  assign n3850 = n3849 ^ n3821;
  assign n3908 = n3872 ^ n3850;
  assign n3913 = n3909 ^ n3908;
  assign n3910 = ~n3908 & ~n3909;
  assign n3875 = n3871 ^ n3760;
  assign n3903 = ~n3875 & n3900;
  assign n3911 = n3910 ^ n3903;
  assign n3702 = n3701 ^ n3640;
  assign n3781 = n3780 ^ n3702;
  assign n3884 = n3781 & n3872;
  assign n3873 = n3872 ^ n3780;
  assign n3879 = n3873 ^ n3848;
  assign n3880 = n3871 ^ n3640;
  assign n3883 = ~n3879 & n3880;
  assign n3885 = n3884 ^ n3883;
  assign n3912 = n3911 ^ n3885;
  assign n3914 = n3913 ^ n3912;
  assign n3881 = n3880 ^ n3879;
  assign n3876 = n3875 ^ n3874;
  assign n3877 = ~n3873 & ~n3876;
  assign n3851 = ~n3797 & ~n3850;
  assign n3878 = n3877 ^ n3851;
  assign n3882 = n3881 ^ n3878;
  assign n3886 = n3885 ^ n3882;
  assign n3894 = n3893 ^ n3872;
  assign n3895 = n3874 & ~n3894;
  assign n3896 = n3895 ^ n3884;
  assign n3892 = n3873 ^ n3702;
  assign n3897 = n3896 ^ n3892;
  assign n3887 = n3849 ^ n3760;
  assign n3888 = n3887 ^ n3880;
  assign n3889 = n3873 ^ n3797;
  assign n3890 = n3888 & n3889;
  assign n3891 = n3890 ^ n3877;
  assign n3898 = n3897 ^ n3891;
  assign n3938 = n3886 & n3898;
  assign n3939 = n3914 & n3938;
  assign n3904 = n3760 & ~n3849;
  assign n3905 = n3904 ^ n3903;
  assign n3901 = n3900 ^ n3875;
  assign n3902 = n3901 ^ n3896;
  assign n3906 = n3905 ^ n3902;
  assign n3907 = n3898 & ~n3906;
  assign n3899 = n3898 ^ n3886;
  assign n3937 = n3907 ^ n3899;
  assign n3940 = n3939 ^ n3937;
  assign n3918 = n3914 ^ n3906;
  assign n3929 = n3918 ^ n3907;
  assign n3927 = ~n3886 & ~n3906;
  assign n3928 = ~n3914 & n3927;
  assign n3930 = n3929 ^ n3928;
  assign n3941 = n3940 ^ n3930;
  assign n3919 = n3907 ^ n3886;
  assign n3920 = ~n3918 & ~n3919;
  assign n3921 = n3920 ^ n3914;
  assign n3915 = n3914 ^ n3907;
  assign n3916 = ~n3899 & n3915;
  assign n3917 = n3916 ^ n3886;
  assign n3922 = n3921 ^ n3917;
  assign n4924 = n3941 ^ n3922;
  assign n4925 = n3874 & ~n4924;
  assign n3924 = n3872 & ~n3922;
  assign n4926 = n4925 ^ n3924;
  assign n4916 = n3888 & ~n3930;
  assign n6838 = n4926 ^ n4916;
  assign n6835 = ~n3894 & ~n4924;
  assign n3923 = n3781 & ~n3922;
  assign n6836 = n6835 ^ n3923;
  assign n4919 = n3889 & ~n3930;
  assign n3931 = n3930 ^ n3921;
  assign n4918 = ~n3876 & ~n3931;
  assign n4920 = n4919 ^ n4918;
  assign n3932 = ~n3873 & ~n3931;
  assign n4921 = n4920 ^ n3932;
  assign n6837 = n6836 ^ n4921;
  assign n6839 = n6838 ^ n6837;
  assign n6942 = n6941 ^ n6839;
  assign n12292 = n10487 ^ n6942;
  assign n12294 = n12293 ^ n12292;
  assign n7009 = ~n6654 & n6694;
  assign n6945 = ~n6653 & ~n6717;
  assign n6946 = n6945 ^ n6859;
  assign n7010 = n7009 ^ n6946;
  assign n7011 = n7010 ^ n6708;
  assign n7007 = n6865 ^ n6722;
  assign n6912 = n6657 & n6720;
  assign n6913 = n6912 ^ n6858;
  assign n7008 = n7007 ^ n6913;
  assign n7012 = n7011 ^ n7008;
  assign n12286 = n9807 ^ n7012;
  assign n6916 = n6685 & ~n6717;
  assign n6915 = ~n6658 & ~n6706;
  assign n6917 = n6916 ^ n6915;
  assign n7036 = n7007 ^ n6917;
  assign n7035 = n6945 ^ n6858;
  assign n7037 = n7036 ^ n7035;
  assign n6826 = n4908 ^ n4897;
  assign n6827 = n4855 & n6826;
  assign n6983 = n6827 ^ n4910;
  assign n6897 = n4844 & n4894;
  assign n6896 = n4872 & n4905;
  assign n6898 = n6897 ^ n6896;
  assign n7031 = n6983 ^ n6898;
  assign n6934 = n4843 & n4905;
  assign n6831 = n4854 & n6826;
  assign n6832 = n6831 ^ n4898;
  assign n7030 = n6934 ^ n6832;
  assign n7032 = n7031 ^ n7030;
  assign n12284 = n7037 ^ n7032;
  assign n7052 = n5768 & ~n5820;
  assign n5810 = n5621 & n5809;
  assign n5817 = n5816 ^ n5810;
  assign n7053 = n7052 ^ n5817;
  assign n6845 = n5769 & ~n5830;
  assign n6843 = n5620 & ~n5820;
  assign n6844 = n6843 ^ n5825;
  assign n6846 = n6845 ^ n6844;
  assign n7054 = n7053 ^ n6846;
  assign n5831 = n5830 ^ n5809;
  assign n6850 = ~n5774 & ~n5831;
  assign n6849 = ~n5762 & ~n5833;
  assign n6851 = n6850 ^ n6849;
  assign n6999 = n6903 ^ n6851;
  assign n5832 = ~n5771 & ~n5831;
  assign n5839 = n5838 ^ n5832;
  assign n7051 = n6999 ^ n5839;
  assign n7055 = n7054 ^ n7051;
  assign n6991 = ~n3850 & n3921;
  assign n4915 = ~n3849 & ~n3940;
  assign n4917 = n4916 ^ n4915;
  assign n6992 = n6991 ^ n4917;
  assign n3934 = ~n3908 & ~n3917;
  assign n3926 = ~n3797 & n3921;
  assign n3933 = n3932 ^ n3926;
  assign n3935 = n3934 ^ n3933;
  assign n6993 = n6992 ^ n3935;
  assign n3944 = n3940 ^ n3917;
  assign n3945 = ~n3875 & n3944;
  assign n3943 = ~n3879 & n3941;
  assign n3946 = n3945 ^ n3943;
  assign n6989 = n6835 ^ n3946;
  assign n4923 = n3900 & n3944;
  assign n4927 = n4926 ^ n4923;
  assign n6990 = n6989 ^ n4927;
  assign n6994 = n6993 ^ n6990;
  assign n12283 = n7055 ^ n6994;
  assign n12285 = n12284 ^ n12283;
  assign n12287 = n12286 ^ n12285;
  assign n12298 = n12294 ^ n12287;
  assign n6947 = n6946 ^ n6866;
  assign n6944 = n6913 ^ n6861;
  assign n6948 = n6947 ^ n6944;
  assign n11351 = n7012 ^ n6948;
  assign n6985 = n4845 & n4882;
  assign n6830 = n4873 & n4886;
  assign n6935 = n6934 ^ n6830;
  assign n6986 = n6985 ^ n6935;
  assign n6987 = n6986 ^ n4896;
  assign n6893 = n4825 & n4906;
  assign n6894 = n6893 ^ n6832;
  assign n6984 = n6983 ^ n6894;
  assign n6988 = n6987 ^ n6984;
  assign n6828 = n6827 ^ n4899;
  assign n6936 = n6935 ^ n6828;
  assign n6823 = n4865 & n4887;
  assign n6933 = n6894 ^ n6823;
  assign n6937 = n6936 ^ n6933;
  assign n10524 = n6988 ^ n6937;
  assign n12274 = n11351 ^ n10524;
  assign n6889 = ~n3909 & ~n3917;
  assign n6965 = n6889 ^ n3926;
  assign n6966 = n6965 ^ n4920;
  assign n6964 = n4926 ^ n4917;
  assign n6967 = n6966 ^ n6964;
  assign n6959 = ~n5772 & ~n5830;
  assign n6960 = n6959 ^ n6843;
  assign n6961 = n6960 ^ n5824;
  assign n6958 = n5838 ^ n5817;
  assign n6962 = n6961 ^ n6958;
  assign n12273 = n6967 ^ n6962;
  assign n12275 = n12274 ^ n12273;
  assign n7060 = n6915 ^ n6695;
  assign n7061 = n7060 ^ n6863;
  assign n7059 = n6946 ^ n6858;
  assign n7062 = n7061 ^ n7059;
  assign n12271 = n9719 ^ n7062;
  assign n12269 = n9708 ^ n7037;
  assign n6918 = n6917 ^ n6702;
  assign n6914 = n6913 ^ n6721;
  assign n6919 = n6918 ^ n6914;
  assign n11346 = n6948 ^ n6919;
  assign n6899 = n6898 ^ n4890;
  assign n6895 = n6894 ^ n4907;
  assign n6900 = n6899 ^ n6895;
  assign n10497 = n6937 ^ n6900;
  assign n12267 = n11346 ^ n10497;
  assign n6888 = n3887 & ~n3940;
  assign n6890 = n6889 ^ n6888;
  assign n7003 = n6989 ^ n6890;
  assign n7002 = n4926 ^ n4915;
  assign n7004 = n7003 ^ n7002;
  assign n6997 = ~n5780 & n5809;
  assign n6998 = n6997 ^ n6959;
  assign n7000 = n6999 ^ n6998;
  assign n6996 = n5838 ^ n5810;
  assign n7001 = n7000 ^ n6996;
  assign n7005 = n7004 ^ n7001;
  assign n12268 = n12267 ^ n7005;
  assign n12270 = n12269 ^ n12268;
  assign n12272 = n12271 ^ n12270;
  assign n12276 = n12275 ^ n12272;
  assign n12299 = n12298 ^ n12276;
  assign n12264 = n9646 ^ n6948;
  assign n6833 = n6832 ^ n6830;
  assign n6822 = n4871 & n4886;
  assign n6824 = n6823 ^ n6822;
  assign n6825 = n6824 ^ n4888;
  assign n6829 = n6828 ^ n6825;
  assign n6834 = n6833 ^ n6829;
  assign n10491 = n6868 ^ n6834;
  assign n6908 = n6836 ^ n4917;
  assign n6907 = n4927 ^ n4918;
  assign n6909 = n6908 ^ n6907;
  assign n6905 = n6904 ^ n5817;
  assign n6902 = n5839 ^ n5822;
  assign n6906 = n6905 ^ n6902;
  assign n6910 = n6909 ^ n6906;
  assign n12263 = n10491 ^ n6910;
  assign n12265 = n12264 ^ n12263;
  assign n6974 = n6946 ^ n6864;
  assign n6975 = n6974 ^ n6913;
  assign n12261 = n9611 ^ n6975;
  assign n11334 = n7062 ^ n6948;
  assign n7046 = n6897 ^ n4889;
  assign n7047 = n7046 ^ n6824;
  assign n7045 = n6935 ^ n6832;
  assign n7048 = n7047 ^ n7045;
  assign n10502 = n7048 ^ n6937;
  assign n12259 = n11334 ^ n10502;
  assign n5827 = n5826 ^ n5817;
  assign n5840 = n5839 ^ n5827;
  assign n4922 = n4921 ^ n4917;
  assign n4928 = n4927 ^ n4922;
  assign n5841 = n5840 ^ n4928;
  assign n12260 = n12259 ^ n5841;
  assign n12262 = n12261 ^ n12260;
  assign n12266 = n12265 ^ n12262;
  assign n12277 = n12276 ^ n12266;
  assign n12337 = n12298 ^ n12277;
  assign n12315 = n12287 ^ n12262;
  assign n12290 = n9839 ^ n6725;
  assign n6970 = n6935 ^ n6825;
  assign n6971 = n6970 ^ n6894;
  assign n10503 = n6975 ^ n6971;
  assign n6848 = n5688 & ~n5833;
  assign n6852 = n6851 ^ n6848;
  assign n6842 = n6841 ^ n5837;
  assign n6847 = n6846 ^ n6842;
  assign n6853 = n6852 ^ n6847;
  assign n3942 = n3880 & n3941;
  assign n3947 = n3946 ^ n3942;
  assign n3925 = n3924 ^ n3923;
  assign n3936 = n3935 ^ n3925;
  assign n3948 = n3947 ^ n3936;
  assign n6854 = n6853 ^ n3948;
  assign n12289 = n10503 ^ n6854;
  assign n12291 = n12290 ^ n12289;
  assign n12305 = n12291 ^ n12287;
  assign n12316 = n12305 ^ n12266;
  assign n12317 = n12315 & ~n12316;
  assign n12300 = n12266 & n12299;
  assign n12318 = n12317 ^ n12300;
  assign n12338 = n12337 ^ n12318;
  assign n12278 = n11346 ^ n6937;
  assign n6891 = n6890 ^ n3933;
  assign n6887 = n4927 ^ n3945;
  assign n6892 = n6891 ^ n6887;
  assign n12279 = n12278 ^ n6892;
  assign n7025 = n6998 ^ n6844;
  assign n7024 = n6850 ^ n5839;
  assign n7026 = n7025 ^ n7024;
  assign n12280 = n12279 ^ n7026;
  assign n12281 = n12280 ^ n9774;
  assign n12282 = n12281 ^ n12277;
  assign n12295 = n12294 ^ n12291;
  assign n12302 = n12295 ^ n12281;
  assign n12333 = n12302 ^ n12270;
  assign n12288 = n12287 ^ n12265;
  assign n12334 = n12333 ^ n12288;
  assign n12335 = n12282 & n12334;
  assign n12309 = n12270 ^ n12265;
  assign n12325 = n12315 ^ n12309;
  assign n12326 = ~n12277 & ~n12325;
  assign n12336 = n12335 ^ n12326;
  assign n12339 = n12338 ^ n12336;
  assign n12296 = n12295 ^ n12277;
  assign n12328 = n12296 ^ n12288;
  assign n12303 = n12302 ^ n12262;
  assign n12324 = ~n12281 & ~n12303;
  assign n12327 = n12326 ^ n12324;
  assign n12329 = n12328 ^ n12327;
  assign n12297 = n12288 & ~n12296;
  assign n12301 = n12300 ^ n12297;
  assign n12330 = n12329 ^ n12301;
  assign n12353 = n12339 ^ n12330;
  assign n12321 = n12270 & ~n12302;
  assign n12306 = n12305 ^ n12276;
  assign n12310 = n12306 & ~n12309;
  assign n12322 = n12321 ^ n12310;
  assign n12319 = n12309 ^ n12306;
  assign n12320 = n12319 ^ n12318;
  assign n12323 = n12322 ^ n12320;
  assign n12340 = ~n12323 & n12339;
  assign n12307 = n12306 ^ n12302;
  assign n12304 = n12303 ^ n12266;
  assign n12313 = n12307 ^ n12304;
  assign n12308 = ~n12304 & ~n12307;
  assign n12311 = n12310 ^ n12308;
  assign n12312 = n12311 ^ n12301;
  assign n12314 = n12313 ^ n12312;
  assign n12362 = n12340 ^ n12314;
  assign n12363 = ~n12353 & n12362;
  assign n12364 = n12363 ^ n12330;
  assign n12341 = n12323 ^ n12314;
  assign n12345 = n12340 ^ n12330;
  assign n12346 = ~n12341 & ~n12345;
  assign n12347 = n12346 ^ n12314;
  assign n12365 = n12364 ^ n12347;
  assign n12960 = n12299 & ~n12365;
  assign n12355 = n12330 & n12339;
  assign n12356 = n12314 & n12355;
  assign n12354 = n12353 ^ n12340;
  assign n12357 = n12356 ^ n12354;
  assign n12342 = n12341 ^ n12340;
  assign n12331 = ~n12323 & ~n12330;
  assign n12332 = ~n12314 & n12331;
  assign n12343 = n12342 ^ n12332;
  assign n12367 = n12357 ^ n12343;
  assign n12368 = n12367 ^ n12365;
  assign n12854 = ~n12316 & ~n12368;
  assign n12961 = n12960 ^ n12854;
  assign n12359 = n12334 & ~n12343;
  assign n12358 = ~n12302 & ~n12357;
  assign n12360 = n12359 ^ n12358;
  assign n12962 = n12961 ^ n12360;
  assign n12371 = n12364 ^ n12357;
  assign n12372 = n12306 & n12371;
  assign n12369 = n12315 & ~n12368;
  assign n12366 = n12266 & ~n12365;
  assign n12370 = n12369 ^ n12366;
  assign n12373 = n12372 ^ n12370;
  assign n12348 = n12347 ^ n12343;
  assign n12349 = ~n12325 & ~n12348;
  assign n12959 = n12373 ^ n12349;
  assign n12963 = n12962 ^ n12959;
  assign n12969 = n12968 ^ n12963;
  assign n12974 = n12973 ^ n12969;
  assign n12989 = n12988 ^ n12974;
  assign n12897 = n12681 & ~n12712;
  assign n12735 = ~n12703 & ~n12726;
  assign n12898 = n12897 ^ n12735;
  assign n12743 = n12726 ^ n12712;
  assign n12894 = ~n12662 & n12743;
  assign n12893 = ~n12672 & n12729;
  assign n12895 = n12894 ^ n12893;
  assign n12896 = n12895 ^ n12747;
  assign n12899 = n12898 ^ n12896;
  assign n12713 = ~n12640 & ~n12712;
  assign n12892 = n12732 ^ n12713;
  assign n12900 = n12899 ^ n12892;
  assign n12919 = n12918 ^ n12900;
  assign n12888 = n12601 ^ n12582;
  assign n12885 = n12555 & n12581;
  assign n12604 = ~n12536 & ~n12596;
  assign n12886 = n12885 ^ n12604;
  assign n12874 = n12543 & n12590;
  assign n12873 = n12538 & ~n12612;
  assign n12875 = n12874 ^ n12873;
  assign n12876 = n12875 ^ n12616;
  assign n12887 = n12886 ^ n12876;
  assign n12889 = n12888 ^ n12887;
  assign n12881 = n12512 & ~n12593;
  assign n12882 = n12881 ^ n12589;
  assign n12879 = n12518 & ~n12596;
  assign n12603 = n12496 & ~n12593;
  assign n12878 = n12622 ^ n12603;
  assign n12880 = n12879 ^ n12878;
  assign n12883 = n12882 ^ n12880;
  assign n12877 = n12876 ^ n12614;
  assign n12884 = n12883 ^ n12877;
  assign n12890 = n12889 ^ n12884;
  assign n12868 = n12420 & n12464;
  assign n12869 = n12868 ^ n12477;
  assign n12866 = n12421 & n12482;
  assign n12864 = n12398 & n12464;
  assign n12468 = n12394 & n12465;
  assign n12865 = n12864 ^ n12468;
  assign n12867 = n12866 ^ n12865;
  assign n12870 = n12869 ^ n12867;
  assign n12859 = n12413 & n12479;
  assign n12858 = n12426 & n12488;
  assign n12860 = n12859 ^ n12858;
  assign n12862 = n12861 ^ n12860;
  assign n12863 = n12862 ^ n12490;
  assign n12871 = n12870 ^ n12863;
  assign n12852 = ~n12296 & n12367;
  assign n12851 = ~n12309 & n12371;
  assign n12853 = n12852 ^ n12851;
  assign n12855 = n12854 ^ n12853;
  assign n12856 = n12855 ^ n12373;
  assign n12848 = ~n12303 & n12347;
  assign n12849 = n12848 ^ n12360;
  assign n12846 = ~n12304 & ~n12364;
  assign n12844 = ~n12281 & n12347;
  assign n12351 = ~n12277 & ~n12348;
  assign n12845 = n12844 ^ n12351;
  assign n12847 = n12846 ^ n12845;
  assign n12850 = n12849 ^ n12847;
  assign n12857 = n12856 ^ n12850;
  assign n12872 = n12871 ^ n12857;
  assign n12891 = n12890 ^ n12872;
  assign n12920 = n12919 ^ n12891;
  assign n12992 = n12989 ^ n12920;
  assign n13068 = n12671 & n12729;
  assign n13069 = n13068 ^ n12895;
  assign n13066 = n12748 ^ n12728;
  assign n13009 = ~n12704 & ~n12726;
  assign n12734 = ~n12639 & n12723;
  assign n12943 = n12942 ^ n12734;
  assign n13010 = n13009 ^ n12943;
  assign n13067 = n13066 ^ n13010;
  assign n13070 = n13069 ^ n13067;
  assign n13078 = n13077 ^ n13070;
  assign n13039 = ~n12541 & n12590;
  assign n13040 = n13039 ^ n12875;
  assign n13037 = n12617 ^ n12600;
  assign n13038 = n13037 ^ n12880;
  assign n13041 = n13040 ^ n13038;
  assign n13064 = n13041 ^ n12972;
  assign n13061 = n12370 ^ n12359;
  assign n12344 = n12282 & ~n12343;
  assign n12350 = n12349 ^ n12344;
  assign n12352 = n12351 ^ n12350;
  assign n13060 = n12961 ^ n12352;
  assign n13062 = n13061 ^ n13060;
  assign n13058 = n12487 ^ n12476;
  assign n12461 = n12399 & n12460;
  assign n12467 = n12466 ^ n12461;
  assign n12469 = n12468 ^ n12467;
  assign n13057 = n12966 ^ n12469;
  assign n13059 = n13058 ^ n13057;
  assign n13063 = n13062 ^ n13059;
  assign n13065 = n13064 ^ n13063;
  assign n13079 = n13078 ^ n13065;
  assign n13083 = n13079 ^ n12920;
  assign n13007 = ~n12645 & n12723;
  assign n12720 = n12719 ^ n12713;
  assign n13008 = n13007 ^ n12720;
  assign n13011 = n13010 ^ n13008;
  assign n12744 = n12694 & n12743;
  assign n12745 = n12744 ^ n12732;
  assign n13006 = n12896 ^ n12745;
  assign n13012 = n13011 ^ n13006;
  assign n12750 = n12749 ^ n12720;
  assign n12746 = n12745 ^ n12738;
  assign n12751 = n12750 ^ n12746;
  assign n13013 = n13012 ^ n12751;
  assign n13022 = n13021 ^ n13013;
  assign n13004 = n12884 ^ n12620;
  assign n12605 = n12604 ^ n12603;
  assign n12610 = n12609 ^ n12605;
  assign n12602 = n12601 ^ n12589;
  assign n12611 = n12610 ^ n12602;
  assign n13005 = n13004 ^ n12611;
  assign n13023 = n13022 ^ n13005;
  assign n12922 = n12424 & n12482;
  assign n12999 = n12922 ^ n12864;
  assign n13000 = n12999 ^ n12467;
  assign n12998 = n12487 ^ n12477;
  assign n13001 = n13000 ^ n12998;
  assign n12996 = n12370 ^ n12360;
  assign n12928 = ~n12307 & ~n12364;
  assign n12994 = n12928 ^ n12844;
  assign n12995 = n12994 ^ n12350;
  assign n12997 = n12996 ^ n12995;
  assign n13002 = n13001 ^ n12997;
  assign n12944 = n12943 ^ n12898;
  assign n12941 = n12894 ^ n12745;
  assign n12945 = n12944 ^ n12941;
  assign n12946 = n12945 ^ n12751;
  assign n12957 = n12956 ^ n12946;
  assign n12936 = n12886 ^ n12878;
  assign n12935 = n12873 ^ n12614;
  assign n12937 = n12936 ^ n12935;
  assign n12938 = n12937 ^ n12620;
  assign n12939 = n12938 ^ n12889;
  assign n12932 = n12370 ^ n12358;
  assign n12929 = n12333 & ~n12357;
  assign n12930 = n12929 ^ n12928;
  assign n12931 = n12930 ^ n12855;
  assign n12933 = n12932 ^ n12931;
  assign n12926 = n12487 ^ n12475;
  assign n12923 = n12450 & n12474;
  assign n12924 = n12923 ^ n12922;
  assign n12925 = n12924 ^ n12862;
  assign n12927 = n12926 ^ n12925;
  assign n12934 = n12933 ^ n12927;
  assign n12940 = n12939 ^ n12934;
  assign n12958 = n12957 ^ n12940;
  assign n13003 = n13002 ^ n12958;
  assign n13024 = n13023 ^ n13003;
  assign n12736 = n12735 ^ n12734;
  assign n12741 = n12740 ^ n12736;
  assign n12733 = n12732 ^ n12720;
  assign n12742 = n12741 ^ n12733;
  assign n12752 = n12751 ^ n12742;
  assign n12842 = n12841 ^ n12752;
  assign n12624 = n12623 ^ n12589;
  assign n12625 = n12624 ^ n12614;
  assign n12621 = n12620 ^ n12611;
  assign n12626 = n12625 ^ n12621;
  assign n12478 = n12477 ^ n12469;
  assign n12491 = n12490 ^ n12478;
  assign n12361 = n12360 ^ n12352;
  assign n12374 = n12373 ^ n12361;
  assign n12492 = n12491 ^ n12374;
  assign n12627 = n12626 ^ n12492;
  assign n12843 = n12842 ^ n12627;
  assign n12993 = n12989 ^ n12843;
  assign n13025 = n13024 ^ n12993;
  assign n13136 = n13083 ^ n13025;
  assign n12921 = n12920 ^ n12843;
  assign n13044 = n12975 ^ n12720;
  assign n13045 = n13044 ^ n12745;
  assign n13055 = n13054 ^ n13045;
  assign n13042 = n13041 ^ n12625;
  assign n13033 = n12404 & n12479;
  assign n13034 = n13033 ^ n12860;
  assign n13031 = n12965 ^ n12486;
  assign n13032 = n13031 ^ n12867;
  assign n13035 = n13034 ^ n13032;
  assign n13028 = n12288 & n12367;
  assign n13029 = n13028 ^ n12853;
  assign n13026 = n12960 ^ n12366;
  assign n13027 = n13026 ^ n12847;
  assign n13030 = n13029 ^ n13027;
  assign n13036 = n13035 ^ n13030;
  assign n13043 = n13042 ^ n13036;
  assign n13056 = n13055 ^ n13043;
  assign n13107 = n13056 ^ n12920;
  assign n13116 = n13107 ^ n12993;
  assign n13117 = n12921 & n13116;
  assign n13084 = n13083 ^ n13024;
  assign n13085 = n12993 & n13084;
  assign n13118 = n13117 ^ n13085;
  assign n13137 = n13136 ^ n13118;
  assign n13102 = n13101 ^ n12751;
  assign n13091 = n12924 ^ n12865;
  assign n13090 = n12858 ^ n12490;
  assign n13092 = n13091 ^ n13090;
  assign n13088 = n12930 ^ n12845;
  assign n13087 = n12851 ^ n12373;
  assign n13089 = n13088 ^ n13087;
  assign n13093 = n13092 ^ n13089;
  assign n13094 = n13093 ^ n12938;
  assign n13103 = n13102 ^ n13094;
  assign n13080 = n13079 ^ n13056;
  assign n13104 = n13103 ^ n13080;
  assign n13131 = n13104 ^ n12958;
  assign n13132 = n13131 ^ n12992;
  assign n13133 = n13103 ^ n13025;
  assign n13134 = n13132 & n13133;
  assign n12990 = n12989 ^ n12958;
  assign n12991 = n12990 ^ n12921;
  assign n13126 = n12991 & n13025;
  assign n13135 = n13134 ^ n13126;
  assign n13138 = n13137 ^ n13135;
  assign n13081 = n13080 ^ n13025;
  assign n13128 = n13081 ^ n12992;
  assign n13105 = n13104 ^ n12843;
  assign n13125 = n13103 & n13105;
  assign n13127 = n13126 ^ n13125;
  assign n13129 = n13128 ^ n13127;
  assign n13082 = n12992 & n13081;
  assign n13086 = n13085 ^ n13082;
  assign n13130 = n13129 ^ n13086;
  assign n13149 = n13138 ^ n13130;
  assign n13121 = ~n12958 & n13104;
  assign n13108 = n13107 ^ n13024;
  assign n13111 = n12990 & n13108;
  assign n13122 = n13121 ^ n13111;
  assign n13119 = n13108 ^ n12990;
  assign n13120 = n13119 ^ n13118;
  assign n13123 = n13122 ^ n13120;
  assign n13139 = n13123 & n13138;
  assign n13155 = n13149 ^ n13139;
  assign n13109 = n13108 ^ n13104;
  assign n13106 = n13105 ^ n12993;
  assign n13114 = n13109 ^ n13106;
  assign n13110 = n13106 & n13109;
  assign n13112 = n13111 ^ n13110;
  assign n13113 = n13112 ^ n13086;
  assign n13115 = n13114 ^ n13113;
  assign n13153 = ~n13130 & n13138;
  assign n13154 = n13115 & n13153;
  assign n13156 = n13155 ^ n13154;
  assign n13124 = n13123 ^ n13115;
  assign n13145 = n13139 ^ n13124;
  assign n13143 = n13123 & n13130;
  assign n13144 = ~n13115 & n13143;
  assign n13146 = n13145 ^ n13144;
  assign n13160 = n13156 ^ n13146;
  assign n13488 = n12992 & n13160;
  assign n13367 = n13081 & n13160;
  assign n13150 = n13139 ^ n13115;
  assign n13151 = n13149 & n13150;
  assign n13152 = n13151 ^ n13130;
  assign n13157 = n13156 ^ n13152;
  assign n13366 = n12990 & n13157;
  assign n13368 = n13367 ^ n13366;
  assign n13489 = n13488 ^ n13368;
  assign n13140 = n13139 ^ n13130;
  assign n13141 = n13124 & n13140;
  assign n13142 = n13141 ^ n13115;
  assign n13159 = n13152 ^ n13142;
  assign n13168 = n13084 & n13159;
  assign n13163 = n12993 & n13159;
  assign n13486 = n13168 ^ n13163;
  assign n13484 = n13106 & n13152;
  assign n13414 = n13103 & n13142;
  assign n13147 = n13146 ^ n13142;
  assign n13314 = n13025 & n13147;
  assign n13436 = n13414 ^ n13314;
  assign n13485 = n13484 ^ n13436;
  assign n13487 = n13486 ^ n13485;
  assign n13490 = n13489 ^ n13487;
  assign n17276 = n15369 ^ n13490;
  assign n10820 = n9785 ^ n9678;
  assign n10822 = n10821 ^ n10820;
  assign n10819 = n10818 ^ n9696;
  assign n10823 = n10822 ^ n10819;
  assign n10764 = n9855 ^ n9820;
  assign n10766 = n10765 ^ n10764;
  assign n10763 = n10762 ^ n9832;
  assign n10767 = n10766 ^ n10763;
  assign n10824 = n10823 ^ n10767;
  assign n10793 = n10792 ^ n9733;
  assign n9753 = n9752 ^ n9287;
  assign n10791 = n10790 ^ n9753;
  assign n10794 = n10793 ^ n10791;
  assign n10782 = n10781 ^ n9678;
  assign n10784 = n10783 ^ n10782;
  assign n9667 = n9666 ^ n9287;
  assign n10780 = n10779 ^ n9667;
  assign n10785 = n10784 ^ n10780;
  assign n10787 = n10786 ^ n10785;
  assign n10795 = n10794 ^ n10787;
  assign n10825 = n10824 ^ n10795;
  assign n10839 = n10838 ^ n10781;
  assign n10837 = n10836 ^ n9287;
  assign n10840 = n10839 ^ n10837;
  assign n10772 = n9820 ^ n9401;
  assign n10774 = n10773 ^ n10772;
  assign n10771 = n10770 ^ n9524;
  assign n10775 = n10774 ^ n10771;
  assign n10776 = n10775 ^ n10767;
  assign n10841 = n10840 ^ n10776;
  assign n10874 = ~n10785 & n10841;
  assign n10830 = n10823 ^ n10775;
  assign n10831 = n10830 ^ n10795;
  assign n10809 = n9855 ^ n9630;
  assign n10811 = n10810 ^ n10809;
  assign n10808 = n10807 ^ n9623;
  assign n10812 = n10811 ^ n10808;
  assign n10832 = n10812 ^ n10785;
  assign n10833 = n10831 & n10832;
  assign n10875 = n10874 ^ n10833;
  assign n10872 = n10832 ^ n10831;
  assign n10801 = n10800 ^ n9401;
  assign n10803 = n10802 ^ n10801;
  assign n9288 = n9287 ^ n9278;
  assign n10799 = n10798 ^ n9288;
  assign n10804 = n10803 ^ n10799;
  assign n10850 = n10823 ^ n10804;
  assign n10813 = n10812 ^ n10804;
  assign n10859 = n10830 ^ n10813;
  assign n10860 = n10850 & n10859;
  assign n10826 = n10813 & n10825;
  assign n10861 = n10860 ^ n10826;
  assign n10873 = n10872 ^ n10861;
  assign n10876 = n10875 ^ n10873;
  assign n10843 = n10841 ^ n10804;
  assign n10844 = n10843 ^ n10813;
  assign n10842 = n10841 ^ n10831;
  assign n10848 = n10844 ^ n10842;
  assign n10845 = n10842 & n10844;
  assign n10846 = n10845 ^ n10833;
  assign n10814 = n10813 ^ n10795;
  assign n10815 = n10814 ^ n10776;
  assign n10827 = n10823 ^ n10812;
  assign n10828 = n10815 & n10827;
  assign n10829 = n10828 ^ n10826;
  assign n10847 = n10846 ^ n10829;
  assign n10849 = n10848 ^ n10847;
  assign n10882 = n10876 ^ n10849;
  assign n10858 = n10824 ^ n10814;
  assign n10862 = n10861 ^ n10858;
  assign n10853 = n10840 ^ n10814;
  assign n10854 = n10841 ^ n10785;
  assign n10855 = n10854 ^ n10827;
  assign n10856 = n10853 & n10855;
  assign n10851 = n10850 ^ n10832;
  assign n10852 = n10814 & n10851;
  assign n10857 = n10856 ^ n10852;
  assign n10863 = n10862 ^ n10857;
  assign n10877 = n10863 & n10876;
  assign n10866 = n10827 ^ n10815;
  assign n10864 = n10840 & n10843;
  assign n10865 = n10864 ^ n10852;
  assign n10867 = n10866 ^ n10865;
  assign n10868 = n10867 ^ n10829;
  assign n10893 = n10877 ^ n10868;
  assign n10894 = n10882 & n10893;
  assign n10895 = n10894 ^ n10849;
  assign n10871 = n10868 ^ n10863;
  assign n10887 = n10877 ^ n10849;
  assign n10888 = n10871 & n10887;
  assign n10889 = n10888 ^ n10868;
  assign n10896 = n10895 ^ n10889;
  assign n11056 = n10825 & n10896;
  assign n10883 = n10882 ^ n10877;
  assign n10880 = n10868 & n10876;
  assign n10881 = ~n10849 & n10880;
  assign n10884 = n10883 ^ n10881;
  assign n10878 = n10877 ^ n10871;
  assign n10869 = n10863 & ~n10868;
  assign n10870 = n10849 & n10869;
  assign n10879 = n10878 ^ n10870;
  assign n10885 = n10884 ^ n10879;
  assign n10897 = n10896 ^ n10885;
  assign n10898 = n10859 & n10897;
  assign n11130 = n11056 ^ n10898;
  assign n10907 = n10855 & n10884;
  assign n10906 = n10841 & n10879;
  assign n10908 = n10907 ^ n10906;
  assign n11131 = n11130 ^ n10908;
  assign n10913 = n10895 ^ n10884;
  assign n11101 = n10851 & n10913;
  assign n10890 = n10889 ^ n10879;
  assign n10903 = n10831 & n10890;
  assign n10901 = n10813 & n10896;
  assign n10900 = n10850 & n10897;
  assign n10902 = n10901 ^ n10900;
  assign n10904 = n10903 ^ n10902;
  assign n11129 = n11101 ^ n10904;
  assign n11132 = n11131 ^ n11129;
  assign n11138 = n11137 ^ n11132;
  assign n10656 = n9808 ^ n7891;
  assign n10654 = n7973 ^ n7904;
  assign n10653 = n7953 ^ n7875;
  assign n10655 = n10654 ^ n10653;
  assign n10657 = n10656 ^ n10655;
  assign n10613 = n9863 ^ n8001;
  assign n10611 = n8012 ^ n7786;
  assign n7836 = n7835 ^ n7824;
  assign n10612 = n10611 ^ n7836;
  assign n10614 = n10613 ^ n10612;
  assign n10666 = n10657 ^ n10614;
  assign n10641 = n7978 ^ n7553;
  assign n7965 = n7897 ^ n7413;
  assign n10640 = n10639 ^ n7965;
  assign n10642 = n10641 ^ n10640;
  assign n10637 = n9720 ^ n7921;
  assign n10635 = n9709 ^ n7953;
  assign n7934 = n7933 ^ n7413;
  assign n10633 = n10632 ^ n7934;
  assign n10631 = n7946 ^ n7884;
  assign n10634 = n10633 ^ n10631;
  assign n10636 = n10635 ^ n10634;
  assign n10638 = n10637 ^ n10636;
  assign n10643 = n10642 ^ n10638;
  assign n10667 = n10666 ^ n10643;
  assign n10617 = n9840 ^ n7824;
  assign n10615 = n8007 ^ n7848;
  assign n7407 = n7406 ^ n7278;
  assign n10616 = n10615 ^ n7407;
  assign n10618 = n10617 ^ n10616;
  assign n10678 = n10657 ^ n10618;
  assign n10685 = n10678 ^ n10643;
  assign n10646 = n10632 ^ n7413;
  assign n10647 = n10646 ^ n7939;
  assign n10648 = n10647 ^ n7985;
  assign n10649 = n10648 ^ n9775;
  assign n10619 = n10618 ^ n10614;
  assign n10650 = n10649 ^ n10619;
  assign n10695 = n10685 ^ n10650;
  assign n10628 = n9612 ^ n7278;
  assign n7420 = n7419 ^ n7413;
  assign n10626 = n10625 ^ n7420;
  assign n10624 = n7851 ^ n7687;
  assign n10627 = n10626 ^ n10624;
  assign n10629 = n10628 ^ n10627;
  assign n10651 = n10650 ^ n10629;
  assign n10622 = n9647 ^ n7800;
  assign n10620 = n7792 ^ n7545;
  assign n8002 = n8001 ^ n7780;
  assign n10621 = n10620 ^ n8002;
  assign n10623 = n10622 ^ n10621;
  assign n10630 = n10629 ^ n10623;
  assign n10694 = n10651 ^ n10630;
  assign n10699 = n10695 ^ n10694;
  assign n10696 = ~n10694 & ~n10695;
  assign n10659 = n10636 ^ n10623;
  assign n10689 = ~n10659 & n10685;
  assign n10697 = n10696 ^ n10689;
  assign n10644 = n10643 ^ n10630;
  assign n10645 = n10644 ^ n10619;
  assign n10663 = n10657 ^ n10623;
  assign n10669 = ~n10645 & n10663;
  assign n10668 = n10630 & n10667;
  assign n10670 = n10669 ^ n10668;
  assign n10698 = n10697 ^ n10670;
  assign n10700 = n10699 ^ n10698;
  assign n10688 = n10636 & ~n10650;
  assign n10690 = n10689 ^ n10688;
  assign n10686 = n10685 ^ n10659;
  assign n10658 = n10657 ^ n10629;
  assign n10679 = n10678 ^ n10630;
  assign n10680 = n10658 & ~n10679;
  assign n10681 = n10680 ^ n10668;
  assign n10687 = n10686 ^ n10681;
  assign n10691 = n10690 ^ n10687;
  assign n10706 = n10700 ^ n10691;
  assign n10677 = n10666 ^ n10644;
  assign n10682 = n10681 ^ n10677;
  assign n10672 = n10650 ^ n10636;
  assign n10673 = n10672 ^ n10663;
  assign n10674 = n10649 ^ n10644;
  assign n10675 = n10673 & n10674;
  assign n10660 = n10659 ^ n10658;
  assign n10661 = ~n10644 & ~n10660;
  assign n10676 = n10675 ^ n10661;
  assign n10683 = n10682 ^ n10676;
  assign n10692 = n10683 & ~n10691;
  assign n10664 = n10663 ^ n10645;
  assign n10652 = ~n10649 & ~n10651;
  assign n10662 = n10661 ^ n10652;
  assign n10665 = n10664 ^ n10662;
  assign n10671 = n10670 ^ n10665;
  assign n10717 = n10692 ^ n10671;
  assign n10718 = ~n10706 & ~n10717;
  assign n10719 = n10718 ^ n10700;
  assign n10684 = n10683 ^ n10671;
  assign n10711 = n10700 ^ n10692;
  assign n10712 = ~n10684 & n10711;
  assign n10713 = n10712 ^ n10671;
  assign n10720 = n10719 ^ n10713;
  assign n11042 = n10667 & ~n10720;
  assign n10707 = n10706 ^ n10692;
  assign n10704 = ~n10671 & ~n10691;
  assign n10705 = ~n10700 & n10704;
  assign n10708 = n10707 ^ n10705;
  assign n10701 = n10671 & n10683;
  assign n10702 = n10700 & n10701;
  assign n10693 = n10692 ^ n10684;
  assign n10703 = n10702 ^ n10693;
  assign n10709 = n10708 ^ n10703;
  assign n10721 = n10720 ^ n10709;
  assign n10722 = ~n10679 & ~n10721;
  assign n11124 = n11042 ^ n10722;
  assign n10731 = n10673 & ~n10708;
  assign n10730 = ~n10650 & ~n10703;
  assign n10732 = n10731 ^ n10730;
  assign n11125 = n11124 ^ n10732;
  assign n10737 = n10719 ^ n10708;
  assign n11072 = ~n10660 & ~n10737;
  assign n10714 = n10713 ^ n10703;
  assign n10727 = n10685 & n10714;
  assign n10725 = n10658 & ~n10721;
  assign n10724 = n10630 & ~n10720;
  assign n10726 = n10725 ^ n10724;
  assign n10728 = n10727 ^ n10726;
  assign n11123 = n11072 ^ n10728;
  assign n11126 = n11125 ^ n11123;
  assign n7033 = n7032 ^ n7004;
  assign n10529 = n7033 ^ n7012;
  assign n10530 = n10529 ^ n6988;
  assign n10531 = n10530 ^ n7055;
  assign n10532 = n10531 ^ n7913;
  assign n4914 = n4913 ^ n3948;
  assign n10492 = n10491 ^ n4914;
  assign n10493 = n10492 ^ n6941;
  assign n10494 = n10493 ^ n8018;
  assign n10542 = n10532 ^ n10494;
  assign n10525 = n10524 ^ n7048;
  assign n7057 = n6994 ^ n6909;
  assign n10523 = n7057 ^ n6962;
  assign n10526 = n10525 ^ n10523;
  assign n10521 = n7928 ^ n7062;
  assign n10519 = n7960 ^ n7037;
  assign n10517 = n10497 ^ n7032;
  assign n7028 = n6909 ^ n6892;
  assign n10516 = n7028 ^ n7001;
  assign n10518 = n10517 ^ n10516;
  assign n10520 = n10519 ^ n10518;
  assign n10522 = n10521 ^ n10520;
  assign n10527 = n10526 ^ n10522;
  assign n10543 = n10542 ^ n10527;
  assign n10488 = n10487 ^ n6853;
  assign n6972 = n6971 ^ n4928;
  assign n10489 = n10488 ^ n6972;
  assign n10490 = n10489 ^ n7867;
  assign n10554 = n10532 ^ n10490;
  assign n10561 = n10554 ^ n10527;
  assign n10499 = n7995 ^ n6919;
  assign n10496 = n7026 ^ n6909;
  assign n10498 = n10497 ^ n10496;
  assign n10500 = n10499 ^ n10498;
  assign n10495 = n10494 ^ n10490;
  assign n10501 = n10500 ^ n10495;
  assign n10571 = n10561 ^ n10501;
  assign n10513 = n7808 ^ n6948;
  assign n10511 = n6937 ^ n6834;
  assign n10510 = n6906 ^ n6839;
  assign n10512 = n10511 ^ n10510;
  assign n10514 = n10513 ^ n10512;
  assign n10504 = n10503 ^ n10502;
  assign n6968 = n6967 ^ n6909;
  assign n10505 = n10504 ^ n6968;
  assign n10506 = n10505 ^ n5840;
  assign n10507 = n10506 ^ n7775;
  assign n10515 = n10514 ^ n10507;
  assign n10508 = n10507 ^ n10501;
  assign n10570 = n10515 ^ n10508;
  assign n10575 = n10571 ^ n10570;
  assign n10572 = ~n10570 & ~n10571;
  assign n10534 = n10520 ^ n10514;
  assign n10565 = ~n10534 & n10561;
  assign n10573 = n10572 ^ n10565;
  assign n10528 = n10527 ^ n10515;
  assign n10538 = n10528 ^ n10495;
  assign n10539 = n10532 ^ n10514;
  assign n10545 = ~n10538 & n10539;
  assign n10544 = n10515 & n10543;
  assign n10546 = n10545 ^ n10544;
  assign n10574 = n10573 ^ n10546;
  assign n10576 = n10575 ^ n10574;
  assign n10564 = ~n10501 & n10520;
  assign n10566 = n10565 ^ n10564;
  assign n10562 = n10561 ^ n10534;
  assign n10533 = n10532 ^ n10507;
  assign n10555 = n10554 ^ n10515;
  assign n10556 = n10533 & ~n10555;
  assign n10557 = n10556 ^ n10544;
  assign n10563 = n10562 ^ n10557;
  assign n10567 = n10566 ^ n10563;
  assign n10584 = n10576 ^ n10567;
  assign n10553 = n10542 ^ n10528;
  assign n10558 = n10557 ^ n10553;
  assign n10548 = n10520 ^ n10501;
  assign n10549 = n10548 ^ n10539;
  assign n10550 = n10528 ^ n10500;
  assign n10551 = n10549 & n10550;
  assign n10535 = n10534 ^ n10533;
  assign n10536 = ~n10528 & ~n10535;
  assign n10552 = n10551 ^ n10536;
  assign n10559 = n10558 ^ n10552;
  assign n10568 = n10559 & ~n10567;
  assign n10540 = n10539 ^ n10538;
  assign n10509 = ~n10500 & ~n10508;
  assign n10537 = n10536 ^ n10509;
  assign n10541 = n10540 ^ n10537;
  assign n10547 = n10546 ^ n10541;
  assign n10585 = n10568 ^ n10547;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = n10586 ^ n10576;
  assign n10560 = n10559 ^ n10547;
  assign n10581 = n10576 ^ n10568;
  assign n10582 = ~n10560 & n10581;
  assign n10583 = n10582 ^ n10547;
  assign n10588 = n10587 ^ n10583;
  assign n11048 = n10543 & ~n10588;
  assign n10592 = n10584 ^ n10568;
  assign n10590 = ~n10547 & ~n10567;
  assign n10591 = ~n10576 & n10590;
  assign n10593 = n10592 ^ n10591;
  assign n10577 = n10547 & n10559;
  assign n10578 = n10576 & n10577;
  assign n10569 = n10568 ^ n10560;
  assign n10579 = n10578 ^ n10569;
  assign n10594 = n10593 ^ n10579;
  assign n10595 = n10594 ^ n10588;
  assign n10603 = ~n10555 & ~n10595;
  assign n11095 = n11048 ^ n10603;
  assign n10747 = n10549 & ~n10593;
  assign n10580 = ~n10501 & ~n10579;
  assign n10748 = n10747 ^ n10580;
  assign n11096 = n11095 ^ n10748;
  assign n10752 = n10593 ^ n10587;
  assign n11036 = ~n10535 & ~n10752;
  assign n10600 = n10583 ^ n10579;
  assign n10743 = n10561 & n10600;
  assign n10596 = n10533 & ~n10595;
  assign n10589 = n10515 & ~n10588;
  assign n10597 = n10596 ^ n10589;
  assign n10744 = n10743 ^ n10597;
  assign n11094 = n11036 ^ n10744;
  assign n11097 = n11096 ^ n11094;
  assign n11127 = n11126 ^ n11097;
  assign n11120 = n10747 ^ n10597;
  assign n11035 = n10550 & ~n10593;
  assign n11037 = n11036 ^ n11035;
  assign n10753 = ~n10528 & ~n10752;
  assign n11038 = n11037 ^ n10753;
  assign n11119 = n11095 ^ n11038;
  assign n11121 = n11120 ^ n11119;
  assign n10394 = n8925 ^ n6928;
  assign n10392 = n8886 ^ n8815;
  assign n8812 = n8811 ^ n8803;
  assign n10393 = n10392 ^ n8812;
  assign n10395 = n10394 ^ n10393;
  assign n10389 = n8874 ^ n6882;
  assign n10387 = n8763 ^ n8456;
  assign n10388 = n10387 ^ n8712;
  assign n10390 = n10389 ^ n10388;
  assign n10385 = n8248 ^ n6818;
  assign n10383 = n8898 ^ n8749;
  assign n10384 = n10383 ^ n8777;
  assign n10386 = n10385 ^ n10384;
  assign n10391 = n10390 ^ n10386;
  assign n10396 = n10395 ^ n10391;
  assign n10375 = n8832 ^ n7041;
  assign n8822 = n8821 ^ n8815;
  assign n10373 = n10372 ^ n8822;
  assign n10374 = n10373 ^ n8921;
  assign n10376 = n10375 ^ n10374;
  assign n10430 = n10396 ^ n10376;
  assign n10402 = n8947 ^ n7019;
  assign n10400 = n8917 ^ n8851;
  assign n8869 = n8868 ^ n8860;
  assign n10401 = n10400 ^ n8869;
  assign n10403 = n10402 ^ n10401;
  assign n10370 = n8785 ^ n6954;
  assign n10368 = n8593 ^ n8469;
  assign n8887 = n8886 ^ n8883;
  assign n10369 = n10368 ^ n8887;
  assign n10371 = n10370 ^ n10369;
  assign n10416 = n10403 ^ n10371;
  assign n10431 = n10430 ^ n10416;
  assign n10451 = n10376 & ~n10396;
  assign n10377 = n10376 ^ n10371;
  assign n10408 = n8906 ^ n7067;
  assign n8955 = n8848 ^ n8815;
  assign n10407 = n10406 ^ n8955;
  assign n10409 = n10408 ^ n10407;
  assign n8941 = n8940 ^ n8936;
  assign n10405 = n10376 ^ n8941;
  assign n10410 = n10409 ^ n10405;
  assign n10404 = n10403 ^ n10386;
  assign n10411 = n10410 ^ n10404;
  assign n10414 = ~n10377 & n10411;
  assign n10452 = n10451 ^ n10414;
  assign n10449 = n10411 ^ n10377;
  assign n10381 = n8728 ^ n6978;
  assign n8895 = n8894 ^ n8815;
  assign n10379 = n10378 ^ n8895;
  assign n10380 = n10379 ^ n8901;
  assign n10382 = n10381 ^ n10380;
  assign n10427 = n10403 ^ n10382;
  assign n10398 = n10382 ^ n10371;
  assign n10436 = n10404 ^ n10398;
  assign n10437 = ~n10427 & ~n10436;
  assign n10420 = n10403 ^ n10390;
  assign n10421 = n10420 ^ n10410;
  assign n10422 = n10398 & n10421;
  assign n10438 = n10437 ^ n10422;
  assign n10450 = n10449 ^ n10438;
  assign n10453 = n10452 ^ n10450;
  assign n10412 = n10411 ^ n10396;
  assign n10397 = n10396 ^ n10382;
  assign n10399 = n10398 ^ n10397;
  assign n10425 = n10412 ^ n10399;
  assign n10417 = n10410 ^ n10398;
  assign n10418 = n10417 ^ n10391;
  assign n10419 = ~n10416 & ~n10418;
  assign n10423 = n10422 ^ n10419;
  assign n10413 = ~n10399 & ~n10412;
  assign n10415 = n10414 ^ n10413;
  assign n10424 = n10423 ^ n10415;
  assign n10426 = n10425 ^ n10424;
  assign n10464 = n10453 ^ n10426;
  assign n10435 = n10420 ^ n10417;
  assign n10439 = n10438 ^ n10435;
  assign n10432 = n10417 ^ n10395;
  assign n10433 = ~n10431 & n10432;
  assign n10428 = n10427 ^ n10377;
  assign n10429 = ~n10417 & n10428;
  assign n10434 = n10433 ^ n10429;
  assign n10440 = n10439 ^ n10434;
  assign n10454 = n10440 & ~n10453;
  assign n10465 = n10464 ^ n10454;
  assign n10443 = n10418 ^ n10416;
  assign n10441 = ~n10395 & ~n10397;
  assign n10442 = n10441 ^ n10429;
  assign n10444 = n10443 ^ n10442;
  assign n10445 = n10444 ^ n10423;
  assign n10462 = n10445 & ~n10453;
  assign n10463 = ~n10426 & n10462;
  assign n10466 = n10465 ^ n10463;
  assign n11029 = ~n10431 & ~n10466;
  assign n10470 = n10454 ^ n10445;
  assign n10471 = ~n10464 & n10470;
  assign n10472 = n10471 ^ n10426;
  assign n10448 = n10445 ^ n10440;
  assign n10457 = n10454 ^ n10426;
  assign n10458 = n10448 & n10457;
  assign n10459 = n10458 ^ n10445;
  assign n10473 = n10472 ^ n10459;
  assign n10482 = n10398 & n10473;
  assign n10455 = n10454 ^ n10448;
  assign n10446 = n10440 & ~n10445;
  assign n10447 = n10426 & n10446;
  assign n10456 = n10455 ^ n10447;
  assign n10467 = n10466 ^ n10456;
  assign n10474 = n10473 ^ n10467;
  assign n10481 = ~n10427 & ~n10474;
  assign n10483 = n10482 ^ n10481;
  assign n11117 = n11029 ^ n10483;
  assign n11085 = n10421 & n10473;
  assign n10475 = ~n10436 & ~n10474;
  assign n11086 = n11085 ^ n10475;
  assign n11024 = n10472 ^ n10466;
  assign n11027 = ~n10417 & ~n11024;
  assign n11025 = n10428 & ~n11024;
  assign n11023 = n10432 & ~n10466;
  assign n11026 = n11025 ^ n11023;
  assign n11028 = n11027 ^ n11026;
  assign n11116 = n11086 ^ n11028;
  assign n11118 = n11117 ^ n11116;
  assign n11122 = n11121 ^ n11118;
  assign n11128 = n11127 ^ n11122;
  assign n11139 = n11138 ^ n11128;
  assign n10914 = n10814 & n10913;
  assign n10912 = n10840 & n10895;
  assign n10915 = n10914 ^ n10912;
  assign n10911 = n10844 & n10889;
  assign n10916 = n10915 ^ n10911;
  assign n10909 = n10843 & n10895;
  assign n10910 = n10909 ^ n10908;
  assign n10917 = n10916 ^ n10910;
  assign n10891 = n10832 & n10890;
  assign n10886 = n10815 & n10885;
  assign n10892 = n10891 ^ n10886;
  assign n10899 = n10898 ^ n10892;
  assign n10905 = n10904 ^ n10899;
  assign n10918 = n10917 ^ n10905;
  assign n11021 = n11020 ^ n10918;
  assign n10751 = ~n10500 & n10587;
  assign n10754 = n10753 ^ n10751;
  assign n10750 = ~n10570 & ~n10583;
  assign n10755 = n10754 ^ n10750;
  assign n10746 = ~n10508 & n10587;
  assign n10749 = n10748 ^ n10746;
  assign n10756 = n10755 ^ n10749;
  assign n10601 = ~n10534 & n10600;
  assign n10599 = ~n10538 & n10594;
  assign n10602 = n10601 ^ n10599;
  assign n10604 = n10603 ^ n10602;
  assign n10745 = n10744 ^ n10604;
  assign n10757 = n10756 ^ n10745;
  assign n10738 = ~n10644 & ~n10737;
  assign n10736 = ~n10649 & n10719;
  assign n10739 = n10738 ^ n10736;
  assign n10735 = ~n10694 & ~n10713;
  assign n10740 = n10739 ^ n10735;
  assign n10733 = ~n10651 & n10719;
  assign n10734 = n10733 ^ n10732;
  assign n10741 = n10740 ^ n10734;
  assign n10715 = ~n10659 & n10714;
  assign n10710 = ~n10645 & n10709;
  assign n10716 = n10715 ^ n10710;
  assign n10723 = n10722 ^ n10716;
  assign n10729 = n10728 ^ n10723;
  assign n10742 = n10741 ^ n10729;
  assign n10758 = n10757 ^ n10742;
  assign n10606 = n10548 & ~n10579;
  assign n10605 = ~n10571 & ~n10583;
  assign n10607 = n10606 ^ n10605;
  assign n10608 = n10607 ^ n10604;
  assign n10598 = n10597 ^ n10580;
  assign n10609 = n10608 ^ n10598;
  assign n10484 = ~n10396 & n10456;
  assign n10485 = n10484 ^ n10483;
  assign n10478 = ~n10412 & n10459;
  assign n10477 = n10430 & n10456;
  assign n10479 = n10478 ^ n10477;
  assign n10468 = ~n10418 & ~n10467;
  assign n10460 = n10459 ^ n10456;
  assign n10461 = ~n10377 & n10460;
  assign n10469 = n10468 ^ n10461;
  assign n10476 = n10475 ^ n10469;
  assign n10480 = n10479 ^ n10476;
  assign n10486 = n10485 ^ n10480;
  assign n10610 = n10609 ^ n10486;
  assign n10759 = n10758 ^ n10610;
  assign n11022 = n11021 ^ n10759;
  assign n11142 = n11139 ^ n11022;
  assign n11161 = n10842 & n10889;
  assign n11232 = n11161 ^ n10912;
  assign n11102 = n10853 & n10884;
  assign n11103 = n11102 ^ n11101;
  assign n11233 = n11232 ^ n11103;
  assign n11231 = n10908 ^ n10902;
  assign n11234 = n11233 ^ n11231;
  assign n11240 = n11239 ^ n11234;
  assign n11229 = n11097 ^ n10757;
  assign n11224 = ~n10397 & n10472;
  assign n11030 = n11029 ^ n10484;
  assign n11225 = n11224 ^ n11030;
  assign n11176 = ~n10399 & n10459;
  assign n11080 = ~n10395 & n10472;
  assign n11151 = n11080 ^ n11027;
  assign n11177 = n11176 ^ n11151;
  assign n11226 = n11225 ^ n11177;
  assign n11032 = n10411 & n10460;
  assign n11033 = n11032 ^ n10483;
  assign n11223 = n11033 ^ n10476;
  assign n11227 = n11226 ^ n11223;
  assign n11087 = n11086 ^ n11030;
  assign n11084 = n11033 ^ n11025;
  assign n11088 = n11087 ^ n11084;
  assign n11228 = n11227 ^ n11088;
  assign n11230 = n11229 ^ n11228;
  assign n11241 = n11240 ^ n11230;
  assign n11145 = ~n10695 & ~n10713;
  assign n11218 = n11145 ^ n10736;
  assign n11073 = n10674 & ~n10708;
  assign n11074 = n11073 ^ n11072;
  assign n11219 = n11218 ^ n11074;
  assign n11217 = n10732 ^ n10726;
  assign n11220 = n11219 ^ n11217;
  assign n11091 = n10751 ^ n10605;
  assign n11092 = n11091 ^ n11037;
  assign n11090 = n10748 ^ n10597;
  assign n11093 = n11092 ^ n11090;
  assign n11221 = n11220 ^ n11093;
  assign n11165 = n10906 ^ n10902;
  assign n11162 = n10854 & n10879;
  assign n11163 = n11162 ^ n11161;
  assign n11164 = n11163 ^ n10899;
  assign n11166 = n11165 ^ n11164;
  assign n11174 = n11173 ^ n11166;
  assign n11156 = n10754 ^ n10607;
  assign n11155 = n10744 ^ n10601;
  assign n11157 = n11156 ^ n11155;
  assign n11158 = n11157 ^ n11097;
  assign n11152 = n11151 ^ n10479;
  assign n11150 = n11033 ^ n10461;
  assign n11153 = n11152 ^ n11150;
  assign n11154 = n11153 ^ n11088;
  assign n11159 = n11158 ^ n11154;
  assign n11144 = n10672 & ~n10703;
  assign n11146 = n11145 ^ n11144;
  assign n11147 = n11146 ^ n10723;
  assign n11143 = n10730 ^ n10726;
  assign n11148 = n11147 ^ n11143;
  assign n11149 = n11148 ^ n10609;
  assign n11160 = n11159 ^ n11149;
  assign n11175 = n11174 ^ n11160;
  assign n11222 = n11221 ^ n11175;
  assign n11242 = n11241 ^ n11222;
  assign n11059 = n10827 & n10885;
  assign n11060 = n11059 ^ n10892;
  assign n11057 = n11056 ^ n10901;
  assign n11058 = n11057 ^ n10916;
  assign n11061 = n11060 ^ n11058;
  assign n11069 = n11068 ^ n11061;
  assign n11051 = n10539 & n10594;
  assign n11052 = n11051 ^ n10602;
  assign n11049 = n11048 ^ n10589;
  assign n11050 = n11049 ^ n10755;
  assign n11053 = n11052 ^ n11050;
  assign n11045 = n10663 & n10709;
  assign n11046 = n11045 ^ n10716;
  assign n11043 = n11042 ^ n10724;
  assign n11044 = n11043 ^ n10740;
  assign n11047 = n11046 ^ n11044;
  assign n11054 = n11053 ^ n11047;
  assign n11039 = n11038 ^ n10748;
  assign n11040 = n11039 ^ n10744;
  assign n11031 = n11030 ^ n11028;
  assign n11034 = n11033 ^ n11031;
  assign n11041 = n11040 ^ n11034;
  assign n11055 = n11054 ^ n11041;
  assign n11070 = n11069 ^ n11055;
  assign n11071 = n11070 ^ n11022;
  assign n11269 = n11242 ^ n11071;
  assign n11206 = n11163 ^ n10915;
  assign n11205 = n10904 ^ n10891;
  assign n11207 = n11206 ^ n11205;
  assign n11212 = n11211 ^ n11207;
  assign n11201 = n11146 ^ n10739;
  assign n11200 = n10728 ^ n10715;
  assign n11202 = n11201 ^ n11200;
  assign n11203 = n11202 ^ n11157;
  assign n11199 = n11097 ^ n11088;
  assign n11204 = n11203 ^ n11199;
  assign n11213 = n11212 ^ n11204;
  assign n11190 = n10907 ^ n10902;
  assign n11104 = n11103 ^ n10914;
  assign n11189 = n11130 ^ n11104;
  assign n11191 = n11190 ^ n11189;
  assign n11196 = n11195 ^ n11191;
  assign n11185 = n10731 ^ n10726;
  assign n11075 = n11074 ^ n10738;
  assign n11184 = n11124 ^ n11075;
  assign n11186 = n11185 ^ n11184;
  assign n11187 = n11186 ^ n11121;
  assign n11180 = ~n10416 & ~n10467;
  assign n11181 = n11180 ^ n10469;
  assign n11178 = n11085 ^ n10482;
  assign n11179 = n11178 ^ n11177;
  assign n11182 = n11181 ^ n11179;
  assign n11183 = n11182 ^ n11053;
  assign n11188 = n11187 ^ n11183;
  assign n11197 = n11196 ^ n11188;
  assign n11198 = n11197 ^ n11070;
  assign n11214 = n11213 ^ n11198;
  assign n11278 = n11269 ^ n11214;
  assign n11105 = n11104 ^ n10908;
  assign n11106 = n11105 ^ n10904;
  assign n11114 = n11113 ^ n11106;
  assign n11098 = n11097 ^ n11093;
  assign n11081 = n11080 ^ n10478;
  assign n11082 = n11081 ^ n11026;
  assign n11079 = n11030 ^ n10483;
  assign n11083 = n11082 ^ n11079;
  assign n11089 = n11088 ^ n11083;
  assign n11099 = n11098 ^ n11089;
  assign n11076 = n11075 ^ n10732;
  assign n11077 = n11076 ^ n10728;
  assign n11078 = n11077 ^ n11040;
  assign n11100 = n11099 ^ n11078;
  assign n11115 = n11114 ^ n11100;
  assign n11259 = n11214 ^ n11115;
  assign n11140 = n11139 ^ n11115;
  assign n11277 = n11259 ^ n11140;
  assign n11282 = n11278 ^ n11277;
  assign n11279 = n11277 & ~n11278;
  assign n11247 = n11175 ^ n11139;
  assign n11273 = n11247 & ~n11269;
  assign n11280 = n11279 ^ n11273;
  assign n11243 = n11242 ^ n11140;
  assign n11262 = n11243 ^ n11198;
  assign n11265 = ~n11142 & ~n11262;
  assign n11251 = n11197 ^ n11022;
  assign n11254 = n11251 ^ n11242;
  assign n11255 = n11140 & ~n11254;
  assign n11266 = n11265 ^ n11255;
  assign n11281 = n11280 ^ n11266;
  assign n11283 = n11282 ^ n11281;
  assign n11263 = n11262 ^ n11142;
  assign n11260 = n11213 & n11259;
  assign n11246 = n11115 ^ n11022;
  assign n11248 = n11247 ^ n11246;
  assign n11249 = ~n11243 & ~n11248;
  assign n11261 = n11260 ^ n11249;
  assign n11264 = n11263 ^ n11261;
  assign n11267 = n11266 ^ n11264;
  assign n11272 = ~n11175 & n11214;
  assign n11274 = n11273 ^ n11272;
  assign n11270 = n11269 ^ n11247;
  assign n11141 = n11140 ^ n11071;
  assign n11253 = n11141 & ~n11246;
  assign n11256 = n11255 ^ n11253;
  assign n11271 = n11270 ^ n11256;
  assign n11275 = n11274 ^ n11271;
  assign n11297 = n11267 & ~n11275;
  assign n11298 = n11283 & n11297;
  assign n11287 = n11283 ^ n11275;
  assign n11252 = n11251 ^ n11243;
  assign n11257 = n11256 ^ n11252;
  assign n11215 = n11214 ^ n11175;
  assign n11216 = n11215 ^ n11142;
  assign n11244 = n11243 ^ n11213;
  assign n11245 = ~n11216 & ~n11244;
  assign n11250 = n11249 ^ n11245;
  assign n11258 = n11257 ^ n11250;
  assign n11276 = ~n11258 & ~n11275;
  assign n11296 = n11287 ^ n11276;
  assign n11299 = n11298 ^ n11296;
  assign n11268 = n11267 ^ n11258;
  assign n11294 = n11276 ^ n11268;
  assign n11292 = ~n11258 & ~n11267;
  assign n11293 = ~n11283 & n11292;
  assign n11295 = n11294 ^ n11293;
  assign n11300 = n11299 ^ n11295;
  assign n13454 = ~n11142 & ~n11300;
  assign n13401 = ~n11262 & ~n11300;
  assign n11284 = n11283 ^ n11276;
  assign n11285 = ~n11268 & ~n11284;
  assign n11286 = n11285 ^ n11267;
  assign n13286 = n11295 ^ n11286;
  assign n13336 = n11247 & ~n13286;
  assign n13402 = n13401 ^ n13336;
  assign n13455 = n13454 ^ n13402;
  assign n11288 = n11276 ^ n11267;
  assign n11289 = n11287 & n11288;
  assign n11290 = n11289 ^ n11283;
  assign n11291 = n11290 ^ n11286;
  assign n11312 = n11140 & ~n11291;
  assign n11303 = ~n11254 & ~n11291;
  assign n13452 = n11312 ^ n11303;
  assign n13407 = n11277 & n11286;
  assign n13296 = n11213 & ~n11290;
  assign n11305 = n11299 ^ n11290;
  assign n11306 = ~n11243 & ~n11305;
  assign n13340 = n13296 ^ n11306;
  assign n13408 = n13407 ^ n13340;
  assign n13453 = n13452 ^ n13408;
  assign n13456 = n13455 ^ n13453;
  assign n11315 = ~n11216 & n11299;
  assign n11301 = n11300 ^ n11291;
  assign n11313 = ~n11246 & n11301;
  assign n11314 = n11313 ^ n11312;
  assign n11316 = n11315 ^ n11314;
  assign n11308 = ~n11244 & n11299;
  assign n11307 = ~n11248 & ~n11305;
  assign n11309 = n11308 ^ n11307;
  assign n11310 = n11309 ^ n11306;
  assign n11302 = n11141 & n11301;
  assign n11304 = n11303 ^ n11302;
  assign n11311 = n11310 ^ n11304;
  assign n11317 = n11316 ^ n11311;
  assign n17274 = n13456 ^ n11317;
  assign n11786 = n9645 ^ n8785;
  assign n11784 = n8874 ^ n8711;
  assign n11785 = n11784 ^ n10392;
  assign n11787 = n11786 ^ n11785;
  assign n11781 = n9806 ^ n8947;
  assign n11779 = n8920 ^ n8832;
  assign n11778 = n8868 ^ n8848;
  assign n11780 = n11779 ^ n11778;
  assign n11782 = n11781 ^ n11780;
  assign n11788 = n11787 ^ n11782;
  assign n11794 = n9707 ^ n8832;
  assign n8926 = n8925 ^ n8785;
  assign n11792 = n11791 ^ n8926;
  assign n11793 = n11792 ^ n10400;
  assign n11795 = n11794 ^ n11793;
  assign n11821 = n9773 ^ n8925;
  assign n11818 = n8821 ^ n8811;
  assign n11820 = n11819 ^ n11818;
  assign n11822 = n11821 ^ n11820;
  assign n11809 = n9861 ^ n8874;
  assign n11808 = n11807 ^ n10368;
  assign n11810 = n11809 ^ n11808;
  assign n11805 = n9838 ^ n8248;
  assign n11804 = n11803 ^ n10387;
  assign n11806 = n11805 ^ n11804;
  assign n11811 = n11810 ^ n11806;
  assign n11823 = n11822 ^ n11811;
  assign n11841 = ~n11795 & n11823;
  assign n11826 = n11806 ^ n11782;
  assign n11799 = n8936 ^ n8894;
  assign n8948 = n8947 ^ n8785;
  assign n11798 = n11797 ^ n8948;
  assign n11800 = n11799 ^ n11798;
  assign n11790 = n9718 ^ n8906;
  assign n11796 = n11795 ^ n11790;
  assign n11801 = n11800 ^ n11796;
  assign n11827 = n11826 ^ n11801;
  assign n11830 = n11795 ^ n11787;
  assign n11831 = n11827 & n11830;
  assign n11842 = n11841 ^ n11831;
  assign n11839 = n11830 ^ n11827;
  assign n11776 = n9610 ^ n8728;
  assign n8907 = n8906 ^ n8785;
  assign n11774 = n11773 ^ n8907;
  assign n11775 = n11774 ^ n10383;
  assign n11777 = n11776 ^ n11775;
  assign n11783 = n11782 ^ n11777;
  assign n11789 = n11787 ^ n11777;
  assign n11836 = n11826 ^ n11789;
  assign n11837 = n11783 & n11836;
  assign n11814 = n11810 ^ n11782;
  assign n11815 = n11814 ^ n11801;
  assign n11816 = n11789 & n11815;
  assign n11838 = n11837 ^ n11816;
  assign n11840 = n11839 ^ n11838;
  assign n11843 = n11842 ^ n11840;
  assign n11802 = n11801 ^ n11789;
  assign n11857 = n11814 ^ n11802;
  assign n11858 = n11857 ^ n11838;
  assign n11852 = n11823 ^ n11795;
  assign n11853 = n11852 ^ n11788;
  assign n11854 = n11822 ^ n11802;
  assign n11855 = n11853 & n11854;
  assign n11846 = n11830 ^ n11783;
  assign n11847 = n11802 & n11846;
  assign n11856 = n11855 ^ n11847;
  assign n11859 = n11858 ^ n11856;
  assign n11860 = n11843 & n11859;
  assign n11828 = n11827 ^ n11823;
  assign n11824 = n11823 ^ n11777;
  assign n11825 = n11824 ^ n11789;
  assign n11834 = n11828 ^ n11825;
  assign n11829 = n11825 & n11828;
  assign n11832 = n11831 ^ n11829;
  assign n11812 = n11811 ^ n11802;
  assign n11813 = n11788 & n11812;
  assign n11817 = n11816 ^ n11813;
  assign n11833 = n11832 ^ n11817;
  assign n11835 = n11834 ^ n11833;
  assign n11844 = n11843 ^ n11835;
  assign n11875 = n11860 ^ n11844;
  assign n11849 = n11812 ^ n11788;
  assign n11845 = n11822 & n11824;
  assign n11848 = n11847 ^ n11845;
  assign n11850 = n11849 ^ n11848;
  assign n11851 = n11850 ^ n11817;
  assign n11873 = n11843 & n11851;
  assign n11874 = ~n11835 & n11873;
  assign n11876 = n11875 ^ n11874;
  assign n11864 = n11859 ^ n11851;
  assign n11871 = n11864 ^ n11860;
  assign n11869 = ~n11851 & n11859;
  assign n11870 = n11835 & n11869;
  assign n11872 = n11871 ^ n11870;
  assign n11877 = n11876 ^ n11872;
  assign n12141 = n11788 & n11877;
  assign n11950 = n11812 & n11877;
  assign n11865 = n11860 ^ n11835;
  assign n11866 = n11864 & n11865;
  assign n11867 = n11866 ^ n11851;
  assign n11882 = n11872 ^ n11867;
  assign n11885 = n11830 & n11882;
  assign n11951 = n11950 ^ n11885;
  assign n12142 = n12141 ^ n11951;
  assign n11861 = n11860 ^ n11851;
  assign n11862 = n11844 & n11861;
  assign n11863 = n11862 ^ n11835;
  assign n11868 = n11867 ^ n11863;
  assign n11899 = n11815 & n11868;
  assign n11880 = n11789 & n11868;
  assign n12139 = n11899 ^ n11880;
  assign n11956 = n11825 & n11867;
  assign n11891 = n11876 ^ n11863;
  assign n11892 = n11802 & n11891;
  assign n11890 = n11822 & n11863;
  assign n11893 = n11892 ^ n11890;
  assign n11957 = n11956 ^ n11893;
  assign n12140 = n12139 ^ n11957;
  assign n12143 = n12142 ^ n12140;
  assign n11357 = n7055 ^ n7001;
  assign n6995 = n6994 ^ n6988;
  assign n11358 = n11357 ^ n6995;
  assign n11356 = n10816 ^ n7037;
  assign n11359 = n11358 ^ n11356;
  assign n11340 = n6941 ^ n6906;
  assign n6938 = n6937 ^ n6909;
  assign n11341 = n11340 ^ n6938;
  assign n11339 = n10805 ^ n6868;
  assign n11342 = n11341 ^ n11339;
  assign n11366 = n11359 ^ n11342;
  assign n11324 = n10768 ^ n6975;
  assign n11322 = n6853 ^ n5840;
  assign n11323 = n11322 ^ n4914;
  assign n11325 = n11324 ^ n11323;
  assign n11381 = n11359 ^ n11325;
  assign n11352 = n11351 ^ n10788;
  assign n7056 = n7055 ^ n6906;
  assign n11350 = n7056 ^ n6962;
  assign n11353 = n11352 ^ n11350;
  assign n11347 = n11346 ^ n10777;
  assign n7027 = n7026 ^ n6906;
  assign n11344 = n7027 ^ n7001;
  assign n11345 = n11344 ^ n7033;
  assign n11348 = n11347 ^ n11345;
  assign n7049 = n7048 ^ n6967;
  assign n11349 = n11348 ^ n7049;
  assign n11354 = n11353 ^ n11349;
  assign n11388 = n11381 ^ n11354;
  assign n11327 = n6941 ^ n6853;
  assign n6840 = n6839 ^ n6834;
  assign n11328 = n11327 ^ n6840;
  assign n11326 = n10760 ^ n6725;
  assign n11329 = n11328 ^ n11326;
  assign n11330 = n11329 ^ n11325;
  assign n6901 = n6900 ^ n6892;
  assign n11320 = n7027 ^ n6901;
  assign n11319 = n10834 ^ n6948;
  assign n11321 = n11320 ^ n11319;
  assign n11331 = n11330 ^ n11321;
  assign n11398 = n11388 ^ n11331;
  assign n11335 = n11334 ^ n10796;
  assign n6963 = n6962 ^ n6906;
  assign n11332 = n6963 ^ n5840;
  assign n11333 = n11332 ^ n6972;
  assign n11336 = n11335 ^ n11333;
  assign n11343 = n11342 ^ n11336;
  assign n11337 = n11336 ^ n11331;
  assign n11397 = n11343 ^ n11337;
  assign n11402 = n11398 ^ n11397;
  assign n11399 = ~n11397 & ~n11398;
  assign n11361 = n11348 ^ n11342;
  assign n11391 = ~n11361 & n11388;
  assign n11400 = n11399 ^ n11391;
  assign n11370 = n11359 ^ n11329;
  assign n11371 = n11370 ^ n11354;
  assign n11372 = n11343 & n11371;
  assign n11355 = n11354 ^ n11343;
  assign n11365 = n11355 ^ n11330;
  assign n11369 = ~n11365 & n11366;
  assign n11373 = n11372 ^ n11369;
  assign n11401 = n11400 ^ n11373;
  assign n11403 = n11402 ^ n11401;
  assign n11392 = ~n11331 & n11348;
  assign n11393 = n11392 ^ n11391;
  assign n11389 = n11388 ^ n11361;
  assign n11360 = n11359 ^ n11336;
  assign n11382 = n11381 ^ n11343;
  assign n11383 = n11360 & ~n11382;
  assign n11384 = n11383 ^ n11372;
  assign n11390 = n11389 ^ n11384;
  assign n11394 = n11393 ^ n11390;
  assign n11410 = n11403 ^ n11394;
  assign n11380 = n11370 ^ n11355;
  assign n11385 = n11384 ^ n11380;
  assign n11375 = n11348 ^ n11331;
  assign n11376 = n11375 ^ n11366;
  assign n11377 = n11355 ^ n11321;
  assign n11378 = n11376 & n11377;
  assign n11362 = n11361 ^ n11360;
  assign n11363 = ~n11355 & ~n11362;
  assign n11379 = n11378 ^ n11363;
  assign n11386 = n11385 ^ n11379;
  assign n11395 = n11386 & ~n11394;
  assign n11411 = n11410 ^ n11395;
  assign n11367 = n11366 ^ n11365;
  assign n11338 = ~n11321 & ~n11337;
  assign n11364 = n11363 ^ n11338;
  assign n11368 = n11367 ^ n11364;
  assign n11374 = n11373 ^ n11368;
  assign n11408 = ~n11374 & ~n11394;
  assign n11409 = ~n11403 & n11408;
  assign n11412 = n11411 ^ n11409;
  assign n11404 = n11374 & n11386;
  assign n11405 = n11403 & n11404;
  assign n11387 = n11386 ^ n11374;
  assign n11396 = n11395 ^ n11387;
  assign n11406 = n11405 ^ n11396;
  assign n11422 = n11412 ^ n11406;
  assign n12041 = n11366 & n11422;
  assign n11928 = ~n11365 & n11422;
  assign n11418 = n11403 ^ n11395;
  assign n11419 = ~n11387 & n11418;
  assign n11420 = n11419 ^ n11374;
  assign n11907 = n11420 ^ n11406;
  assign n11910 = ~n11361 & n11907;
  assign n11929 = n11928 ^ n11910;
  assign n12042 = n12041 ^ n11929;
  assign n11415 = n11395 ^ n11374;
  assign n11416 = ~n11410 & ~n11415;
  assign n11417 = n11416 ^ n11403;
  assign n11421 = n11420 ^ n11417;
  assign n11920 = n11371 & ~n11421;
  assign n11425 = n11343 & ~n11421;
  assign n12039 = n11920 ^ n11425;
  assign n11964 = ~n11397 & ~n11420;
  assign n11432 = n11417 ^ n11412;
  assign n11914 = ~n11355 & ~n11432;
  assign n11429 = ~n11321 & n11417;
  assign n11915 = n11914 ^ n11429;
  assign n11965 = n11964 ^ n11915;
  assign n12040 = n12039 ^ n11965;
  assign n12043 = n12042 ^ n12040;
  assign n12144 = n12143 ^ n12043;
  assign n11679 = n11678 ^ n7953;
  assign n7940 = n7939 ^ n7545;
  assign n11676 = n11675 ^ n7940;
  assign n11677 = n11676 ^ n7885;
  assign n11680 = n11679 ^ n11677;
  assign n11657 = n11656 ^ n8001;
  assign n11655 = n11654 ^ n10615;
  assign n11658 = n11657 ^ n11655;
  assign n11652 = n11651 ^ n7824;
  assign n11650 = n10624 ^ n8008;
  assign n11653 = n11652 ^ n11650;
  assign n11659 = n11658 ^ n11653;
  assign n11648 = n11647 ^ n7990;
  assign n11646 = n11645 ^ n10620;
  assign n11649 = n11648 ^ n11646;
  assign n11660 = n11659 ^ n11649;
  assign n11710 = n11680 ^ n11660;
  assign n11693 = n11692 ^ n7891;
  assign n11691 = n11690 ^ n10631;
  assign n11694 = n11693 ^ n11691;
  assign n11672 = n11671 ^ n7800;
  assign n11670 = n11669 ^ n10611;
  assign n11673 = n11672 ^ n11670;
  assign n11701 = n11694 ^ n11673;
  assign n11711 = n11710 ^ n11701;
  assign n11665 = n11664 ^ n7278;
  assign n7554 = n7553 ^ n7545;
  assign n11662 = n11661 ^ n7554;
  assign n11663 = n11662 ^ n7852;
  assign n11666 = n11665 ^ n11663;
  assign n11674 = n11673 ^ n11666;
  assign n11667 = n11666 ^ n11660;
  assign n11733 = n11674 ^ n11667;
  assign n11716 = n11694 ^ n11653;
  assign n11686 = n11685 ^ n7921;
  assign n7974 = n7973 ^ n7545;
  assign n11684 = n11683 ^ n7974;
  assign n11687 = n11686 ^ n11684;
  assign n11682 = n11681 ^ n11680;
  assign n11688 = n11687 ^ n11682;
  assign n11723 = n11716 ^ n11688;
  assign n11732 = n11723 ^ n11660;
  assign n11737 = n11733 ^ n11732;
  assign n11734 = ~n11732 & ~n11733;
  assign n11696 = n11680 ^ n11673;
  assign n11726 = n11696 & n11723;
  assign n11735 = n11734 ^ n11726;
  assign n11705 = n11694 ^ n11658;
  assign n11706 = n11705 ^ n11688;
  assign n11707 = n11674 & n11706;
  assign n11689 = n11688 ^ n11674;
  assign n11700 = n11689 ^ n11659;
  assign n11704 = n11700 & ~n11701;
  assign n11708 = n11707 ^ n11704;
  assign n11736 = n11735 ^ n11708;
  assign n11738 = n11737 ^ n11736;
  assign n11727 = ~n11660 & ~n11680;
  assign n11728 = n11727 ^ n11726;
  assign n11724 = n11723 ^ n11696;
  assign n11695 = n11694 ^ n11666;
  assign n11717 = n11716 ^ n11674;
  assign n11718 = ~n11695 & n11717;
  assign n11719 = n11718 ^ n11707;
  assign n11725 = n11724 ^ n11719;
  assign n11729 = n11728 ^ n11725;
  assign n11746 = n11738 ^ n11729;
  assign n11715 = n11705 ^ n11689;
  assign n11720 = n11719 ^ n11715;
  assign n11712 = n11689 ^ n11649;
  assign n11713 = n11711 & ~n11712;
  assign n11697 = n11696 ^ n11695;
  assign n11698 = n11689 & ~n11697;
  assign n11714 = n11713 ^ n11698;
  assign n11721 = n11720 ^ n11714;
  assign n11730 = n11721 & n11729;
  assign n11754 = n11746 ^ n11730;
  assign n11702 = n11701 ^ n11700;
  assign n11668 = ~n11649 & ~n11667;
  assign n11699 = n11698 ^ n11668;
  assign n11703 = n11702 ^ n11699;
  assign n11709 = n11708 ^ n11703;
  assign n11752 = ~n11709 & n11729;
  assign n11753 = ~n11738 & n11752;
  assign n11755 = n11754 ^ n11753;
  assign n11981 = n11711 & n11755;
  assign n11739 = n11709 & n11721;
  assign n11740 = n11738 & n11739;
  assign n11722 = n11721 ^ n11709;
  assign n11731 = n11730 ^ n11722;
  assign n11741 = n11740 ^ n11731;
  assign n11756 = n11755 ^ n11741;
  assign n11747 = n11730 ^ n11709;
  assign n11748 = n11746 & ~n11747;
  assign n11749 = n11748 ^ n11738;
  assign n11743 = n11738 ^ n11730;
  assign n11744 = ~n11722 & n11743;
  assign n11745 = n11744 ^ n11709;
  assign n11750 = n11749 ^ n11745;
  assign n11757 = n11756 ^ n11750;
  assign n11758 = ~n11695 & n11757;
  assign n11751 = n11674 & ~n11750;
  assign n11759 = n11758 ^ n11751;
  assign n12136 = n11981 ^ n11759;
  assign n12060 = n11706 & ~n11750;
  assign n11765 = n11717 & n11757;
  assign n12134 = n12060 ^ n11765;
  assign n11986 = n11755 ^ n11749;
  assign n12019 = n11689 & n11986;
  assign n11988 = ~n11712 & n11755;
  assign n11987 = ~n11697 & n11986;
  assign n11989 = n11988 ^ n11987;
  assign n12096 = n12019 ^ n11989;
  assign n12135 = n12134 ^ n12096;
  assign n12137 = n12136 ^ n12135;
  assign n11573 = n10937 ^ n9666;
  assign n11571 = n9767 ^ n9636;
  assign n9659 = n9658 ^ n9162;
  assign n11572 = n11571 ^ n9659;
  assign n11574 = n11573 ^ n11572;
  assign n9624 = n9623 ^ n9620;
  assign n11559 = n10773 ^ n9624;
  assign n11560 = n11559 ^ n9855;
  assign n11561 = n11560 ^ n10935;
  assign n9849 = n9848 ^ n9832;
  assign n11556 = n9849 ^ n9820;
  assign n11557 = n11556 ^ n10802;
  assign n11558 = n11557 ^ n10919;
  assign n11562 = n11561 ^ n11558;
  assign n11575 = n11574 ^ n11562;
  assign n11534 = n10922 ^ n9696;
  assign n11532 = n9796 ^ n9659;
  assign n11531 = n11530 ^ n9678;
  assign n11533 = n11532 ^ n11531;
  assign n11535 = n11534 ^ n11533;
  assign n11588 = n11575 ^ n11535;
  assign n11537 = n10783 ^ n9752;
  assign n11538 = n11537 ^ n9744;
  assign n11539 = n11538 ^ n9785;
  assign n11540 = n11539 ^ n10920;
  assign n11528 = n10926 ^ n9287;
  assign n11526 = n9620 ^ n9162;
  assign n11525 = n9852 ^ n9630;
  assign n11527 = n11526 ^ n11525;
  assign n11529 = n11528 ^ n11527;
  assign n11541 = n11540 ^ n11529;
  assign n11589 = n11588 ^ n11541;
  assign n11609 = ~n11535 & n11575;
  assign n11536 = n11535 ^ n11529;
  assign n11569 = n11558 ^ n11540;
  assign n9745 = n9744 ^ n9162;
  assign n11552 = n9745 ^ n9153;
  assign n11551 = n11550 ^ n9733;
  assign n11553 = n11552 ^ n11551;
  assign n11548 = n10923 ^ n9278;
  assign n11549 = n11548 ^ n11535;
  assign n11554 = n11553 ^ n11549;
  assign n11570 = n11569 ^ n11554;
  assign n11580 = n11536 & n11570;
  assign n11610 = n11609 ^ n11580;
  assign n11607 = n11570 ^ n11536;
  assign n9815 = n9814 ^ n9524;
  assign n9163 = n9162 ^ n9153;
  assign n11542 = n9815 ^ n9163;
  assign n11544 = n11543 ^ n11542;
  assign n11545 = n11544 ^ n9401;
  assign n11546 = n11545 ^ n10927;
  assign n11585 = n11546 ^ n11540;
  assign n11547 = n11546 ^ n11529;
  assign n11594 = n11569 ^ n11547;
  assign n11595 = n11585 & n11594;
  assign n11565 = n11561 ^ n11540;
  assign n11566 = n11565 ^ n11554;
  assign n11567 = n11547 & n11566;
  assign n11596 = n11595 ^ n11567;
  assign n11608 = n11607 ^ n11596;
  assign n11611 = n11610 ^ n11608;
  assign n11577 = n11575 ^ n11546;
  assign n11578 = n11577 ^ n11547;
  assign n11576 = n11575 ^ n11570;
  assign n11583 = n11578 ^ n11576;
  assign n11579 = n11576 & n11578;
  assign n11581 = n11580 ^ n11579;
  assign n11555 = n11554 ^ n11547;
  assign n11563 = n11562 ^ n11555;
  assign n11564 = n11541 & n11563;
  assign n11568 = n11567 ^ n11564;
  assign n11582 = n11581 ^ n11568;
  assign n11584 = n11583 ^ n11582;
  assign n11622 = n11611 ^ n11584;
  assign n11593 = n11565 ^ n11555;
  assign n11597 = n11596 ^ n11593;
  assign n11590 = n11574 ^ n11555;
  assign n11591 = n11589 & n11590;
  assign n11586 = n11585 ^ n11536;
  assign n11587 = n11555 & n11586;
  assign n11592 = n11591 ^ n11587;
  assign n11598 = n11597 ^ n11592;
  assign n11612 = n11598 & n11611;
  assign n11623 = n11622 ^ n11612;
  assign n11601 = n11563 ^ n11541;
  assign n11599 = n11574 & n11577;
  assign n11600 = n11599 ^ n11587;
  assign n11602 = n11601 ^ n11600;
  assign n11603 = n11602 ^ n11568;
  assign n11620 = n11603 & n11611;
  assign n11621 = ~n11584 & n11620;
  assign n11624 = n11623 ^ n11621;
  assign n11970 = n11589 & n11624;
  assign n11628 = n11612 ^ n11603;
  assign n11629 = n11622 & n11628;
  assign n11630 = n11629 ^ n11584;
  assign n11606 = n11603 ^ n11598;
  assign n11615 = n11612 ^ n11584;
  assign n11616 = n11606 & n11615;
  assign n11617 = n11616 ^ n11603;
  assign n11631 = n11630 ^ n11617;
  assign n11641 = n11547 & n11631;
  assign n11613 = n11612 ^ n11606;
  assign n11604 = n11598 & ~n11603;
  assign n11605 = n11584 & n11604;
  assign n11614 = n11613 ^ n11605;
  assign n11625 = n11624 ^ n11614;
  assign n11632 = n11631 ^ n11625;
  assign n11640 = n11585 & n11632;
  assign n11642 = n11641 ^ n11640;
  assign n12132 = n11970 ^ n11642;
  assign n12054 = n11566 & n11631;
  assign n11633 = n11594 & n11632;
  assign n12130 = n12054 ^ n11633;
  assign n11975 = n11630 ^ n11624;
  assign n12030 = n11555 & n11975;
  assign n11977 = n11590 & n11624;
  assign n11976 = n11586 & n11975;
  assign n11978 = n11977 ^ n11976;
  assign n12099 = n12030 ^ n11978;
  assign n12131 = n12130 ^ n12099;
  assign n12133 = n12132 ^ n12131;
  assign n12138 = n12137 ^ n12133;
  assign n12145 = n12144 ^ n12138;
  assign n11423 = n11422 ^ n11421;
  assign n11424 = n11360 & ~n11423;
  assign n11426 = n11425 ^ n11424;
  assign n11413 = n11376 & ~n11412;
  assign n12120 = n11426 ^ n11413;
  assign n11433 = ~n11362 & ~n11432;
  assign n11431 = n11377 & ~n11412;
  assign n11434 = n11433 ^ n11431;
  assign n12072 = n11914 ^ n11434;
  assign n11919 = ~n11382 & ~n11423;
  assign n11921 = n11920 ^ n11919;
  assign n12119 = n12072 ^ n11921;
  assign n12121 = n12120 ^ n12119;
  assign n12129 = n12128 ^ n12121;
  assign n12146 = n12145 ^ n12129;
  assign n11407 = ~n11331 & ~n11406;
  assign n11414 = n11413 ^ n11407;
  assign n12073 = n12072 ^ n11414;
  assign n11908 = n11388 & n11907;
  assign n11909 = n11908 ^ n11426;
  assign n12074 = n12073 ^ n11909;
  assign n12067 = n11854 & n11876;
  assign n11896 = n11846 & n11891;
  assign n12068 = n12067 ^ n11896;
  assign n12069 = n12068 ^ n11892;
  assign n11902 = n11853 & n11876;
  assign n11901 = n11823 & n11872;
  assign n11903 = n11902 ^ n11901;
  assign n12070 = n12069 ^ n11903;
  assign n11883 = n11827 & n11882;
  assign n11878 = n11877 ^ n11868;
  assign n11879 = n11783 & n11878;
  assign n11881 = n11880 ^ n11879;
  assign n11884 = n11883 ^ n11881;
  assign n12071 = n12070 ^ n11884;
  assign n12075 = n12074 ^ n12071;
  assign n12063 = ~n11701 & ~n11756;
  assign n11763 = n11700 & ~n11756;
  assign n11761 = n11745 ^ n11741;
  assign n11762 = n11696 & n11761;
  assign n11764 = n11763 ^ n11762;
  assign n12064 = n12063 ^ n11764;
  assign n12061 = n12060 ^ n11751;
  assign n12021 = ~n11733 & ~n11745;
  assign n11984 = ~n11649 & n11749;
  assign n12020 = n12019 ^ n11984;
  assign n12022 = n12021 ^ n12020;
  assign n12062 = n12061 ^ n12022;
  assign n12065 = n12064 ^ n12062;
  assign n12057 = n11541 & n11625;
  assign n11626 = n11563 & n11625;
  assign n11618 = n11617 ^ n11614;
  assign n11619 = n11536 & n11618;
  assign n11627 = n11626 ^ n11619;
  assign n12058 = n12057 ^ n11627;
  assign n12055 = n12054 ^ n11641;
  assign n12032 = n11578 & n11617;
  assign n11973 = n11574 & n11630;
  assign n12031 = n12030 ^ n11973;
  assign n12033 = n12032 ^ n12031;
  assign n12056 = n12055 ^ n12033;
  assign n12059 = n12058 ^ n12056;
  assign n12066 = n12065 ^ n12059;
  assign n12076 = n12075 ^ n12066;
  assign n12053 = n12052 ^ n12043;
  assign n12077 = n12076 ^ n12053;
  assign n12147 = n12146 ^ n12077;
  assign n11922 = n11921 ^ n11414;
  assign n11918 = n11909 ^ n11433;
  assign n11923 = n11922 ^ n11918;
  assign n11912 = n11375 & ~n11406;
  assign n11428 = ~n11398 & ~n11420;
  assign n11913 = n11912 ^ n11428;
  assign n11916 = n11915 ^ n11913;
  assign n11911 = n11910 ^ n11909;
  assign n11917 = n11916 ^ n11911;
  assign n11924 = n11923 ^ n11917;
  assign n11898 = n11836 & n11878;
  assign n11900 = n11899 ^ n11898;
  assign n11904 = n11903 ^ n11900;
  assign n11897 = n11896 ^ n11884;
  assign n11905 = n11904 ^ n11897;
  assign n12086 = n11924 ^ n11905;
  assign n11636 = n11576 & n11617;
  assign n11635 = n11588 & n11614;
  assign n11637 = n11636 ^ n11635;
  assign n12084 = n12031 ^ n11637;
  assign n12025 = n11570 & n11618;
  assign n12026 = n12025 ^ n11642;
  assign n12083 = n12026 ^ n11619;
  assign n12085 = n12084 ^ n12083;
  assign n12087 = n12086 ^ n12085;
  assign n11768 = ~n11732 & ~n11745;
  assign n11767 = ~n11710 & ~n11741;
  assign n11769 = n11768 ^ n11767;
  assign n12081 = n12020 ^ n11769;
  assign n12014 = n11723 & n11761;
  assign n12015 = n12014 ^ n11759;
  assign n12080 = n12015 ^ n11762;
  assign n12082 = n12081 ^ n12080;
  assign n12088 = n12087 ^ n12082;
  assign n12095 = n12094 ^ n12088;
  assign n12148 = n12147 ^ n12095;
  assign n11930 = n11929 ^ n11919;
  assign n11931 = n11930 ^ n11913;
  assign n11927 = n11426 ^ n11407;
  assign n11932 = n11931 ^ n11927;
  assign n11947 = n11946 ^ n11932;
  assign n11888 = n11828 & n11867;
  assign n11887 = n11852 & n11872;
  assign n11889 = n11888 ^ n11887;
  assign n11894 = n11893 ^ n11889;
  assign n11886 = n11885 ^ n11884;
  assign n11895 = n11894 ^ n11886;
  assign n11906 = n11905 ^ n11895;
  assign n11925 = n11924 ^ n11906;
  assign n11766 = n11765 ^ n11764;
  assign n11770 = n11769 ^ n11766;
  assign n11742 = ~n11660 & ~n11741;
  assign n11760 = n11759 ^ n11742;
  assign n11771 = n11770 ^ n11760;
  assign n11639 = n11575 & n11614;
  assign n11643 = n11642 ^ n11639;
  assign n11634 = n11633 ^ n11627;
  assign n11638 = n11637 ^ n11634;
  assign n11644 = n11643 ^ n11638;
  assign n11772 = n11771 ^ n11644;
  assign n11926 = n11925 ^ n11772;
  assign n11948 = n11947 ^ n11926;
  assign n12188 = n12148 ^ n11948;
  assign n12166 = n11902 ^ n11881;
  assign n12165 = n12069 ^ n11900;
  assign n12167 = n12166 ^ n12165;
  assign n12168 = n12167 ^ n12121;
  assign n11971 = n11970 ^ n11639;
  assign n12162 = n12130 ^ n11971;
  assign n12161 = n12026 ^ n11976;
  assign n12163 = n12162 ^ n12161;
  assign n11982 = n11981 ^ n11742;
  assign n12159 = n12134 ^ n11982;
  assign n12158 = n12015 ^ n11987;
  assign n12160 = n12159 ^ n12158;
  assign n12164 = n12163 ^ n12160;
  assign n12169 = n12168 ^ n12164;
  assign n12157 = n12156 ^ n11923;
  assign n12170 = n12169 ^ n12157;
  assign n12028 = n11577 & n11630;
  assign n12029 = n12028 ^ n11971;
  assign n12034 = n12033 ^ n12029;
  assign n12027 = n12026 ^ n11634;
  assign n12035 = n12034 ^ n12027;
  assign n12017 = ~n11667 & n11749;
  assign n12018 = n12017 ^ n11982;
  assign n12023 = n12022 ^ n12018;
  assign n12016 = n12015 ^ n11766;
  assign n12024 = n12023 ^ n12016;
  assign n12036 = n12035 ^ n12024;
  assign n12011 = n11901 ^ n11881;
  assign n11952 = n11951 ^ n11898;
  assign n12010 = n11952 ^ n11889;
  assign n12012 = n12011 ^ n12010;
  assign n12013 = n12012 ^ n11932;
  assign n12037 = n12036 ^ n12013;
  assign n11962 = ~n11337 & n11417;
  assign n11963 = n11962 ^ n11414;
  assign n11966 = n11965 ^ n11963;
  assign n11961 = n11930 ^ n11909;
  assign n11967 = n11966 ^ n11961;
  assign n12009 = n12008 ^ n11967;
  assign n12038 = n12037 ^ n12009;
  assign n12179 = n12170 ^ n12038;
  assign n12189 = n12188 ^ n12179;
  assign n12078 = n12077 ^ n12038;
  assign n11985 = n11984 ^ n11768;
  assign n11990 = n11989 ^ n11985;
  assign n11983 = n11982 ^ n11759;
  assign n11991 = n11990 ^ n11983;
  assign n11974 = n11973 ^ n11636;
  assign n11979 = n11978 ^ n11974;
  assign n11972 = n11971 ^ n11642;
  assign n11980 = n11979 ^ n11972;
  assign n11992 = n11991 ^ n11980;
  assign n11968 = n11967 ^ n11923;
  assign n11954 = n11824 & n11863;
  assign n11955 = n11954 ^ n11903;
  assign n11958 = n11957 ^ n11955;
  assign n11953 = n11952 ^ n11884;
  assign n11959 = n11958 ^ n11953;
  assign n11960 = n11959 ^ n11905;
  assign n11969 = n11968 ^ n11960;
  assign n11993 = n11992 ^ n11969;
  assign n11430 = n11429 ^ n11428;
  assign n11435 = n11434 ^ n11430;
  assign n11427 = n11426 ^ n11414;
  assign n11436 = n11435 ^ n11427;
  assign n11524 = n11523 ^ n11436;
  assign n11949 = n11948 ^ n11524;
  assign n11994 = n11993 ^ n11949;
  assign n12079 = n12078 ^ n11994;
  assign n12208 = n12148 ^ n12079;
  assign n12117 = n12116 ^ n12074;
  assign n12108 = n11923 ^ n11436;
  assign n12104 = n11890 ^ n11888;
  assign n12105 = n12104 ^ n12068;
  assign n12103 = n11903 ^ n11881;
  assign n12106 = n12105 ^ n12103;
  assign n12107 = n12106 ^ n11905;
  assign n12109 = n12108 ^ n12107;
  assign n12100 = n12099 ^ n11971;
  assign n12101 = n12100 ^ n12026;
  assign n12097 = n12096 ^ n11982;
  assign n12098 = n12097 ^ n12015;
  assign n12102 = n12101 ^ n12098;
  assign n12110 = n12109 ^ n12102;
  assign n12118 = n12117 ^ n12110;
  assign n12171 = n12170 ^ n12118;
  assign n12149 = n12148 ^ n12118;
  assign n12207 = n12171 ^ n12149;
  assign n12212 = n12208 ^ n12207;
  assign n12209 = ~n12207 & ~n12208;
  assign n12174 = n12170 ^ n11948;
  assign n12202 = n12079 & ~n12174;
  assign n12210 = n12209 ^ n12202;
  assign n12183 = n12146 ^ n12038;
  assign n12184 = n12183 ^ n11994;
  assign n12185 = n12171 & n12184;
  assign n12172 = n12171 ^ n11994;
  assign n12178 = n12172 ^ n12147;
  assign n12182 = ~n12178 & n12179;
  assign n12186 = n12185 ^ n12182;
  assign n12211 = n12210 ^ n12186;
  assign n12213 = n12212 ^ n12211;
  assign n12203 = n11948 & ~n12148;
  assign n12204 = n12203 ^ n12202;
  assign n12200 = n12174 ^ n12079;
  assign n12173 = n12118 ^ n12038;
  assign n12194 = n12171 ^ n12078;
  assign n12195 = n12173 & ~n12194;
  assign n12196 = n12195 ^ n12185;
  assign n12201 = n12200 ^ n12196;
  assign n12205 = n12204 ^ n12201;
  assign n12223 = n12213 ^ n12205;
  assign n12193 = n12183 ^ n12172;
  assign n12197 = n12196 ^ n12193;
  assign n12190 = n12172 ^ n12095;
  assign n12191 = n12189 & n12190;
  assign n12175 = n12174 ^ n12173;
  assign n12176 = ~n12172 & ~n12175;
  assign n12192 = n12191 ^ n12176;
  assign n12198 = n12197 ^ n12192;
  assign n12206 = n12198 & ~n12205;
  assign n12231 = n12223 ^ n12206;
  assign n12180 = n12179 ^ n12178;
  assign n12150 = ~n12095 & ~n12149;
  assign n12177 = n12176 ^ n12150;
  assign n12181 = n12180 ^ n12177;
  assign n12187 = n12186 ^ n12181;
  assign n12229 = ~n12187 & ~n12205;
  assign n12230 = ~n12213 & n12229;
  assign n12232 = n12231 ^ n12230;
  assign n12242 = n12189 & ~n12232;
  assign n12218 = n12187 & n12198;
  assign n12219 = n12213 & n12218;
  assign n12199 = n12198 ^ n12187;
  assign n12217 = n12206 ^ n12199;
  assign n12220 = n12219 ^ n12217;
  assign n12233 = n12232 ^ n12220;
  assign n12224 = n12206 ^ n12187;
  assign n12225 = ~n12223 & ~n12224;
  assign n12226 = n12225 ^ n12213;
  assign n12214 = n12213 ^ n12206;
  assign n12215 = ~n12199 & n12214;
  assign n12216 = n12215 ^ n12187;
  assign n12227 = n12226 ^ n12216;
  assign n12234 = n12233 ^ n12227;
  assign n12235 = n12173 & ~n12234;
  assign n12228 = n12171 & ~n12227;
  assign n12236 = n12235 ^ n12228;
  assign n13459 = n12242 ^ n12236;
  assign n12238 = n12232 ^ n12226;
  assign n13306 = ~n12172 & ~n12238;
  assign n13304 = n12190 & ~n12232;
  assign n12239 = ~n12175 & ~n12238;
  assign n13305 = n13304 ^ n12239;
  assign n13307 = n13306 ^ n13305;
  assign n12245 = n12184 & ~n12227;
  assign n12244 = ~n12194 & ~n12234;
  assign n12246 = n12245 ^ n12244;
  assign n13458 = n13307 ^ n12246;
  assign n13460 = n13459 ^ n13458;
  assign n8911 = n8910 ^ n8907;
  assign n8896 = n8895 ^ n8749;
  assign n8902 = n8901 ^ n8896;
  assign n8912 = n8911 ^ n8902;
  assign n8880 = n8815 ^ n8469;
  assign n8888 = n8887 ^ n8880;
  assign n8879 = n8878 ^ n8874;
  assign n8889 = n8888 ^ n8879;
  assign n8913 = n8912 ^ n8889;
  assign n8956 = n8955 ^ n8894;
  assign n8954 = n8953 ^ n8948;
  assign n8957 = n8956 ^ n8954;
  assign n8931 = n8930 ^ n8926;
  assign n8914 = n8851 ^ n8822;
  assign n8922 = n8921 ^ n8914;
  assign n8932 = n8931 ^ n8922;
  assign n8942 = n8941 ^ n8932;
  assign n8958 = n8957 ^ n8942;
  assign n8959 = n8958 ^ n8913;
  assign n8750 = n8749 ^ n8456;
  assign n8778 = n8777 ^ n8750;
  assign n8743 = n8742 ^ n8728;
  assign n8779 = n8778 ^ n8743;
  assign n8470 = n8469 ^ n8456;
  assign n8713 = n8712 ^ n8470;
  assign n8342 = n8341 ^ n8248;
  assign n8714 = n8713 ^ n8342;
  assign n8780 = n8779 ^ n8714;
  assign n8960 = n8959 ^ n8780;
  assign n8852 = n8851 ^ n8848;
  assign n8870 = n8869 ^ n8852;
  assign n8842 = n8841 ^ n8832;
  assign n8871 = n8870 ^ n8842;
  assign n8890 = n8889 ^ n8871;
  assign n8994 = n8960 ^ n8890;
  assign n8823 = n8822 ^ n8812;
  assign n8795 = n8794 ^ n8785;
  assign n8824 = n8823 ^ n8795;
  assign n8825 = n8824 ^ n8780;
  assign n8966 = n8912 ^ n8825;
  assign n8992 = n8824 & n8966;
  assign n8978 = n8912 ^ n8871;
  assign n8972 = n8932 ^ n8889;
  assign n8979 = n8978 ^ n8972;
  assign n8980 = n8959 & n8979;
  assign n8993 = n8992 ^ n8980;
  assign n8995 = n8994 ^ n8993;
  assign n8962 = n8871 ^ n8714;
  assign n8963 = n8962 ^ n8958;
  assign n8964 = n8913 & n8963;
  assign n8961 = n8890 & n8960;
  assign n8965 = n8964 ^ n8961;
  assign n8996 = n8995 ^ n8965;
  assign n8968 = n8871 ^ n8779;
  assign n8987 = n8968 ^ n8913;
  assign n8988 = n8978 & n8987;
  assign n8989 = n8988 ^ n8964;
  assign n8986 = n8962 ^ n8959;
  assign n8990 = n8989 ^ n8986;
  assign n8981 = n8932 ^ n8825;
  assign n8982 = n8981 ^ n8890;
  assign n8983 = n8959 ^ n8824;
  assign n8984 = n8982 & n8983;
  assign n8985 = n8984 ^ n8980;
  assign n8991 = n8990 ^ n8985;
  assign n8999 = n8996 ^ n8991;
  assign n9002 = n8825 & ~n8932;
  assign n8969 = n8968 ^ n8958;
  assign n8973 = n8969 & n8972;
  assign n9003 = n9002 ^ n8973;
  assign n9000 = n8972 ^ n8969;
  assign n9001 = n9000 ^ n8989;
  assign n9004 = n9003 ^ n9001;
  assign n9005 = n8991 & n9004;
  assign n8970 = n8969 ^ n8825;
  assign n8967 = n8966 ^ n8913;
  assign n8976 = n8970 ^ n8967;
  assign n8971 = n8967 & n8970;
  assign n8974 = n8973 ^ n8971;
  assign n8975 = n8974 ^ n8965;
  assign n8977 = n8976 ^ n8975;
  assign n9027 = n9005 ^ n8977;
  assign n9028 = n8999 & n9027;
  assign n9029 = n9028 ^ n8996;
  assign n9011 = n9004 ^ n8977;
  assign n9016 = n9005 ^ n8996;
  assign n9017 = n9011 & n9016;
  assign n9018 = n9017 ^ n8977;
  assign n9030 = n9029 ^ n9018;
  assign n9033 = n8913 & n9030;
  assign n9012 = n9011 ^ n9005;
  assign n9009 = n8996 & n9004;
  assign n9010 = ~n8977 & n9009;
  assign n9013 = n9012 ^ n9010;
  assign n9006 = n9005 ^ n8999;
  assign n8997 = n8991 & ~n8996;
  assign n8998 = n8977 & n8997;
  assign n9007 = n9006 ^ n8998;
  assign n9026 = n9013 ^ n9007;
  assign n9031 = n9030 ^ n9026;
  assign n9032 = n8978 & n9031;
  assign n9034 = n9033 ^ n9032;
  assign n9014 = n8982 & n9013;
  assign n10252 = n9034 ^ n9014;
  assign n10071 = n8987 & n9031;
  assign n10070 = n8963 & n9030;
  assign n10072 = n10071 ^ n10070;
  assign n9019 = n9018 ^ n9013;
  assign n9023 = n8959 & n9019;
  assign n9021 = n8983 & n9013;
  assign n9020 = n8979 & n9019;
  assign n9022 = n9021 ^ n9020;
  assign n9024 = n9023 ^ n9022;
  assign n10251 = n10072 ^ n9024;
  assign n10253 = n10252 ^ n10251;
  assign n9649 = n9648 ^ n9287;
  assign n9638 = n9637 ^ n9624;
  assign n9650 = n9649 ^ n9638;
  assign n9614 = n9613 ^ n9524;
  assign n9289 = n9288 ^ n9163;
  assign n9520 = n9519 ^ n9289;
  assign n9615 = n9614 ^ n9520;
  assign n9651 = n9650 ^ n9615;
  assign n9865 = n9864 ^ n9623;
  assign n9857 = n9856 ^ n9849;
  assign n9866 = n9865 ^ n9857;
  assign n9810 = n9809 ^ n9752;
  assign n9797 = n9796 ^ n9696;
  assign n9793 = n9792 ^ n9785;
  assign n9798 = n9797 ^ n9793;
  assign n9811 = n9810 ^ n9798;
  assign n9870 = n9866 ^ n9811;
  assign n9754 = n9753 ^ n9745;
  assign n9734 = n9733 ^ n9728;
  assign n9755 = n9754 ^ n9734;
  assign n9722 = n9721 ^ n9278;
  assign n9711 = n9710 ^ n9696;
  assign n9668 = n9667 ^ n9659;
  assign n9690 = n9689 ^ n9668;
  assign n9712 = n9711 ^ n9690;
  assign n9723 = n9722 ^ n9712;
  assign n9756 = n9755 ^ n9723;
  assign n9757 = n9756 ^ n9651;
  assign n9909 = n9870 ^ n9757;
  assign n9887 = n9811 ^ n9615;
  assign n9842 = n9841 ^ n9832;
  assign n9827 = n9826 ^ n9815;
  assign n9843 = n9842 ^ n9827;
  assign n9877 = n9843 ^ n9811;
  assign n9888 = n9877 ^ n9651;
  assign n9889 = n9887 & n9888;
  assign n9871 = n9870 ^ n9756;
  assign n9872 = n9651 & n9871;
  assign n9890 = n9889 ^ n9872;
  assign n9910 = n9909 ^ n9890;
  assign n9758 = n9667 ^ n9162;
  assign n9763 = n9762 ^ n9758;
  assign n9768 = n9767 ^ n9763;
  assign n9777 = n9776 ^ n9768;
  assign n9778 = n9777 ^ n9757;
  assign n9867 = n9866 ^ n9843;
  assign n9874 = n9867 ^ n9777;
  assign n9905 = n9874 ^ n9712;
  assign n9812 = n9811 ^ n9650;
  assign n9906 = n9905 ^ n9812;
  assign n9907 = n9778 & n9906;
  assign n9881 = n9712 ^ n9650;
  assign n9897 = n9887 ^ n9881;
  assign n9898 = n9757 & n9897;
  assign n9908 = n9907 ^ n9898;
  assign n9911 = n9910 ^ n9908;
  assign n9868 = n9867 ^ n9757;
  assign n9900 = n9868 ^ n9812;
  assign n9875 = n9874 ^ n9615;
  assign n9896 = n9777 & n9875;
  assign n9899 = n9898 ^ n9896;
  assign n9901 = n9900 ^ n9899;
  assign n9869 = n9812 & n9868;
  assign n9873 = n9872 ^ n9869;
  assign n9902 = n9901 ^ n9873;
  assign n9927 = n9911 ^ n9902;
  assign n9893 = ~n9712 & n9874;
  assign n9878 = n9877 ^ n9756;
  assign n9882 = n9878 & n9881;
  assign n9894 = n9893 ^ n9882;
  assign n9891 = n9881 ^ n9878;
  assign n9892 = n9891 ^ n9890;
  assign n9895 = n9894 ^ n9892;
  assign n9912 = n9895 & n9911;
  assign n9879 = n9878 ^ n9874;
  assign n9876 = n9875 ^ n9651;
  assign n9885 = n9879 ^ n9876;
  assign n9880 = n9876 & n9879;
  assign n9883 = n9882 ^ n9880;
  assign n9884 = n9883 ^ n9873;
  assign n9886 = n9885 ^ n9884;
  assign n9935 = n9912 ^ n9886;
  assign n9936 = n9927 & n9935;
  assign n9937 = n9936 ^ n9902;
  assign n9913 = n9895 ^ n9886;
  assign n9917 = n9912 ^ n9902;
  assign n9918 = n9913 & n9917;
  assign n9919 = n9918 ^ n9886;
  assign n9938 = n9937 ^ n9919;
  assign n9941 = n9651 & n9938;
  assign n9928 = n9927 ^ n9912;
  assign n9925 = ~n9902 & n9911;
  assign n9926 = n9886 & n9925;
  assign n9929 = n9928 ^ n9926;
  assign n9914 = n9913 ^ n9912;
  assign n9903 = n9895 & n9902;
  assign n9904 = ~n9886 & n9903;
  assign n9915 = n9914 ^ n9904;
  assign n9934 = n9929 ^ n9915;
  assign n9939 = n9938 ^ n9934;
  assign n9940 = n9887 & n9939;
  assign n9942 = n9941 ^ n9940;
  assign n9931 = n9906 & n9915;
  assign n10065 = n9942 ^ n9931;
  assign n9956 = n9871 & n9938;
  assign n9955 = n9888 & n9939;
  assign n9957 = n9956 ^ n9955;
  assign n9920 = n9919 ^ n9915;
  assign n9923 = n9757 & n9920;
  assign n9921 = n9897 & n9920;
  assign n9916 = n9778 & n9915;
  assign n9922 = n9921 ^ n9916;
  assign n9924 = n9923 ^ n9922;
  assign n10064 = n9957 ^ n9924;
  assign n10066 = n10065 ^ n10064;
  assign n10254 = n10253 ^ n10066;
  assign n7892 = n7891 ^ n7885;
  assign n7898 = n7897 ^ n7892;
  assign n7905 = n7904 ^ n7898;
  assign n7915 = n7914 ^ n7905;
  assign n7810 = n7809 ^ n7800;
  assign n7793 = n7792 ^ n7786;
  assign n7781 = n7780 ^ n7413;
  assign n7794 = n7793 ^ n7781;
  assign n7811 = n7810 ^ n7794;
  assign n8035 = n7915 ^ n7811;
  assign n8009 = n8008 ^ n8002;
  assign n8013 = n8012 ^ n8009;
  assign n8020 = n8019 ^ n8013;
  assign n7849 = n7848 ^ n7836;
  assign n7853 = n7852 ^ n7849;
  assign n7869 = n7868 ^ n7853;
  assign n8021 = n8020 ^ n7869;
  assign n7997 = n7996 ^ n7990;
  assign n7986 = n7985 ^ n7545;
  assign n7987 = n7986 ^ n7934;
  assign n7998 = n7997 ^ n7987;
  assign n8022 = n8021 ^ n7998;
  assign n7421 = n7420 ^ n7407;
  assign n7555 = n7554 ^ n7421;
  assign n7688 = n7687 ^ n7555;
  assign n7777 = n7776 ^ n7688;
  assign n8024 = n8022 ^ n7777;
  assign n7812 = n7811 ^ n7777;
  assign n8025 = n8024 ^ n7812;
  assign n7979 = n7978 ^ n7974;
  assign n7966 = n7965 ^ n7419;
  assign n7980 = n7979 ^ n7966;
  assign n7962 = n7961 ^ n7953;
  assign n7947 = n7946 ^ n7940;
  assign n7935 = n7934 ^ n7875;
  assign n7948 = n7947 ^ n7935;
  assign n7963 = n7962 ^ n7948;
  assign n7930 = n7929 ^ n7921;
  assign n7964 = n7963 ^ n7930;
  assign n7981 = n7980 ^ n7964;
  assign n7916 = n7915 ^ n7869;
  assign n7982 = n7981 ^ n7916;
  assign n8023 = n8022 ^ n7982;
  assign n8039 = n8025 ^ n8023;
  assign n8033 = n7981 ^ n7812;
  assign n8034 = n8033 ^ n8021;
  assign n8036 = ~n8034 & n8035;
  assign n8030 = n8020 ^ n7915;
  assign n8031 = n8030 ^ n7981;
  assign n8032 = n7812 & n8031;
  assign n8037 = n8036 ^ n8032;
  assign n8027 = n7963 ^ n7811;
  assign n8028 = n7982 & ~n8027;
  assign n8026 = ~n8023 & ~n8025;
  assign n8029 = n8028 ^ n8026;
  assign n8038 = n8037 ^ n8029;
  assign n8040 = n8039 ^ n8038;
  assign n8058 = n8033 ^ n8030;
  assign n8042 = n7915 ^ n7777;
  assign n8043 = n7916 ^ n7812;
  assign n8044 = n8042 & ~n8043;
  assign n8045 = n8044 ^ n8032;
  assign n8059 = n8058 ^ n8045;
  assign n8055 = n8042 ^ n8027;
  assign n8056 = ~n8033 & ~n8055;
  assign n8051 = n8033 ^ n7998;
  assign n8052 = n8022 ^ n7963;
  assign n8053 = n8052 ^ n8035;
  assign n8054 = n8051 & n8053;
  assign n8057 = n8056 ^ n8054;
  assign n8060 = n8059 ^ n8057;
  assign n8064 = n8035 ^ n8034;
  assign n8062 = ~n7998 & ~n8024;
  assign n8063 = n8062 ^ n8056;
  assign n8065 = n8064 ^ n8063;
  assign n8066 = n8065 ^ n8037;
  assign n8081 = n8060 & n8066;
  assign n8082 = n8040 & n8081;
  assign n8070 = n8066 ^ n8060;
  assign n8047 = n7963 & ~n8022;
  assign n8048 = n8047 ^ n8028;
  assign n8041 = n8027 ^ n7982;
  assign n8046 = n8045 ^ n8041;
  assign n8049 = n8048 ^ n8046;
  assign n8061 = ~n8049 & n8060;
  assign n8080 = n8070 ^ n8061;
  assign n8083 = n8082 ^ n8080;
  assign n8050 = n8049 ^ n8040;
  assign n8078 = n8061 ^ n8050;
  assign n8076 = ~n8049 & ~n8066;
  assign n8077 = ~n8040 & n8076;
  assign n8079 = n8078 ^ n8077;
  assign n8084 = n8083 ^ n8079;
  assign n10247 = n8035 & n8084;
  assign n10164 = ~n8034 & n8084;
  assign n8071 = n8061 ^ n8040;
  assign n8072 = ~n8070 & n8071;
  assign n8073 = n8072 ^ n8066;
  assign n8101 = n8083 ^ n8073;
  assign n10111 = ~n8027 & n8101;
  assign n10165 = n10164 ^ n10111;
  assign n10248 = n10247 ^ n10165;
  assign n8067 = n8066 ^ n8061;
  assign n8068 = ~n8050 & ~n8067;
  assign n8069 = n8068 ^ n8040;
  assign n8074 = n8073 ^ n8069;
  assign n8106 = n8031 & ~n8074;
  assign n8075 = n7812 & ~n8074;
  assign n10245 = n8106 ^ n8075;
  assign n10170 = ~n8025 & ~n8073;
  assign n8096 = n8079 ^ n8069;
  assign n10058 = ~n8033 & ~n8096;
  assign n8093 = ~n7998 & n8069;
  assign n10115 = n10058 ^ n8093;
  assign n10171 = n10170 ^ n10115;
  assign n10246 = n10245 ^ n10171;
  assign n10249 = n10248 ^ n10246;
  assign n10226 = n9812 & n9934;
  assign n9943 = n9937 ^ n9929;
  assign n10121 = n9881 & n9943;
  assign n10120 = n9868 & n9934;
  assign n10122 = n10121 ^ n10120;
  assign n10227 = n10226 ^ n10122;
  assign n10224 = n9956 ^ n9941;
  assign n10179 = n9876 & n9937;
  assign n9950 = n9777 & n9919;
  assign n10130 = n9950 ^ n9923;
  assign n10180 = n10179 ^ n10130;
  assign n10225 = n10224 ^ n10180;
  assign n10228 = n10227 ^ n10225;
  assign n10250 = n10249 ^ n10228;
  assign n10255 = n10254 ^ n10250;
  assign n7021 = n7020 ^ n7012;
  assign n7006 = n7005 ^ n6995;
  assign n7022 = n7021 ^ n7006;
  assign n6980 = n6979 ^ n6975;
  assign n6969 = n6968 ^ n6963;
  assign n6973 = n6972 ^ n6969;
  assign n6981 = n6980 ^ n6973;
  assign n7091 = n7022 ^ n6981;
  assign n6820 = n6819 ^ n6725;
  assign n5842 = n5841 ^ n4914;
  assign n6821 = n6820 ^ n5842;
  assign n7079 = n7022 ^ n6821;
  assign n7069 = n7068 ^ n7062;
  assign n7058 = n7057 ^ n7056;
  assign n7070 = n7069 ^ n7058;
  assign n7043 = n7042 ^ n7037;
  assign n7029 = n7028 ^ n7027;
  assign n7034 = n7033 ^ n7029;
  assign n7044 = n7043 ^ n7034;
  assign n7050 = n7049 ^ n7044;
  assign n7071 = n7070 ^ n7050;
  assign n7080 = n7079 ^ n7071;
  assign n6930 = n6929 ^ n6919;
  assign n6911 = n6910 ^ n6901;
  assign n6931 = n6930 ^ n6911;
  assign n6884 = n6883 ^ n6868;
  assign n6855 = n6854 ^ n6840;
  assign n6885 = n6884 ^ n6855;
  assign n6886 = n6885 ^ n6821;
  assign n6932 = n6931 ^ n6886;
  assign n7085 = n7080 ^ n6932;
  assign n7083 = n6981 ^ n6932;
  assign n6956 = n6955 ^ n6948;
  assign n6943 = n6942 ^ n6938;
  assign n6957 = n6956 ^ n6943;
  assign n6982 = n6981 ^ n6957;
  assign n7084 = n7083 ^ n6982;
  assign n7089 = n7085 ^ n7084;
  assign n7086 = n7084 & ~n7085;
  assign n7081 = n7044 ^ n6957;
  assign n7082 = ~n7080 & ~n7081;
  assign n7087 = n7086 ^ n7082;
  assign n7074 = n7022 ^ n6957;
  assign n7075 = n7071 ^ n6982;
  assign n7076 = n7075 ^ n6886;
  assign n7077 = ~n7074 & ~n7076;
  assign n7023 = n7022 ^ n6885;
  assign n7072 = n7071 ^ n7023;
  assign n7073 = n6982 & ~n7072;
  assign n7078 = n7077 ^ n7073;
  assign n7088 = n7087 ^ n7078;
  assign n7090 = n7089 ^ n7088;
  assign n7096 = n7076 ^ n7074;
  assign n7094 = n6931 & n7083;
  assign n7092 = n7091 ^ n7081;
  assign n7093 = ~n7075 & n7092;
  assign n7095 = n7094 ^ n7093;
  assign n7097 = n7096 ^ n7095;
  assign n7098 = n7097 ^ n7078;
  assign n7115 = n6932 & n7044;
  assign n7116 = n7115 ^ n7082;
  assign n7113 = n7081 ^ n7080;
  assign n7105 = n7079 ^ n6982;
  assign n7106 = ~n7091 & n7105;
  assign n7107 = n7106 ^ n7073;
  assign n7114 = n7113 ^ n7107;
  assign n7117 = n7116 ^ n7114;
  assign n7124 = n7098 & n7117;
  assign n7125 = n7090 & n7124;
  assign n7122 = n7117 ^ n7090;
  assign n7104 = n7075 ^ n7023;
  assign n7108 = n7107 ^ n7104;
  assign n7099 = n7044 ^ n6932;
  assign n7100 = n7099 ^ n7074;
  assign n7101 = n7075 ^ n6931;
  assign n7102 = n7100 & ~n7101;
  assign n7103 = n7102 ^ n7093;
  assign n7109 = n7108 ^ n7103;
  assign n7118 = ~n7109 & n7117;
  assign n7123 = n7122 ^ n7118;
  assign n7126 = n7125 ^ n7123;
  assign n7112 = n7109 ^ n7098;
  assign n7119 = n7118 ^ n7112;
  assign n7110 = ~n7098 & ~n7109;
  assign n7111 = ~n7090 & n7110;
  assign n7120 = n7119 ^ n7111;
  assign n7144 = n7126 ^ n7120;
  assign n7139 = n7118 ^ n7090;
  assign n7140 = ~n7112 & ~n7139;
  assign n7141 = n7140 ^ n7098;
  assign n7129 = n7118 ^ n7098;
  assign n7130 = ~n7122 & n7129;
  assign n7131 = n7130 ^ n7090;
  assign n7142 = n7141 ^ n7131;
  assign n7145 = n7144 ^ n7142;
  assign n7146 = ~n7091 & ~n7145;
  assign n7143 = n6982 & ~n7142;
  assign n7147 = n7146 ^ n7143;
  assign n7127 = n7100 & ~n7126;
  assign n10243 = n7147 ^ n7127;
  assign n10054 = n7105 & ~n7145;
  assign n10053 = ~n7072 & ~n7142;
  assign n10055 = n10054 ^ n10053;
  assign n7132 = n7131 ^ n7126;
  assign n7136 = ~n7075 & n7132;
  assign n7134 = ~n7101 & ~n7126;
  assign n7133 = n7092 & n7132;
  assign n7135 = n7134 ^ n7133;
  assign n7137 = n7136 ^ n7135;
  assign n10242 = n10055 ^ n7137;
  assign n10244 = n10243 ^ n10242;
  assign n10256 = n10255 ^ n10244;
  assign n10262 = n10261 ^ n10256;
  assign n10221 = n8890 & n9026;
  assign n9035 = n9029 ^ n9007;
  assign n10137 = n8972 & n9035;
  assign n10136 = n8960 & n9026;
  assign n10138 = n10137 ^ n10136;
  assign n10222 = n10221 ^ n10138;
  assign n10219 = n10070 ^ n9033;
  assign n10217 = n8967 & n9029;
  assign n10088 = n8824 & n9018;
  assign n10195 = n10088 ^ n9023;
  assign n10218 = n10217 ^ n10195;
  assign n10220 = n10219 ^ n10218;
  assign n10223 = n10222 ^ n10220;
  assign n10229 = n10228 ^ n10223;
  assign n10214 = n10053 ^ n7143;
  assign n10212 = n7084 & n7141;
  assign n10160 = n6931 & ~n7131;
  assign n10189 = n10160 ^ n7136;
  assign n10213 = n10212 ^ n10189;
  assign n10215 = n10214 ^ n10213;
  assign n10210 = ~n7074 & n7144;
  assign n7148 = n7141 ^ n7120;
  assign n10102 = ~n7081 & ~n7148;
  assign n10101 = ~n7076 & n7144;
  assign n10103 = n10102 ^ n10101;
  assign n10211 = n10210 ^ n10103;
  assign n10216 = n10215 ^ n10211;
  assign n10230 = n10229 ^ n10216;
  assign n8097 = ~n8055 & ~n8096;
  assign n8095 = n8051 & ~n8079;
  assign n8098 = n8097 ^ n8095;
  assign n10059 = n10058 ^ n8098;
  assign n8089 = n8053 & ~n8079;
  assign n8088 = ~n8022 & ~n8083;
  assign n8090 = n8089 ^ n8088;
  assign n10207 = n10059 ^ n8090;
  assign n8102 = n7982 & n8101;
  assign n8085 = n8084 ^ n8074;
  assign n8086 = n8042 & ~n8085;
  assign n8087 = n8086 ^ n8075;
  assign n8103 = n8102 ^ n8087;
  assign n10208 = n10207 ^ n8103;
  assign n9944 = n9878 & n9943;
  assign n9945 = n9944 ^ n9942;
  assign n9930 = n9874 & n9929;
  assign n9932 = n9931 ^ n9930;
  assign n9933 = n9932 ^ n9924;
  assign n9946 = n9945 ^ n9933;
  assign n10209 = n10208 ^ n9946;
  assign n10231 = n10230 ^ n10209;
  assign n10241 = n10240 ^ n10231;
  assign n10263 = n10262 ^ n10241;
  assign n10140 = n8981 & n9007;
  assign n10087 = n8970 & n9029;
  assign n10141 = n10140 ^ n10087;
  assign n10196 = n10195 ^ n10141;
  assign n9036 = n8969 & n9035;
  assign n9037 = n9036 ^ n9034;
  assign n10194 = n10137 ^ n9037;
  assign n10197 = n10196 ^ n10194;
  assign n10204 = n10203 ^ n10197;
  assign n10106 = ~n7085 & n7141;
  assign n10105 = ~n7099 & ~n7120;
  assign n10107 = n10106 ^ n10105;
  assign n10190 = n10189 ^ n10107;
  assign n7149 = ~n7080 & ~n7148;
  assign n7150 = n7149 ^ n7147;
  assign n10188 = n10102 ^ n7150;
  assign n10191 = n10190 ^ n10188;
  assign n8105 = ~n8043 & ~n8085;
  assign n8107 = n8106 ^ n8105;
  assign n8108 = n8107 ^ n8090;
  assign n8104 = n8103 ^ n8097;
  assign n8109 = n8108 ^ n8104;
  assign n10192 = n10191 ^ n8109;
  assign n10124 = n9905 & n9929;
  assign n9949 = n9879 & n9937;
  assign n10125 = n10124 ^ n9949;
  assign n10131 = n10130 ^ n10125;
  assign n10129 = n10121 ^ n9945;
  assign n10132 = n10131 ^ n10129;
  assign n9958 = n9957 ^ n9932;
  assign n9954 = n9945 ^ n9921;
  assign n9959 = n9958 ^ n9954;
  assign n10133 = n10132 ^ n9959;
  assign n10193 = n10192 ^ n10133;
  assign n10205 = n10204 ^ n10193;
  assign n10264 = n10263 ^ n10205;
  assign n9008 = n8825 & n9007;
  assign n10143 = n9034 ^ n9008;
  assign n10139 = n10138 ^ n10071;
  assign n10142 = n10141 ^ n10139;
  assign n10144 = n10143 ^ n10142;
  assign n10156 = n10155 ^ n10144;
  assign n10127 = n9942 ^ n9930;
  assign n10123 = n10122 ^ n9955;
  assign n10126 = n10125 ^ n10123;
  assign n10128 = n10127 ^ n10126;
  assign n10134 = n10133 ^ n10128;
  assign n10113 = n8052 & ~n8083;
  assign n8092 = ~n8023 & ~n8073;
  assign n10114 = n10113 ^ n8092;
  assign n10116 = n10115 ^ n10114;
  assign n10112 = n10111 ^ n8103;
  assign n10117 = n10116 ^ n10112;
  assign n10118 = n10117 ^ n8109;
  assign n7121 = n6932 & ~n7120;
  assign n10109 = n7147 ^ n7121;
  assign n10104 = n10103 ^ n10054;
  assign n10108 = n10107 ^ n10104;
  assign n10110 = n10109 ^ n10108;
  assign n10119 = n10118 ^ n10110;
  assign n10135 = n10134 ^ n10119;
  assign n10157 = n10156 ^ n10135;
  assign n10328 = n10264 ^ n10157;
  assign n10277 = n8966 & n9018;
  assign n9015 = n9014 ^ n9008;
  assign n10278 = n10277 ^ n9015;
  assign n10279 = n10278 ^ n10218;
  assign n10276 = n10139 ^ n9037;
  assign n10280 = n10279 ^ n10276;
  assign n10166 = n10165 ^ n8105;
  assign n10273 = n10166 ^ n10114;
  assign n10272 = n8088 ^ n8087;
  assign n10274 = n10273 ^ n10272;
  assign n10275 = n10274 ^ n10128;
  assign n10281 = n10280 ^ n10275;
  assign n10177 = n9875 & n9919;
  assign n10178 = n10177 ^ n9932;
  assign n10181 = n10180 ^ n10178;
  assign n10176 = n10123 ^ n9945;
  assign n10182 = n10181 ^ n10176;
  assign n10282 = n10281 ^ n10182;
  assign n10268 = n7083 & ~n7131;
  assign n7128 = n7127 ^ n7121;
  assign n10269 = n10268 ^ n7128;
  assign n10270 = n10269 ^ n10213;
  assign n10267 = n10104 ^ n7150;
  assign n10271 = n10270 ^ n10267;
  assign n10283 = n10282 ^ n10271;
  assign n10291 = n10290 ^ n10283;
  assign n10073 = n10072 ^ n9015;
  assign n10069 = n9037 ^ n9020;
  assign n10074 = n10073 ^ n10069;
  assign n10083 = n10082 ^ n10074;
  assign n10067 = n10066 ^ n9959;
  assign n10061 = n8089 ^ n8087;
  assign n10060 = n10059 ^ n8107;
  assign n10062 = n10061 ^ n10060;
  assign n10056 = n10055 ^ n7128;
  assign n10052 = n7150 ^ n7133;
  assign n10057 = n10056 ^ n10052;
  assign n10063 = n10062 ^ n10057;
  assign n10068 = n10067 ^ n10063;
  assign n10084 = n10083 ^ n10068;
  assign n10299 = n10291 ^ n10084;
  assign n10329 = n10328 ^ n10299;
  assign n10315 = n10157 & ~n10264;
  assign n10292 = n10291 ^ n10241;
  assign n10183 = n10182 ^ n9959;
  assign n9951 = n9950 ^ n9949;
  assign n9952 = n9951 ^ n9922;
  assign n9948 = n9942 ^ n9932;
  assign n9953 = n9952 ^ n9948;
  assign n10184 = n10183 ^ n9953;
  assign n10168 = ~n8024 & n8069;
  assign n10169 = n10168 ^ n8090;
  assign n10172 = n10171 ^ n10169;
  assign n10167 = n10166 ^ n8103;
  assign n10173 = n10172 ^ n10167;
  assign n10174 = n10173 ^ n8109;
  assign n10161 = n10160 ^ n10106;
  assign n10162 = n10161 ^ n7135;
  assign n10159 = n7147 ^ n7128;
  assign n10163 = n10162 ^ n10159;
  assign n10175 = n10174 ^ n10163;
  assign n10185 = n10184 ^ n10175;
  assign n10089 = n10088 ^ n10087;
  assign n10090 = n10089 ^ n9022;
  assign n10086 = n9034 ^ n9015;
  assign n10091 = n10090 ^ n10086;
  assign n10100 = n10099 ^ n10091;
  assign n10158 = n10157 ^ n10100;
  assign n10186 = n10185 ^ n10158;
  assign n10293 = n10292 ^ n10186;
  assign n10296 = n10157 ^ n10084;
  assign n10297 = n10293 & ~n10296;
  assign n10316 = n10315 ^ n10297;
  assign n10313 = n10296 ^ n10293;
  assign n9960 = n9959 ^ n9953;
  assign n9025 = n9024 ^ n9015;
  assign n9038 = n9037 ^ n9025;
  assign n9947 = n9946 ^ n9038;
  assign n9961 = n9960 ^ n9947;
  assign n8094 = n8093 ^ n8092;
  assign n8099 = n8098 ^ n8094;
  assign n8091 = n8090 ^ n8087;
  assign n8100 = n8099 ^ n8091;
  assign n8110 = n8109 ^ n8100;
  assign n9962 = n9961 ^ n8110;
  assign n7138 = n7137 ^ n7128;
  assign n7151 = n7150 ^ n7138;
  assign n9963 = n9962 ^ n7151;
  assign n10051 = n10050 ^ n9963;
  assign n10309 = n10291 ^ n10051;
  assign n10085 = n10084 ^ n10051;
  assign n10310 = n10292 ^ n10085;
  assign n10311 = n10309 & ~n10310;
  assign n10302 = n10291 ^ n10262;
  assign n10303 = n10302 ^ n10186;
  assign n10304 = n10085 & n10303;
  assign n10312 = n10311 ^ n10304;
  assign n10314 = n10313 ^ n10312;
  assign n10317 = n10316 ^ n10314;
  assign n10187 = n10186 ^ n10085;
  assign n10332 = n10302 ^ n10187;
  assign n10333 = n10332 ^ n10312;
  assign n10206 = n10205 ^ n10187;
  assign n10330 = n10206 & n10329;
  assign n10319 = n10309 ^ n10296;
  assign n10320 = ~n10187 & ~n10319;
  assign n10331 = n10330 ^ n10320;
  assign n10334 = n10333 ^ n10331;
  assign n10335 = ~n10317 & n10334;
  assign n10294 = n10293 ^ n10264;
  assign n10265 = n10264 ^ n10051;
  assign n10266 = n10265 ^ n10085;
  assign n10307 = n10294 ^ n10266;
  assign n10300 = n10263 ^ n10187;
  assign n10301 = n10299 & ~n10300;
  assign n10305 = n10304 ^ n10301;
  assign n10295 = ~n10266 & ~n10294;
  assign n10298 = n10297 ^ n10295;
  assign n10306 = n10305 ^ n10298;
  assign n10308 = n10307 ^ n10306;
  assign n10327 = n10317 ^ n10308;
  assign n10336 = n10335 ^ n10327;
  assign n10322 = n10300 ^ n10299;
  assign n10318 = ~n10205 & ~n10265;
  assign n10321 = n10320 ^ n10318;
  assign n10323 = n10322 ^ n10321;
  assign n10324 = n10323 ^ n10305;
  assign n10325 = ~n10317 & ~n10324;
  assign n10326 = ~n10308 & n10325;
  assign n10337 = n10336 ^ n10326;
  assign n10365 = n10329 & ~n10337;
  assign n10353 = n10324 & n10334;
  assign n10354 = n10308 & n10353;
  assign n10347 = n10334 ^ n10324;
  assign n10352 = n10347 ^ n10335;
  assign n10355 = n10354 ^ n10352;
  assign n10356 = n10355 ^ n10337;
  assign n10348 = n10335 ^ n10308;
  assign n10349 = ~n10347 & n10348;
  assign n10350 = n10349 ^ n10324;
  assign n10339 = n10335 ^ n10324;
  assign n10340 = ~n10327 & ~n10339;
  assign n10341 = n10340 ^ n10308;
  assign n10351 = n10350 ^ n10341;
  assign n10357 = n10356 ^ n10351;
  assign n10363 = n10309 & ~n10357;
  assign n10362 = n10085 & ~n10351;
  assign n10364 = n10363 ^ n10362;
  assign n10366 = n10365 ^ n10364;
  assign n10359 = n10303 & ~n10351;
  assign n10358 = ~n10310 & ~n10357;
  assign n10360 = n10359 ^ n10358;
  assign n10342 = n10341 ^ n10337;
  assign n10345 = ~n10187 & ~n10342;
  assign n10343 = ~n10319 & ~n10342;
  assign n10338 = n10206 & ~n10337;
  assign n10344 = n10343 ^ n10338;
  assign n10346 = n10345 ^ n10344;
  assign n10361 = n10360 ^ n10346;
  assign n10367 = n10366 ^ n10361;
  assign n13461 = n13460 ^ n10367;
  assign n17275 = n17274 ^ n13461;
  assign n17277 = n17276 ^ n17275;
  assign n13312 = n13133 & n13146;
  assign n13148 = n12991 & n13147;
  assign n13313 = n13312 ^ n13148;
  assign n13315 = n13314 ^ n13313;
  assign n13171 = n13104 & n13156;
  assign n13170 = n13132 & n13146;
  assign n13172 = n13171 ^ n13170;
  assign n13316 = n13315 ^ n13172;
  assign n13161 = n13160 ^ n13159;
  assign n13162 = n12921 & n13161;
  assign n13164 = n13163 ^ n13162;
  assign n13158 = n13108 & n13157;
  assign n13165 = n13164 ^ n13158;
  assign n13317 = n13316 ^ n13165;
  assign n17272 = n15333 ^ n13317;
  assign n13290 = n11214 & ~n11295;
  assign n13291 = n13290 ^ n11315;
  assign n13472 = n13291 ^ n11310;
  assign n13287 = ~n11269 & ~n13286;
  assign n13288 = n13287 ^ n11314;
  assign n13473 = n13472 ^ n13288;
  assign n17270 = n13473 ^ n13456;
  assign n13479 = n12179 & n12233;
  assign n13349 = ~n12178 & n12233;
  assign n12221 = n12220 ^ n12216;
  assign n13348 = ~n12174 & n12221;
  assign n13350 = n13349 ^ n13348;
  assign n13480 = n13479 ^ n13350;
  assign n13476 = ~n12207 & ~n12216;
  assign n13386 = ~n12095 & n12226;
  assign n13430 = n13386 ^ n13306;
  assign n13477 = n13476 ^ n13430;
  assign n13475 = n12245 ^ n12228;
  assign n13478 = n13477 ^ n13475;
  assign n13481 = n13480 ^ n13478;
  assign n13449 = n10299 & n10356;
  assign n13356 = ~n10300 & n10356;
  assign n12249 = n10355 ^ n10350;
  assign n13328 = ~n10296 & n12249;
  assign n13357 = n13356 ^ n13328;
  assign n13450 = n13449 ^ n13357;
  assign n13447 = n10362 ^ n10359;
  assign n13394 = ~n10266 & ~n10350;
  assign n13281 = ~n10205 & n10341;
  assign n13332 = n13281 ^ n10345;
  assign n13395 = n13394 ^ n13332;
  assign n13448 = n13447 ^ n13395;
  assign n13451 = n13450 ^ n13448;
  assign n13482 = n13481 ^ n13451;
  assign n17271 = n17270 ^ n13482;
  assign n17273 = n17272 ^ n17271;
  assign n17278 = n17277 ^ n17273;
  assign n13167 = n13116 & n13161;
  assign n13169 = n13168 ^ n13167;
  assign n13173 = n13172 ^ n13169;
  assign n13166 = n13165 ^ n13148;
  assign n13174 = n13173 ^ n13166;
  assign n17262 = n15317 ^ n13174;
  assign n13346 = n12188 & ~n12220;
  assign n13345 = ~n12208 & ~n12216;
  assign n13347 = n13346 ^ n13345;
  assign n13431 = n13430 ^ n13347;
  assign n12222 = n12079 & n12221;
  assign n12237 = n12236 ^ n12222;
  assign n13429 = n13348 ^ n12237;
  assign n13432 = n13431 ^ n13429;
  assign n13330 = n10328 & ~n10355;
  assign n13280 = ~n10294 & ~n10350;
  assign n13331 = n13330 ^ n13280;
  assign n13333 = n13332 ^ n13331;
  assign n12250 = n10293 & n12249;
  assign n12251 = n12250 ^ n10364;
  assign n13329 = n13328 ^ n12251;
  assign n13334 = n13333 ^ n13329;
  assign n13433 = n13432 ^ n13334;
  assign n13338 = n11215 & ~n11295;
  assign n13295 = ~n11278 & n11286;
  assign n13339 = n13338 ^ n13295;
  assign n13341 = n13340 ^ n13339;
  assign n13337 = n13336 ^ n13288;
  assign n13342 = n13341 ^ n13337;
  assign n13292 = n13291 ^ n11304;
  assign n13289 = n13288 ^ n11307;
  assign n13293 = n13292 ^ n13289;
  assign n13343 = n13342 ^ n13293;
  assign n17261 = n13433 ^ n13343;
  assign n17263 = n17262 ^ n17261;
  assign n17287 = n17278 ^ n17263;
  assign n13363 = n13109 & n13152;
  assign n13415 = n13414 ^ n13363;
  assign n13416 = n13415 ^ n13313;
  assign n13413 = n13172 ^ n13164;
  assign n13417 = n13416 ^ n13413;
  assign n17241 = n13417 ^ n13174;
  assign n17242 = n17241 ^ n15281;
  assign n13297 = n13296 ^ n13295;
  assign n13298 = n13297 ^ n11309;
  assign n13294 = n13291 ^ n11314;
  assign n13299 = n13298 ^ n13294;
  assign n13300 = n13299 ^ n13293;
  assign n17239 = n13473 ^ n13300;
  assign n12241 = ~n12148 & ~n12220;
  assign n12243 = n12242 ^ n12241;
  assign n13308 = n13307 ^ n12243;
  assign n13309 = n13308 ^ n12237;
  assign n12253 = ~n10264 & ~n10355;
  assign n12254 = n12253 ^ n10365;
  assign n13302 = n12254 ^ n10346;
  assign n13303 = n13302 ^ n12251;
  assign n13310 = n13309 ^ n13303;
  assign n17240 = n17239 ^ n13310;
  assign n17243 = n17242 ^ n17240;
  assign n17289 = n17287 ^ n17243;
  assign n13364 = n13131 & n13156;
  assign n13365 = n13364 ^ n13363;
  assign n13437 = n13436 ^ n13365;
  assign n13435 = n13366 ^ n13165;
  assign n13438 = n13437 ^ n13435;
  assign n17251 = n13438 ^ n13174;
  assign n17252 = n17251 ^ n14782;
  assign n13403 = n13402 ^ n11302;
  assign n13505 = n13403 ^ n13339;
  assign n13504 = n13290 ^ n11314;
  assign n13506 = n13505 ^ n13504;
  assign n17249 = n13506 ^ n13343;
  assign n13358 = n13357 ^ n10358;
  assign n13359 = n13358 ^ n13331;
  assign n13355 = n12253 ^ n10364;
  assign n13360 = n13359 ^ n13355;
  assign n13353 = n12241 ^ n12236;
  assign n13351 = n13350 ^ n12244;
  assign n13352 = n13351 ^ n13347;
  assign n13354 = n13353 ^ n13352;
  assign n13361 = n13360 ^ n13354;
  assign n17250 = n17249 ^ n13361;
  assign n17253 = n17252 ^ n17250;
  assign n17304 = ~n17253 & n17287;
  assign n13371 = n13171 ^ n13164;
  assign n13369 = n13368 ^ n13167;
  assign n13370 = n13369 ^ n13365;
  assign n13372 = n13371 ^ n13370;
  assign n17267 = n15408 ^ n13372;
  assign n13405 = n11259 & ~n11290;
  assign n13406 = n13405 ^ n13291;
  assign n13409 = n13408 ^ n13406;
  assign n13404 = n13403 ^ n13288;
  assign n13410 = n13409 ^ n13404;
  assign n17265 = n13506 ^ n13410;
  assign n13511 = n13351 ^ n12237;
  assign n13508 = ~n12149 & n12226;
  assign n13509 = n13508 ^ n12243;
  assign n13510 = n13509 ^ n13477;
  assign n13512 = n13511 ^ n13510;
  assign n13396 = ~n10265 & n10341;
  assign n13397 = n13396 ^ n12254;
  assign n13398 = n13397 ^ n13395;
  assign n13393 = n13358 ^ n12251;
  assign n13399 = n13398 ^ n13393;
  assign n13513 = n13512 ^ n13399;
  assign n17266 = n17265 ^ n13513;
  assign n17268 = n17267 ^ n17266;
  assign n17285 = n17273 ^ n17268;
  assign n13516 = n13105 & n13142;
  assign n13517 = n13516 ^ n13172;
  assign n13518 = n13517 ^ n13485;
  assign n13515 = n13369 ^ n13165;
  assign n13519 = n13518 ^ n13515;
  assign n17256 = n13519 ^ n13174;
  assign n17257 = n17256 ^ n15252;
  assign n13411 = n13410 ^ n13293;
  assign n17255 = n13411 ^ n13299;
  assign n17258 = n17257 ^ n17255;
  assign n13389 = n12243 ^ n12236;
  assign n13387 = n13386 ^ n13345;
  assign n13388 = n13387 ^ n13305;
  assign n13390 = n13389 ^ n13388;
  assign n13282 = n13281 ^ n13280;
  assign n13283 = n13282 ^ n10344;
  assign n13279 = n12254 ^ n10364;
  assign n13284 = n13283 ^ n13279;
  assign n13391 = n13390 ^ n13284;
  assign n17254 = n17253 ^ n13391;
  assign n17259 = n17258 ^ n17254;
  assign n17286 = n17285 ^ n17259;
  assign n13464 = n13170 ^ n13164;
  assign n13463 = n13315 ^ n13169;
  assign n13465 = n13464 ^ n13463;
  assign n17246 = n15211 ^ n13465;
  assign n17244 = n13293 ^ n11317;
  assign n12255 = n12254 ^ n10360;
  assign n12252 = n12251 ^ n10343;
  assign n12256 = n12255 ^ n12252;
  assign n12247 = n12246 ^ n12243;
  assign n12240 = n12239 ^ n12237;
  assign n12248 = n12247 ^ n12240;
  assign n12257 = n12256 ^ n12248;
  assign n17245 = n17244 ^ n12257;
  assign n17247 = n17246 ^ n17245;
  assign n17292 = n17253 ^ n17247;
  assign n17293 = n17286 & n17292;
  assign n17305 = n17304 ^ n17293;
  assign n17302 = n17292 ^ n17286;
  assign n17298 = n17268 ^ n17243;
  assign n17248 = n17247 ^ n17243;
  assign n17299 = n17285 ^ n17248;
  assign n17300 = n17298 & n17299;
  assign n17281 = n17277 ^ n17268;
  assign n17282 = n17281 ^ n17259;
  assign n17283 = n17248 & n17282;
  assign n17301 = n17300 ^ n17283;
  assign n17303 = n17302 ^ n17301;
  assign n17306 = n17305 ^ n17303;
  assign n17290 = n17289 ^ n17248;
  assign n17288 = n17287 ^ n17286;
  assign n17296 = n17290 ^ n17288;
  assign n17291 = n17288 & n17290;
  assign n17294 = n17293 ^ n17291;
  assign n17269 = n17268 ^ n17247;
  assign n17260 = n17259 ^ n17248;
  assign n17279 = n17278 ^ n17260;
  assign n17280 = n17269 & n17279;
  assign n17284 = n17283 ^ n17280;
  assign n17295 = n17294 ^ n17284;
  assign n17297 = n17296 ^ n17295;
  assign n17324 = n17306 ^ n17297;
  assign n17320 = n17281 ^ n17260;
  assign n17321 = n17320 ^ n17301;
  assign n17264 = n17263 ^ n17260;
  assign n17316 = n17287 ^ n17253;
  assign n17317 = n17316 ^ n17269;
  assign n17318 = n17264 & n17317;
  assign n17308 = n17298 ^ n17292;
  assign n17309 = n17260 & n17308;
  assign n17319 = n17318 ^ n17309;
  assign n17322 = n17321 ^ n17319;
  assign n17323 = n17306 & n17322;
  assign n17311 = n17279 ^ n17269;
  assign n17307 = n17263 & n17289;
  assign n17310 = n17309 ^ n17307;
  assign n17312 = n17311 ^ n17310;
  assign n17313 = n17312 ^ n17284;
  assign n17328 = n17323 ^ n17313;
  assign n17329 = n17324 & n17328;
  assign n17330 = n17329 ^ n17297;
  assign n17678 = n17289 & n17330;
  assign n17338 = n17322 ^ n17313;
  assign n17339 = n17338 ^ n17323;
  assign n17336 = ~n17313 & n17322;
  assign n17337 = n17297 & n17336;
  assign n17340 = n17339 ^ n17337;
  assign n17514 = n17287 & n17340;
  assign n17325 = n17324 ^ n17323;
  assign n17314 = n17306 & n17313;
  assign n17315 = ~n17297 & n17314;
  assign n17326 = n17325 ^ n17315;
  assign n17354 = n17317 & n17326;
  assign n17515 = n17514 ^ n17354;
  assign n17679 = n17678 ^ n17515;
  assign n17342 = n17323 ^ n17297;
  assign n17343 = n17338 & n17342;
  assign n17344 = n17343 ^ n17313;
  assign n17581 = n17290 & n17344;
  assign n17509 = n17263 & n17330;
  assign n17331 = n17330 ^ n17326;
  assign n17334 = n17260 & n17331;
  assign n17510 = n17509 ^ n17334;
  assign n17582 = n17581 ^ n17510;
  assign n17680 = n17679 ^ n17582;
  assign n17341 = n17340 ^ n17326;
  assign n17585 = n17279 & n17341;
  assign n17501 = n17344 ^ n17340;
  assign n17502 = n17292 & n17501;
  assign n17586 = n17585 ^ n17502;
  assign n17345 = n17344 ^ n17330;
  assign n17346 = n17345 ^ n17341;
  assign n17347 = n17299 & n17346;
  assign n17676 = n17586 ^ n17347;
  assign n17503 = n17286 & n17501;
  assign n17352 = n17248 & n17345;
  assign n17351 = n17298 & n17346;
  assign n17353 = n17352 ^ n17351;
  assign n17504 = n17503 ^ n17353;
  assign n17677 = n17676 ^ n17504;
  assign n17681 = n17680 ^ n17677;
  assign n17348 = n17282 & n17345;
  assign n17349 = n17348 ^ n17347;
  assign n17516 = n17515 ^ n17349;
  assign n17332 = n17308 & n17331;
  assign n17513 = n17504 ^ n17332;
  assign n17517 = n17516 ^ n17513;
  assign n17682 = n17681 ^ n17517;
  assign n17689 = n17688 ^ n17682;
  assign n13772 = n11154 ^ n10486;
  assign n13773 = n13772 ^ n11149;
  assign n13770 = n11207 ^ n11132;
  assign n13771 = n13770 ^ n12953;
  assign n13774 = n13773 ^ n13771;
  assign n13764 = n13074 ^ n11061;
  assign n13762 = n11182 ^ n11118;
  assign n13763 = n13762 ^ n11187;
  assign n13765 = n13764 ^ n13763;
  assign n13745 = n13051 ^ n11106;
  assign n13743 = n11182 ^ n11034;
  assign n13744 = n13743 ^ n11054;
  assign n13746 = n13745 ^ n13744;
  assign n13766 = n13765 ^ n13746;
  assign n13760 = n13098 ^ n11132;
  assign n13759 = n11203 ^ n11154;
  assign n13761 = n13760 ^ n13759;
  assign n13767 = n13766 ^ n13761;
  assign n13797 = n13774 ^ n13767;
  assign n13755 = n12984 ^ n11191;
  assign n13753 = n11118 ^ n11088;
  assign n13754 = n13753 ^ n11127;
  assign n13756 = n13755 ^ n13754;
  assign n13741 = n12915 ^ n11166;
  assign n13739 = n11227 ^ n10486;
  assign n13740 = n13739 ^ n10758;
  assign n13742 = n13741 ^ n13740;
  assign n13787 = n13756 ^ n13742;
  assign n13798 = n13797 ^ n13787;
  assign n13778 = n11228 ^ n11083;
  assign n13776 = n11132 ^ n10918;
  assign n13777 = n13776 ^ n13018;
  assign n13779 = n13778 ^ n13777;
  assign n13775 = n13774 ^ n11221;
  assign n13780 = n13779 ^ n13775;
  assign n13747 = n13746 ^ n13742;
  assign n13808 = n13780 ^ n13747;
  assign n13817 = n13808 ^ n13767;
  assign n13750 = n11089 ^ n11034;
  assign n13751 = n13750 ^ n11078;
  assign n13748 = n11234 ^ n11132;
  assign n13749 = n13748 ^ n12838;
  assign n13752 = n13751 ^ n13749;
  assign n13768 = n13767 ^ n13752;
  assign n13757 = n13756 ^ n13752;
  assign n13816 = n13768 ^ n13757;
  assign n13821 = n13817 ^ n13816;
  assign n13818 = ~n13816 & ~n13817;
  assign n13783 = n13774 ^ n13756;
  assign n13812 = ~n13783 & n13808;
  assign n13819 = n13818 ^ n13812;
  assign n13792 = n13765 ^ n13742;
  assign n13793 = n13792 ^ n13780;
  assign n13794 = n13757 & n13793;
  assign n13781 = n13780 ^ n13757;
  assign n13788 = n13781 ^ n13766;
  assign n13791 = n13787 & ~n13788;
  assign n13795 = n13794 ^ n13791;
  assign n13820 = n13819 ^ n13795;
  assign n13822 = n13821 ^ n13820;
  assign n13811 = ~n13767 & n13774;
  assign n13813 = n13812 ^ n13811;
  assign n13809 = n13808 ^ n13783;
  assign n13758 = n13757 ^ n13747;
  assign n13782 = n13752 ^ n13742;
  assign n13803 = ~n13758 & n13782;
  assign n13804 = n13803 ^ n13794;
  assign n13810 = n13809 ^ n13804;
  assign n13814 = n13813 ^ n13810;
  assign n13826 = n13822 ^ n13814;
  assign n13802 = n13792 ^ n13781;
  assign n13805 = n13804 ^ n13802;
  assign n13799 = n13781 ^ n13761;
  assign n13800 = n13798 & n13799;
  assign n13784 = n13783 ^ n13782;
  assign n13785 = ~n13781 & ~n13784;
  assign n13801 = n13800 ^ n13785;
  assign n13806 = n13805 ^ n13801;
  assign n13815 = n13806 & ~n13814;
  assign n13837 = n13826 ^ n13815;
  assign n13789 = n13788 ^ n13787;
  assign n13769 = ~n13761 & ~n13768;
  assign n13786 = n13785 ^ n13769;
  assign n13790 = n13789 ^ n13786;
  assign n13796 = n13795 ^ n13790;
  assign n13835 = ~n13796 & ~n13814;
  assign n13836 = ~n13822 & n13835;
  assign n13838 = n13837 ^ n13836;
  assign n13854 = n13798 & ~n13838;
  assign n13832 = n13796 & n13806;
  assign n13833 = n13822 & n13832;
  assign n13807 = n13806 ^ n13796;
  assign n13831 = n13815 ^ n13807;
  assign n13834 = n13833 ^ n13831;
  assign n13839 = n13838 ^ n13834;
  assign n13827 = n13815 ^ n13796;
  assign n13828 = ~n13826 & ~n13827;
  assign n13829 = n13828 ^ n13822;
  assign n13823 = n13822 ^ n13815;
  assign n13824 = ~n13807 & n13823;
  assign n13825 = n13824 ^ n13796;
  assign n13830 = n13829 ^ n13825;
  assign n13840 = n13839 ^ n13830;
  assign n13852 = n13782 & ~n13840;
  assign n13851 = n13757 & ~n13830;
  assign n13853 = n13852 ^ n13851;
  assign n13855 = n13854 ^ n13853;
  assign n13844 = n13838 ^ n13829;
  assign n13848 = ~n13781 & ~n13844;
  assign n13846 = n13799 & ~n13838;
  assign n13845 = ~n13784 & ~n13844;
  assign n13847 = n13846 ^ n13845;
  assign n13849 = n13848 ^ n13847;
  assign n13842 = n13793 & ~n13830;
  assign n13841 = ~n13758 & ~n13840;
  assign n13843 = n13842 ^ n13841;
  assign n13850 = n13849 ^ n13843;
  assign n13856 = n13855 ^ n13850;
  assign n17141 = n17140 ^ n13856;
  assign n14041 = n14040 ^ n10280;
  assign n14038 = n10274 ^ n10110;
  assign n14037 = n10182 ^ n10173;
  assign n14039 = n14038 ^ n14037;
  assign n14042 = n14041 ^ n14039;
  assign n14006 = n14005 ^ n10074;
  assign n14003 = n10244 ^ n10062;
  assign n14002 = n9959 ^ n8109;
  assign n14004 = n14003 ^ n14002;
  assign n14007 = n14006 ^ n14004;
  assign n14043 = n14042 ^ n14007;
  assign n14033 = n14032 ^ n10223;
  assign n14030 = n10208 ^ n7151;
  assign n14031 = n14030 ^ n10250;
  assign n14034 = n14033 ^ n14031;
  assign n14058 = n14042 ^ n14034;
  assign n14020 = n14019 ^ n10091;
  assign n14017 = n10271 ^ n10057;
  assign n14018 = n14017 ^ n10174;
  assign n14021 = n14020 ^ n14018;
  assign n14014 = n14013 ^ n10144;
  assign n14010 = n10191 ^ n10057;
  assign n14011 = n14010 ^ n10118;
  assign n14012 = n14011 ^ n10275;
  assign n14015 = n14014 ^ n14012;
  assign n14009 = n9953 ^ n8100;
  assign n14016 = n14015 ^ n14009;
  assign n14022 = n14021 ^ n14016;
  assign n14059 = n14058 ^ n14022;
  assign n14053 = n14052 ^ n10197;
  assign n14050 = n10057 ^ n8109;
  assign n14049 = n10132 ^ n10117;
  assign n14051 = n14050 ^ n14049;
  assign n14054 = n14053 ^ n14051;
  assign n14028 = n14027 ^ n10253;
  assign n14025 = n10249 ^ n10216;
  assign n14024 = n10066 ^ n10062;
  assign n14026 = n14025 ^ n14024;
  assign n14029 = n14028 ^ n14026;
  assign n14035 = n14034 ^ n14029;
  assign n14055 = n14054 ^ n14035;
  assign n14060 = n14059 ^ n14055;
  assign n14000 = n13999 ^ n9038;
  assign n13996 = n10163 ^ n10057;
  assign n13997 = n13996 ^ n8110;
  assign n13998 = n13997 ^ n10209;
  assign n14001 = n14000 ^ n13998;
  assign n14056 = n14055 ^ n14001;
  assign n14008 = n14007 ^ n14001;
  assign n14057 = n14056 ^ n14008;
  assign n14066 = n14060 ^ n14057;
  assign n14062 = n14015 ^ n14007;
  assign n14063 = n14059 & n14062;
  assign n14061 = ~n14057 & ~n14060;
  assign n14064 = n14063 ^ n14061;
  assign n14045 = n14042 ^ n14029;
  assign n14046 = n14045 ^ n14022;
  assign n14047 = n14008 & n14046;
  assign n14023 = n14022 ^ n14008;
  assign n14036 = n14035 ^ n14023;
  assign n14044 = ~n14036 & n14043;
  assign n14048 = n14047 ^ n14044;
  assign n14065 = n14064 ^ n14048;
  assign n14067 = n14066 ^ n14065;
  assign n14081 = n14043 ^ n14036;
  assign n14068 = n14042 ^ n14001;
  assign n14078 = n14068 ^ n14062;
  assign n14079 = ~n14023 & n14078;
  assign n14077 = ~n14054 & ~n14056;
  assign n14080 = n14079 ^ n14077;
  assign n14082 = n14081 ^ n14080;
  assign n14083 = n14082 ^ n14048;
  assign n14091 = n14045 ^ n14023;
  assign n14069 = n14058 ^ n14008;
  assign n14070 = n14068 & ~n14069;
  assign n14071 = n14070 ^ n14047;
  assign n14092 = n14091 ^ n14071;
  assign n14086 = n14055 ^ n14015;
  assign n14087 = n14086 ^ n14043;
  assign n14088 = n14054 ^ n14023;
  assign n14089 = ~n14087 & n14088;
  assign n14090 = n14089 ^ n14079;
  assign n14093 = n14092 ^ n14090;
  assign n14114 = n14083 & n14093;
  assign n14115 = n14067 & n14114;
  assign n14107 = n14093 ^ n14083;
  assign n14074 = ~n14015 & ~n14055;
  assign n14075 = n14074 ^ n14063;
  assign n14072 = n14062 ^ n14059;
  assign n14073 = n14072 ^ n14071;
  assign n14076 = n14075 ^ n14073;
  assign n14094 = n14076 & n14093;
  assign n14113 = n14107 ^ n14094;
  assign n14116 = n14115 ^ n14113;
  assign n14095 = n14076 ^ n14067;
  assign n14096 = n14095 ^ n14094;
  assign n14084 = n14076 & ~n14083;
  assign n14085 = ~n14067 & n14084;
  assign n14097 = n14096 ^ n14085;
  assign n14117 = n14116 ^ n14097;
  assign n14240 = n14043 & ~n14117;
  assign n14238 = ~n14036 & ~n14117;
  assign n14108 = n14094 ^ n14067;
  assign n14109 = ~n14107 & n14108;
  assign n14110 = n14109 ^ n14083;
  assign n14236 = n14116 ^ n14110;
  assign n14237 = n14062 & n14236;
  assign n14239 = n14238 ^ n14237;
  assign n14241 = n14240 ^ n14239;
  assign n14098 = n14094 ^ n14083;
  assign n14099 = n14095 & ~n14098;
  assign n14100 = n14099 ^ n14067;
  assign n14111 = n14110 ^ n14100;
  assign n14122 = n14008 & ~n14111;
  assign n14112 = n14046 & ~n14111;
  assign n14234 = n14122 ^ n14112;
  assign n14232 = ~n14057 & ~n14110;
  assign n14230 = ~n14054 & n14100;
  assign n14101 = n14100 ^ n14097;
  assign n14102 = ~n14023 & n14101;
  assign n14231 = n14230 ^ n14102;
  assign n14233 = n14232 ^ n14231;
  assign n14235 = n14234 ^ n14233;
  assign n14242 = n14241 ^ n14235;
  assign n13898 = n12012 ^ n11644;
  assign n13899 = n13898 ^ n11967;
  assign n13900 = n13899 ^ n11959;
  assign n13901 = n13900 ^ n12024;
  assign n13902 = n13901 ^ n13177;
  assign n13893 = n12167 ^ n11905;
  assign n13892 = n12160 ^ n12133;
  assign n13894 = n13893 ^ n13892;
  assign n13891 = n13186 ^ n11923;
  assign n13895 = n13894 ^ n13891;
  assign n13903 = n13902 ^ n13895;
  assign n13872 = n12144 ^ n12065;
  assign n13871 = n12101 ^ n12071;
  assign n13873 = n13872 ^ n13871;
  assign n13874 = n13873 ^ n13175;
  assign n13938 = n13902 ^ n13874;
  assign n13914 = n12106 ^ n11960;
  assign n13912 = n12163 ^ n12035;
  assign n13913 = n13912 ^ n11991;
  assign n13915 = n13914 ^ n13913;
  assign n13908 = n12012 ^ n11906;
  assign n13906 = n12163 ^ n12085;
  assign n13907 = n13906 ^ n11771;
  assign n13909 = n13908 ^ n13907;
  assign n13905 = n13180 ^ n11932;
  assign n13910 = n13909 ^ n13905;
  assign n13904 = n13182 ^ n11436;
  assign n13911 = n13910 ^ n13904;
  assign n13916 = n13915 ^ n13911;
  assign n13946 = n13938 ^ n13916;
  assign n13881 = n12163 ^ n12082;
  assign n13882 = n13881 ^ n11906;
  assign n13880 = n13197 ^ n11917;
  assign n13883 = n13882 ^ n13880;
  assign n13875 = n12143 ^ n12059;
  assign n13876 = n13875 ^ n12168;
  assign n13877 = n13876 ^ n12137;
  assign n13878 = n13877 ^ n13199;
  assign n13879 = n13878 ^ n13874;
  assign n13884 = n13883 ^ n13879;
  assign n13947 = n13946 ^ n13884;
  assign n13886 = n12107 ^ n12075;
  assign n13885 = n12163 ^ n11980;
  assign n13887 = n13886 ^ n13885;
  assign n13888 = n13887 ^ n12098;
  assign n13889 = n13888 ^ n13188;
  assign n13896 = n13895 ^ n13889;
  assign n13890 = n13889 ^ n13884;
  assign n13897 = n13896 ^ n13890;
  assign n13952 = n13947 ^ n13897;
  assign n13925 = n13910 ^ n13895;
  assign n13949 = ~n13925 & n13946;
  assign n13948 = ~n13897 & ~n13947;
  assign n13950 = n13949 ^ n13948;
  assign n13920 = n13902 ^ n13878;
  assign n13921 = n13920 ^ n13916;
  assign n13922 = n13896 & n13921;
  assign n13917 = n13916 ^ n13896;
  assign n13918 = n13917 ^ n13879;
  assign n13919 = n13903 & ~n13918;
  assign n13923 = n13922 ^ n13919;
  assign n13951 = n13950 ^ n13923;
  assign n13953 = n13952 ^ n13951;
  assign n13930 = n13918 ^ n13903;
  assign n13926 = n13902 ^ n13889;
  assign n13927 = n13926 ^ n13925;
  assign n13928 = ~n13917 & ~n13927;
  assign n13924 = ~n13883 & ~n13890;
  assign n13929 = n13928 ^ n13924;
  assign n13931 = n13930 ^ n13929;
  assign n13932 = n13931 ^ n13923;
  assign n13942 = n13920 ^ n13917;
  assign n13939 = n13938 ^ n13896;
  assign n13940 = n13926 & ~n13939;
  assign n13941 = n13940 ^ n13922;
  assign n13943 = n13942 ^ n13941;
  assign n13933 = n13910 ^ n13884;
  assign n13934 = n13933 ^ n13903;
  assign n13935 = n13917 ^ n13883;
  assign n13936 = n13934 & n13935;
  assign n13937 = n13936 ^ n13928;
  assign n13944 = n13943 ^ n13937;
  assign n13983 = n13932 & n13944;
  assign n13984 = n13953 & n13983;
  assign n13956 = ~n13884 & n13910;
  assign n13957 = n13956 ^ n13949;
  assign n13954 = n13946 ^ n13925;
  assign n13955 = n13954 ^ n13941;
  assign n13958 = n13957 ^ n13955;
  assign n13959 = n13944 & ~n13958;
  assign n13945 = n13944 ^ n13932;
  assign n13982 = n13959 ^ n13945;
  assign n13985 = n13984 ^ n13982;
  assign n13966 = n13958 ^ n13953;
  assign n13967 = n13966 ^ n13959;
  assign n13964 = ~n13932 & ~n13958;
  assign n13965 = ~n13953 & n13964;
  assign n13968 = n13967 ^ n13965;
  assign n13986 = n13985 ^ n13968;
  assign n13991 = n13903 & n13986;
  assign n13960 = n13959 ^ n13953;
  assign n13961 = ~n13945 & n13960;
  assign n13962 = n13961 ^ n13932;
  assign n13988 = n13985 ^ n13962;
  assign n13989 = ~n13925 & n13988;
  assign n13987 = ~n13918 & n13986;
  assign n13990 = n13989 ^ n13987;
  assign n13992 = n13991 ^ n13990;
  assign n13969 = n13959 ^ n13932;
  assign n13970 = ~n13966 & ~n13969;
  assign n13971 = n13970 ^ n13953;
  assign n13977 = n13971 ^ n13962;
  assign n13979 = n13921 & ~n13977;
  assign n13978 = n13896 & ~n13977;
  assign n13980 = n13979 ^ n13978;
  assign n13974 = ~n13883 & n13971;
  assign n13972 = n13971 ^ n13968;
  assign n13973 = ~n13917 & ~n13972;
  assign n13975 = n13974 ^ n13973;
  assign n13963 = ~n13897 & ~n13962;
  assign n13976 = n13975 ^ n13963;
  assign n13981 = n13980 ^ n13976;
  assign n13993 = n13992 ^ n13981;
  assign n17138 = n14242 ^ n13993;
  assign n14252 = n13986 ^ n13977;
  assign n14253 = n13926 & ~n14252;
  assign n14254 = n14253 ^ n13978;
  assign n14249 = n13934 & ~n13968;
  assign n14398 = n14254 ^ n14249;
  assign n14311 = ~n13939 & ~n14252;
  assign n14312 = n14311 ^ n13979;
  assign n14245 = ~n13927 & ~n13972;
  assign n14244 = n13935 & ~n13968;
  assign n14246 = n14245 ^ n14244;
  assign n14247 = n14246 ^ n13973;
  assign n14397 = n14312 ^ n14247;
  assign n14399 = n14398 ^ n14397;
  assign n13664 = n12963 ^ n12946;
  assign n13665 = n13664 ^ n13092;
  assign n13666 = n13665 ^ n12937;
  assign n13668 = n13667 ^ n13666;
  assign n13637 = n13059 ^ n12972;
  assign n13636 = n13070 ^ n13030;
  assign n13638 = n13637 ^ n13636;
  assign n13635 = n13634 ^ n12978;
  assign n13639 = n13638 ^ n13635;
  assign n13614 = n13041 ^ n13035;
  assign n13613 = n13045 ^ n12374;
  assign n13615 = n13614 ^ n13613;
  assign n13612 = n13611 ^ n13070;
  assign n13616 = n13615 ^ n13612;
  assign n13640 = n13639 ^ n13616;
  assign n13669 = n13668 ^ n13640;
  assign n13646 = n13089 ^ n12963;
  assign n13647 = n13646 ^ n12946;
  assign n13645 = n12927 ^ n12889;
  assign n13648 = n13647 ^ n13645;
  assign n13644 = n13643 ^ n12900;
  assign n13649 = n13648 ^ n13644;
  assign n13683 = n13669 ^ n13649;
  assign n13621 = n12968 ^ n12620;
  assign n13620 = n13062 ^ n12978;
  assign n13622 = n13621 ^ n13620;
  assign n13619 = n13618 ^ n12751;
  assign n13623 = n13622 ^ n13619;
  assign n13608 = n12933 ^ n12900;
  assign n13607 = n12884 ^ n12871;
  assign n13609 = n13608 ^ n13607;
  assign n13606 = n13605 ^ n13012;
  assign n13610 = n13609 ^ n13606;
  assign n13633 = n13623 ^ n13610;
  assign n13684 = n13683 ^ n13633;
  assign n13703 = ~n13649 & n13669;
  assign n13653 = n13001 ^ n12611;
  assign n13651 = n12963 ^ n12857;
  assign n13652 = n13651 ^ n13013;
  assign n13654 = n13653 ^ n13652;
  assign n13642 = n13641 ^ n12742;
  assign n13650 = n13649 ^ n13642;
  assign n13655 = n13654 ^ n13650;
  assign n13617 = n13616 ^ n13610;
  assign n13663 = n13655 ^ n13617;
  assign n13674 = n13649 ^ n13623;
  assign n13675 = n13663 & n13674;
  assign n13704 = n13703 ^ n13675;
  assign n13701 = n13674 ^ n13663;
  assign n13627 = n12997 ^ n12963;
  assign n13628 = n13627 ^ n12752;
  assign n13626 = n12625 ^ n12491;
  assign n13629 = n13628 ^ n13626;
  assign n13625 = n13624 ^ n13045;
  assign n13630 = n13629 ^ n13625;
  assign n13631 = n13630 ^ n13623;
  assign n13632 = n13631 ^ n13617;
  assign n13680 = n13630 ^ n13610;
  assign n13689 = n13632 & n13680;
  assign n13659 = n13639 ^ n13610;
  assign n13660 = n13659 ^ n13655;
  assign n13661 = n13631 & n13660;
  assign n13690 = n13689 ^ n13661;
  assign n13702 = n13701 ^ n13690;
  assign n13705 = n13704 ^ n13702;
  assign n13671 = n13669 ^ n13630;
  assign n13672 = n13671 ^ n13631;
  assign n13670 = n13669 ^ n13663;
  assign n13678 = n13672 ^ n13670;
  assign n13673 = n13670 & n13672;
  assign n13676 = n13675 ^ n13673;
  assign n13656 = n13655 ^ n13631;
  assign n13657 = n13656 ^ n13640;
  assign n13658 = n13633 & n13657;
  assign n13662 = n13661 ^ n13658;
  assign n13677 = n13676 ^ n13662;
  assign n13679 = n13678 ^ n13677;
  assign n13711 = n13705 ^ n13679;
  assign n13688 = n13659 ^ n13656;
  assign n13691 = n13690 ^ n13688;
  assign n13685 = n13668 ^ n13656;
  assign n13686 = n13684 & n13685;
  assign n13681 = n13680 ^ n13674;
  assign n13682 = n13656 & n13681;
  assign n13687 = n13686 ^ n13682;
  assign n13692 = n13691 ^ n13687;
  assign n13706 = n13692 & n13705;
  assign n13712 = n13711 ^ n13706;
  assign n13695 = n13657 ^ n13633;
  assign n13693 = n13668 & n13671;
  assign n13694 = n13693 ^ n13682;
  assign n13696 = n13695 ^ n13694;
  assign n13697 = n13696 ^ n13662;
  assign n13709 = n13697 & n13705;
  assign n13710 = ~n13679 & n13709;
  assign n13713 = n13712 ^ n13710;
  assign n13736 = n13684 & n13713;
  assign n13718 = n13706 ^ n13697;
  assign n13719 = n13711 & n13718;
  assign n13720 = n13719 ^ n13679;
  assign n13700 = n13697 ^ n13692;
  assign n13715 = n13706 ^ n13679;
  assign n13716 = n13700 & n13715;
  assign n13717 = n13716 ^ n13697;
  assign n13721 = n13720 ^ n13717;
  assign n13734 = n13631 & n13721;
  assign n13707 = n13706 ^ n13700;
  assign n13698 = n13692 & ~n13697;
  assign n13699 = n13679 & n13698;
  assign n13708 = n13707 ^ n13699;
  assign n13714 = n13713 ^ n13708;
  assign n13722 = n13721 ^ n13714;
  assign n13733 = n13680 & n13722;
  assign n13735 = n13734 ^ n13733;
  assign n13737 = n13736 ^ n13735;
  assign n13726 = n13720 ^ n13713;
  assign n13730 = n13656 & n13726;
  assign n13728 = n13685 & n13713;
  assign n13727 = n13681 & n13726;
  assign n13729 = n13728 ^ n13727;
  assign n13731 = n13730 ^ n13729;
  assign n13724 = n13660 & n13721;
  assign n13723 = n13632 & n13722;
  assign n13725 = n13724 ^ n13723;
  assign n13732 = n13731 ^ n13725;
  assign n13738 = n13737 ^ n13732;
  assign n17137 = n14399 ^ n13738;
  assign n17139 = n17138 ^ n17137;
  assign n17142 = n17141 ^ n17139;
  assign n14226 = n13787 & n13839;
  assign n14223 = n13834 ^ n13825;
  assign n14224 = ~n13783 & n14223;
  assign n14222 = ~n13788 & n13839;
  assign n14225 = n14224 ^ n14222;
  assign n14227 = n14226 ^ n14225;
  assign n14220 = n13851 ^ n13842;
  assign n14217 = ~n13761 & n13829;
  assign n14218 = n14217 ^ n13848;
  assign n14216 = ~n13816 & ~n13825;
  assign n14219 = n14218 ^ n14216;
  assign n14221 = n14220 ^ n14219;
  assign n14228 = n14227 ^ n14221;
  assign n17135 = n17134 ^ n14228;
  assign n14336 = ~n14055 & ~n14116;
  assign n14125 = ~n14087 & n14097;
  assign n14383 = n14336 ^ n14125;
  assign n14104 = n14088 & n14097;
  assign n14103 = n14078 & n14101;
  assign n14105 = n14104 ^ n14103;
  assign n14106 = n14105 ^ n14102;
  assign n14459 = n14383 ^ n14106;
  assign n14302 = n14059 & n14236;
  assign n14118 = n14117 ^ n14111;
  assign n14123 = n14068 & n14118;
  assign n14124 = n14123 ^ n14122;
  assign n14303 = n14302 ^ n14124;
  assign n14460 = n14459 ^ n14303;
  assign n14255 = n13946 & n13988;
  assign n14256 = n14255 ^ n14254;
  assign n14248 = ~n13884 & ~n13985;
  assign n14250 = n14249 ^ n14248;
  assign n14251 = n14250 ^ n14247;
  assign n14257 = n14256 ^ n14251;
  assign n17132 = n14460 ^ n14257;
  assign n13868 = n13633 & n13714;
  assign n13865 = n13717 ^ n13708;
  assign n13866 = n13674 & n13865;
  assign n13864 = n13657 & n13714;
  assign n13867 = n13866 ^ n13864;
  assign n13869 = n13868 ^ n13867;
  assign n13862 = n13734 ^ n13724;
  assign n13859 = n13668 & n13720;
  assign n13860 = n13859 ^ n13730;
  assign n13858 = n13672 & n13717;
  assign n13861 = n13860 ^ n13858;
  assign n13863 = n13862 ^ n13861;
  assign n13870 = n13869 ^ n13863;
  assign n13994 = n13993 ^ n13870;
  assign n17133 = n17132 ^ n13994;
  assign n17136 = n17135 ^ n17133;
  assign n17143 = n17142 ^ n17136;
  assign n14287 = ~n13817 & ~n13825;
  assign n14286 = n13797 & ~n13834;
  assign n14288 = n14287 ^ n14286;
  assign n14289 = n14288 ^ n14218;
  assign n14283 = n13808 & n14223;
  assign n14284 = n14283 ^ n13853;
  assign n14285 = n14284 ^ n14224;
  assign n14290 = n14289 ^ n14285;
  assign n17129 = n17128 ^ n14290;
  assign n14119 = ~n14069 & n14118;
  assign n14120 = n14119 ^ n14112;
  assign n14401 = n14383 ^ n14120;
  assign n14400 = n14303 ^ n14103;
  assign n14402 = n14401 ^ n14400;
  assign n14313 = n14312 ^ n14250;
  assign n14310 = n14256 ^ n14245;
  assign n14314 = n14313 ^ n14310;
  assign n17126 = n14402 ^ n14314;
  assign n14331 = ~n13947 & ~n13962;
  assign n14330 = n13933 & ~n13985;
  assign n14332 = n14331 ^ n14330;
  assign n14333 = n14332 ^ n13975;
  assign n14329 = n14256 ^ n13989;
  assign n14334 = n14333 ^ n14329;
  assign n14321 = n13683 & n13708;
  assign n14320 = n13670 & n13717;
  assign n14322 = n14321 ^ n14320;
  assign n14323 = n14322 ^ n13860;
  assign n14258 = n13663 & n13865;
  assign n14259 = n14258 ^ n13735;
  assign n14319 = n14259 ^ n13866;
  assign n14324 = n14323 ^ n14319;
  assign n17125 = n14334 ^ n14324;
  assign n17127 = n17126 ^ n17125;
  assign n17130 = n17129 ^ n17127;
  assign n17144 = n17143 ^ n17130;
  assign n14348 = ~n13767 & ~n13834;
  assign n14370 = n14348 ^ n13854;
  assign n14448 = n14370 ^ n13849;
  assign n14449 = n14448 ^ n14284;
  assign n17121 = n17120 ^ n14449;
  assign n14306 = ~n14060 & ~n14110;
  assign n14436 = n14306 ^ n14230;
  assign n14437 = n14436 ^ n14105;
  assign n14435 = n14383 ^ n14124;
  assign n14438 = n14437 ^ n14435;
  assign n17117 = n14438 ^ n14402;
  assign n14454 = n14331 ^ n13974;
  assign n14455 = n14454 ^ n14246;
  assign n14453 = n14254 ^ n14250;
  assign n14456 = n14455 ^ n14453;
  assign n14457 = n14456 ^ n14314;
  assign n17118 = n17117 ^ n14457;
  assign n14260 = n13669 & n13708;
  assign n14261 = n14260 ^ n13736;
  assign n14262 = n14261 ^ n13731;
  assign n14263 = n14262 ^ n14259;
  assign n14264 = n14263 ^ n14257;
  assign n17119 = n17118 ^ n14264;
  assign n17122 = n17121 ^ n17119;
  assign n17181 = n17144 ^ n17122;
  assign n14364 = n14311 ^ n13990;
  assign n14365 = n14364 ^ n14332;
  assign n14363 = n14254 ^ n14248;
  assign n14366 = n14365 ^ n14363;
  assign n14338 = n14239 ^ n14119;
  assign n14305 = ~n14086 & ~n14116;
  assign n14307 = n14306 ^ n14305;
  assign n14339 = n14338 ^ n14307;
  assign n14337 = n14336 ^ n14124;
  assign n14340 = n14339 ^ n14337;
  assign n17149 = n14366 ^ n14340;
  assign n14430 = ~n13890 & n13971;
  assign n14431 = n14430 ^ n14250;
  assign n14432 = n14431 ^ n13976;
  assign n14429 = n14364 ^ n14256;
  assign n14433 = n14432 ^ n14429;
  assign n14376 = n13671 & n13720;
  assign n14377 = n14376 ^ n14261;
  assign n14378 = n14377 ^ n13861;
  assign n14342 = n13867 ^ n13723;
  assign n14375 = n14342 ^ n14259;
  assign n14379 = n14378 ^ n14375;
  assign n17148 = n14433 ^ n14379;
  assign n17150 = n17149 ^ n17148;
  assign n14369 = ~n13768 & n13829;
  assign n14371 = n14370 ^ n14369;
  assign n14372 = n14371 ^ n14219;
  assign n14350 = n14225 ^ n13841;
  assign n14368 = n14350 ^ n14284;
  assign n14373 = n14372 ^ n14368;
  assign n17147 = n17146 ^ n14373;
  assign n17151 = n17150 ^ n17147;
  assign n17152 = n17151 ^ n17136;
  assign n14418 = n14287 ^ n14217;
  assign n14419 = n14418 ^ n13847;
  assign n14417 = n14370 ^ n13853;
  assign n14420 = n14419 ^ n14417;
  assign n17108 = n17107 ^ n14420;
  assign n14382 = ~n14056 & n14100;
  assign n14384 = n14383 ^ n14382;
  assign n14385 = n14384 ^ n14233;
  assign n14381 = n14338 ^ n14303;
  assign n14386 = n14385 ^ n14381;
  assign n17105 = n14402 ^ n14386;
  assign n14434 = n14433 ^ n14314;
  assign n17106 = n17105 ^ n14434;
  assign n17109 = n17108 ^ n17106;
  assign n14351 = n14350 ^ n14288;
  assign n14349 = n14348 ^ n13853;
  assign n14352 = n14351 ^ n14349;
  assign n17102 = n17101 ^ n14352;
  assign n14308 = n14307 ^ n14231;
  assign n14304 = n14303 ^ n14237;
  assign n14309 = n14308 ^ n14304;
  assign n17098 = n14402 ^ n14309;
  assign n14335 = n14334 ^ n14314;
  assign n17099 = n17098 ^ n14335;
  assign n14344 = n14260 ^ n13735;
  assign n14343 = n14342 ^ n14322;
  assign n14345 = n14344 ^ n14343;
  assign n14367 = n14366 ^ n14345;
  assign n17100 = n17099 ^ n14367;
  assign n17103 = n17102 ^ n17100;
  assign n14442 = n14320 ^ n13859;
  assign n14443 = n14442 ^ n13729;
  assign n14441 = n14261 ^ n13735;
  assign n14444 = n14443 ^ n14441;
  assign n17097 = n14456 ^ n14444;
  assign n17104 = n17103 ^ n17097;
  assign n17110 = n17109 ^ n17104;
  assign n17153 = n17152 ^ n17110;
  assign n17183 = n17153 ^ n17144;
  assign n14407 = n14370 ^ n13843;
  assign n14406 = n14284 ^ n13845;
  assign n14408 = n14407 ^ n14406;
  assign n17115 = n17114 ^ n14408;
  assign n14126 = n14125 ^ n14124;
  assign n14121 = n14120 ^ n14106;
  assign n14127 = n14126 ^ n14121;
  assign n17112 = n14399 ^ n14127;
  assign n14317 = n14261 ^ n13725;
  assign n14316 = n14259 ^ n13727;
  assign n14318 = n14317 ^ n14316;
  assign n17111 = n14318 ^ n14314;
  assign n17113 = n17112 ^ n17111;
  assign n17116 = n17115 ^ n17113;
  assign n17123 = n17122 ^ n17116;
  assign n17182 = n17181 ^ n17123;
  assign n17187 = n17183 ^ n17182;
  assign n17184 = ~n17182 & n17183;
  assign n17154 = n17116 ^ n17103;
  assign n17155 = ~n17153 & n17154;
  assign n17185 = n17184 ^ n17155;
  assign n17168 = n17151 ^ n17116;
  assign n17124 = n17123 ^ n17110;
  assign n17178 = n17143 ^ n17124;
  assign n17179 = ~n17168 & ~n17178;
  assign n17160 = n17151 ^ n17142;
  assign n17161 = n17160 ^ n17110;
  assign n17162 = ~n17123 & ~n17161;
  assign n17180 = n17179 ^ n17162;
  assign n17186 = n17185 ^ n17180;
  assign n17188 = n17187 ^ n17186;
  assign n17164 = n17154 ^ n17153;
  assign n17157 = n17151 ^ n17122;
  assign n17158 = n17152 ^ n17123;
  assign n17159 = n17157 & n17158;
  assign n17163 = n17162 ^ n17159;
  assign n17165 = n17164 ^ n17163;
  assign n17145 = ~n17103 & ~n17144;
  assign n17156 = n17155 ^ n17145;
  assign n17166 = n17165 ^ n17156;
  assign n17189 = n17188 ^ n17166;
  assign n17193 = n17178 ^ n17168;
  assign n17191 = ~n17130 & n17181;
  assign n17171 = n17157 ^ n17154;
  assign n17172 = ~n17124 & n17171;
  assign n17192 = n17191 ^ n17172;
  assign n17194 = n17193 ^ n17192;
  assign n17195 = n17194 ^ n17180;
  assign n17174 = n17160 ^ n17124;
  assign n17175 = n17174 ^ n17163;
  assign n17131 = n17130 ^ n17124;
  assign n17167 = n17144 ^ n17103;
  assign n17169 = n17168 ^ n17167;
  assign n17170 = n17131 & n17169;
  assign n17173 = n17172 ^ n17170;
  assign n17176 = n17175 ^ n17173;
  assign n17177 = ~n17166 & n17176;
  assign n17200 = n17195 ^ n17177;
  assign n17201 = n17189 & n17200;
  assign n17202 = n17201 ^ n17188;
  assign n17670 = n17181 & ~n17202;
  assign n17208 = n17195 ^ n17176;
  assign n17216 = n17208 ^ n17177;
  assign n17214 = n17176 & ~n17195;
  assign n17215 = ~n17188 & n17214;
  assign n17217 = n17216 ^ n17215;
  assign n17233 = ~n17144 & n17217;
  assign n17196 = ~n17166 & n17195;
  assign n17197 = n17188 & n17196;
  assign n17190 = n17189 ^ n17177;
  assign n17198 = n17197 ^ n17190;
  assign n17226 = n17169 & n17198;
  assign n17234 = n17233 ^ n17226;
  assign n17671 = n17670 ^ n17234;
  assign n17209 = n17188 ^ n17177;
  assign n17210 = n17208 & ~n17209;
  assign n17211 = n17210 ^ n17195;
  assign n17574 = ~n17182 & n17211;
  assign n17494 = ~n17130 & ~n17202;
  assign n17203 = n17202 ^ n17198;
  assign n17206 = ~n17124 & ~n17203;
  assign n17495 = n17494 ^ n17206;
  assign n17575 = n17574 ^ n17495;
  assign n17672 = n17671 ^ n17575;
  assign n17229 = n17217 ^ n17211;
  assign n17487 = n17154 & n17229;
  assign n17218 = n17217 ^ n17198;
  assign n17486 = ~n17178 & n17218;
  assign n17488 = n17487 ^ n17486;
  assign n17212 = n17211 ^ n17202;
  assign n17219 = n17218 ^ n17212;
  assign n17220 = n17158 & ~n17219;
  assign n17489 = n17488 ^ n17220;
  assign n17230 = ~n17153 & n17229;
  assign n17224 = n17157 & ~n17219;
  assign n17223 = ~n17123 & ~n17212;
  assign n17225 = n17224 ^ n17223;
  assign n17231 = n17230 ^ n17225;
  assign n17669 = n17489 ^ n17231;
  assign n17673 = n17672 ^ n17669;
  assign n17213 = ~n17161 & ~n17212;
  assign n17221 = n17220 ^ n17213;
  assign n17235 = n17234 ^ n17221;
  assign n17204 = n17171 & ~n17203;
  assign n17232 = n17231 ^ n17204;
  assign n17236 = n17235 ^ n17232;
  assign n17674 = n17673 ^ n17236;
  assign n17484 = n17183 & n17211;
  assign n17639 = n17494 ^ n17484;
  assign n17199 = n17131 & n17198;
  assign n17205 = n17204 ^ n17199;
  assign n17640 = n17639 ^ n17205;
  assign n17638 = n17234 ^ n17225;
  assign n17641 = n17640 ^ n17638;
  assign n17675 = n17674 ^ n17641;
  assign n17690 = n17689 ^ n17675;
  assign n15066 = n12155 ^ n10074;
  assign n15065 = n14050 ^ n10254;
  assign n15067 = n15066 ^ n15065;
  assign n15063 = n12007 ^ n10280;
  assign n15061 = n10144 ^ n10128;
  assign n15060 = n10271 ^ n10173;
  assign n15062 = n15061 ^ n15060;
  assign n15064 = n15063 ^ n15062;
  assign n15068 = n15067 ^ n15064;
  assign n15057 = n11945 ^ n10144;
  assign n15042 = n10197 ^ n10074;
  assign n15055 = n15042 ^ n10133;
  assign n15056 = n15055 ^ n14038;
  assign n15058 = n15057 ^ n15056;
  assign n15051 = n12127 ^ n10253;
  assign n15050 = n14003 ^ n10229;
  assign n15052 = n15051 ^ n15050;
  assign n15048 = n12051 ^ n10223;
  assign n15047 = n14025 ^ n9947;
  assign n15049 = n15048 ^ n15047;
  assign n15053 = n15052 ^ n15049;
  assign n15043 = n15042 ^ n9959;
  assign n15044 = n15043 ^ n10117;
  assign n15045 = n15044 ^ n10191;
  assign n15046 = n15045 ^ n12093;
  assign n15054 = n15053 ^ n15046;
  assign n15059 = n15058 ^ n15054;
  assign n15069 = n15068 ^ n15059;
  assign n15091 = n15064 ^ n15049;
  assign n15073 = n10280 ^ n10074;
  assign n15074 = n15073 ^ n10183;
  assign n15072 = n10163 ^ n8100;
  assign n15075 = n15074 ^ n15072;
  assign n15070 = n11522 ^ n10091;
  assign n15071 = n15070 ^ n15058;
  assign n15076 = n15075 ^ n15071;
  assign n15101 = n15091 ^ n15076;
  assign n15121 = n15101 ^ n15054;
  assign n15080 = n12115 ^ n9038;
  assign n15077 = n10091 ^ n10074;
  assign n15078 = n15077 ^ n9960;
  assign n15079 = n15078 ^ n14030;
  assign n15081 = n15080 ^ n15079;
  assign n15109 = n15081 ^ n15054;
  assign n15082 = n15081 ^ n15067;
  assign n15120 = n15109 ^ n15082;
  assign n15125 = n15121 ^ n15120;
  assign n15122 = ~n15120 & ~n15121;
  assign n15087 = n15067 ^ n15058;
  assign n15105 = ~n15087 & n15101;
  assign n15123 = n15122 ^ n15105;
  assign n15083 = n15082 ^ n15076;
  assign n15112 = n15083 ^ n15053;
  assign n15115 = n15068 & ~n15112;
  assign n15094 = n15064 ^ n15052;
  assign n15095 = n15094 ^ n15076;
  assign n15096 = n15082 & n15095;
  assign n15116 = n15115 ^ n15096;
  assign n15124 = n15123 ^ n15116;
  assign n15126 = n15125 ^ n15124;
  assign n15104 = ~n15054 & n15058;
  assign n15106 = n15105 ^ n15104;
  assign n15102 = n15101 ^ n15087;
  assign n15086 = n15081 ^ n15064;
  assign n15092 = n15091 ^ n15082;
  assign n15093 = n15086 & ~n15092;
  assign n15097 = n15096 ^ n15093;
  assign n15103 = n15102 ^ n15097;
  assign n15107 = n15106 ^ n15103;
  assign n15131 = n15126 ^ n15107;
  assign n15098 = n15094 ^ n15083;
  assign n15099 = n15098 ^ n15097;
  assign n15088 = n15087 ^ n15086;
  assign n15089 = ~n15083 & ~n15088;
  assign n15084 = n15083 ^ n15046;
  assign n15085 = n15069 & n15084;
  assign n15090 = n15089 ^ n15085;
  assign n15100 = n15099 ^ n15090;
  assign n15108 = n15100 & ~n15107;
  assign n15142 = n15131 ^ n15108;
  assign n15113 = n15112 ^ n15068;
  assign n15110 = ~n15046 & ~n15109;
  assign n15111 = n15110 ^ n15089;
  assign n15114 = n15113 ^ n15111;
  assign n15117 = n15116 ^ n15114;
  assign n15140 = ~n15107 & ~n15117;
  assign n15141 = ~n15126 & n15140;
  assign n15143 = n15142 ^ n15141;
  assign n15181 = n15069 & ~n15143;
  assign n15127 = n15100 & n15117;
  assign n15128 = n15126 & n15127;
  assign n15118 = n15117 ^ n15100;
  assign n15119 = n15118 ^ n15108;
  assign n15129 = n15128 ^ n15119;
  assign n15130 = ~n15054 & ~n15129;
  assign n15182 = n15181 ^ n15130;
  assign n15135 = n15126 ^ n15108;
  assign n15136 = ~n15118 & n15135;
  assign n15137 = n15136 ^ n15117;
  assign n15132 = n15117 ^ n15108;
  assign n15133 = ~n15131 & ~n15132;
  assign n15134 = n15133 ^ n15126;
  assign n15138 = n15137 ^ n15134;
  assign n15179 = n15095 & ~n15138;
  assign n15144 = n15143 ^ n15129;
  assign n15145 = n15144 ^ n15138;
  assign n15152 = ~n15092 & ~n15145;
  assign n15180 = n15179 ^ n15152;
  assign n15183 = n15182 ^ n15180;
  assign n15176 = n15143 ^ n15134;
  assign n15177 = ~n15088 & ~n15176;
  assign n15153 = n15137 ^ n15129;
  assign n15174 = n15101 & n15153;
  assign n15146 = n15086 & ~n15145;
  assign n15139 = n15082 & ~n15138;
  assign n15147 = n15146 ^ n15139;
  assign n15175 = n15174 ^ n15147;
  assign n15178 = n15177 ^ n15175;
  assign n15184 = n15183 ^ n15178;
  assign n14588 = n12137 ^ n12065;
  assign n14587 = n12167 ^ n12133;
  assign n14589 = n14588 ^ n14587;
  assign n14586 = n13076 ^ n12043;
  assign n14590 = n14589 ^ n14586;
  assign n14570 = n12098 ^ n12065;
  assign n14571 = n14570 ^ n13875;
  assign n14569 = n13053 ^ n12074;
  assign n14572 = n14571 ^ n14569;
  assign n14600 = n14590 ^ n14572;
  assign n14597 = n12085 ^ n11895;
  assign n14559 = n12160 ^ n12082;
  assign n14598 = n14597 ^ n14559;
  assign n14596 = n13100 ^ n11923;
  assign n14599 = n14598 ^ n14596;
  assign n14601 = n14600 ^ n14599;
  assign n14560 = n14559 ^ n11771;
  assign n14561 = n14560 ^ n13898;
  assign n14558 = n12955 ^ n11924;
  assign n14562 = n14561 ^ n14558;
  assign n14620 = n14601 ^ n14562;
  assign n14566 = n12024 ^ n11771;
  assign n14565 = n12035 ^ n11959;
  assign n14567 = n14566 ^ n14565;
  assign n14564 = n12917 ^ n11932;
  assign n14568 = n14567 ^ n14564;
  assign n14554 = n12160 ^ n12137;
  assign n14553 = n12163 ^ n11905;
  assign n14555 = n14554 ^ n14553;
  assign n14552 = n12986 ^ n12121;
  assign n14556 = n14555 ^ n14552;
  assign n14608 = n14568 ^ n14556;
  assign n14621 = n14620 ^ n14608;
  assign n14563 = n14562 ^ n14556;
  assign n14577 = n12160 ^ n12024;
  assign n14578 = n14577 ^ n11991;
  assign n14576 = n13020 ^ n11968;
  assign n14579 = n14578 ^ n14576;
  assign n14574 = n12106 ^ n11980;
  assign n14575 = n14574 ^ n14562;
  assign n14580 = n14579 ^ n14575;
  assign n14573 = n14572 ^ n14568;
  assign n14581 = n14580 ^ n14573;
  assign n14603 = ~n14563 & n14581;
  assign n14602 = n14562 & ~n14601;
  assign n14604 = n14603 ^ n14602;
  assign n14548 = n12160 ^ n11991;
  assign n14549 = n14548 ^ n12098;
  assign n14550 = n14549 ^ n13871;
  assign n14547 = n12840 ^ n12108;
  assign n14551 = n14550 ^ n14547;
  assign n14557 = n14556 ^ n14551;
  assign n14591 = n14590 ^ n14568;
  assign n14592 = n14591 ^ n14580;
  assign n14593 = n14557 & n14592;
  assign n14583 = n14568 ^ n14551;
  assign n14584 = n14573 ^ n14557;
  assign n14585 = n14583 & ~n14584;
  assign n14594 = n14593 ^ n14585;
  assign n14582 = n14581 ^ n14563;
  assign n14595 = n14594 ^ n14582;
  assign n14605 = n14604 ^ n14595;
  assign n14606 = n14580 ^ n14557;
  assign n14627 = n14606 ^ n14591;
  assign n14628 = n14627 ^ n14594;
  assign n14624 = n14583 ^ n14563;
  assign n14625 = ~n14606 & ~n14624;
  assign n14622 = n14606 ^ n14599;
  assign n14623 = n14621 & n14622;
  assign n14626 = n14625 ^ n14623;
  assign n14629 = n14628 ^ n14626;
  assign n14630 = ~n14605 & n14629;
  assign n14613 = n14601 ^ n14581;
  assign n14611 = n14601 ^ n14551;
  assign n14612 = n14611 ^ n14557;
  assign n14617 = n14613 ^ n14612;
  assign n14614 = ~n14612 & ~n14613;
  assign n14615 = n14614 ^ n14603;
  assign n14607 = n14606 ^ n14600;
  assign n14609 = ~n14607 & n14608;
  assign n14610 = n14609 ^ n14593;
  assign n14616 = n14615 ^ n14610;
  assign n14618 = n14617 ^ n14616;
  assign n14619 = n14618 ^ n14605;
  assign n14647 = n14630 ^ n14619;
  assign n14633 = n14608 ^ n14607;
  assign n14631 = ~n14599 & ~n14611;
  assign n14632 = n14631 ^ n14625;
  assign n14634 = n14633 ^ n14632;
  assign n14635 = n14634 ^ n14610;
  assign n14645 = ~n14605 & ~n14635;
  assign n14646 = ~n14618 & n14645;
  assign n14648 = n14647 ^ n14646;
  assign n14677 = n14621 & ~n14648;
  assign n14650 = n14629 & n14635;
  assign n14651 = n14618 & n14650;
  assign n14639 = n14635 ^ n14629;
  assign n14649 = n14639 ^ n14630;
  assign n14652 = n14651 ^ n14649;
  assign n14676 = ~n14601 & ~n14652;
  assign n14678 = n14677 ^ n14676;
  assign n14653 = n14652 ^ n14648;
  assign n14640 = n14630 ^ n14618;
  assign n14641 = ~n14639 & n14640;
  assign n14642 = n14641 ^ n14635;
  assign n14636 = n14635 ^ n14630;
  assign n14637 = ~n14619 & ~n14636;
  assign n14638 = n14637 ^ n14618;
  assign n14643 = n14642 ^ n14638;
  assign n14654 = n14653 ^ n14643;
  assign n14674 = ~n14584 & ~n14654;
  assign n14673 = n14592 & ~n14643;
  assign n14675 = n14674 ^ n14673;
  assign n14679 = n14678 ^ n14675;
  assign n14666 = n14648 ^ n14638;
  assign n14671 = ~n14624 & ~n14666;
  assign n14657 = n14652 ^ n14642;
  assign n14658 = n14581 & n14657;
  assign n14655 = n14583 & ~n14654;
  assign n14644 = n14557 & ~n14643;
  assign n14656 = n14655 ^ n14644;
  assign n14659 = n14658 ^ n14656;
  assign n14672 = n14671 ^ n14659;
  assign n14680 = n14679 ^ n14672;
  assign n14667 = ~n14606 & ~n14666;
  assign n14665 = ~n14599 & n14638;
  assign n14668 = n14667 ^ n14665;
  assign n14663 = n14620 & ~n14652;
  assign n14662 = ~n14613 & ~n14642;
  assign n14664 = n14663 ^ n14662;
  assign n14669 = n14668 ^ n14664;
  assign n14660 = ~n14563 & n14657;
  assign n14661 = n14660 ^ n14659;
  assign n14670 = n14669 ^ n14661;
  assign n14681 = n14680 ^ n14670;
  assign n17017 = n15184 ^ n14681;
  assign n14957 = n11229 ^ n11083;
  assign n14955 = n11126 ^ n10742;
  assign n14956 = n14955 ^ n11220;
  assign n14958 = n14957 ^ n14956;
  assign n14952 = n11166 ^ n10154;
  assign n14950 = n11158 ^ n10486;
  assign n14931 = n11202 ^ n11126;
  assign n14949 = n14931 ^ n11148;
  assign n14951 = n14950 ^ n14949;
  assign n14953 = n14952 ^ n14951;
  assign n14948 = n11234 ^ n10098;
  assign n14954 = n14953 ^ n14948;
  assign n14959 = n14958 ^ n14954;
  assign n14925 = n11220 ^ n11126;
  assign n14924 = n11106 ^ n11077;
  assign n14926 = n14925 ^ n14924;
  assign n14927 = n14926 ^ n11098;
  assign n14928 = n14927 ^ n11034;
  assign n14929 = n14928 ^ n10049;
  assign n14921 = n11187 ^ n11088;
  assign n14920 = n11132 ^ n11126;
  assign n14922 = n14921 ^ n14920;
  assign n14923 = n14922 ^ n10081;
  assign n14930 = n14929 ^ n14923;
  assign n14960 = n14959 ^ n14930;
  assign n14961 = n11149 ^ n10918;
  assign n14962 = n14961 ^ n10742;
  assign n14963 = n14962 ^ n11227;
  assign n14964 = n14963 ^ n10289;
  assign n14940 = n11061 ^ n11047;
  assign n14941 = n14940 ^ n11182;
  assign n14942 = n14941 ^ n11078;
  assign n14943 = n14942 ^ n10239;
  assign n14986 = n14964 ^ n14943;
  assign n14993 = n14986 ^ n14959;
  assign n14938 = n11191 ^ n10260;
  assign n14936 = n11118 ^ n11054;
  assign n14937 = n14936 ^ n11186;
  assign n14939 = n14938 ^ n14937;
  assign n14944 = n14943 ^ n14939;
  assign n14934 = n11207 ^ n10202;
  assign n14932 = n11153 ^ n11097;
  assign n14933 = n14932 ^ n14931;
  assign n14935 = n14934 ^ n14933;
  assign n14945 = n14944 ^ n14935;
  assign n15002 = n14993 ^ n14945;
  assign n14946 = n14945 ^ n14929;
  assign n15001 = n14946 ^ n14930;
  assign n15006 = n15002 ^ n15001;
  assign n15003 = ~n15001 & ~n15002;
  assign n14966 = n14953 ^ n14923;
  assign n14996 = ~n14966 & n14993;
  assign n15004 = n15003 ^ n14996;
  assign n14975 = n14964 ^ n14939;
  assign n14976 = n14975 ^ n14959;
  assign n14977 = n14930 & n14976;
  assign n14970 = n14960 ^ n14944;
  assign n14971 = n14964 ^ n14923;
  assign n14974 = ~n14970 & n14971;
  assign n14978 = n14977 ^ n14974;
  assign n15005 = n15004 ^ n14978;
  assign n15007 = n15006 ^ n15005;
  assign n14997 = ~n14945 & n14953;
  assign n14998 = n14997 ^ n14996;
  assign n14994 = n14993 ^ n14966;
  assign n14965 = n14964 ^ n14929;
  assign n14987 = n14986 ^ n14930;
  assign n14988 = n14965 & ~n14987;
  assign n14989 = n14988 ^ n14977;
  assign n14995 = n14994 ^ n14989;
  assign n14999 = n14998 ^ n14995;
  assign n15011 = n15007 ^ n14999;
  assign n14985 = n14975 ^ n14960;
  assign n14990 = n14989 ^ n14985;
  assign n14980 = n14953 ^ n14945;
  assign n14981 = n14980 ^ n14971;
  assign n14982 = n14960 ^ n14935;
  assign n14983 = n14981 & n14982;
  assign n14967 = n14966 ^ n14965;
  assign n14968 = ~n14960 & ~n14967;
  assign n14984 = n14983 ^ n14968;
  assign n14991 = n14990 ^ n14984;
  assign n15000 = n14991 & ~n14999;
  assign n15023 = n15011 ^ n15000;
  assign n14972 = n14971 ^ n14970;
  assign n14947 = ~n14935 & ~n14946;
  assign n14969 = n14968 ^ n14947;
  assign n14973 = n14972 ^ n14969;
  assign n14979 = n14978 ^ n14973;
  assign n15021 = ~n14979 & ~n14999;
  assign n15022 = ~n15007 & n15021;
  assign n15024 = n15023 ^ n15022;
  assign n15012 = n15000 ^ n14979;
  assign n15013 = ~n15011 & ~n15012;
  assign n15014 = n15013 ^ n15007;
  assign n15163 = n15024 ^ n15014;
  assign n15290 = ~n14960 & ~n15163;
  assign n15228 = ~n14935 & n15014;
  assign n15304 = n15290 ^ n15228;
  assign n14992 = n14991 ^ n14979;
  assign n15008 = n15007 ^ n15000;
  assign n15009 = ~n14992 & n15008;
  assign n15010 = n15009 ^ n14979;
  assign n15032 = ~n15002 & ~n15010;
  assign n15018 = n14979 & n14991;
  assign n15019 = n15007 & n15018;
  assign n15017 = n15000 ^ n14992;
  assign n15020 = n15019 ^ n15017;
  assign n15031 = n14980 & ~n15020;
  assign n15033 = n15032 ^ n15031;
  assign n15305 = n15304 ^ n15033;
  assign n15036 = n15020 ^ n15010;
  assign n15165 = n14993 & n15036;
  assign n15025 = n15024 ^ n15020;
  assign n15015 = n15014 ^ n15010;
  assign n15026 = n15025 ^ n15015;
  assign n15027 = n14965 & ~n15026;
  assign n15016 = n14930 & ~n15015;
  assign n15028 = n15027 ^ n15016;
  assign n15166 = n15165 ^ n15028;
  assign n15037 = ~n14966 & n15036;
  assign n15303 = n15166 ^ n15037;
  assign n15306 = n15305 ^ n15303;
  assign n17018 = n17017 ^ n15306;
  assign n14832 = n13621 ^ n13093;
  assign n14831 = n14712 ^ n12945;
  assign n14833 = n14832 ^ n14831;
  assign n14820 = n14693 ^ n12978;
  assign n14819 = n13614 ^ n13063;
  assign n14821 = n14820 ^ n14819;
  assign n14807 = n14703 ^ n13070;
  assign n14806 = n13626 ^ n13036;
  assign n14808 = n14807 ^ n14806;
  assign n14830 = n14821 ^ n14808;
  assign n14834 = n14833 ^ n14830;
  assign n14813 = n14696 ^ n12742;
  assign n14811 = n12968 ^ n12871;
  assign n14812 = n14811 ^ n13004;
  assign n14814 = n14813 ^ n14812;
  assign n14802 = n14685 ^ n12900;
  assign n14799 = n13092 ^ n12968;
  assign n14800 = n14799 ^ n12938;
  assign n14801 = n14800 ^ n12934;
  assign n14803 = n14802 ^ n14801;
  assign n14810 = n14803 ^ n13002;
  assign n14815 = n14814 ^ n14810;
  assign n14788 = n14691 ^ n13012;
  assign n14787 = n13645 ^ n12872;
  assign n14789 = n14788 ^ n14787;
  assign n14809 = n14808 ^ n14789;
  assign n14816 = n14815 ^ n14809;
  assign n14852 = n14834 ^ n14816;
  assign n14793 = n14688 ^ n13045;
  assign n14790 = n13001 ^ n12968;
  assign n14791 = n14790 ^ n12621;
  assign n14792 = n14791 ^ n12492;
  assign n14794 = n14793 ^ n14792;
  assign n14850 = n14834 ^ n14794;
  assign n14797 = n13637 ^ n12969;
  assign n14796 = n14683 ^ n12751;
  assign n14798 = n14797 ^ n14796;
  assign n14818 = n14798 ^ n14794;
  assign n14851 = n14850 ^ n14818;
  assign n14859 = n14852 ^ n14851;
  assign n14839 = n14798 ^ n14789;
  assign n14841 = n14818 ^ n14815;
  assign n14855 = n14841 ^ n14830;
  assign n14856 = n14839 & ~n14855;
  assign n14822 = n14821 ^ n14789;
  assign n14823 = n14822 ^ n14815;
  assign n14824 = n14818 & ~n14823;
  assign n14857 = n14856 ^ n14824;
  assign n14853 = n14851 & ~n14852;
  assign n14804 = n14803 ^ n14798;
  assign n14829 = n14804 & ~n14816;
  assign n14854 = n14853 ^ n14829;
  assign n14858 = n14857 ^ n14854;
  assign n14860 = n14859 ^ n14858;
  assign n14835 = ~n14803 & n14834;
  assign n14836 = n14835 ^ n14829;
  assign n14795 = n14794 ^ n14789;
  assign n14825 = n14818 ^ n14809;
  assign n14826 = n14795 & n14825;
  assign n14827 = n14826 ^ n14824;
  assign n14817 = n14816 ^ n14804;
  assign n14828 = n14827 ^ n14817;
  assign n14837 = n14836 ^ n14828;
  assign n14861 = n14860 ^ n14837;
  assign n14865 = n14855 ^ n14839;
  assign n14863 = n14833 & n14850;
  assign n14805 = n14804 ^ n14795;
  assign n14844 = n14805 & ~n14841;
  assign n14864 = n14863 ^ n14844;
  assign n14866 = n14865 ^ n14864;
  assign n14867 = n14866 ^ n14857;
  assign n14846 = n14841 ^ n14822;
  assign n14847 = n14846 ^ n14827;
  assign n14838 = n14834 ^ n14803;
  assign n14840 = n14839 ^ n14838;
  assign n14842 = n14841 ^ n14833;
  assign n14843 = n14840 & ~n14842;
  assign n14845 = n14844 ^ n14843;
  assign n14848 = n14847 ^ n14845;
  assign n14849 = ~n14837 & ~n14848;
  assign n14871 = n14867 ^ n14849;
  assign n14872 = n14861 & ~n14871;
  assign n14873 = n14872 ^ n14860;
  assign n14908 = n14833 & ~n14873;
  assign n14868 = ~n14837 & ~n14867;
  assign n14869 = n14860 & n14868;
  assign n14862 = n14861 ^ n14849;
  assign n14870 = n14869 ^ n14862;
  assign n14874 = n14873 ^ n14870;
  assign n14907 = ~n14841 & ~n14874;
  assign n14909 = n14908 ^ n14907;
  assign n14876 = n14867 ^ n14848;
  assign n14877 = n14860 ^ n14849;
  assign n14878 = n14876 & ~n14877;
  assign n14879 = n14878 ^ n14867;
  assign n14905 = ~n14852 & ~n14879;
  assign n14883 = n14876 ^ n14849;
  assign n14881 = ~n14848 & n14867;
  assign n14882 = ~n14860 & n14881;
  assign n14884 = n14883 ^ n14882;
  assign n14904 = n14838 & n14884;
  assign n14906 = n14905 ^ n14904;
  assign n14910 = n14909 ^ n14906;
  assign n14890 = n14884 ^ n14879;
  assign n14902 = n14804 & ~n14890;
  assign n14891 = ~n14816 & ~n14890;
  assign n14880 = n14879 ^ n14873;
  assign n14888 = n14818 & n14880;
  assign n14885 = n14884 ^ n14870;
  assign n14886 = n14885 ^ n14880;
  assign n14887 = n14795 & n14886;
  assign n14889 = n14888 ^ n14887;
  assign n14892 = n14891 ^ n14889;
  assign n14903 = n14902 ^ n14892;
  assign n14911 = n14910 ^ n14903;
  assign n17019 = n17018 ^ n14911;
  assign n17021 = n17020 ^ n17019;
  assign n15198 = n14677 ^ n14656;
  assign n15194 = n14622 & ~n14648;
  assign n15195 = n15194 ^ n14671;
  assign n15196 = n15195 ^ n14667;
  assign n15197 = n15196 ^ n14675;
  assign n15199 = n15198 ^ n15197;
  assign n17014 = n17013 ^ n15199;
  assign n15170 = n14981 & ~n15024;
  assign n15379 = n15170 ^ n15028;
  assign n15226 = n14982 & ~n15024;
  assign n15164 = ~n14967 & ~n15163;
  assign n15227 = n15226 ^ n15164;
  assign n15291 = n15290 ^ n15227;
  assign n15168 = n14976 & ~n15015;
  assign n15034 = ~n14987 & ~n15026;
  assign n15169 = n15168 ^ n15034;
  assign n15378 = n15291 ^ n15169;
  assign n15380 = n15379 ^ n15378;
  assign n14897 = n14840 & n14870;
  assign n15190 = n14897 ^ n14889;
  assign n15186 = ~n14842 & n14870;
  assign n14875 = n14805 & ~n14874;
  assign n15187 = n15186 ^ n14875;
  assign n15188 = n15187 ^ n14907;
  assign n14895 = n14825 & n14886;
  assign n14894 = ~n14823 & n14880;
  assign n14896 = n14895 ^ n14894;
  assign n15189 = n15188 ^ n14896;
  assign n15191 = n15190 ^ n15189;
  assign n17011 = n15380 ^ n15191;
  assign n15363 = n14608 & n14653;
  assign n15239 = ~n14607 & n14653;
  assign n15240 = n15239 ^ n14660;
  assign n15364 = n15363 ^ n15240;
  assign n15361 = n14673 ^ n14644;
  assign n15234 = ~n14612 & ~n14642;
  assign n15235 = n15234 ^ n14668;
  assign n15362 = n15361 ^ n15235;
  assign n15365 = n15364 ^ n15362;
  assign n15348 = n15068 & n15144;
  assign n15155 = ~n15112 & n15144;
  assign n15154 = ~n15087 & n15153;
  assign n15156 = n15155 ^ n15154;
  assign n15349 = n15348 ^ n15156;
  assign n15345 = ~n15120 & ~n15137;
  assign n15294 = ~n15083 & ~n15176;
  assign n15219 = ~n15046 & n15134;
  assign n15308 = n15294 ^ n15219;
  assign n15346 = n15345 ^ n15308;
  assign n15344 = n15179 ^ n15139;
  assign n15347 = n15346 ^ n15344;
  assign n15350 = n15349 ^ n15347;
  assign n17010 = n15365 ^ n15350;
  assign n17012 = n17011 ^ n17010;
  assign n17015 = n17014 ^ n17012;
  assign n15355 = n14971 & n15025;
  assign n15035 = ~n14970 & n15025;
  assign n15038 = n15037 ^ n15035;
  assign n15356 = n15355 ^ n15038;
  assign n15352 = ~n15001 & ~n15010;
  assign n15353 = n15352 ^ n15304;
  assign n15351 = n15168 ^ n15016;
  assign n15354 = n15353 ^ n15351;
  assign n15357 = n15356 ^ n15354;
  assign n15340 = n14839 & n14885;
  assign n14913 = ~n14855 & n14885;
  assign n14914 = n14913 ^ n14902;
  assign n15341 = n15340 ^ n14914;
  assign n15338 = n14894 ^ n14888;
  assign n15258 = n14851 & ~n14879;
  assign n15259 = n15258 ^ n14909;
  assign n15339 = n15338 ^ n15259;
  assign n15342 = n15341 ^ n15339;
  assign n16979 = n15357 ^ n15342;
  assign n15324 = n15196 ^ n14678;
  assign n15325 = n15324 ^ n14659;
  assign n15221 = n15084 & ~n15143;
  assign n15222 = n15221 ^ n15177;
  assign n15295 = n15294 ^ n15222;
  assign n15296 = n15295 ^ n15182;
  assign n15297 = n15296 ^ n15175;
  assign n16978 = n15325 ^ n15297;
  assign n16980 = n16979 ^ n16978;
  assign n16977 = n16976 ^ n15365;
  assign n16981 = n16980 ^ n16977;
  assign n17016 = n17015 ^ n16981;
  assign n17022 = n17021 ^ n17016;
  assign n17001 = n17000 ^ n15325;
  assign n15149 = ~n15121 & ~n15137;
  assign n15220 = n15219 ^ n15149;
  assign n15223 = n15222 ^ n15220;
  assign n15218 = n15182 ^ n15147;
  assign n15224 = n15223 ^ n15218;
  assign n16997 = n15224 ^ n15184;
  assign n15274 = n14678 ^ n14656;
  assign n15272 = n14665 ^ n14662;
  assign n15273 = n15272 ^ n15195;
  assign n15275 = n15274 ^ n15273;
  assign n15276 = n15275 ^ n14680;
  assign n16998 = n16997 ^ n15276;
  assign n15029 = ~n14945 & ~n15020;
  assign n15171 = n15170 ^ n15029;
  assign n15292 = n15291 ^ n15171;
  assign n15293 = n15292 ^ n15166;
  assign n14898 = n14834 & n14884;
  assign n14899 = n14898 ^ n14897;
  assign n15287 = n15188 ^ n14899;
  assign n15288 = n15287 ^ n14892;
  assign n16996 = n15293 ^ n15288;
  assign n16999 = n16998 ^ n16996;
  assign n17002 = n17001 ^ n16999;
  assign n17044 = n17022 ^ n17002;
  assign n16994 = n16993 ^ n14680;
  assign n15172 = n15171 ^ n15169;
  assign n15167 = n15166 ^ n15164;
  assign n15173 = n15172 ^ n15167;
  assign n14900 = n14899 ^ n14896;
  assign n14893 = n14892 ^ n14875;
  assign n14901 = n14900 ^ n14893;
  assign n16991 = n15173 ^ n14901;
  assign n15376 = n15181 ^ n15147;
  assign n15375 = n15295 ^ n15180;
  assign n15377 = n15376 ^ n15375;
  assign n16990 = n15377 ^ n15199;
  assign n16992 = n16991 ^ n16990;
  assign n16995 = n16994 ^ n16992;
  assign n17003 = n17002 ^ n16995;
  assign n17056 = n17044 ^ n17003;
  assign n15241 = n15240 ^ n14674;
  assign n15242 = n15241 ^ n14659;
  assign n15236 = ~n14611 & n14638;
  assign n15237 = n15236 ^ n14678;
  assign n15238 = n15237 ^ n15235;
  assign n15243 = n15242 ^ n15238;
  assign n16986 = n16985 ^ n15243;
  assign n15401 = n14676 ^ n14656;
  assign n15400 = n15241 ^ n14664;
  assign n15402 = n15401 ^ n15400;
  assign n15157 = n15156 ^ n15152;
  assign n15150 = n15059 & ~n15129;
  assign n15151 = n15150 ^ n15149;
  assign n15158 = n15157 ^ n15151;
  assign n15148 = n15147 ^ n15130;
  assign n15159 = n15158 ^ n15148;
  assign n16983 = n15402 ^ n15159;
  assign n15393 = ~n14946 & n15014;
  assign n15394 = n15393 ^ n15171;
  assign n15395 = n15394 ^ n15353;
  assign n15039 = n15038 ^ n15034;
  assign n15392 = n15166 ^ n15039;
  assign n15396 = n15395 ^ n15392;
  assign n15260 = n14850 & ~n14873;
  assign n15261 = n15260 ^ n14899;
  assign n15262 = n15261 ^ n15259;
  assign n14915 = n14914 ^ n14895;
  assign n15257 = n14915 ^ n14892;
  assign n15263 = n15262 ^ n15257;
  assign n16982 = n15396 ^ n15263;
  assign n16984 = n16983 ^ n16982;
  assign n16987 = n16986 ^ n16984;
  assign n16988 = n16987 ^ n16981;
  assign n15266 = n14908 ^ n14905;
  assign n15267 = n15266 ^ n15187;
  assign n15265 = n14899 ^ n14889;
  assign n15268 = n15267 ^ n15265;
  assign n15229 = n15228 ^ n15032;
  assign n15230 = n15229 ^ n15227;
  assign n15225 = n15171 ^ n15028;
  assign n15231 = n15230 ^ n15225;
  assign n16973 = n15268 ^ n15231;
  assign n15388 = ~n15109 & n15134;
  assign n15389 = n15388 ^ n15182;
  assign n15390 = n15389 ^ n15346;
  assign n15387 = n15175 ^ n15157;
  assign n15391 = n15390 ^ n15387;
  assign n16971 = n15391 ^ n15184;
  assign n15244 = n15243 ^ n14680;
  assign n16972 = n16971 ^ n15244;
  assign n16974 = n16973 ^ n16972;
  assign n16969 = n16968 ^ n15275;
  assign n16966 = n16965 ^ n15402;
  assign n15309 = n15308 ^ n15151;
  assign n15307 = n15175 ^ n15154;
  assign n15310 = n15309 ^ n15307;
  assign n16962 = n15310 ^ n15184;
  assign n16963 = n16962 ^ n14681;
  assign n15040 = n15039 ^ n15033;
  assign n15030 = n15029 ^ n15028;
  assign n15041 = n15040 ^ n15030;
  assign n14917 = n14898 ^ n14889;
  assign n14916 = n14915 ^ n14906;
  assign n14918 = n14917 ^ n14916;
  assign n16961 = n15041 ^ n14918;
  assign n16964 = n16963 ^ n16961;
  assign n16967 = n16966 ^ n16964;
  assign n16970 = n16969 ^ n16967;
  assign n16975 = n16974 ^ n16970;
  assign n16989 = n16988 ^ n16975;
  assign n17055 = n17022 ^ n16989;
  assign n17060 = n17056 ^ n17055;
  assign n17057 = ~n17055 & ~n17056;
  assign n17005 = n16995 ^ n16967;
  assign n17040 = n16989 & ~n17005;
  assign n17058 = n17057 ^ n17040;
  assign n17009 = n16995 ^ n16987;
  assign n17004 = n17003 ^ n16975;
  assign n17047 = n17016 ^ n17004;
  assign n17050 = n17009 & ~n17047;
  assign n17028 = n17015 ^ n16987;
  assign n17030 = n17028 ^ n16975;
  assign n17031 = n17003 & n17030;
  assign n17051 = n17050 ^ n17031;
  assign n17059 = n17058 ^ n17051;
  assign n17061 = n17060 ^ n17059;
  assign n17039 = n16967 & ~n17022;
  assign n17041 = n17040 ^ n17039;
  assign n17037 = n17005 ^ n16989;
  assign n17006 = n17002 ^ n16987;
  assign n17032 = n17003 ^ n16988;
  assign n17033 = n17006 & ~n17032;
  assign n17034 = n17033 ^ n17031;
  assign n17038 = n17037 ^ n17034;
  assign n17042 = n17041 ^ n17038;
  assign n17070 = n17061 ^ n17042;
  assign n17048 = n17047 ^ n17009;
  assign n17045 = ~n17021 & ~n17044;
  assign n17007 = n17006 ^ n17005;
  assign n17008 = ~n17004 & ~n17007;
  assign n17046 = n17045 ^ n17008;
  assign n17049 = n17048 ^ n17046;
  assign n17052 = n17051 ^ n17049;
  assign n17029 = n17028 ^ n17004;
  assign n17035 = n17034 ^ n17029;
  assign n17023 = n17022 ^ n16967;
  assign n17024 = n17023 ^ n17009;
  assign n17025 = n17021 ^ n17004;
  assign n17026 = n17024 & n17025;
  assign n17027 = n17026 ^ n17008;
  assign n17036 = n17035 ^ n17027;
  assign n17043 = n17036 & ~n17042;
  assign n17071 = n17052 ^ n17043;
  assign n17072 = ~n17070 & ~n17071;
  assign n17073 = n17072 ^ n17061;
  assign n17536 = ~n17021 & n17073;
  assign n17053 = n17052 ^ n17036;
  assign n17065 = n17061 ^ n17043;
  assign n17066 = ~n17053 & n17065;
  assign n17067 = n17066 ^ n17052;
  assign n17478 = ~n17055 & ~n17067;
  assign n17664 = n17536 ^ n17478;
  assign n17078 = n17070 ^ n17043;
  assign n17076 = ~n17042 & ~n17052;
  assign n17077 = ~n17061 & n17076;
  assign n17079 = n17078 ^ n17077;
  assign n17558 = n17025 & ~n17079;
  assign n17085 = n17079 ^ n17073;
  assign n17086 = ~n17007 & ~n17085;
  assign n17559 = n17558 ^ n17086;
  assign n17665 = n17664 ^ n17559;
  assign n17062 = n17036 & n17052;
  assign n17063 = n17061 & n17062;
  assign n17054 = n17053 ^ n17043;
  assign n17064 = n17063 ^ n17054;
  assign n17092 = ~n17022 & ~n17064;
  assign n17091 = n17024 & ~n17079;
  assign n17093 = n17092 ^ n17091;
  assign n17080 = n17079 ^ n17064;
  assign n17074 = n17073 ^ n17067;
  assign n17081 = n17080 ^ n17074;
  assign n17082 = n17006 & ~n17081;
  assign n17075 = n17003 & ~n17074;
  assign n17083 = n17082 ^ n17075;
  assign n17663 = n17093 ^ n17083;
  assign n17666 = n17665 ^ n17663;
  assign n15981 = n13012 ^ n12934;
  assign n15982 = n15981 ^ n12857;
  assign n15983 = n15982 ^ n12884;
  assign n15984 = n15983 ^ n13178;
  assign n15966 = n13620 ^ n13036;
  assign n15967 = n15966 ^ n12972;
  assign n15968 = n15967 ^ n13200;
  assign n16014 = n15984 ^ n15968;
  assign n15989 = n14811 ^ n12611;
  assign n15988 = n13651 ^ n12997;
  assign n15990 = n15989 ^ n15988;
  assign n15986 = n13183 ^ n12742;
  assign n15978 = n13181 ^ n12900;
  assign n15976 = n14799 ^ n12889;
  assign n15975 = n13646 ^ n12933;
  assign n15977 = n15976 ^ n15975;
  assign n15979 = n15978 ^ n15977;
  assign n15987 = n15986 ^ n15979;
  assign n15991 = n15990 ^ n15987;
  assign n16015 = n16014 ^ n15991;
  assign n15971 = n12968 ^ n12937;
  assign n15972 = n15971 ^ n13646;
  assign n15970 = n13198 ^ n12945;
  assign n15973 = n15972 ^ n15970;
  assign n15963 = n13636 ^ n13041;
  assign n15964 = n15963 ^ n12492;
  assign n15965 = n15964 ^ n13176;
  assign n15969 = n15968 ^ n15965;
  assign n15974 = n15973 ^ n15969;
  assign n16043 = n15974 & ~n15979;
  assign n15985 = n15984 ^ n15965;
  assign n15992 = n15991 ^ n15985;
  assign n16001 = n13062 ^ n12963;
  assign n16000 = n13059 ^ n12620;
  assign n16002 = n16001 ^ n16000;
  assign n15999 = n13187 ^ n12751;
  assign n16003 = n16002 ^ n15999;
  assign n16007 = n16003 ^ n15979;
  assign n16008 = n15992 & n16007;
  assign n16044 = n16043 ^ n16008;
  assign n16041 = n16007 ^ n15992;
  assign n15994 = n13627 ^ n13613;
  assign n15995 = n15994 ^ n14790;
  assign n15996 = n15995 ^ n12625;
  assign n15997 = n15996 ^ n13189;
  assign n16021 = n15997 ^ n15984;
  assign n16004 = n16003 ^ n15997;
  assign n16028 = n16004 ^ n15985;
  assign n16029 = n16021 & n16028;
  assign n16016 = n16004 & n16015;
  assign n16030 = n16029 ^ n16016;
  assign n16042 = n16041 ^ n16030;
  assign n16045 = n16044 ^ n16042;
  assign n15998 = n15997 ^ n15974;
  assign n16005 = n16004 ^ n15998;
  assign n15993 = n15992 ^ n15974;
  assign n16019 = n16005 ^ n15993;
  assign n16010 = n16003 ^ n15984;
  assign n16011 = n16004 ^ n15991;
  assign n16012 = n16011 ^ n15969;
  assign n16013 = n16010 & n16012;
  assign n16017 = n16016 ^ n16013;
  assign n16006 = n15993 & n16005;
  assign n16009 = n16008 ^ n16006;
  assign n16018 = n16017 ^ n16009;
  assign n16020 = n16019 ^ n16018;
  assign n16056 = n16045 ^ n16020;
  assign n16031 = n16014 ^ n16011;
  assign n16032 = n16031 ^ n16030;
  assign n16024 = n16011 ^ n15973;
  assign n15980 = n15979 ^ n15974;
  assign n16025 = n16010 ^ n15980;
  assign n16026 = n16024 & n16025;
  assign n16022 = n16021 ^ n16007;
  assign n16023 = n16011 & n16022;
  assign n16027 = n16026 ^ n16023;
  assign n16033 = n16032 ^ n16027;
  assign n16046 = n16033 & n16045;
  assign n16036 = n16012 ^ n16010;
  assign n16034 = n15973 & n15998;
  assign n16035 = n16034 ^ n16023;
  assign n16037 = n16036 ^ n16035;
  assign n16038 = n16037 ^ n16017;
  assign n16057 = n16046 ^ n16038;
  assign n16058 = n16056 & n16057;
  assign n16059 = n16058 ^ n16020;
  assign n16047 = n16038 ^ n16033;
  assign n16051 = n16046 ^ n16020;
  assign n16052 = n16047 & n16051;
  assign n16053 = n16052 ^ n16038;
  assign n16060 = n16059 ^ n16053;
  assign n16200 = n16015 & n16060;
  assign n16063 = n16056 ^ n16046;
  assign n16061 = n16038 & n16045;
  assign n16062 = ~n16020 & n16061;
  assign n16064 = n16063 ^ n16062;
  assign n16048 = n16047 ^ n16046;
  assign n16039 = n16033 & ~n16038;
  assign n16040 = n16020 & n16039;
  assign n16049 = n16048 ^ n16040;
  assign n16065 = n16064 ^ n16049;
  assign n16066 = n16065 ^ n16060;
  assign n16067 = n16028 & n16066;
  assign n16274 = n16200 ^ n16067;
  assign n16136 = n16025 & n16064;
  assign n16077 = n15974 & n16049;
  assign n16137 = n16136 ^ n16077;
  assign n16309 = n16274 ^ n16137;
  assign n16068 = n16053 ^ n16049;
  assign n16154 = n15992 & n16068;
  assign n16075 = n16004 & n16060;
  assign n16074 = n16021 & n16066;
  assign n16076 = n16075 ^ n16074;
  assign n16155 = n16154 ^ n16076;
  assign n16141 = n16064 ^ n16059;
  assign n16142 = n16022 & n16141;
  assign n16308 = n16155 ^ n16142;
  assign n16310 = n16309 ^ n16308;
  assign n15879 = n14577 ^ n13912;
  assign n15878 = n14695 ^ n11436;
  assign n15880 = n15879 ^ n15878;
  assign n15875 = n14684 ^ n11932;
  assign n15873 = n14559 ^ n13906;
  assign n15874 = n15873 ^ n13898;
  assign n15876 = n15875 ^ n15874;
  assign n15877 = n15876 ^ n14574;
  assign n15881 = n15880 ^ n15877;
  assign n15870 = n14553 ^ n12138;
  assign n15869 = n14682 ^ n11923;
  assign n15871 = n15870 ^ n15869;
  assign n15865 = n14687 ^ n12074;
  assign n15863 = n14548 ^ n13885;
  assign n15864 = n15863 ^ n13871;
  assign n15866 = n15865 ^ n15864;
  assign n15872 = n15871 ^ n15866;
  assign n15882 = n15881 ^ n15872;
  assign n15884 = n14565 ^ n11772;
  assign n15883 = n14690 ^ n11967;
  assign n15885 = n15884 ^ n15883;
  assign n15856 = n13875 ^ n12102;
  assign n15855 = n14702 ^ n12043;
  assign n15857 = n15856 ^ n15855;
  assign n15907 = n15885 ^ n15857;
  assign n15914 = n15907 ^ n15881;
  assign n15859 = n14587 ^ n12066;
  assign n15858 = n14692 ^ n12121;
  assign n15860 = n15859 ^ n15858;
  assign n15861 = n15860 ^ n15857;
  assign n15853 = n14597 ^ n12164;
  assign n15852 = n14711 ^ n11917;
  assign n15854 = n15853 ^ n15852;
  assign n15862 = n15861 ^ n15854;
  assign n15924 = n15914 ^ n15862;
  assign n15867 = n15866 ^ n15862;
  assign n15923 = n15872 ^ n15867;
  assign n15928 = n15924 ^ n15923;
  assign n15925 = ~n15923 & ~n15924;
  assign n15887 = n15876 ^ n15871;
  assign n15917 = ~n15887 & n15914;
  assign n15926 = n15925 ^ n15917;
  assign n15896 = n15885 ^ n15860;
  assign n15897 = n15896 ^ n15881;
  assign n15898 = n15872 & n15897;
  assign n15891 = n15882 ^ n15861;
  assign n15892 = n15885 ^ n15871;
  assign n15895 = n15891 & ~n15892;
  assign n15899 = n15898 ^ n15895;
  assign n15927 = n15926 ^ n15899;
  assign n15929 = n15928 ^ n15927;
  assign n15918 = ~n15862 & n15876;
  assign n15919 = n15918 ^ n15917;
  assign n15915 = n15914 ^ n15887;
  assign n15886 = n15885 ^ n15866;
  assign n15908 = n15907 ^ n15872;
  assign n15909 = ~n15886 & n15908;
  assign n15910 = n15909 ^ n15898;
  assign n15916 = n15915 ^ n15910;
  assign n15920 = n15919 ^ n15916;
  assign n15937 = n15929 ^ n15920;
  assign n15906 = n15896 ^ n15882;
  assign n15911 = n15910 ^ n15906;
  assign n15901 = n15876 ^ n15862;
  assign n15902 = n15901 ^ n15892;
  assign n15903 = n15882 ^ n15854;
  assign n15904 = ~n15902 & ~n15903;
  assign n15888 = n15887 ^ n15886;
  assign n15889 = n15882 & n15888;
  assign n15905 = n15904 ^ n15889;
  assign n15912 = n15911 ^ n15905;
  assign n15921 = n15912 & ~n15920;
  assign n15945 = n15937 ^ n15921;
  assign n15893 = n15892 ^ n15891;
  assign n15868 = ~n15854 & ~n15867;
  assign n15890 = n15889 ^ n15868;
  assign n15894 = n15893 ^ n15890;
  assign n15900 = n15899 ^ n15894;
  assign n15943 = ~n15900 & ~n15920;
  assign n15944 = ~n15929 & n15943;
  assign n15946 = n15945 ^ n15944;
  assign n15938 = n15921 ^ n15900;
  assign n15939 = ~n15937 & ~n15938;
  assign n15940 = n15939 ^ n15929;
  assign n16130 = n15946 ^ n15940;
  assign n16170 = n15882 & ~n16130;
  assign n16128 = ~n15854 & n15940;
  assign n16171 = n16170 ^ n16128;
  assign n15913 = n15912 ^ n15900;
  assign n15934 = n15929 ^ n15921;
  assign n15935 = ~n15913 & n15934;
  assign n15936 = n15935 ^ n15900;
  assign n15959 = ~n15924 & ~n15936;
  assign n15930 = n15900 & n15912;
  assign n15931 = n15929 & n15930;
  assign n15922 = n15921 ^ n15913;
  assign n15932 = n15931 ^ n15922;
  assign n15958 = n15901 & ~n15932;
  assign n15960 = n15959 ^ n15958;
  assign n16264 = n16171 ^ n15960;
  assign n15952 = n15936 ^ n15932;
  assign n16165 = n15914 & n15952;
  assign n15947 = n15946 ^ n15932;
  assign n15941 = n15940 ^ n15936;
  assign n15948 = n15947 ^ n15941;
  assign n15949 = ~n15886 & ~n15948;
  assign n15942 = n15872 & ~n15941;
  assign n15950 = n15949 ^ n15942;
  assign n16166 = n16165 ^ n15950;
  assign n15953 = ~n15887 & n15952;
  assign n16263 = n16166 ^ n15953;
  assign n16265 = n16264 ^ n16263;
  assign n16886 = n16310 ^ n16265;
  assign n15760 = n12154 ^ n11132;
  assign n15758 = n11191 ^ n11186;
  assign n15759 = n15758 ^ n11199;
  assign n15761 = n15760 ^ n15759;
  assign n15749 = n12114 ^ n11106;
  assign n15747 = n14925 ^ n13748;
  assign n15748 = n15747 ^ n11041;
  assign n15750 = n15749 ^ n15748;
  assign n15762 = n15761 ^ n15750;
  assign n15739 = n12050 ^ n11061;
  assign n15738 = n14924 ^ n11183;
  assign n15740 = n15739 ^ n15738;
  assign n15736 = n12006 ^ n10918;
  assign n15734 = n11227 ^ n10757;
  assign n15733 = n11166 ^ n11148;
  assign n15735 = n15734 ^ n15733;
  assign n15737 = n15736 ^ n15735;
  assign n15741 = n15740 ^ n15737;
  assign n15785 = n15762 ^ n15741;
  assign n15752 = n12126 ^ n11191;
  assign n15751 = n14940 ^ n11122;
  assign n15753 = n15752 ^ n15751;
  assign n15754 = n15753 ^ n15740;
  assign n15745 = n12092 ^ n11207;
  assign n15743 = n11157 ^ n11153;
  assign n15744 = n15743 ^ n14920;
  assign n15746 = n15745 ^ n15744;
  assign n15755 = n15754 ^ n15746;
  assign n15730 = n11093 ^ n11083;
  assign n15729 = n14955 ^ n13776;
  assign n15731 = n15730 ^ n15729;
  assign n15726 = n11944 ^ n11166;
  assign n15724 = n14931 ^ n13770;
  assign n15725 = n15724 ^ n10610;
  assign n15727 = n15726 ^ n15725;
  assign n15723 = n11521 ^ n11234;
  assign n15728 = n15727 ^ n15723;
  assign n15732 = n15731 ^ n15728;
  assign n15742 = n15741 ^ n15732;
  assign n15799 = n15755 ^ n15742;
  assign n15756 = n15755 ^ n15750;
  assign n15798 = n15762 ^ n15756;
  assign n15803 = n15799 ^ n15798;
  assign n15800 = ~n15798 & ~n15799;
  assign n15765 = n15761 ^ n15727;
  assign n15793 = n15742 & ~n15765;
  assign n15801 = n15800 ^ n15793;
  assign n15774 = n15753 ^ n15737;
  assign n15775 = n15774 ^ n15732;
  assign n15776 = n15762 & n15775;
  assign n15763 = n15762 ^ n15732;
  assign n15769 = n15763 ^ n15754;
  assign n15770 = n15761 ^ n15737;
  assign n15773 = ~n15769 & n15770;
  assign n15777 = n15776 ^ n15773;
  assign n15802 = n15801 ^ n15777;
  assign n15804 = n15803 ^ n15802;
  assign n15794 = n15727 & ~n15755;
  assign n15795 = n15794 ^ n15793;
  assign n15791 = n15765 ^ n15742;
  assign n15764 = n15750 ^ n15737;
  assign n15786 = n15764 & ~n15785;
  assign n15787 = n15786 ^ n15776;
  assign n15792 = n15791 ^ n15787;
  assign n15796 = n15795 ^ n15792;
  assign n15814 = n15804 ^ n15796;
  assign n15784 = n15774 ^ n15763;
  assign n15788 = n15787 ^ n15784;
  assign n15779 = n15755 ^ n15727;
  assign n15780 = n15779 ^ n15770;
  assign n15781 = n15763 ^ n15746;
  assign n15782 = n15780 & n15781;
  assign n15766 = n15765 ^ n15764;
  assign n15767 = ~n15763 & ~n15766;
  assign n15783 = n15782 ^ n15767;
  assign n15789 = n15788 ^ n15783;
  assign n15797 = n15789 & ~n15796;
  assign n15822 = n15814 ^ n15797;
  assign n15771 = n15770 ^ n15769;
  assign n15757 = ~n15746 & ~n15756;
  assign n15768 = n15767 ^ n15757;
  assign n15772 = n15771 ^ n15768;
  assign n15778 = n15777 ^ n15772;
  assign n15820 = ~n15778 & ~n15796;
  assign n15821 = ~n15804 & n15820;
  assign n15823 = n15822 ^ n15821;
  assign n15809 = n15778 & n15789;
  assign n15810 = n15804 & n15809;
  assign n15790 = n15789 ^ n15778;
  assign n15808 = n15797 ^ n15790;
  assign n15811 = n15810 ^ n15808;
  assign n15824 = n15823 ^ n15811;
  assign n15815 = n15797 ^ n15778;
  assign n15816 = ~n15814 & ~n15815;
  assign n15817 = n15816 ^ n15804;
  assign n15805 = n15804 ^ n15797;
  assign n15806 = ~n15790 & n15805;
  assign n15807 = n15806 ^ n15778;
  assign n15818 = n15817 ^ n15807;
  assign n15825 = n15824 ^ n15818;
  assign n15846 = ~n15785 & ~n15825;
  assign n15845 = n15775 & ~n15818;
  assign n15847 = n15846 ^ n15845;
  assign n15843 = n15780 & ~n15823;
  assign n15842 = ~n15755 & ~n15811;
  assign n15844 = n15843 ^ n15842;
  assign n15848 = n15847 ^ n15844;
  assign n15835 = n15823 ^ n15817;
  assign n15840 = ~n15766 & ~n15835;
  assign n15826 = n15764 & ~n15825;
  assign n15819 = n15762 & ~n15818;
  assign n15827 = n15826 ^ n15819;
  assign n15812 = n15811 ^ n15807;
  assign n15813 = n15742 & n15812;
  assign n15828 = n15827 ^ n15813;
  assign n15841 = n15840 ^ n15828;
  assign n15849 = n15848 ^ n15841;
  assign n15836 = ~n15763 & ~n15835;
  assign n15834 = ~n15746 & n15817;
  assign n15837 = n15836 ^ n15834;
  assign n15832 = ~n15799 & ~n15807;
  assign n15831 = n15779 & ~n15811;
  assign n15833 = n15832 ^ n15831;
  assign n15838 = n15837 ^ n15833;
  assign n15829 = ~n15765 & n15812;
  assign n15830 = n15829 ^ n15828;
  assign n15839 = n15838 ^ n15830;
  assign n15850 = n15849 ^ n15839;
  assign n16887 = n16886 ^ n15850;
  assign n15532 = n15073 ^ n13019;
  assign n15531 = n14017 ^ n10163;
  assign n15533 = n15532 ^ n15531;
  assign n15528 = n15042 ^ n12954;
  assign n15526 = n14010 ^ n10110;
  assign n15527 = n15526 ^ n10275;
  assign n15529 = n15528 ^ n15527;
  assign n15530 = n15529 ^ n14009;
  assign n15534 = n15533 ^ n15530;
  assign n15523 = n12985 ^ n10253;
  assign n15521 = n10244 ^ n10057;
  assign n15522 = n15521 ^ n14002;
  assign n15524 = n15523 ^ n15522;
  assign n15517 = n15077 ^ n12839;
  assign n15515 = n13996 ^ n7151;
  assign n15516 = n15515 ^ n10209;
  assign n15518 = n15517 ^ n15516;
  assign n15525 = n15524 ^ n15518;
  assign n15535 = n15534 ^ n15525;
  assign n15538 = n12916 ^ n10144;
  assign n15536 = n10271 ^ n10110;
  assign n15537 = n15536 ^ n14037;
  assign n15539 = n15538 ^ n15537;
  assign n15507 = n13052 ^ n9038;
  assign n15505 = n10216 ^ n7151;
  assign n15506 = n15505 ^ n10250;
  assign n15508 = n15507 ^ n15506;
  assign n15561 = n15539 ^ n15508;
  assign n15568 = n15561 ^ n15534;
  assign n15511 = n13075 ^ n10223;
  assign n15509 = n10244 ^ n10216;
  assign n15510 = n15509 ^ n14024;
  assign n15512 = n15511 ^ n15510;
  assign n15513 = n15512 ^ n15508;
  assign n15503 = n13099 ^ n10074;
  assign n15502 = n14049 ^ n14010;
  assign n15504 = n15503 ^ n15502;
  assign n15514 = n15513 ^ n15504;
  assign n15578 = n15568 ^ n15514;
  assign n15519 = n15518 ^ n15514;
  assign n15577 = n15525 ^ n15519;
  assign n15582 = n15578 ^ n15577;
  assign n15579 = ~n15577 & ~n15578;
  assign n15541 = n15529 ^ n15524;
  assign n15571 = ~n15541 & n15568;
  assign n15580 = n15579 ^ n15571;
  assign n15550 = n15539 ^ n15512;
  assign n15551 = n15550 ^ n15534;
  assign n15552 = n15525 & n15551;
  assign n15545 = n15535 ^ n15513;
  assign n15546 = n15539 ^ n15524;
  assign n15549 = ~n15545 & n15546;
  assign n15553 = n15552 ^ n15549;
  assign n15581 = n15580 ^ n15553;
  assign n15583 = n15582 ^ n15581;
  assign n15572 = ~n15514 & n15529;
  assign n15573 = n15572 ^ n15571;
  assign n15569 = n15568 ^ n15541;
  assign n15540 = n15539 ^ n15518;
  assign n15562 = n15561 ^ n15525;
  assign n15563 = n15540 & ~n15562;
  assign n15564 = n15563 ^ n15552;
  assign n15570 = n15569 ^ n15564;
  assign n15574 = n15573 ^ n15570;
  assign n15590 = n15583 ^ n15574;
  assign n15560 = n15550 ^ n15535;
  assign n15565 = n15564 ^ n15560;
  assign n15555 = n15529 ^ n15514;
  assign n15556 = n15555 ^ n15546;
  assign n15557 = n15535 ^ n15504;
  assign n15558 = n15556 & n15557;
  assign n15542 = n15541 ^ n15540;
  assign n15543 = ~n15535 & ~n15542;
  assign n15559 = n15558 ^ n15543;
  assign n15566 = n15565 ^ n15559;
  assign n15575 = n15566 & ~n15574;
  assign n15547 = n15546 ^ n15545;
  assign n15520 = ~n15504 & ~n15519;
  assign n15544 = n15543 ^ n15520;
  assign n15548 = n15547 ^ n15544;
  assign n15554 = n15553 ^ n15548;
  assign n15598 = n15575 ^ n15554;
  assign n15599 = ~n15590 & ~n15598;
  assign n15600 = n15599 ^ n15583;
  assign n15591 = n15590 ^ n15575;
  assign n15588 = ~n15554 & ~n15574;
  assign n15589 = ~n15583 & n15588;
  assign n15592 = n15591 ^ n15589;
  assign n15611 = n15600 ^ n15592;
  assign n15718 = ~n15535 & ~n15611;
  assign n15609 = ~n15504 & n15600;
  assign n15719 = n15718 ^ n15609;
  assign n15584 = n15554 & n15566;
  assign n15585 = n15583 & n15584;
  assign n15567 = n15566 ^ n15554;
  assign n15576 = n15575 ^ n15567;
  assign n15586 = n15585 ^ n15576;
  assign n15716 = n15555 & ~n15586;
  assign n15595 = n15583 ^ n15575;
  assign n15596 = ~n15567 & n15595;
  assign n15597 = n15596 ^ n15554;
  assign n15608 = ~n15578 & ~n15597;
  assign n15717 = n15716 ^ n15608;
  assign n15720 = n15719 ^ n15717;
  assign n15705 = n15597 ^ n15586;
  assign n15714 = ~n15541 & n15705;
  assign n15706 = n15568 & n15705;
  assign n15603 = n15592 ^ n15586;
  assign n15601 = n15600 ^ n15597;
  assign n15604 = n15603 ^ n15601;
  assign n15605 = n15540 & ~n15604;
  assign n15602 = n15525 & ~n15601;
  assign n15606 = n15605 ^ n15602;
  assign n15707 = n15706 ^ n15606;
  assign n15715 = n15714 ^ n15707;
  assign n15721 = n15720 ^ n15715;
  assign n16885 = n16884 ^ n15721;
  assign n16888 = n16887 ^ n16885;
  assign n16083 = ~n15545 & n15603;
  assign n16084 = n16083 ^ n15714;
  assign n15710 = ~n15562 & ~n15604;
  assign n16085 = n16084 ^ n15710;
  assign n16086 = n16085 ^ n15717;
  assign n15587 = ~n15514 & ~n15586;
  assign n16082 = n15606 ^ n15587;
  assign n16087 = n16086 ^ n16082;
  assign n16834 = n16833 ^ n16087;
  assign n16159 = n16011 & n16141;
  assign n16139 = n15973 & n16059;
  assign n16160 = n16159 ^ n16139;
  assign n16054 = n15993 & n16053;
  assign n16050 = n15980 & n16049;
  assign n16055 = n16054 ^ n16050;
  assign n16260 = n16160 ^ n16055;
  assign n16069 = n16007 & n16068;
  assign n16259 = n16155 ^ n16069;
  assign n16261 = n16260 ^ n16259;
  assign n16830 = n16310 ^ n16261;
  assign n15956 = n15908 & ~n15948;
  assign n15954 = n15891 & n15947;
  assign n15955 = n15954 ^ n15953;
  assign n15957 = n15956 ^ n15955;
  assign n15961 = n15960 ^ n15957;
  assign n15933 = ~n15862 & ~n15932;
  assign n15951 = n15950 ^ n15933;
  assign n15962 = n15961 ^ n15951;
  assign n16831 = n16830 ^ n15962;
  assign n16113 = ~n15769 & n15824;
  assign n16114 = n16113 ^ n15829;
  assign n16115 = n16114 ^ n15846;
  assign n16151 = n16115 ^ n15833;
  assign n16150 = n15842 ^ n15827;
  assign n16152 = n16151 ^ n16150;
  assign n16829 = n16152 ^ n15850;
  assign n16832 = n16831 ^ n16829;
  assign n16835 = n16834 ^ n16832;
  assign n16285 = n15770 & n15824;
  assign n16286 = n16285 ^ n16114;
  assign n16283 = n15845 ^ n15819;
  assign n16119 = ~n15798 & ~n15807;
  assign n16120 = n16119 ^ n15837;
  assign n16284 = n16283 ^ n16120;
  assign n16287 = n16286 ^ n16284;
  assign n16203 = n16010 & n16065;
  assign n16070 = n16012 & n16065;
  assign n16071 = n16070 ^ n16069;
  assign n16204 = n16203 ^ n16071;
  assign n16201 = n16200 ^ n16075;
  assign n16161 = n16005 & n16053;
  assign n16162 = n16161 ^ n16160;
  assign n16202 = n16201 ^ n16162;
  assign n16205 = n16204 ^ n16202;
  assign n16872 = n16287 ^ n16205;
  assign n16313 = n15843 ^ n15827;
  assign n16210 = n15781 & ~n15823;
  assign n16211 = n16210 ^ n15840;
  assign n16212 = n16211 ^ n15836;
  assign n16312 = n16212 ^ n15847;
  assign n16314 = n16313 ^ n16312;
  assign n15593 = n15556 & ~n15592;
  assign n16291 = n15606 ^ n15593;
  assign n15613 = n15557 & ~n15592;
  assign n15612 = ~n15542 & ~n15611;
  assign n15614 = n15613 ^ n15612;
  assign n16207 = n15718 ^ n15614;
  assign n15709 = n15551 & ~n15601;
  assign n15711 = n15710 ^ n15709;
  assign n16290 = n16207 ^ n15711;
  assign n16292 = n16291 ^ n16290;
  assign n16315 = n16314 ^ n16292;
  assign n16873 = n16872 ^ n16315;
  assign n16125 = ~n15902 & ~n15946;
  assign n16280 = n16125 ^ n15950;
  assign n16194 = n15897 & ~n15941;
  assign n16278 = n16194 ^ n15956;
  assign n16132 = ~n15903 & ~n15946;
  assign n16131 = n15888 & ~n16130;
  assign n16133 = n16132 ^ n16131;
  assign n16242 = n16170 ^ n16133;
  assign n16279 = n16278 ^ n16242;
  assign n16281 = n16280 ^ n16279;
  assign n16874 = n16873 ^ n16281;
  assign n16876 = n16875 ^ n16874;
  assign n16219 = n15546 & n15603;
  assign n16220 = n16219 ^ n16084;
  assign n16217 = n15709 ^ n15602;
  assign n16108 = ~n15577 & ~n15597;
  assign n16109 = n16108 ^ n15719;
  assign n16218 = n16217 ^ n16109;
  assign n16221 = n16220 ^ n16218;
  assign n16288 = n16287 ^ n16221;
  assign n16197 = ~n15892 & n15947;
  assign n16198 = n16197 ^ n15955;
  assign n16195 = n16194 ^ n15942;
  assign n16172 = ~n15923 & ~n15936;
  assign n16173 = n16172 ^ n16171;
  assign n16196 = n16195 ^ n16173;
  assign n16199 = n16198 ^ n16196;
  assign n16851 = n16288 ^ n16199;
  assign n16143 = n16024 & n16064;
  assign n16144 = n16143 ^ n16142;
  assign n16245 = n16159 ^ n16144;
  assign n16246 = n16245 ^ n16137;
  assign n16247 = n16246 ^ n16155;
  assign n16213 = n16212 ^ n15844;
  assign n16214 = n16213 ^ n15828;
  assign n16850 = n16247 ^ n16214;
  assign n16852 = n16851 ^ n16850;
  assign n16854 = n16853 ^ n16852;
  assign n16877 = n16876 ^ n16854;
  assign n16889 = n16888 ^ n16877;
  assign n16922 = ~n16835 & n16889;
  assign n16078 = n16077 ^ n16076;
  assign n16072 = n16071 ^ n16067;
  assign n16073 = n16072 ^ n16055;
  assign n16079 = n16078 ^ n16073;
  assign n16844 = n16152 ^ n16079;
  assign n16106 = ~n15519 & n15600;
  assign n15594 = n15593 ^ n15587;
  assign n16107 = n16106 ^ n15594;
  assign n16110 = n16109 ^ n16107;
  assign n16105 = n16085 ^ n15707;
  assign n16111 = n16110 ^ n16105;
  assign n16845 = n16844 ^ n16111;
  assign n16117 = ~n15756 & n15817;
  assign n16118 = n16117 ^ n15844;
  assign n16121 = n16120 ^ n16118;
  assign n16116 = n16115 ^ n15828;
  assign n16122 = n16121 ^ n16116;
  assign n16846 = n16845 ^ n16122;
  assign n16168 = ~n15867 & n15940;
  assign n16126 = n16125 ^ n15933;
  assign n16169 = n16168 ^ n16126;
  assign n16174 = n16173 ^ n16169;
  assign n16167 = n16166 ^ n15957;
  assign n16175 = n16174 ^ n16167;
  assign n16847 = n16846 ^ n16175;
  assign n16849 = n16848 ^ n16847;
  assign n16855 = n16854 ^ n16849;
  assign n16157 = n15998 & n16059;
  assign n16158 = n16157 ^ n16137;
  assign n16163 = n16162 ^ n16158;
  assign n16156 = n16155 ^ n16072;
  assign n16164 = n16163 ^ n16156;
  assign n16840 = n16310 ^ n16164;
  assign n16129 = n16128 ^ n15959;
  assign n16134 = n16133 ^ n16129;
  assign n16127 = n16126 ^ n15950;
  assign n16135 = n16134 ^ n16127;
  assign n16841 = n16840 ^ n16135;
  assign n16237 = n15834 ^ n15832;
  assign n16238 = n16237 ^ n16211;
  assign n16236 = n15844 ^ n15827;
  assign n16239 = n16238 ^ n16236;
  assign n16123 = n16122 ^ n15849;
  assign n16839 = n16239 ^ n16123;
  assign n16842 = n16841 ^ n16839;
  assign n15610 = n15609 ^ n15608;
  assign n15615 = n15614 ^ n15610;
  assign n15607 = n15606 ^ n15594;
  assign n15616 = n15615 ^ n15607;
  assign n16837 = n16836 ^ n15616;
  assign n16838 = n16837 ^ n16835;
  assign n16843 = n16842 ^ n16838;
  assign n16856 = n16855 ^ n16843;
  assign n15712 = n15711 ^ n15594;
  assign n15708 = n15707 ^ n15612;
  assign n15713 = n15712 ^ n15708;
  assign n16861 = n16860 ^ n15713;
  assign n16306 = n16278 ^ n16126;
  assign n16305 = n16166 ^ n16131;
  assign n16307 = n16306 ^ n16305;
  assign n16276 = n16136 ^ n16076;
  assign n16275 = n16274 ^ n16245;
  assign n16277 = n16276 ^ n16275;
  assign n16858 = n16307 ^ n16277;
  assign n16857 = n16314 ^ n15849;
  assign n16859 = n16858 ^ n16857;
  assign n16862 = n16861 ^ n16859;
  assign n16892 = n16862 ^ n16835;
  assign n16915 = n16856 & n16892;
  assign n16923 = n16922 ^ n16915;
  assign n16920 = n16892 ^ n16856;
  assign n16240 = n16239 ^ n15849;
  assign n16208 = n16207 ^ n15594;
  assign n16209 = n16208 ^ n15707;
  assign n16215 = n16214 ^ n16209;
  assign n16865 = n16240 ^ n16215;
  assign n16140 = n16139 ^ n16054;
  assign n16145 = n16144 ^ n16140;
  assign n16138 = n16137 ^ n16076;
  assign n16146 = n16145 ^ n16138;
  assign n16864 = n16310 ^ n16146;
  assign n16866 = n16865 ^ n16864;
  assign n16243 = n16242 ^ n16126;
  assign n16244 = n16243 ^ n16166;
  assign n16867 = n16866 ^ n16244;
  assign n16869 = n16868 ^ n16867;
  assign n16893 = n16869 ^ n16849;
  assign n16870 = n16869 ^ n16862;
  assign n16906 = n16870 ^ n16855;
  assign n16907 = n16893 & n16906;
  assign n16880 = n16876 ^ n16849;
  assign n16881 = n16880 ^ n16843;
  assign n16882 = n16870 & n16881;
  assign n16908 = n16907 ^ n16882;
  assign n16921 = n16920 ^ n16908;
  assign n16924 = n16923 ^ n16921;
  assign n16890 = n16889 ^ n16869;
  assign n16913 = n16890 ^ n16870;
  assign n16912 = n16889 ^ n16856;
  assign n16918 = n16913 ^ n16912;
  assign n16914 = n16912 & n16913;
  assign n16916 = n16915 ^ n16914;
  assign n16863 = n16862 ^ n16849;
  assign n16871 = n16870 ^ n16843;
  assign n16878 = n16877 ^ n16871;
  assign n16879 = n16863 & n16878;
  assign n16883 = n16882 ^ n16879;
  assign n16917 = n16916 ^ n16883;
  assign n16919 = n16918 ^ n16917;
  assign n16937 = n16924 ^ n16919;
  assign n16905 = n16880 ^ n16871;
  assign n16909 = n16908 ^ n16905;
  assign n16900 = n16888 ^ n16871;
  assign n16901 = n16889 ^ n16835;
  assign n16902 = n16901 ^ n16863;
  assign n16903 = n16900 & n16902;
  assign n16894 = n16893 ^ n16892;
  assign n16895 = n16871 & n16894;
  assign n16904 = n16903 ^ n16895;
  assign n16910 = n16909 ^ n16904;
  assign n16925 = n16910 & n16924;
  assign n16897 = n16878 ^ n16863;
  assign n16891 = n16888 & n16890;
  assign n16896 = n16895 ^ n16891;
  assign n16898 = n16897 ^ n16896;
  assign n16899 = n16898 ^ n16883;
  assign n16941 = n16925 ^ n16899;
  assign n16942 = n16937 & n16941;
  assign n16943 = n16942 ^ n16919;
  assign n17542 = n16888 & n16943;
  assign n16911 = n16910 ^ n16899;
  assign n16926 = n16925 ^ n16919;
  assign n16927 = n16911 & n16926;
  assign n16928 = n16927 ^ n16899;
  assign n17463 = n16912 & n16928;
  assign n17660 = n17542 ^ n17463;
  assign n16938 = n16937 ^ n16925;
  assign n16935 = n16899 & n16924;
  assign n16936 = ~n16919 & n16935;
  assign n16939 = n16938 ^ n16936;
  assign n17564 = n16900 & n16939;
  assign n16950 = n16943 ^ n16939;
  assign n16951 = n16894 & n16950;
  assign n17565 = n17564 ^ n16951;
  assign n17661 = n17660 ^ n17565;
  assign n16931 = n16925 ^ n16911;
  assign n16929 = ~n16899 & n16910;
  assign n16930 = n16919 & n16929;
  assign n16932 = n16931 ^ n16930;
  assign n16957 = n16889 & n16932;
  assign n16956 = n16902 & n16939;
  assign n16958 = n16957 ^ n16956;
  assign n16944 = n16943 ^ n16928;
  assign n16947 = n16870 & n16944;
  assign n16940 = n16939 ^ n16932;
  assign n16945 = n16944 ^ n16940;
  assign n16946 = n16893 & n16945;
  assign n16948 = n16947 ^ n16946;
  assign n17659 = n16958 ^ n16948;
  assign n17662 = n17661 ^ n17659;
  assign n17667 = n17666 ^ n17662;
  assign n17507 = n17288 & n17344;
  assign n17506 = n17316 & n17340;
  assign n17508 = n17507 ^ n17506;
  assign n17511 = n17510 ^ n17508;
  assign n17505 = n17504 ^ n17502;
  assign n17512 = n17511 ^ n17505;
  assign n17518 = n17517 ^ n17512;
  assign n17531 = n17530 ^ n17518;
  assign n17483 = ~n17167 & n17217;
  assign n17485 = n17484 ^ n17483;
  assign n17496 = n17495 ^ n17485;
  assign n17493 = n17487 ^ n17231;
  assign n17497 = n17496 ^ n17493;
  assign n17498 = n17497 ^ n17236;
  assign n17491 = n17233 ^ n17225;
  assign n17490 = n17489 ^ n17485;
  assign n17492 = n17491 ^ n17490;
  assign n17499 = n17498 ^ n17492;
  assign n17477 = n17023 & ~n17064;
  assign n17479 = n17478 ^ n17477;
  assign n17068 = n17067 ^ n17064;
  assign n17474 = ~n17005 & n17068;
  assign n17473 = ~n17047 & n17080;
  assign n17475 = n17474 ^ n17473;
  assign n17089 = ~n17032 & ~n17081;
  assign n17476 = n17475 ^ n17089;
  assign n17480 = n17479 ^ n17476;
  assign n17472 = n17092 ^ n17083;
  assign n17481 = n17480 ^ n17472;
  assign n17470 = n16957 ^ n16948;
  assign n17466 = n16878 & n16940;
  assign n16933 = n16932 ^ n16928;
  assign n17465 = n16892 & n16933;
  assign n17467 = n17466 ^ n17465;
  assign n16954 = n16906 & n16945;
  assign n17468 = n17467 ^ n16954;
  assign n17462 = n16901 & n16932;
  assign n17464 = n17463 ^ n17462;
  assign n17469 = n17468 ^ n17464;
  assign n17471 = n17470 ^ n17469;
  assign n17482 = n17481 ^ n17471;
  assign n17500 = n17499 ^ n17482;
  assign n17532 = n17531 ^ n17500;
  assign n17668 = n17667 ^ n17532;
  assign n17691 = n17690 ^ n17668;
  assign n17646 = n17509 ^ n17507;
  assign n17327 = n17264 & n17326;
  assign n17333 = n17332 ^ n17327;
  assign n17647 = n17646 ^ n17333;
  assign n17645 = n17515 ^ n17353;
  assign n17648 = n17647 ^ n17645;
  assign n17649 = n17648 ^ n17517;
  assign n17654 = n17653 ^ n17649;
  assign n17642 = n17641 ^ n17236;
  assign n17207 = n17206 ^ n17205;
  assign n17614 = n17234 ^ n17207;
  assign n17615 = n17614 ^ n17231;
  assign n17643 = n17642 ^ n17615;
  assign n17541 = n16871 & n16950;
  assign n17566 = n17565 ^ n17541;
  assign n17635 = n17566 ^ n16958;
  assign n16934 = n16856 & n16933;
  assign n16949 = n16948 ^ n16934;
  assign n17636 = n17635 ^ n16949;
  assign n17535 = ~n17004 & ~n17085;
  assign n17560 = n17559 ^ n17535;
  assign n17633 = n17560 ^ n17093;
  assign n17069 = n16989 & n17068;
  assign n17084 = n17083 ^ n17069;
  assign n17634 = n17633 ^ n17084;
  assign n17637 = n17636 ^ n17634;
  assign n17644 = n17643 ^ n17637;
  assign n17655 = n17654 ^ n17644;
  assign n17355 = n17354 ^ n17353;
  assign n17335 = n17334 ^ n17333;
  assign n17350 = n17349 ^ n17335;
  assign n17356 = n17355 ^ n17350;
  assign n17460 = n17459 ^ n17356;
  assign n17227 = n17226 ^ n17225;
  assign n17222 = n17221 ^ n17207;
  assign n17228 = n17227 ^ n17222;
  assign n17237 = n17236 ^ n17228;
  assign n17088 = n17030 & ~n17074;
  assign n17090 = n17089 ^ n17088;
  assign n17094 = n17093 ^ n17090;
  assign n17087 = n17086 ^ n17084;
  assign n17095 = n17094 ^ n17087;
  assign n16953 = n16881 & n16944;
  assign n16955 = n16954 ^ n16953;
  assign n16959 = n16958 ^ n16955;
  assign n16952 = n16951 ^ n16949;
  assign n16960 = n16959 ^ n16952;
  assign n17096 = n17095 ^ n16960;
  assign n17238 = n17237 ^ n17096;
  assign n17461 = n17460 ^ n17238;
  assign n17658 = n17655 ^ n17461;
  assign n17692 = n17691 ^ n17658;
  assign n17556 = n17555 ^ n17517;
  assign n17543 = n17542 ^ n17541;
  assign n17544 = n17543 ^ n17464;
  assign n17540 = n17465 ^ n16949;
  assign n17545 = n17544 ^ n17540;
  assign n17537 = n17536 ^ n17535;
  assign n17538 = n17537 ^ n17479;
  assign n17534 = n17474 ^ n17084;
  assign n17539 = n17538 ^ n17534;
  assign n17546 = n17545 ^ n17539;
  assign n17547 = n17546 ^ n17498;
  assign n17557 = n17556 ^ n17547;
  assign n17734 = n17692 ^ n17557;
  assign n17707 = n17514 ^ n17353;
  assign n17706 = n17676 ^ n17508;
  assign n17708 = n17707 ^ n17706;
  assign n17716 = n17715 ^ n17708;
  assign n17704 = n17673 ^ n17492;
  assign n17699 = n16890 & n16943;
  assign n17700 = n17699 ^ n16958;
  assign n17599 = n16913 & n16928;
  assign n17600 = n17599 ^ n17543;
  assign n17701 = n17700 ^ n17600;
  assign n17698 = n17468 ^ n16949;
  assign n17702 = n17701 ^ n17698;
  assign n17694 = ~n17044 & n17073;
  assign n17695 = n17694 ^ n17093;
  assign n17606 = ~n17056 & ~n17067;
  assign n17607 = n17606 ^ n17537;
  assign n17696 = n17695 ^ n17607;
  assign n17693 = n17476 ^ n17084;
  assign n17697 = n17696 ^ n17693;
  assign n17703 = n17702 ^ n17697;
  assign n17705 = n17704 ^ n17703;
  assign n17717 = n17716 ^ n17705;
  assign n17618 = n17515 ^ n17335;
  assign n17619 = n17618 ^ n17504;
  assign n17629 = n17628 ^ n17619;
  assign n17573 = n17223 ^ n17213;
  assign n17576 = n17575 ^ n17573;
  assign n17571 = ~n17168 & n17218;
  assign n17572 = n17571 ^ n17488;
  assign n17577 = n17576 ^ n17572;
  assign n17616 = n17615 ^ n17577;
  assign n17610 = n17009 & n17080;
  assign n17611 = n17610 ^ n17475;
  assign n17608 = n17088 ^ n17075;
  assign n17609 = n17608 ^ n17607;
  assign n17612 = n17611 ^ n17609;
  assign n17603 = n16863 & n16940;
  assign n17604 = n17603 ^ n17467;
  assign n17601 = n16953 ^ n16947;
  assign n17602 = n17601 ^ n17600;
  assign n17605 = n17604 ^ n17602;
  assign n17613 = n17612 ^ n17605;
  assign n17617 = n17616 ^ n17613;
  assign n17630 = n17629 ^ n17617;
  assign n17738 = n17717 ^ n17630;
  assign n17745 = n17738 ^ n17691;
  assign n17584 = n17269 & n17341;
  assign n17587 = n17586 ^ n17584;
  assign n17580 = n17352 ^ n17348;
  assign n17583 = n17582 ^ n17580;
  assign n17588 = n17587 ^ n17583;
  assign n17597 = n17596 ^ n17588;
  assign n17578 = n17577 ^ n17228;
  assign n17568 = n16956 ^ n16948;
  assign n17567 = n17566 ^ n16955;
  assign n17569 = n17568 ^ n17567;
  assign n17562 = n17091 ^ n17083;
  assign n17561 = n17560 ^ n17090;
  assign n17563 = n17562 ^ n17561;
  assign n17570 = n17569 ^ n17563;
  assign n17579 = n17578 ^ n17570;
  assign n17598 = n17597 ^ n17579;
  assign n17631 = n17630 ^ n17598;
  assign n17632 = n17631 ^ n17557;
  assign n17754 = n17745 ^ n17632;
  assign n17656 = n17655 ^ n17632;
  assign n17753 = n17658 ^ n17656;
  assign n17758 = n17754 ^ n17753;
  assign n17755 = n17753 & n17754;
  assign n17533 = n17532 ^ n17461;
  assign n17748 = n17533 & n17745;
  assign n17756 = n17755 ^ n17748;
  assign n17727 = n17717 ^ n17598;
  assign n17728 = n17727 ^ n17691;
  assign n17729 = n17658 & n17728;
  assign n17722 = n17692 ^ n17631;
  assign n17723 = n17717 ^ n17461;
  assign n17726 = n17722 & n17723;
  assign n17730 = n17729 ^ n17726;
  assign n17757 = n17756 ^ n17730;
  assign n17759 = n17758 ^ n17757;
  assign n17749 = ~n17532 & n17632;
  assign n17750 = n17749 ^ n17748;
  assign n17746 = n17745 ^ n17533;
  assign n17718 = n17717 ^ n17655;
  assign n17739 = n17738 ^ n17658;
  assign n17740 = n17718 & n17739;
  assign n17741 = n17740 ^ n17729;
  assign n17747 = n17746 ^ n17741;
  assign n17751 = n17750 ^ n17747;
  assign n17771 = n17759 ^ n17751;
  assign n17737 = n17727 ^ n17692;
  assign n17742 = n17741 ^ n17737;
  assign n17732 = n17632 ^ n17532;
  assign n17733 = n17732 ^ n17723;
  assign n17735 = n17733 & n17734;
  assign n17719 = n17718 ^ n17533;
  assign n17720 = n17692 & n17719;
  assign n17736 = n17735 ^ n17720;
  assign n17743 = n17742 ^ n17736;
  assign n17752 = n17743 & n17751;
  assign n17772 = n17771 ^ n17752;
  assign n17724 = n17723 ^ n17722;
  assign n17657 = n17557 & n17656;
  assign n17721 = n17720 ^ n17657;
  assign n17725 = n17724 ^ n17721;
  assign n17731 = n17730 ^ n17725;
  assign n17769 = n17731 & n17751;
  assign n17770 = ~n17759 & n17769;
  assign n17773 = n17772 ^ n17770;
  assign n19760 = n17734 & n17773;
  assign n17775 = n17752 ^ n17731;
  assign n17776 = n17771 & n17775;
  assign n17777 = n17776 ^ n17759;
  assign n17790 = n17777 ^ n17773;
  assign n17795 = n17719 & n17790;
  assign n19761 = n19760 ^ n17795;
  assign n17789 = n17557 & n17777;
  assign n17744 = n17743 ^ n17731;
  assign n17760 = n17759 ^ n17752;
  assign n17761 = n17744 & n17760;
  assign n17762 = n17761 ^ n17731;
  assign n17787 = n17754 & n17762;
  assign n19759 = n17789 ^ n17787;
  assign n19762 = n19761 ^ n19759;
  assign n17801 = n17733 & n17773;
  assign n17765 = n17752 ^ n17744;
  assign n17763 = ~n17731 & n17743;
  assign n17764 = n17759 & n17763;
  assign n17766 = n17765 ^ n17764;
  assign n17800 = n17632 & n17766;
  assign n17802 = n17801 ^ n17800;
  assign n17778 = n17777 ^ n17762;
  assign n17781 = n17658 & n17778;
  assign n17774 = n17773 ^ n17766;
  assign n17779 = n17778 ^ n17774;
  assign n17780 = n17718 & n17779;
  assign n17782 = n17781 ^ n17780;
  assign n19758 = n17802 ^ n17782;
  assign n19763 = n19762 ^ n19758;
  assign n17798 = n17728 & n17778;
  assign n17797 = n17739 & n17779;
  assign n17799 = n17798 ^ n17797;
  assign n17803 = n17802 ^ n17799;
  assign n17767 = n17766 ^ n17762;
  assign n17783 = n17745 & n17767;
  assign n17784 = n17783 ^ n17782;
  assign n17796 = n17795 ^ n17784;
  assign n17804 = n17803 ^ n17796;
  assign n19921 = n19763 ^ n17804;
  assign n25583 = n22718 ^ n19921;
  assign n19137 = n15318 ^ n14408;
  assign n19136 = n17125 ^ n17098;
  assign n19138 = n19137 ^ n19136;
  assign n19133 = n15334 ^ n14449;
  assign n19131 = n14460 ^ n14242;
  assign n19132 = n19131 ^ n13994;
  assign n19134 = n19133 ^ n19132;
  assign n19118 = n15370 ^ n14228;
  assign n19116 = n14242 ^ n14127;
  assign n19117 = n19116 ^ n17137;
  assign n19119 = n19118 ^ n19117;
  assign n19135 = n19134 ^ n19119;
  assign n19139 = n19138 ^ n19135;
  assign n18044 = n14408 ^ n14290;
  assign n19105 = n18044 ^ n14783;
  assign n19103 = n17098 ^ n14340;
  assign n19104 = n19103 ^ n14367;
  assign n19106 = n19105 ^ n19104;
  assign n19170 = n19139 ^ n19106;
  assign n19124 = n15212 ^ n13856;
  assign n19122 = n14402 ^ n14127;
  assign n19123 = n19122 ^ n17111;
  assign n19125 = n19124 ^ n19123;
  assign n19114 = n15409 ^ n14352;
  assign n19112 = n14386 ^ n14340;
  assign n19113 = n19112 ^ n17148;
  assign n19115 = n19114 ^ n19113;
  assign n19149 = n19125 ^ n19115;
  assign n19171 = n19170 ^ n19149;
  assign n19164 = ~n19106 & n19139;
  assign n19142 = n19134 ^ n19115;
  assign n18051 = n14408 ^ n14373;
  assign n19109 = n18051 ^ n15253;
  assign n19108 = n17105 ^ n14438;
  assign n19110 = n19109 ^ n19108;
  assign n19107 = n19106 ^ n17097;
  assign n19111 = n19110 ^ n19107;
  assign n19143 = n19142 ^ n19111;
  assign n19146 = n19125 ^ n19106;
  assign n19147 = n19143 & n19146;
  assign n19165 = n19164 ^ n19147;
  assign n18070 = n14420 ^ n14408;
  assign n19128 = n18070 ^ n15282;
  assign n19126 = n17117 ^ n14460;
  assign n19127 = n19126 ^ n14264;
  assign n19129 = n19128 ^ n19127;
  assign n19130 = n19129 ^ n19125;
  assign n19159 = n19142 ^ n19130;
  assign n19160 = n19129 ^ n19115;
  assign n19161 = n19159 & n19160;
  assign n19120 = n19119 ^ n19115;
  assign n19121 = n19120 ^ n19111;
  assign n19153 = n19121 & n19130;
  assign n19162 = n19161 ^ n19153;
  assign n19158 = n19146 ^ n19143;
  assign n19163 = n19162 ^ n19158;
  assign n19166 = n19165 ^ n19163;
  assign n19150 = n19130 ^ n19111;
  assign n19175 = n19150 ^ n19120;
  assign n19176 = n19175 ^ n19162;
  assign n19172 = n19150 ^ n19138;
  assign n19173 = n19171 & n19172;
  assign n19168 = n19160 ^ n19146;
  assign n19169 = n19150 & n19168;
  assign n19174 = n19173 ^ n19169;
  assign n19177 = n19176 ^ n19174;
  assign n19178 = n19166 & n19177;
  assign n19144 = n19143 ^ n19139;
  assign n19140 = n19139 ^ n19129;
  assign n19141 = n19140 ^ n19130;
  assign n19156 = n19144 ^ n19141;
  assign n19151 = n19150 ^ n19135;
  assign n19152 = n19149 & n19151;
  assign n19154 = n19153 ^ n19152;
  assign n19145 = n19141 & n19144;
  assign n19148 = n19147 ^ n19145;
  assign n19155 = n19154 ^ n19148;
  assign n19157 = n19156 ^ n19155;
  assign n19167 = n19166 ^ n19157;
  assign n19197 = n19178 ^ n19167;
  assign n19181 = n19151 ^ n19149;
  assign n19179 = n19138 & n19140;
  assign n19180 = n19179 ^ n19169;
  assign n19182 = n19181 ^ n19180;
  assign n19183 = n19182 ^ n19154;
  assign n19195 = n19166 & n19183;
  assign n19196 = ~n19157 & n19195;
  assign n19198 = n19197 ^ n19196;
  assign n19358 = n19171 & n19198;
  assign n19187 = n19183 ^ n19177;
  assign n19208 = n19187 ^ n19178;
  assign n19206 = n19177 & ~n19183;
  assign n19207 = n19157 & n19206;
  assign n19209 = n19208 ^ n19207;
  assign n19210 = n19209 ^ n19198;
  assign n19188 = n19178 ^ n19157;
  assign n19189 = n19187 & n19188;
  assign n19190 = n19189 ^ n19183;
  assign n19184 = n19183 ^ n19178;
  assign n19185 = n19167 & n19184;
  assign n19186 = n19185 ^ n19157;
  assign n19191 = n19190 ^ n19186;
  assign n19349 = n19210 ^ n19191;
  assign n19352 = n19160 & n19349;
  assign n19193 = n19130 & n19191;
  assign n19353 = n19352 ^ n19193;
  assign n19474 = n19358 ^ n19353;
  assign n19350 = n19159 & n19349;
  assign n19192 = n19121 & n19191;
  assign n19445 = n19350 ^ n19192;
  assign n19199 = n19198 ^ n19186;
  assign n19415 = n19168 & n19199;
  assign n19414 = n19172 & n19198;
  assign n19416 = n19415 ^ n19414;
  assign n19200 = n19150 & n19199;
  assign n19417 = n19416 ^ n19200;
  assign n19473 = n19445 ^ n19417;
  assign n19475 = n19474 ^ n19473;
  assign n19482 = n19481 ^ n19475;
  assign n18995 = n17357 ^ n16111;
  assign n17951 = n16164 ^ n16122;
  assign n16080 = n16079 ^ n15962;
  assign n18994 = n17951 ^ n16080;
  assign n18996 = n18995 ^ n18994;
  assign n18992 = n17378 ^ n15713;
  assign n17922 = n16310 ^ n15849;
  assign n16282 = n16281 ^ n16277;
  assign n18991 = n17922 ^ n16282;
  assign n18993 = n18992 ^ n18991;
  assign n18997 = n18996 ^ n18993;
  assign n19009 = n17362 ^ n15616;
  assign n17940 = n16307 ^ n16175;
  assign n19008 = n17940 ^ n16840;
  assign n19010 = n19009 ^ n19008;
  assign n18988 = n17364 ^ n16087;
  assign n17933 = n16307 ^ n16265;
  assign n18986 = n17933 ^ n16830;
  assign n18987 = n18986 ^ n16844;
  assign n18989 = n18988 ^ n18987;
  assign n17937 = n16239 ^ n16146;
  assign n19007 = n18989 ^ n17937;
  assign n19011 = n19010 ^ n19007;
  assign n19001 = n17375 ^ n16209;
  assign n17927 = n16307 ^ n16135;
  assign n18999 = n17927 ^ n16864;
  assign n19000 = n18999 ^ n16850;
  assign n19002 = n19001 ^ n19000;
  assign n19004 = n19002 ^ n18993;
  assign n19021 = n19011 ^ n19004;
  assign n18982 = n17368 ^ n16292;
  assign n17956 = n16314 ^ n16277;
  assign n16206 = n16205 ^ n16199;
  assign n18981 = n17956 ^ n16206;
  assign n18983 = n18982 ^ n18981;
  assign n18979 = n17359 ^ n16221;
  assign n16248 = n16247 ^ n16244;
  assign n18978 = n16872 ^ n16248;
  assign n18980 = n18979 ^ n18978;
  assign n18984 = n18983 ^ n18980;
  assign n19022 = n19021 ^ n18984;
  assign n19050 = n19022 ^ n18997;
  assign n18976 = n17371 ^ n15721;
  assign n17945 = n16261 ^ n15839;
  assign n16311 = n16310 ^ n16307;
  assign n18975 = n17945 ^ n16311;
  assign n18977 = n18976 ^ n18975;
  assign n18985 = n18984 ^ n18977;
  assign n19003 = n19002 ^ n18985;
  assign n19048 = ~n18977 & n19003;
  assign n19029 = n19002 ^ n18996;
  assign n19015 = n18993 ^ n18989;
  assign n19040 = n19029 ^ n19015;
  assign n19041 = n19021 & ~n19040;
  assign n19049 = n19048 ^ n19041;
  assign n19051 = n19050 ^ n19049;
  assign n19023 = n18997 & n19022;
  assign n19018 = n18996 ^ n18983;
  assign n19019 = n19018 ^ n19011;
  assign n19020 = ~n19004 & ~n19019;
  assign n19024 = n19023 ^ n19020;
  assign n19052 = n19051 ^ n19024;
  assign n19043 = n19021 ^ n19018;
  assign n19006 = n18996 ^ n18980;
  assign n19030 = n19006 ^ n19004;
  assign n19031 = ~n19029 & ~n19030;
  assign n19032 = n19031 ^ n19020;
  assign n19044 = n19043 ^ n19032;
  assign n18990 = n18989 ^ n18985;
  assign n18998 = n18997 ^ n18990;
  assign n19038 = n19021 ^ n18977;
  assign n19039 = ~n18998 & ~n19038;
  assign n19042 = n19041 ^ n19039;
  assign n19045 = n19044 ^ n19042;
  assign n19059 = n19052 ^ n19045;
  assign n19034 = ~n18985 & ~n18989;
  assign n19012 = n19011 ^ n19006;
  assign n19016 = ~n19012 & n19015;
  assign n19035 = n19034 ^ n19016;
  assign n19028 = n19015 ^ n19012;
  assign n19033 = n19032 ^ n19028;
  assign n19036 = n19035 ^ n19033;
  assign n19046 = ~n19036 & n19045;
  assign n19060 = n19059 ^ n19046;
  assign n19013 = n19012 ^ n18985;
  assign n19005 = n19004 ^ n19003;
  assign n19026 = n19013 ^ n19005;
  assign n19014 = ~n19005 & n19013;
  assign n19017 = n19016 ^ n19014;
  assign n19025 = n19024 ^ n19017;
  assign n19027 = n19026 ^ n19025;
  assign n19057 = n19045 & ~n19052;
  assign n19058 = ~n19027 & n19057;
  assign n19061 = n19060 ^ n19058;
  assign n19053 = ~n19036 & n19052;
  assign n19054 = n19027 & n19053;
  assign n19037 = n19036 ^ n19027;
  assign n19047 = n19046 ^ n19037;
  assign n19055 = n19054 ^ n19047;
  assign n19081 = n19061 ^ n19055;
  assign n19468 = n18997 & n19081;
  assign n19316 = n19022 & n19081;
  assign n19074 = n19046 ^ n19027;
  assign n19075 = n19059 & ~n19074;
  assign n19076 = n19075 ^ n19052;
  assign n19077 = n19076 ^ n19061;
  assign n19315 = n19015 & n19077;
  assign n19317 = n19316 ^ n19315;
  assign n19469 = n19468 ^ n19317;
  assign n19064 = n19052 ^ n19046;
  assign n19065 = n19037 & n19064;
  assign n19066 = n19065 ^ n19027;
  assign n19079 = n19076 ^ n19066;
  assign n19407 = ~n19019 & ~n19079;
  assign n19080 = ~n19004 & ~n19079;
  assign n19466 = n19407 ^ n19080;
  assign n19464 = ~n19005 & n19076;
  assign n19401 = ~n18977 & ~n19066;
  assign n19067 = n19066 ^ n19055;
  assign n19068 = n19021 & ~n19067;
  assign n19463 = n19401 ^ n19068;
  assign n19465 = n19464 ^ n19463;
  assign n19467 = n19466 ^ n19465;
  assign n19470 = n19469 ^ n19467;
  assign n18882 = n16997 ^ n16978;
  assign n17810 = n15231 ^ n15173;
  assign n18883 = n18882 ^ n17810;
  assign n18884 = n18883 ^ n15288;
  assign n18885 = n18884 ^ n18540;
  assign n15381 = n15380 ^ n15377;
  assign n18879 = n15381 ^ n14901;
  assign n18880 = n18879 ^ n15184;
  assign n18878 = n18631 ^ n14680;
  assign n18881 = n18880 ^ n18878;
  assign n18886 = n18885 ^ n18881;
  assign n18866 = n16971 ^ n15224;
  assign n17822 = n15396 ^ n15173;
  assign n18865 = n17822 ^ n15268;
  assign n18867 = n18866 ^ n18865;
  assign n18863 = n18588 ^ n15275;
  assign n18861 = n18573 ^ n15402;
  assign n18859 = n16962 ^ n15159;
  assign n17816 = n15306 ^ n15173;
  assign n18858 = n17816 ^ n14918;
  assign n18860 = n18859 ^ n18858;
  assign n18862 = n18861 ^ n18860;
  assign n18864 = n18863 ^ n18862;
  assign n18868 = n18867 ^ n18864;
  assign n18906 = n18886 ^ n18868;
  assign n18891 = n17010 ^ n15342;
  assign n15298 = n15297 ^ n15293;
  assign n18892 = n18891 ^ n15298;
  assign n18893 = n18892 ^ n18457;
  assign n15358 = n15357 ^ n15350;
  assign n18873 = n16990 ^ n15358;
  assign n18874 = n18873 ^ n15191;
  assign n18875 = n18874 ^ n18388;
  assign n18894 = n18893 ^ n18875;
  assign n18907 = n18906 ^ n18894;
  assign n15160 = n15159 ^ n15041;
  assign n18869 = n15243 ^ n15160;
  assign n18870 = n18869 ^ n15391;
  assign n18871 = n18870 ^ n15263;
  assign n18872 = n18871 ^ n18662;
  assign n18898 = n18893 ^ n18872;
  assign n18899 = n18898 ^ n18868;
  assign n18888 = n15173 ^ n14911;
  assign n18889 = n18888 ^ n16962;
  assign n18887 = n18505 ^ n14670;
  assign n18890 = n18889 ^ n18887;
  assign n18895 = n18894 ^ n18890;
  assign n18900 = n18899 ^ n18895;
  assign n18896 = n18895 ^ n18885;
  assign n18897 = n18896 ^ n18886;
  assign n18912 = n18900 ^ n18897;
  assign n18876 = n18875 ^ n18872;
  assign n18877 = n18876 ^ n18868;
  assign n18909 = n18877 & n18886;
  assign n18905 = n18881 ^ n18872;
  assign n18908 = n18905 & ~n18907;
  assign n18910 = n18909 ^ n18908;
  assign n18902 = n18881 ^ n18862;
  assign n18903 = n18899 & ~n18902;
  assign n18901 = ~n18897 & ~n18900;
  assign n18904 = n18903 ^ n18901;
  assign n18911 = n18910 ^ n18904;
  assign n18913 = n18912 ^ n18911;
  assign n18931 = n18906 ^ n18876;
  assign n18915 = n18885 ^ n18872;
  assign n18916 = n18898 ^ n18886;
  assign n18917 = n18915 & ~n18916;
  assign n18918 = n18917 ^ n18909;
  assign n18932 = n18931 ^ n18918;
  assign n18926 = n18906 ^ n18890;
  assign n18927 = n18895 ^ n18862;
  assign n18928 = n18927 ^ n18905;
  assign n18929 = n18926 & n18928;
  assign n18924 = n18915 ^ n18902;
  assign n18925 = ~n18906 & ~n18924;
  assign n18930 = n18929 ^ n18925;
  assign n18933 = n18932 ^ n18930;
  assign n18937 = n18907 ^ n18905;
  assign n18935 = ~n18890 & ~n18896;
  assign n18936 = n18935 ^ n18925;
  assign n18938 = n18937 ^ n18936;
  assign n18939 = n18938 ^ n18910;
  assign n18963 = n18933 & n18939;
  assign n18964 = n18913 & n18963;
  assign n18943 = n18939 ^ n18933;
  assign n18920 = n18862 & ~n18895;
  assign n18921 = n18920 ^ n18903;
  assign n18914 = n18902 ^ n18899;
  assign n18919 = n18918 ^ n18914;
  assign n18922 = n18921 ^ n18919;
  assign n18934 = ~n18922 & n18933;
  assign n18962 = n18943 ^ n18934;
  assign n18965 = n18964 ^ n18962;
  assign n18923 = n18922 ^ n18913;
  assign n18954 = n18934 ^ n18923;
  assign n18952 = ~n18922 & ~n18939;
  assign n18953 = ~n18913 & n18952;
  assign n18955 = n18954 ^ n18953;
  assign n18966 = n18965 ^ n18955;
  assign n18970 = ~n18907 & n18966;
  assign n18944 = n18934 ^ n18913;
  assign n18945 = ~n18943 & n18944;
  assign n18946 = n18945 ^ n18939;
  assign n18968 = n18965 ^ n18946;
  assign n18969 = ~n18902 & n18968;
  assign n18971 = n18970 ^ n18969;
  assign n18967 = n18905 & n18966;
  assign n18972 = n18971 ^ n18967;
  assign n18959 = ~n18897 & ~n18946;
  assign n18940 = n18939 ^ n18934;
  assign n18941 = ~n18923 & ~n18940;
  assign n18942 = n18941 ^ n18913;
  assign n18956 = n18955 ^ n18942;
  assign n18957 = ~n18906 & ~n18956;
  assign n18951 = ~n18890 & n18942;
  assign n18958 = n18957 ^ n18951;
  assign n18960 = n18959 ^ n18958;
  assign n18947 = n18946 ^ n18942;
  assign n18949 = n18886 & ~n18947;
  assign n18948 = n18877 & ~n18947;
  assign n18950 = n18949 ^ n18948;
  assign n18961 = n18960 ^ n18950;
  assign n18973 = n18972 ^ n18961;
  assign n19471 = n19470 ^ n18973;
  assign n18777 = n16270 ^ n13438;
  assign n18775 = n13342 ^ n13334;
  assign n18205 = n13174 ^ n12248;
  assign n18776 = n18775 ^ n18205;
  assign n18778 = n18777 ^ n18776;
  assign n18772 = n16228 ^ n13490;
  assign n18197 = n13317 ^ n13309;
  assign n13457 = n13456 ^ n13451;
  assign n18771 = n18197 ^ n13457;
  assign n18773 = n18772 ^ n18771;
  assign n18748 = n16297 ^ n13465;
  assign n18172 = n13490 ^ n13481;
  assign n11318 = n11317 ^ n10367;
  assign n18747 = n18172 ^ n11318;
  assign n18749 = n18748 ^ n18747;
  assign n18774 = n18773 ^ n18749;
  assign n18779 = n18778 ^ n18774;
  assign n18753 = n16099 ^ n13372;
  assign n18164 = n13432 ^ n12248;
  assign n18751 = n18164 ^ n17251;
  assign n13507 = n13506 ^ n13360;
  assign n18752 = n18751 ^ n13507;
  assign n18754 = n18753 ^ n18752;
  assign n18808 = n18779 ^ n18754;
  assign n18764 = n16320 ^ n13174;
  assign n18762 = n13465 ^ n13460;
  assign n13428 = n13293 ^ n12256;
  assign n18763 = n18762 ^ n13428;
  assign n18765 = n18764 ^ n18763;
  assign n18745 = n16189 ^ n13519;
  assign n18743 = n13410 ^ n13399;
  assign n18742 = n13372 ^ n13354;
  assign n18744 = n18743 ^ n18742;
  assign n18746 = n18745 ^ n18744;
  assign n18792 = n18765 ^ n18746;
  assign n18809 = n18808 ^ n18792;
  assign n18804 = ~n18754 & n18779;
  assign n18782 = n18773 ^ n18746;
  assign n18758 = n13299 ^ n13284;
  assign n18184 = n13512 ^ n12248;
  assign n18757 = n18184 ^ n17256;
  assign n18759 = n18758 ^ n18757;
  assign n18755 = n15701 ^ n13417;
  assign n18756 = n18755 ^ n18754;
  assign n18760 = n18759 ^ n18756;
  assign n18783 = n18782 ^ n18760;
  assign n18786 = n18765 ^ n18754;
  assign n18787 = n18783 & n18786;
  assign n18805 = n18804 ^ n18787;
  assign n18768 = n16253 ^ n13317;
  assign n18198 = n13390 ^ n12248;
  assign n18766 = n18198 ^ n17241;
  assign n13474 = n13473 ^ n13303;
  assign n18767 = n18766 ^ n13474;
  assign n18769 = n18768 ^ n18767;
  assign n18799 = n18769 ^ n18746;
  assign n18770 = n18769 ^ n18765;
  assign n18800 = n18782 ^ n18770;
  assign n18801 = n18799 & n18800;
  assign n18750 = n18749 ^ n18746;
  assign n18761 = n18760 ^ n18750;
  assign n18789 = n18761 & n18770;
  assign n18802 = n18801 ^ n18789;
  assign n18798 = n18786 ^ n18783;
  assign n18803 = n18802 ^ n18798;
  assign n18806 = n18805 ^ n18803;
  assign n18790 = n18770 ^ n18760;
  assign n18815 = n18790 ^ n18750;
  assign n18816 = n18815 ^ n18802;
  assign n18812 = n18799 ^ n18786;
  assign n18813 = n18790 & n18812;
  assign n18810 = n18790 ^ n18778;
  assign n18811 = n18809 & n18810;
  assign n18814 = n18813 ^ n18811;
  assign n18817 = n18816 ^ n18814;
  assign n18818 = n18806 & n18817;
  assign n18784 = n18783 ^ n18779;
  assign n18780 = n18779 ^ n18769;
  assign n18781 = n18780 ^ n18770;
  assign n18796 = n18784 ^ n18781;
  assign n18791 = n18790 ^ n18774;
  assign n18793 = n18791 & n18792;
  assign n18794 = n18793 ^ n18789;
  assign n18785 = n18781 & n18784;
  assign n18788 = n18787 ^ n18785;
  assign n18795 = n18794 ^ n18788;
  assign n18797 = n18796 ^ n18795;
  assign n18807 = n18806 ^ n18797;
  assign n18837 = n18818 ^ n18807;
  assign n18821 = n18792 ^ n18791;
  assign n18819 = n18778 & n18780;
  assign n18820 = n18819 ^ n18813;
  assign n18822 = n18821 ^ n18820;
  assign n18823 = n18822 ^ n18794;
  assign n18835 = n18806 & n18823;
  assign n18836 = ~n18797 & n18835;
  assign n18838 = n18837 ^ n18836;
  assign n19336 = n18809 & n18838;
  assign n18827 = n18823 ^ n18817;
  assign n18848 = n18827 ^ n18818;
  assign n18846 = n18817 & ~n18823;
  assign n18847 = n18797 & n18846;
  assign n18849 = n18848 ^ n18847;
  assign n18850 = n18849 ^ n18838;
  assign n18828 = n18818 ^ n18797;
  assign n18829 = n18827 & n18828;
  assign n18830 = n18829 ^ n18823;
  assign n18824 = n18823 ^ n18818;
  assign n18825 = n18807 & n18824;
  assign n18826 = n18825 ^ n18797;
  assign n18831 = n18830 ^ n18826;
  assign n19327 = n18850 ^ n18831;
  assign n19330 = n18799 & n19327;
  assign n18833 = n18770 & n18831;
  assign n19331 = n19330 ^ n18833;
  assign n19460 = n19336 ^ n19331;
  assign n19328 = n18800 & n19327;
  assign n18832 = n18761 & n18831;
  assign n19439 = n19328 ^ n18832;
  assign n18839 = n18838 ^ n18826;
  assign n19386 = n18812 & n18839;
  assign n19385 = n18810 & n18838;
  assign n19387 = n19386 ^ n19385;
  assign n18840 = n18790 & n18839;
  assign n19388 = n19387 ^ n18840;
  assign n19459 = n19439 ^ n19388;
  assign n19461 = n19460 ^ n19459;
  assign n19095 = n18966 ^ n18947;
  assign n19096 = n18915 & ~n19095;
  assign n19097 = n19096 ^ n18949;
  assign n19092 = n18928 & ~n18955;
  assign n19432 = n19097 ^ n19092;
  assign n19311 = ~n18916 & ~n19095;
  assign n19397 = n19311 ^ n18948;
  assign n19088 = ~n18924 & ~n18956;
  assign n19087 = n18926 & ~n18955;
  assign n19089 = n19088 ^ n19087;
  assign n19090 = n19089 ^ n18957;
  assign n19431 = n19397 ^ n19090;
  assign n19433 = n19432 ^ n19431;
  assign n19462 = n19461 ^ n19433;
  assign n19472 = n19471 ^ n19462;
  assign n19483 = n19482 ^ n19472;
  assign n19360 = n19140 & n19186;
  assign n19357 = n19139 & n19209;
  assign n19359 = n19358 ^ n19357;
  assign n19361 = n19360 ^ n19359;
  assign n19203 = n19141 & n19190;
  assign n19201 = n19138 & n19186;
  assign n19202 = n19201 ^ n19200;
  assign n19204 = n19203 ^ n19202;
  assign n19362 = n19361 ^ n19204;
  assign n19212 = n19209 ^ n19190;
  assign n19354 = n19143 & n19212;
  assign n19355 = n19354 ^ n19353;
  assign n19214 = n19151 & n19210;
  assign n19213 = n19146 & n19212;
  assign n19215 = n19214 ^ n19213;
  assign n19351 = n19350 ^ n19215;
  assign n19356 = n19355 ^ n19351;
  assign n19363 = n19362 ^ n19356;
  assign n19382 = n19381 ^ n19363;
  assign n19343 = ~n18896 & n18942;
  assign n19091 = ~n18895 & ~n18965;
  assign n19093 = n19092 ^ n19091;
  assign n19344 = n19343 ^ n19093;
  assign n19345 = n19344 ^ n18960;
  assign n19312 = n19311 ^ n18971;
  assign n19098 = n18899 & n18968;
  assign n19099 = n19098 ^ n19097;
  assign n19342 = n19312 ^ n19099;
  assign n19346 = n19345 ^ n19342;
  assign n19338 = n18780 & n18826;
  assign n19335 = n18779 & n18849;
  assign n19337 = n19336 ^ n19335;
  assign n19339 = n19338 ^ n19337;
  assign n18843 = n18781 & n18830;
  assign n18841 = n18778 & n18826;
  assign n18842 = n18841 ^ n18840;
  assign n18844 = n18843 ^ n18842;
  assign n19340 = n19339 ^ n18844;
  assign n18852 = n18849 ^ n18830;
  assign n19332 = n18783 & n18852;
  assign n19333 = n19332 ^ n19331;
  assign n18854 = n18791 & n18850;
  assign n18853 = n18786 & n18852;
  assign n18855 = n18854 ^ n18853;
  assign n19329 = n19328 ^ n18855;
  assign n19334 = n19333 ^ n19329;
  assign n19341 = n19340 ^ n19334;
  assign n19347 = n19346 ^ n19341;
  assign n19082 = n19081 ^ n19079;
  assign n19083 = ~n19029 & ~n19082;
  assign n19084 = n19083 ^ n19080;
  assign n19062 = ~n18985 & n19061;
  assign n19324 = n19084 ^ n19062;
  assign n19321 = ~n18990 & n19061;
  assign n19320 = n19013 & n19076;
  assign n19322 = n19321 ^ n19320;
  assign n19318 = ~n19030 & ~n19082;
  assign n19319 = n19318 ^ n19317;
  assign n19323 = n19322 ^ n19319;
  assign n19325 = n19324 ^ n19323;
  assign n19309 = ~n18900 & ~n18946;
  assign n19308 = n18927 & ~n18965;
  assign n19310 = n19309 ^ n19308;
  assign n19313 = n19312 ^ n19310;
  assign n19307 = n19097 ^ n19091;
  assign n19314 = n19313 ^ n19307;
  assign n19326 = n19325 ^ n19314;
  assign n19348 = n19347 ^ n19326;
  assign n19383 = n19382 ^ n19348;
  assign n19577 = n19483 ^ n19383;
  assign n19499 = n19144 & n19190;
  assign n19554 = n19499 ^ n19201;
  assign n19555 = n19554 ^ n19416;
  assign n19553 = n19359 ^ n19353;
  assign n19556 = n19555 ^ n19553;
  assign n19564 = n19563 ^ n19556;
  assign n19078 = ~n19012 & n19077;
  assign n19085 = n19084 ^ n19078;
  assign n19549 = n19319 ^ n19085;
  assign n19546 = n19003 & ~n19066;
  assign n19056 = ~n18998 & n19055;
  assign n19063 = n19062 ^ n19056;
  assign n19547 = n19546 ^ n19063;
  assign n19548 = n19547 ^ n19465;
  assign n19550 = n19549 ^ n19548;
  assign n19408 = n19407 ^ n19318;
  assign n19409 = n19408 ^ n19063;
  assign n19069 = ~n19040 & ~n19067;
  assign n19406 = n19085 ^ n19069;
  assign n19410 = n19409 ^ n19406;
  assign n19551 = n19550 ^ n19410;
  assign n19398 = n19397 ^ n19093;
  assign n19396 = n19099 ^ n19088;
  assign n19399 = n19398 ^ n19396;
  assign n19545 = n19399 ^ n19346;
  assign n19552 = n19551 ^ n19545;
  assign n19565 = n19564 ^ n19552;
  assign n19488 = n18784 & n18830;
  assign n19540 = n19488 ^ n18841;
  assign n19541 = n19540 ^ n19387;
  assign n19539 = n19337 ^ n19331;
  assign n19542 = n19541 ^ n19539;
  assign n19393 = n19309 ^ n18951;
  assign n19394 = n19393 ^ n19089;
  assign n19392 = n19097 ^ n19093;
  assign n19395 = n19394 ^ n19392;
  assign n19543 = n19542 ^ n19395;
  assign n19529 = n19357 ^ n19353;
  assign n19498 = n19170 & n19209;
  assign n19500 = n19499 ^ n19498;
  assign n19528 = n19500 ^ n19351;
  assign n19530 = n19529 ^ n19528;
  assign n19537 = n19536 ^ n19530;
  assign n19523 = n19463 ^ n19322;
  assign n19522 = n19315 ^ n19085;
  assign n19524 = n19523 ^ n19522;
  assign n19525 = n19524 ^ n19410;
  assign n19493 = n19310 ^ n18958;
  assign n19492 = n19099 ^ n18969;
  assign n19494 = n19493 ^ n19492;
  assign n19521 = n19494 ^ n19399;
  assign n19526 = n19525 ^ n19521;
  assign n19518 = n19335 ^ n19331;
  assign n19487 = n18808 & n18849;
  assign n19489 = n19488 ^ n19487;
  assign n19517 = n19489 ^ n19329;
  assign n19519 = n19518 ^ n19517;
  assign n19520 = n19519 ^ n19314;
  assign n19527 = n19526 ^ n19520;
  assign n19538 = n19537 ^ n19527;
  assign n19544 = n19543 ^ n19538;
  assign n19566 = n19565 ^ n19544;
  assign n19578 = n19577 ^ n19566;
  assign n19446 = n19445 ^ n19359;
  assign n19444 = n19415 ^ n19355;
  assign n19447 = n19446 ^ n19444;
  assign n19455 = n19454 ^ n19447;
  assign n19440 = n19439 ^ n19337;
  assign n19438 = n19386 ^ n19333;
  assign n19441 = n19440 ^ n19438;
  assign n19442 = n19441 ^ n19399;
  assign n19435 = n19084 ^ n19056;
  assign n19070 = ~n19038 & n19055;
  assign n19071 = n19070 ^ n19069;
  assign n19072 = n19071 ^ n19068;
  assign n19434 = n19408 ^ n19072;
  assign n19436 = n19435 ^ n19434;
  assign n19437 = n19436 ^ n19433;
  assign n19443 = n19442 ^ n19437;
  assign n19456 = n19455 ^ n19443;
  assign n19418 = n19417 ^ n19359;
  assign n19419 = n19418 ^ n19355;
  assign n19429 = n19428 ^ n19419;
  assign n19404 = n19084 ^ n19063;
  assign n19402 = n19401 ^ n19320;
  assign n19403 = n19402 ^ n19071;
  assign n19405 = n19404 ^ n19403;
  assign n19411 = n19410 ^ n19405;
  assign n19400 = n19399 ^ n19395;
  assign n19412 = n19411 ^ n19400;
  assign n19389 = n19388 ^ n19337;
  assign n19390 = n19389 ^ n19333;
  assign n19094 = n19093 ^ n19090;
  assign n19100 = n19099 ^ n19094;
  assign n19391 = n19390 ^ n19100;
  assign n19413 = n19412 ^ n19391;
  assign n19430 = n19429 ^ n19413;
  assign n19457 = n19456 ^ n19430;
  assign n19574 = n19566 ^ n19457;
  assign n19211 = n19149 & n19210;
  assign n19216 = n19215 ^ n19211;
  assign n19194 = n19193 ^ n19192;
  assign n19205 = n19204 ^ n19194;
  assign n19217 = n19216 ^ n19205;
  assign n19305 = n19304 ^ n19217;
  assign n19073 = n19072 ^ n19063;
  assign n19086 = n19085 ^ n19073;
  assign n19101 = n19100 ^ n19086;
  assign n18851 = n18792 & n18850;
  assign n18856 = n18855 ^ n18851;
  assign n18834 = n18833 ^ n18832;
  assign n18845 = n18844 ^ n18834;
  assign n18857 = n18856 ^ n18845;
  assign n18974 = n18973 ^ n18857;
  assign n19102 = n19101 ^ n18974;
  assign n19306 = n19305 ^ n19102;
  assign n19484 = n19483 ^ n19306;
  assign n19575 = n19574 ^ n19484;
  assign n19573 = n19456 ^ n19383;
  assign n19606 = n19575 ^ n19573;
  assign n19501 = n19500 ^ n19202;
  assign n19497 = n19355 ^ n19213;
  assign n19502 = n19501 ^ n19497;
  assign n19512 = n19511 ^ n19502;
  assign n19490 = n19489 ^ n18842;
  assign n19486 = n19333 ^ n18853;
  assign n19491 = n19490 ^ n19486;
  assign n19495 = n19494 ^ n19491;
  assign n19485 = n19410 ^ n19399;
  assign n19496 = n19495 ^ n19485;
  assign n19513 = n19512 ^ n19496;
  assign n19514 = n19513 ^ n19484;
  assign n19515 = n19514 ^ n19430;
  assign n19604 = n19513 & n19515;
  assign n19585 = n19430 ^ n19383;
  assign n19570 = n19538 ^ n19456;
  assign n19593 = n19585 ^ n19570;
  assign n19594 = ~n19574 & ~n19593;
  assign n19605 = n19604 ^ n19594;
  assign n19607 = n19606 ^ n19605;
  assign n19579 = ~n19457 & ~n19578;
  assign n19576 = n19573 & n19575;
  assign n19580 = n19579 ^ n19576;
  assign n19608 = n19607 ^ n19580;
  assign n19600 = n19577 ^ n19574;
  assign n19384 = n19383 ^ n19306;
  assign n19458 = n19457 ^ n19384;
  assign n19586 = ~n19458 & ~n19585;
  assign n19587 = n19586 ^ n19579;
  assign n19601 = n19600 ^ n19587;
  assign n19595 = n19574 ^ n19513;
  assign n19596 = n19538 ^ n19514;
  assign n19597 = n19596 ^ n19573;
  assign n19598 = ~n19595 & ~n19597;
  assign n19599 = n19598 ^ n19594;
  assign n19602 = n19601 ^ n19599;
  assign n19612 = n19608 ^ n19602;
  assign n19589 = ~n19514 & ~n19538;
  assign n19567 = n19566 ^ n19384;
  assign n19571 = n19567 & n19570;
  assign n19590 = n19589 ^ n19571;
  assign n19584 = n19570 ^ n19567;
  assign n19588 = n19587 ^ n19584;
  assign n19591 = n19590 ^ n19588;
  assign n19603 = n19591 & n19602;
  assign n19568 = n19567 ^ n19514;
  assign n19516 = n19515 ^ n19457;
  assign n19582 = n19568 ^ n19516;
  assign n19569 = ~n19516 & ~n19568;
  assign n19572 = n19571 ^ n19569;
  assign n19581 = n19580 ^ n19572;
  assign n19583 = n19582 ^ n19581;
  assign n19613 = n19603 ^ n19583;
  assign n19614 = n19612 & n19613;
  assign n19615 = n19614 ^ n19608;
  assign n19592 = n19591 ^ n19583;
  assign n19609 = n19608 ^ n19603;
  assign n19610 = n19592 & n19609;
  assign n19611 = n19610 ^ n19583;
  assign n19616 = n19615 ^ n19611;
  assign n19888 = ~n19578 & n19616;
  assign n19623 = n19612 ^ n19603;
  assign n19621 = n19602 & ~n19608;
  assign n19622 = n19583 & n19621;
  assign n19624 = n19623 ^ n19622;
  assign n19619 = n19603 ^ n19592;
  assign n19617 = n19591 & n19608;
  assign n19618 = ~n19583 & n19617;
  assign n19620 = n19619 ^ n19618;
  assign n19625 = n19624 ^ n19620;
  assign n19626 = n19625 ^ n19616;
  assign n19627 = ~n19458 & n19626;
  assign n19953 = n19888 ^ n19627;
  assign n19813 = ~n19597 & n19620;
  assign n19637 = ~n19514 & n19624;
  assign n19814 = n19813 ^ n19637;
  assign n19954 = n19953 ^ n19814;
  assign n19629 = n19624 ^ n19615;
  assign n19838 = n19567 & n19629;
  assign n19639 = ~n19457 & n19616;
  assign n19638 = ~n19585 & n19626;
  assign n19640 = n19639 ^ n19638;
  assign n19839 = n19838 ^ n19640;
  assign n19819 = n19620 ^ n19611;
  assign n19820 = ~n19593 & n19819;
  assign n19952 = n19839 ^ n19820;
  assign n19955 = n19954 ^ n19952;
  assign n19818 = ~n19595 & n19620;
  assign n19821 = n19820 ^ n19818;
  assign n19816 = n19513 & n19611;
  assign n19634 = ~n19568 & n19615;
  assign n19817 = n19816 ^ n19634;
  assign n19822 = n19821 ^ n19817;
  assign n19815 = n19814 ^ n19640;
  assign n19823 = n19822 ^ n19815;
  assign n24272 = n19955 ^ n19823;
  assign n19843 = ~n19574 & n19819;
  assign n19926 = n19843 ^ n19821;
  assign n19927 = n19926 ^ n19814;
  assign n19928 = n19927 ^ n19839;
  assign n25581 = n24272 ^ n19928;
  assign n17965 = n16209 ^ n15335;
  assign n17963 = n16244 ^ n16199;
  assign n17964 = n17963 ^ n16872;
  assign n17966 = n17965 ^ n17964;
  assign n17958 = n16221 ^ n15371;
  assign n17955 = n16281 ^ n16199;
  assign n17957 = n17956 ^ n17955;
  assign n17959 = n17958 ^ n17957;
  assign n17967 = n17966 ^ n17959;
  assign n17947 = n15713 ^ n15319;
  assign n17946 = n17945 ^ n17933;
  assign n17948 = n17947 ^ n17946;
  assign n17976 = n17967 ^ n17948;
  assign n17953 = n16087 ^ n15410;
  assign n17950 = n16175 ^ n15962;
  assign n17952 = n17951 ^ n17950;
  assign n17954 = n17953 ^ n17952;
  assign n17960 = n17959 ^ n17954;
  assign n17941 = n17940 ^ n16135;
  assign n16112 = n16111 ^ n15713;
  assign n17939 = n16112 ^ n15254;
  assign n17942 = n17941 ^ n17939;
  assign n17934 = n17933 ^ n15962;
  assign n17935 = n17934 ^ n16844;
  assign n15722 = n15721 ^ n15713;
  assign n17932 = n15722 ^ n14784;
  assign n17936 = n17935 ^ n17932;
  assign n17938 = n17937 ^ n17936;
  assign n17943 = n17942 ^ n17938;
  assign n17928 = n17927 ^ n16244;
  assign n17929 = n17928 ^ n16850;
  assign n16235 = n15713 ^ n15616;
  assign n17926 = n16235 ^ n15283;
  assign n17930 = n17929 ^ n17926;
  assign n17924 = n16292 ^ n15213;
  assign n17921 = n16307 ^ n16281;
  assign n17923 = n17922 ^ n17921;
  assign n17925 = n17924 ^ n17923;
  assign n17931 = n17930 ^ n17925;
  assign n17944 = n17943 ^ n17931;
  assign n18007 = n17960 ^ n17944;
  assign n17985 = n17954 ^ n17930;
  assign n17972 = n17966 ^ n17954;
  assign n17986 = n17972 ^ n17931;
  assign n17987 = n17985 & n17986;
  assign n17961 = n17960 ^ n17943;
  assign n17962 = n17931 & n17961;
  assign n17988 = n17987 ^ n17962;
  assign n18008 = n18007 ^ n17988;
  assign n17949 = n17948 ^ n17944;
  assign n18003 = n17976 ^ n17936;
  assign n17969 = n17954 ^ n17925;
  assign n18004 = n18003 ^ n17969;
  assign n18005 = n17949 & n18004;
  assign n17974 = n17936 ^ n17925;
  assign n17995 = n17985 ^ n17974;
  assign n17996 = n17944 & n17995;
  assign n18006 = n18005 ^ n17996;
  assign n18009 = n18008 ^ n18006;
  assign n17968 = n17967 ^ n17944;
  assign n17998 = n17969 ^ n17968;
  assign n17978 = n17976 ^ n17930;
  assign n17994 = n17948 & n17978;
  assign n17997 = n17996 ^ n17994;
  assign n17999 = n17998 ^ n17997;
  assign n17970 = n17968 & n17969;
  assign n17971 = n17970 ^ n17962;
  assign n18000 = n17999 ^ n17971;
  assign n18023 = n18009 ^ n18000;
  assign n17991 = ~n17936 & n17976;
  assign n17973 = n17972 ^ n17943;
  assign n17975 = n17973 & n17974;
  assign n17992 = n17991 ^ n17975;
  assign n17989 = n17974 ^ n17973;
  assign n17990 = n17989 ^ n17988;
  assign n17993 = n17992 ^ n17990;
  assign n18010 = n17993 & n18009;
  assign n18031 = n18023 ^ n18010;
  assign n17979 = n17978 ^ n17931;
  assign n17977 = n17976 ^ n17973;
  assign n17983 = n17979 ^ n17977;
  assign n17980 = n17977 & n17979;
  assign n17981 = n17980 ^ n17975;
  assign n17982 = n17981 ^ n17971;
  assign n17984 = n17983 ^ n17982;
  assign n18029 = ~n18000 & n18009;
  assign n18030 = n17984 & n18029;
  assign n18032 = n18031 ^ n18030;
  assign n18520 = n17976 & n18032;
  assign n18011 = n17993 ^ n17984;
  assign n18012 = n18011 ^ n18010;
  assign n18001 = n17993 & n18000;
  assign n18002 = ~n17984 & n18001;
  assign n18013 = n18012 ^ n18002;
  assign n18041 = n18004 & n18013;
  assign n18521 = n18520 ^ n18041;
  assign n18033 = n18032 ^ n18013;
  assign n18024 = n18010 ^ n17984;
  assign n18025 = n18023 & n18024;
  assign n18026 = n18025 ^ n18000;
  assign n18015 = n18010 ^ n18000;
  assign n18016 = n18011 & n18015;
  assign n18017 = n18016 ^ n17984;
  assign n18027 = n18026 ^ n18017;
  assign n18034 = n18033 ^ n18027;
  assign n18035 = n17986 & n18034;
  assign n18028 = n17961 & n18027;
  assign n18036 = n18035 ^ n18028;
  assign n18623 = n18521 ^ n18036;
  assign n18432 = n18032 ^ n18026;
  assign n18486 = n17973 & n18432;
  assign n18039 = n17931 & n18027;
  assign n18038 = n17985 & n18034;
  assign n18040 = n18039 ^ n18038;
  assign n18487 = n18486 ^ n18040;
  assign n18018 = n18017 ^ n18013;
  assign n18019 = n17995 & n18018;
  assign n18622 = n18487 ^ n18019;
  assign n18624 = n18623 ^ n18622;
  assign n18633 = n18632 ^ n18624;
  assign n18199 = n18198 ^ n18197;
  assign n13285 = n13284 ^ n12256;
  assign n18200 = n18199 ^ n13285;
  assign n18201 = n18200 ^ n13473;
  assign n18202 = n18201 ^ n14464;
  assign n18168 = n13519 ^ n13361;
  assign n18169 = n18168 ^ n13512;
  assign n18170 = n18169 ^ n13410;
  assign n18171 = n18170 ^ n14394;
  assign n18226 = n18202 ^ n18171;
  assign n18192 = n14213 ^ n13465;
  assign n18190 = n13482 ^ n11317;
  assign n18191 = n18190 ^ n13460;
  assign n18193 = n18192 ^ n18191;
  assign n18218 = n18193 ^ n18171;
  assign n18204 = n13461 ^ n13293;
  assign n18206 = n18205 ^ n18204;
  assign n18207 = n18206 ^ n14412;
  assign n18208 = n18207 ^ n18202;
  assign n13400 = n13399 ^ n12256;
  assign n18186 = n13400 ^ n13299;
  assign n18185 = n18184 ^ n13390;
  assign n18187 = n18186 ^ n18185;
  assign n18182 = n14425 ^ n13417;
  assign n18180 = n14358 ^ n13372;
  assign n13335 = n13334 ^ n12256;
  assign n18178 = n13506 ^ n13335;
  assign n18177 = n18164 ^ n13354;
  assign n18179 = n18178 ^ n18177;
  assign n18181 = n18180 ^ n18179;
  assign n18183 = n18182 ^ n18181;
  assign n18188 = n18187 ^ n18183;
  assign n18215 = n18208 ^ n18188;
  assign n18247 = n18218 ^ n18215;
  assign n18173 = n18172 ^ n13456;
  assign n18174 = n18173 ^ n13310;
  assign n18175 = n18174 ^ n14279;
  assign n18176 = n18175 ^ n18171;
  assign n18227 = n18208 ^ n18176;
  assign n18228 = n18226 & n18227;
  assign n18219 = n18218 ^ n18188;
  assign n18220 = n18208 & n18219;
  assign n18229 = n18228 ^ n18220;
  assign n18248 = n18247 ^ n18229;
  assign n18166 = n14299 ^ n13438;
  assign n18163 = n13342 ^ n12256;
  assign n18165 = n18164 ^ n18163;
  assign n18167 = n18166 ^ n18165;
  assign n18242 = n18215 ^ n18167;
  assign n18194 = n18193 ^ n18175;
  assign n18195 = n18194 ^ n18167;
  assign n18243 = n18195 ^ n18181;
  assign n18214 = n18207 ^ n18171;
  assign n18244 = n18243 ^ n18214;
  assign n18245 = n18242 & n18244;
  assign n18211 = n18207 ^ n18181;
  assign n18236 = n18226 ^ n18211;
  assign n18237 = n18215 & n18236;
  assign n18246 = n18245 ^ n18237;
  assign n18249 = n18248 ^ n18246;
  assign n18216 = n18215 ^ n18194;
  assign n18239 = n18216 ^ n18214;
  assign n18203 = n18202 ^ n18195;
  assign n18235 = n18167 & n18203;
  assign n18238 = n18237 ^ n18235;
  assign n18240 = n18239 ^ n18238;
  assign n18217 = n18214 & n18216;
  assign n18221 = n18220 ^ n18217;
  assign n18241 = n18240 ^ n18221;
  assign n18262 = n18249 ^ n18241;
  assign n18231 = ~n18181 & n18195;
  assign n18189 = n18188 ^ n18176;
  assign n18212 = n18189 & n18211;
  assign n18232 = n18231 ^ n18212;
  assign n18225 = n18211 ^ n18189;
  assign n18230 = n18229 ^ n18225;
  assign n18233 = n18232 ^ n18230;
  assign n18250 = n18233 & n18249;
  assign n18275 = n18262 ^ n18250;
  assign n18209 = n18208 ^ n18203;
  assign n18196 = n18195 ^ n18189;
  assign n18223 = n18209 ^ n18196;
  assign n18210 = n18196 & n18209;
  assign n18213 = n18212 ^ n18210;
  assign n18222 = n18221 ^ n18213;
  assign n18224 = n18223 ^ n18222;
  assign n18273 = ~n18241 & n18249;
  assign n18274 = n18224 & n18273;
  assign n18276 = n18275 ^ n18274;
  assign n18234 = n18233 ^ n18224;
  assign n18257 = n18250 ^ n18234;
  assign n18255 = n18233 & n18241;
  assign n18256 = ~n18224 & n18255;
  assign n18258 = n18257 ^ n18256;
  assign n18277 = n18276 ^ n18258;
  assign n18263 = n18250 ^ n18224;
  assign n18264 = n18262 & n18263;
  assign n18265 = n18264 ^ n18241;
  assign n18251 = n18250 ^ n18241;
  assign n18252 = n18234 & n18251;
  assign n18253 = n18252 ^ n18224;
  assign n18268 = n18265 ^ n18253;
  assign n18400 = n18277 ^ n18268;
  assign n18401 = n18226 & n18400;
  assign n18270 = n18208 & n18268;
  assign n18402 = n18401 ^ n18270;
  assign n18391 = n18244 & n18258;
  assign n18617 = n18402 ^ n18391;
  assign n18480 = n18227 & n18400;
  assign n18269 = n18219 & n18268;
  assign n18481 = n18480 ^ n18269;
  assign n18395 = n18242 & n18258;
  assign n18259 = n18258 ^ n18253;
  assign n18394 = n18236 & n18259;
  assign n18396 = n18395 ^ n18394;
  assign n18260 = n18215 & n18259;
  assign n18397 = n18396 ^ n18260;
  assign n18616 = n18481 ^ n18397;
  assign n18618 = n18617 ^ n18616;
  assign n18073 = n16254 ^ n14449;
  assign n14451 = n14444 ^ n14318;
  assign n18071 = n18070 ^ n14451;
  assign n18072 = n18071 ^ n17132;
  assign n18074 = n18073 ^ n18072;
  assign n18067 = n16321 ^ n14408;
  assign n13857 = n13856 ^ n13738;
  assign n18066 = n17126 ^ n13857;
  assign n18068 = n18067 ^ n18066;
  assign n18075 = n18074 ^ n18068;
  assign n18047 = n16100 ^ n14352;
  assign n14325 = n14324 ^ n14318;
  assign n18045 = n18044 ^ n14325;
  assign n18046 = n18045 ^ n17149;
  assign n18048 = n18047 ^ n18046;
  assign n18085 = n18044 ^ n14318;
  assign n18086 = n18085 ^ n14334;
  assign n18087 = n18086 ^ n14309;
  assign n18088 = n18087 ^ n16271;
  assign n18078 = n16229 ^ n14228;
  assign n14450 = n14449 ^ n14263;
  assign n18077 = n17138 ^ n14450;
  assign n18079 = n18078 ^ n18077;
  assign n18062 = n16298 ^ n13856;
  assign n14229 = n14228 ^ n13870;
  assign n18061 = n17112 ^ n14229;
  assign n18063 = n18062 ^ n18061;
  assign n18080 = n18079 ^ n18063;
  assign n18089 = n18088 ^ n18080;
  assign n18124 = ~n18048 & n18089;
  assign n18092 = n18068 ^ n18048;
  assign n18059 = n16190 ^ n14373;
  assign n18057 = n14352 ^ n14345;
  assign n18056 = n14433 ^ n14386;
  assign n18058 = n18057 ^ n18056;
  assign n18060 = n18059 ^ n18058;
  assign n18105 = n18079 ^ n18060;
  assign n18053 = n14456 ^ n14438;
  assign n14440 = n14379 ^ n14318;
  assign n18052 = n18051 ^ n14440;
  assign n18054 = n18053 ^ n18052;
  assign n18049 = n15702 ^ n14420;
  assign n18050 = n18049 ^ n18048;
  assign n18055 = n18054 ^ n18050;
  assign n18113 = n18105 ^ n18055;
  assign n18117 = n18092 & n18113;
  assign n18125 = n18124 ^ n18117;
  assign n18122 = n18113 ^ n18092;
  assign n18093 = n18074 ^ n18060;
  assign n18106 = n18105 ^ n18075;
  assign n18107 = n18093 & n18106;
  assign n18064 = n18063 ^ n18060;
  assign n18065 = n18064 ^ n18055;
  assign n18083 = n18065 & n18075;
  assign n18108 = n18107 ^ n18083;
  assign n18123 = n18122 ^ n18108;
  assign n18126 = n18125 ^ n18123;
  assign n18090 = n18089 ^ n18074;
  assign n18115 = n18090 ^ n18075;
  assign n18114 = n18113 ^ n18089;
  assign n18120 = n18115 ^ n18114;
  assign n18116 = n18114 & n18115;
  assign n18118 = n18117 ^ n18116;
  assign n18069 = n18068 ^ n18060;
  assign n18076 = n18075 ^ n18055;
  assign n18081 = n18080 ^ n18076;
  assign n18082 = n18069 & n18081;
  assign n18084 = n18083 ^ n18082;
  assign n18119 = n18118 ^ n18084;
  assign n18121 = n18120 ^ n18119;
  assign n18131 = n18126 ^ n18121;
  assign n18109 = n18076 ^ n18064;
  assign n18110 = n18109 ^ n18108;
  assign n18100 = n18088 ^ n18076;
  assign n18101 = n18089 ^ n18048;
  assign n18102 = n18101 ^ n18069;
  assign n18103 = n18100 & n18102;
  assign n18094 = n18093 ^ n18092;
  assign n18095 = n18076 & n18094;
  assign n18104 = n18103 ^ n18095;
  assign n18111 = n18110 ^ n18104;
  assign n18127 = n18111 & n18126;
  assign n18097 = n18081 ^ n18069;
  assign n18091 = n18088 & n18090;
  assign n18096 = n18095 ^ n18091;
  assign n18098 = n18097 ^ n18096;
  assign n18099 = n18098 ^ n18084;
  assign n18132 = n18127 ^ n18099;
  assign n18133 = n18131 & n18132;
  assign n18134 = n18133 ^ n18121;
  assign n18112 = n18111 ^ n18099;
  assign n18128 = n18127 ^ n18121;
  assign n18129 = n18112 & n18128;
  assign n18130 = n18129 ^ n18099;
  assign n18135 = n18134 ^ n18130;
  assign n18158 = n18075 & n18135;
  assign n18143 = n18127 ^ n18112;
  assign n18141 = ~n18099 & n18111;
  assign n18142 = n18121 & n18141;
  assign n18144 = n18143 ^ n18142;
  assign n18139 = n18131 ^ n18127;
  assign n18137 = n18099 & n18126;
  assign n18138 = ~n18121 & n18137;
  assign n18140 = n18139 ^ n18138;
  assign n18145 = n18144 ^ n18140;
  assign n18146 = n18145 ^ n18135;
  assign n18157 = n18093 & n18146;
  assign n18159 = n18158 ^ n18157;
  assign n18156 = n18102 & n18140;
  assign n18160 = n18159 ^ n18156;
  assign n18149 = n18140 ^ n18134;
  assign n18153 = n18076 & n18149;
  assign n18151 = n18100 & n18140;
  assign n18150 = n18094 & n18149;
  assign n18152 = n18151 ^ n18150;
  assign n18154 = n18153 ^ n18152;
  assign n18147 = n18106 & n18146;
  assign n18136 = n18065 & n18135;
  assign n18148 = n18147 ^ n18136;
  assign n18155 = n18154 ^ n18148;
  assign n18161 = n18160 ^ n18155;
  assign n18619 = n18618 ^ n18161;
  assign n17836 = n16979 ^ n15381;
  assign n17835 = n17369 ^ n15199;
  assign n17837 = n17836 ^ n17835;
  assign n17833 = n16996 ^ n15358;
  assign n17832 = n17360 ^ n15365;
  assign n17834 = n17833 ^ n17832;
  assign n17838 = n17837 ^ n17834;
  assign n17829 = n17372 ^ n14670;
  assign n15311 = n15310 ^ n15306;
  assign n17828 = n16991 ^ n15311;
  assign n17830 = n17829 ^ n17828;
  assign n17839 = n17838 ^ n17830;
  assign n17843 = n17358 ^ n15243;
  assign n15397 = n15396 ^ n15391;
  assign n17842 = n16961 ^ n15397;
  assign n17844 = n17843 ^ n17842;
  assign n17855 = n17844 ^ n17837;
  assign n17824 = n17363 ^ n15275;
  assign n15264 = n15263 ^ n14901;
  assign n17823 = n17822 ^ n15264;
  assign n17825 = n17824 ^ n17823;
  assign n17819 = n17365 ^ n15402;
  assign n14912 = n14911 ^ n14901;
  assign n17817 = n17816 ^ n14912;
  assign n17818 = n17817 ^ n15160;
  assign n17820 = n17819 ^ n17818;
  assign n15232 = n15231 ^ n15224;
  assign n17821 = n17820 ^ n15232;
  assign n17826 = n17825 ^ n17821;
  assign n17813 = n17376 ^ n15325;
  assign n15286 = n15268 ^ n14901;
  assign n17811 = n17810 ^ n15286;
  assign n17812 = n17811 ^ n15298;
  assign n17814 = n17813 ^ n17812;
  assign n17808 = n17379 ^ n14680;
  assign n15185 = n15184 ^ n15173;
  assign n17807 = n17011 ^ n15185;
  assign n17809 = n17808 ^ n17807;
  assign n17815 = n17814 ^ n17809;
  assign n17827 = n17826 ^ n17815;
  assign n17884 = n17855 ^ n17827;
  assign n17862 = n17844 ^ n17814;
  assign n17845 = n17844 ^ n17834;
  assign n17863 = n17845 ^ n17815;
  assign n17864 = ~n17862 & n17863;
  assign n17856 = n17855 ^ n17826;
  assign n17857 = ~n17815 & n17856;
  assign n17865 = n17864 ^ n17857;
  assign n17885 = n17884 ^ n17865;
  assign n17831 = n17830 ^ n17827;
  assign n17880 = n17839 ^ n17820;
  assign n17852 = n17844 ^ n17809;
  assign n17881 = n17880 ^ n17852;
  assign n17882 = n17831 & ~n17881;
  assign n17849 = n17820 ^ n17809;
  assign n17872 = n17862 ^ n17849;
  assign n17873 = n17827 & n17872;
  assign n17883 = n17882 ^ n17873;
  assign n17886 = n17885 ^ n17883;
  assign n17853 = n17838 ^ n17827;
  assign n17875 = n17853 ^ n17852;
  assign n17840 = n17839 ^ n17814;
  assign n17871 = n17830 & ~n17840;
  assign n17874 = n17873 ^ n17871;
  assign n17876 = n17875 ^ n17874;
  assign n17854 = n17852 & n17853;
  assign n17858 = n17857 ^ n17854;
  assign n17877 = n17876 ^ n17858;
  assign n17900 = n17886 ^ n17877;
  assign n17868 = n17820 & n17839;
  assign n17846 = n17845 ^ n17826;
  assign n17850 = n17846 & ~n17849;
  assign n17869 = n17868 ^ n17850;
  assign n17866 = n17849 ^ n17846;
  assign n17867 = n17866 ^ n17865;
  assign n17870 = n17869 ^ n17867;
  assign n17887 = ~n17870 & ~n17886;
  assign n17908 = n17900 ^ n17887;
  assign n17847 = n17846 ^ n17839;
  assign n17841 = n17840 ^ n17815;
  assign n17860 = n17847 ^ n17841;
  assign n17848 = n17841 & n17847;
  assign n17851 = n17850 ^ n17848;
  assign n17859 = n17858 ^ n17851;
  assign n17861 = n17860 ^ n17859;
  assign n17906 = ~n17877 & ~n17886;
  assign n17907 = n17861 & n17906;
  assign n17909 = n17908 ^ n17907;
  assign n18510 = n17839 & ~n17909;
  assign n17888 = n17870 ^ n17861;
  assign n17889 = n17888 ^ n17887;
  assign n17878 = ~n17870 & n17877;
  assign n17879 = ~n17861 & n17878;
  assign n17890 = n17889 ^ n17879;
  assign n17918 = ~n17881 & ~n17890;
  assign n18511 = n18510 ^ n17918;
  assign n17910 = n17909 ^ n17890;
  assign n17901 = n17887 ^ n17861;
  assign n17902 = ~n17900 & n17901;
  assign n17903 = n17902 ^ n17877;
  assign n17892 = n17887 ^ n17877;
  assign n17893 = ~n17888 & n17892;
  assign n17894 = n17893 ^ n17861;
  assign n17904 = n17903 ^ n17894;
  assign n17911 = n17910 ^ n17904;
  assign n17912 = n17863 & n17911;
  assign n17905 = n17856 & n17904;
  assign n17913 = n17912 ^ n17905;
  assign n18614 = n18511 ^ n17913;
  assign n18419 = n17909 ^ n17903;
  assign n18471 = n17846 & ~n18419;
  assign n17916 = ~n17815 & n17904;
  assign n17915 = ~n17862 & n17911;
  assign n17917 = n17916 ^ n17915;
  assign n18472 = n18471 ^ n17917;
  assign n17895 = n17894 ^ n17890;
  assign n17896 = n17872 & ~n17895;
  assign n18613 = n18472 ^ n17896;
  assign n18615 = n18614 ^ n18613;
  assign n18620 = n18619 ^ n18615;
  assign n18405 = n18089 & n18144;
  assign n18406 = n18405 ^ n18156;
  assign n18468 = n18406 ^ n18148;
  assign n18292 = n18144 ^ n18130;
  assign n18408 = n18113 & n18292;
  assign n18409 = n18408 ^ n18159;
  assign n18467 = n18409 ^ n18150;
  assign n18469 = n18468 ^ n18467;
  assign n18621 = n18620 ^ n18469;
  assign n18634 = n18633 ^ n18621;
  assign n18463 = n18114 & n18130;
  assign n18286 = n18088 & n18134;
  assign n18526 = n18463 ^ n18286;
  assign n18527 = n18526 ^ n18152;
  assign n18525 = n18406 ^ n18159;
  assign n18528 = n18527 ^ n18525;
  assign n18529 = n18528 ^ n18469;
  assign n18021 = n17944 & n18018;
  assign n18014 = n17949 & n18013;
  assign n18020 = n18019 ^ n18014;
  assign n18022 = n18021 ^ n18020;
  assign n18522 = n18521 ^ n18022;
  assign n18523 = n18522 ^ n18487;
  assign n18407 = n18406 ^ n18154;
  assign n18410 = n18409 ^ n18407;
  assign n18524 = n18523 ^ n18410;
  assign n18530 = n18529 ^ n18524;
  assign n18515 = n18196 & n18265;
  assign n18254 = n18167 & n18253;
  assign n18516 = n18515 ^ n18254;
  assign n18517 = n18516 ^ n18396;
  assign n18392 = n18195 & n18276;
  assign n18393 = n18392 ^ n18391;
  assign n18514 = n18402 ^ n18393;
  assign n18518 = n18517 ^ n18514;
  assign n18482 = n18481 ^ n18393;
  assign n18279 = n18276 ^ n18265;
  assign n18399 = n18189 & n18279;
  assign n18403 = n18402 ^ n18399;
  assign n18479 = n18403 ^ n18394;
  assign n18483 = n18482 ^ n18479;
  assign n18519 = n18518 ^ n18483;
  assign n18531 = n18530 ^ n18519;
  assign n17898 = n17827 & ~n17895;
  assign n17891 = n17831 & ~n17890;
  assign n17897 = n17896 ^ n17891;
  assign n17899 = n17898 ^ n17897;
  assign n18512 = n18511 ^ n17899;
  assign n18513 = n18512 ^ n18472;
  assign n18532 = n18531 ^ n18513;
  assign n18542 = n18541 ^ n18532;
  assign n18635 = n18634 ^ n18542;
  assign n18605 = n18090 & n18134;
  assign n18606 = n18605 ^ n18406;
  assign n18288 = n18115 & n18130;
  assign n18287 = n18286 ^ n18153;
  assign n18289 = n18288 ^ n18287;
  assign n18607 = n18606 ^ n18289;
  assign n18294 = n18081 & n18145;
  assign n18293 = n18092 & n18292;
  assign n18295 = n18294 ^ n18293;
  assign n18556 = n18295 ^ n18147;
  assign n18604 = n18556 ^ n18409;
  assign n18608 = n18607 ^ n18604;
  assign n18609 = n18608 ^ n18469;
  assign n18610 = n18609 ^ n18528;
  assign n18598 = n18203 & n18253;
  assign n18599 = n18598 ^ n18393;
  assign n18266 = n18209 & n18265;
  assign n18261 = n18260 ^ n18254;
  assign n18267 = n18266 ^ n18261;
  assign n18600 = n18599 ^ n18267;
  assign n18281 = n18216 & n18277;
  assign n18280 = n18211 & n18279;
  assign n18282 = n18281 ^ n18280;
  assign n18596 = n18480 ^ n18282;
  assign n18597 = n18596 ^ n18403;
  assign n18601 = n18600 ^ n18597;
  assign n18602 = n18601 ^ n18483;
  assign n18475 = n17847 & n17903;
  assign n18413 = n17830 & n17894;
  assign n18593 = n18475 ^ n18413;
  assign n18594 = n18593 ^ n17897;
  assign n18592 = n18511 ^ n17917;
  assign n18595 = n18594 ^ n18592;
  assign n18603 = n18602 ^ n18595;
  assign n18611 = n18610 ^ n18603;
  assign n18489 = n17977 & n18026;
  assign n18426 = n17948 & n18017;
  assign n18578 = n18489 ^ n18426;
  assign n18579 = n18578 ^ n18020;
  assign n18577 = n18521 ^ n18040;
  assign n18580 = n18579 ^ n18577;
  assign n18590 = n18589 ^ n18580;
  assign n18564 = n18520 ^ n18040;
  assign n18434 = n17968 & n18033;
  assign n18433 = n17974 & n18432;
  assign n18435 = n18434 ^ n18433;
  assign n18562 = n18435 ^ n18035;
  assign n18490 = n18003 & n18032;
  assign n18491 = n18490 ^ n18489;
  assign n18563 = n18562 ^ n18491;
  assign n18565 = n18564 ^ n18563;
  assign n18575 = n18574 ^ n18565;
  assign n18558 = n18405 ^ n18159;
  assign n18462 = n18101 & n18144;
  assign n18464 = n18463 ^ n18462;
  assign n18557 = n18556 ^ n18464;
  assign n18559 = n18558 ^ n18557;
  assign n18465 = n18464 ^ n18287;
  assign n18461 = n18409 ^ n18293;
  assign n18466 = n18465 ^ n18461;
  assign n18470 = n18469 ^ n18466;
  assign n18560 = n18559 ^ n18470;
  assign n18550 = n18243 & n18276;
  assign n18551 = n18550 ^ n18515;
  assign n18552 = n18551 ^ n18261;
  assign n18549 = n18403 ^ n18280;
  assign n18553 = n18552 ^ n18549;
  assign n18554 = n18553 ^ n18483;
  assign n18547 = n18510 ^ n17917;
  assign n18421 = n17853 & n17910;
  assign n18420 = ~n17849 & ~n18419;
  assign n18422 = n18421 ^ n18420;
  assign n18545 = n18422 ^ n17912;
  assign n18474 = ~n17880 & ~n17909;
  assign n18476 = n18475 ^ n18474;
  assign n18546 = n18545 ^ n18476;
  assign n18548 = n18547 ^ n18546;
  assign n18555 = n18554 ^ n18548;
  assign n18561 = n18560 ^ n18555;
  assign n18576 = n18575 ^ n18561;
  assign n18591 = n18590 ^ n18576;
  assign n18612 = n18611 ^ n18591;
  assign n18636 = n18635 ^ n18612;
  assign n18648 = n18402 ^ n18392;
  assign n18647 = n18596 ^ n18551;
  assign n18649 = n18648 ^ n18647;
  assign n18650 = n18649 ^ n18559;
  assign n18643 = n17978 & n18017;
  assign n18644 = n18643 ^ n18521;
  assign n18428 = n17979 & n18026;
  assign n18427 = n18426 ^ n18021;
  assign n18429 = n18428 ^ n18427;
  assign n18645 = n18644 ^ n18429;
  assign n18642 = n18562 ^ n18487;
  assign n18646 = n18645 ^ n18642;
  assign n18651 = n18650 ^ n18646;
  assign n18652 = n18651 ^ n18608;
  assign n18638 = ~n17840 & n17894;
  assign n18639 = n18638 ^ n18511;
  assign n18415 = n17841 & n17903;
  assign n18414 = n18413 ^ n17898;
  assign n18416 = n18415 ^ n18414;
  assign n18640 = n18639 ^ n18416;
  assign n18637 = n18545 ^ n18472;
  assign n18641 = n18640 ^ n18637;
  assign n18653 = n18652 ^ n18641;
  assign n18664 = n18663 ^ n18653;
  assign n18431 = n17969 & n18033;
  assign n18436 = n18435 ^ n18431;
  assign n18425 = n18039 ^ n18028;
  assign n18430 = n18429 ^ n18425;
  assign n18437 = n18436 ^ n18430;
  assign n18291 = n18069 & n18145;
  assign n18296 = n18295 ^ n18291;
  assign n18285 = n18158 ^ n18136;
  assign n18290 = n18289 ^ n18285;
  assign n18297 = n18296 ^ n18290;
  assign n18438 = n18437 ^ n18297;
  assign n18418 = n17852 & n17910;
  assign n18423 = n18422 ^ n18418;
  assign n18412 = n17916 ^ n17905;
  assign n18417 = n18416 ^ n18412;
  assign n18424 = n18423 ^ n18417;
  assign n18439 = n18438 ^ n18424;
  assign n18398 = n18397 ^ n18393;
  assign n18404 = n18403 ^ n18398;
  assign n18411 = n18410 ^ n18404;
  assign n18440 = n18439 ^ n18411;
  assign n18459 = n18458 ^ n18440;
  assign n18686 = n18664 ^ n18459;
  assign n18693 = n18686 ^ n18612;
  assign n18492 = n18491 ^ n18427;
  assign n18488 = n18487 ^ n18433;
  assign n18493 = n18492 ^ n18488;
  assign n18507 = n18506 ^ n18493;
  assign n18477 = n18476 ^ n18414;
  assign n18473 = n18472 ^ n18420;
  assign n18478 = n18477 ^ n18473;
  assign n18484 = n18483 ^ n18478;
  assign n18485 = n18484 ^ n18470;
  assign n18508 = n18507 ^ n18485;
  assign n18278 = n18214 & n18277;
  assign n18283 = n18282 ^ n18278;
  assign n18271 = n18270 ^ n18269;
  assign n18272 = n18271 ^ n18267;
  assign n18284 = n18283 ^ n18272;
  assign n18298 = n18297 ^ n18284;
  assign n18042 = n18041 ^ n18040;
  assign n18037 = n18036 ^ n18022;
  assign n18043 = n18042 ^ n18037;
  assign n18162 = n18161 ^ n18043;
  assign n18299 = n18298 ^ n18162;
  assign n17919 = n17918 ^ n17917;
  assign n17914 = n17913 ^ n17899;
  assign n17920 = n17919 ^ n17914;
  assign n18300 = n18299 ^ n17920;
  assign n18390 = n18389 ^ n18300;
  assign n18460 = n18459 ^ n18390;
  assign n18509 = n18508 ^ n18460;
  assign n18703 = n18693 ^ n18509;
  assign n18543 = n18542 ^ n18509;
  assign n18702 = n18635 ^ n18543;
  assign n18707 = n18703 ^ n18702;
  assign n18704 = ~n18702 & ~n18703;
  assign n18666 = n18634 ^ n18576;
  assign n18697 = ~n18666 & n18693;
  assign n18705 = n18704 ^ n18697;
  assign n18675 = n18664 ^ n18390;
  assign n18676 = n18675 ^ n18612;
  assign n18677 = n18635 & n18676;
  assign n18670 = n18636 ^ n18460;
  assign n18671 = n18664 ^ n18634;
  assign n18674 = ~n18670 & n18671;
  assign n18678 = n18677 ^ n18674;
  assign n18706 = n18705 ^ n18678;
  assign n18708 = n18707 ^ n18706;
  assign n18696 = ~n18509 & n18576;
  assign n18698 = n18697 ^ n18696;
  assign n18694 = n18693 ^ n18666;
  assign n18665 = n18664 ^ n18542;
  assign n18687 = n18686 ^ n18635;
  assign n18688 = n18665 & ~n18687;
  assign n18689 = n18688 ^ n18677;
  assign n18695 = n18694 ^ n18689;
  assign n18699 = n18698 ^ n18695;
  assign n18713 = n18708 ^ n18699;
  assign n18685 = n18675 ^ n18636;
  assign n18690 = n18689 ^ n18685;
  assign n18680 = n18576 ^ n18509;
  assign n18681 = n18680 ^ n18671;
  assign n18682 = n18636 ^ n18508;
  assign n18683 = n18681 & n18682;
  assign n18667 = n18666 ^ n18665;
  assign n18668 = ~n18636 & ~n18667;
  assign n18684 = n18683 ^ n18668;
  assign n18691 = n18690 ^ n18684;
  assign n18700 = n18691 & ~n18699;
  assign n18723 = n18713 ^ n18700;
  assign n18672 = n18671 ^ n18670;
  assign n18544 = ~n18508 & ~n18543;
  assign n18669 = n18668 ^ n18544;
  assign n18673 = n18672 ^ n18669;
  assign n18679 = n18678 ^ n18673;
  assign n18721 = ~n18679 & ~n18699;
  assign n18722 = ~n18708 & n18721;
  assign n18724 = n18723 ^ n18722;
  assign n18714 = n18700 ^ n18679;
  assign n18715 = ~n18713 & ~n18714;
  assign n18716 = n18715 ^ n18708;
  assign n19807 = n18724 ^ n18716;
  assign n19832 = ~n18636 & ~n19807;
  assign n19809 = n18682 & ~n18724;
  assign n19808 = ~n18667 & ~n19807;
  assign n19810 = n19809 ^ n19808;
  assign n19923 = n19832 ^ n19810;
  assign n19802 = n18681 & ~n18724;
  assign n18709 = n18679 & n18691;
  assign n18710 = n18708 & n18709;
  assign n18692 = n18691 ^ n18679;
  assign n18701 = n18700 ^ n18692;
  assign n18711 = n18710 ^ n18701;
  assign n18712 = ~n18509 & ~n18711;
  assign n19803 = n19802 ^ n18712;
  assign n19924 = n19923 ^ n19803;
  assign n18717 = n18708 ^ n18700;
  assign n18718 = ~n18692 & n18717;
  assign n18719 = n18718 ^ n18679;
  assign n18733 = n18719 ^ n18711;
  assign n19827 = n18693 & n18733;
  assign n18720 = n18719 ^ n18716;
  assign n18728 = n18635 & ~n18720;
  assign n18725 = n18724 ^ n18711;
  assign n18726 = n18725 ^ n18720;
  assign n18727 = n18665 & ~n18726;
  assign n18729 = n18728 ^ n18727;
  assign n19828 = n19827 ^ n18729;
  assign n19925 = n19924 ^ n19828;
  assign n15374 = n15342 ^ n15191;
  assign n15382 = n15381 ^ n15374;
  assign n15373 = n15372 ^ n15365;
  assign n15383 = n15382 ^ n15373;
  assign n15343 = n15342 ^ n15288;
  assign n15359 = n15358 ^ n15343;
  assign n15337 = n15336 ^ n15325;
  assign n15360 = n15359 ^ n15337;
  assign n15384 = n15383 ^ n15360;
  assign n15321 = n15320 ^ n14680;
  assign n15312 = n15311 ^ n14912;
  assign n15322 = n15321 ^ n15312;
  assign n15385 = n15384 ^ n15322;
  assign n15412 = n15411 ^ n15402;
  assign n15398 = n15263 ^ n14918;
  assign n15399 = n15398 ^ n15397;
  assign n15413 = n15412 ^ n15399;
  assign n15421 = n15413 ^ n15360;
  assign n15269 = n15268 ^ n15264;
  assign n15256 = n15255 ^ n15244;
  assign n15270 = n15269 ^ n15256;
  assign n14919 = n14918 ^ n14912;
  assign n15161 = n15160 ^ n14919;
  assign n14786 = n14785 ^ n14681;
  assign n15162 = n15161 ^ n14786;
  assign n15233 = n15232 ^ n15162;
  assign n15271 = n15270 ^ n15233;
  assign n15441 = n15421 ^ n15271;
  assign n15450 = n15441 ^ n15385;
  assign n15289 = n15288 ^ n15286;
  assign n15299 = n15298 ^ n15289;
  assign n15285 = n15284 ^ n15276;
  assign n15300 = n15299 ^ n15285;
  assign n15431 = n15385 ^ n15300;
  assign n15215 = n15214 ^ n15199;
  assign n15192 = n15191 ^ n14901;
  assign n15193 = n15192 ^ n15185;
  assign n15216 = n15215 ^ n15193;
  assign n15301 = n15300 ^ n15216;
  assign n15449 = n15431 ^ n15301;
  assign n15454 = n15450 ^ n15449;
  assign n15451 = ~n15449 & ~n15450;
  assign n15217 = n15216 ^ n15162;
  assign n15445 = ~n15217 & n15441;
  assign n15452 = n15451 ^ n15445;
  assign n15414 = n15413 ^ n15216;
  assign n15302 = n15301 ^ n15271;
  assign n15434 = n15384 ^ n15302;
  assign n15437 = n15414 & ~n15434;
  assign n15424 = n15413 ^ n15383;
  assign n15425 = n15424 ^ n15271;
  assign n15426 = n15301 & n15425;
  assign n15438 = n15437 ^ n15426;
  assign n15453 = n15452 ^ n15438;
  assign n15455 = n15454 ^ n15453;
  assign n15428 = n15424 ^ n15302;
  assign n15417 = n15413 ^ n15300;
  assign n15422 = n15421 ^ n15301;
  assign n15423 = n15417 & ~n15422;
  assign n15427 = n15426 ^ n15423;
  assign n15429 = n15428 ^ n15427;
  assign n15418 = n15417 ^ n15217;
  assign n15419 = ~n15302 & ~n15418;
  assign n15323 = n15322 ^ n15302;
  assign n15386 = n15385 ^ n15162;
  assign n15415 = n15414 ^ n15386;
  assign n15416 = n15323 & n15415;
  assign n15420 = n15419 ^ n15416;
  assign n15430 = n15429 ^ n15420;
  assign n15435 = n15434 ^ n15414;
  assign n15432 = ~n15322 & ~n15431;
  assign n15433 = n15432 ^ n15419;
  assign n15436 = n15435 ^ n15433;
  assign n15439 = n15438 ^ n15436;
  assign n15460 = n15430 & n15439;
  assign n15461 = n15455 & n15460;
  assign n15444 = n15162 & ~n15385;
  assign n15446 = n15445 ^ n15444;
  assign n15442 = n15441 ^ n15217;
  assign n15443 = n15442 ^ n15427;
  assign n15447 = n15446 ^ n15443;
  assign n15448 = n15430 & ~n15447;
  assign n15440 = n15439 ^ n15430;
  assign n15459 = n15448 ^ n15440;
  assign n15462 = n15461 ^ n15459;
  assign n15497 = ~n15385 & ~n15462;
  assign n15465 = n15455 ^ n15447;
  assign n15473 = n15465 ^ n15448;
  assign n15471 = ~n15439 & ~n15447;
  assign n15472 = ~n15455 & n15471;
  assign n15474 = n15473 ^ n15472;
  assign n15496 = n15415 & ~n15474;
  assign n15498 = n15497 ^ n15496;
  assign n15475 = n15474 ^ n15462;
  assign n15466 = n15448 ^ n15439;
  assign n15467 = ~n15465 & ~n15466;
  assign n15468 = n15467 ^ n15455;
  assign n15456 = n15455 ^ n15448;
  assign n15457 = ~n15440 & n15456;
  assign n15458 = n15457 ^ n15439;
  assign n15469 = n15468 ^ n15458;
  assign n15476 = n15475 ^ n15469;
  assign n15494 = ~n15422 & ~n15476;
  assign n15493 = n15425 & ~n15469;
  assign n15495 = n15494 ^ n15493;
  assign n15499 = n15498 ^ n15495;
  assign n15486 = n15474 ^ n15468;
  assign n15491 = ~n15418 & ~n15486;
  assign n15463 = n15462 ^ n15458;
  assign n15479 = n15441 & n15463;
  assign n15477 = n15417 & ~n15476;
  assign n15470 = n15301 & ~n15469;
  assign n15478 = n15477 ^ n15470;
  assign n15480 = n15479 ^ n15478;
  assign n15492 = n15491 ^ n15480;
  assign n15500 = n15499 ^ n15492;
  assign n16738 = n16737 ^ n15500;
  assign n16300 = n16299 ^ n16292;
  assign n16289 = n16288 ^ n16282;
  assign n16301 = n16300 ^ n16289;
  assign n16231 = n16230 ^ n16221;
  assign n16216 = n16215 ^ n16206;
  assign n16232 = n16231 ^ n16216;
  assign n16302 = n16301 ^ n16232;
  assign n16258 = n15849 ^ n15722;
  assign n16262 = n16261 ^ n16258;
  assign n16266 = n16265 ^ n16262;
  assign n16273 = n16272 ^ n16266;
  assign n16303 = n16302 ^ n16273;
  assign n16102 = n16101 ^ n16087;
  assign n15851 = n15850 ^ n15722;
  assign n16081 = n16080 ^ n15851;
  assign n16103 = n16102 ^ n16081;
  assign n16346 = n16303 ^ n16103;
  assign n16323 = n16322 ^ n15713;
  assign n16316 = n16315 ^ n16311;
  assign n16324 = n16323 ^ n16316;
  assign n16192 = n16191 ^ n16111;
  assign n16176 = n16175 ^ n16164;
  assign n16153 = n16152 ^ n16087;
  assign n16177 = n16176 ^ n16153;
  assign n16193 = n16192 ^ n16177;
  assign n16332 = n16324 ^ n16193;
  assign n16347 = n16346 ^ n16332;
  assign n16367 = ~n16103 & n16303;
  assign n16233 = n16232 ^ n16193;
  assign n16147 = n16146 ^ n16135;
  assign n16124 = n16123 ^ n16112;
  assign n16148 = n16147 ^ n16124;
  assign n15704 = n15703 ^ n15616;
  assign n16104 = n16103 ^ n15704;
  assign n16149 = n16148 ^ n16104;
  assign n16234 = n16233 ^ n16149;
  assign n16329 = n16324 ^ n16103;
  assign n16330 = n16234 & n16329;
  assign n16368 = n16367 ^ n16330;
  assign n16365 = n16329 ^ n16234;
  assign n16256 = n16255 ^ n16209;
  assign n16241 = n16240 ^ n16235;
  assign n16249 = n16248 ^ n16241;
  assign n16257 = n16256 ^ n16249;
  assign n16343 = n16257 ^ n16193;
  assign n16325 = n16324 ^ n16257;
  assign n16352 = n16325 ^ n16233;
  assign n16353 = n16343 & n16352;
  assign n16336 = n16301 ^ n16193;
  assign n16337 = n16336 ^ n16149;
  assign n16338 = n16325 & n16337;
  assign n16354 = n16353 ^ n16338;
  assign n16366 = n16365 ^ n16354;
  assign n16369 = n16368 ^ n16366;
  assign n16327 = n16303 ^ n16234;
  assign n16304 = n16303 ^ n16257;
  assign n16326 = n16325 ^ n16304;
  assign n16341 = n16327 ^ n16326;
  assign n16333 = n16325 ^ n16149;
  assign n16334 = n16333 ^ n16302;
  assign n16335 = n16332 & n16334;
  assign n16339 = n16338 ^ n16335;
  assign n16328 = n16326 & n16327;
  assign n16331 = n16330 ^ n16328;
  assign n16340 = n16339 ^ n16331;
  assign n16342 = n16341 ^ n16340;
  assign n16380 = n16369 ^ n16342;
  assign n16351 = n16336 ^ n16333;
  assign n16355 = n16354 ^ n16351;
  assign n16348 = n16333 ^ n16273;
  assign n16349 = n16347 & n16348;
  assign n16344 = n16343 ^ n16329;
  assign n16345 = n16333 & n16344;
  assign n16350 = n16349 ^ n16345;
  assign n16356 = n16355 ^ n16350;
  assign n16370 = n16356 & n16369;
  assign n16381 = n16380 ^ n16370;
  assign n16359 = n16334 ^ n16332;
  assign n16357 = n16273 & n16304;
  assign n16358 = n16357 ^ n16345;
  assign n16360 = n16359 ^ n16358;
  assign n16361 = n16360 ^ n16339;
  assign n16378 = n16361 & n16369;
  assign n16379 = ~n16342 & n16378;
  assign n16382 = n16381 ^ n16379;
  assign n16407 = n16347 & n16382;
  assign n16384 = n16370 ^ n16361;
  assign n16385 = n16380 & n16384;
  assign n16386 = n16385 ^ n16342;
  assign n16364 = n16361 ^ n16356;
  assign n16373 = n16370 ^ n16342;
  assign n16374 = n16364 & n16373;
  assign n16375 = n16374 ^ n16361;
  assign n16387 = n16386 ^ n16375;
  assign n16390 = n16325 & n16387;
  assign n16371 = n16370 ^ n16364;
  assign n16362 = n16356 & ~n16361;
  assign n16363 = n16342 & n16362;
  assign n16372 = n16371 ^ n16363;
  assign n16383 = n16382 ^ n16372;
  assign n16388 = n16387 ^ n16383;
  assign n16389 = n16343 & n16388;
  assign n16391 = n16390 ^ n16389;
  assign n16730 = n16407 ^ n16391;
  assign n16596 = n16348 & n16382;
  assign n16396 = n16386 ^ n16382;
  assign n16404 = n16344 & n16396;
  assign n16597 = n16596 ^ n16404;
  assign n16397 = n16333 & n16396;
  assign n16598 = n16597 ^ n16397;
  assign n16410 = n16337 & n16387;
  assign n16409 = n16352 & n16388;
  assign n16411 = n16410 ^ n16409;
  assign n16729 = n16598 ^ n16411;
  assign n16731 = n16730 ^ n16729;
  assign n16709 = n15496 ^ n15478;
  assign n16512 = n15323 & ~n15474;
  assign n16513 = n16512 ^ n15491;
  assign n15487 = ~n15302 & ~n15486;
  assign n16601 = n16513 ^ n15487;
  assign n16708 = n16601 ^ n15495;
  assign n16710 = n16709 ^ n16708;
  assign n16732 = n16731 ^ n16710;
  assign n14374 = n14373 ^ n14367;
  assign n14380 = n14379 ^ n14374;
  assign n14387 = n14386 ^ n14380;
  assign n14396 = n14395 ^ n14387;
  assign n13995 = n13994 ^ n13857;
  assign n14128 = n14127 ^ n13995;
  assign n14215 = n14214 ^ n14128;
  assign n14471 = n14396 ^ n14215;
  assign n14445 = n14444 ^ n14440;
  assign n14439 = n14438 ^ n14434;
  assign n14446 = n14445 ^ n14439;
  assign n14427 = n14426 ^ n14420;
  assign n14360 = n14359 ^ n14352;
  assign n14346 = n14345 ^ n14325;
  assign n14341 = n14340 ^ n14335;
  assign n14347 = n14346 ^ n14341;
  assign n14361 = n14360 ^ n14347;
  assign n14428 = n14427 ^ n14361;
  assign n14447 = n14446 ^ n14428;
  assign n14472 = n14471 ^ n14447;
  assign n14315 = n14314 ^ n14309;
  assign n14326 = n14325 ^ n14315;
  assign n14301 = n14300 ^ n14290;
  assign n14327 = n14326 ^ n14301;
  assign n14243 = n14242 ^ n14229;
  assign n14265 = n14264 ^ n14243;
  assign n14281 = n14280 ^ n14265;
  assign n14282 = n14281 ^ n14215;
  assign n14328 = n14327 ^ n14282;
  assign n14510 = n14328 & ~n14361;
  assign n14475 = n14396 ^ n14281;
  assign n14476 = n14475 ^ n14447;
  assign n14414 = n14413 ^ n14408;
  assign n14404 = n14318 ^ n13738;
  assign n14403 = n14402 ^ n14399;
  assign n14405 = n14404 ^ n14403;
  assign n14415 = n14414 ^ n14405;
  assign n14481 = n14415 ^ n14361;
  assign n14482 = n14476 & n14481;
  assign n14511 = n14510 ^ n14482;
  assign n14508 = n14481 ^ n14476;
  assign n14452 = n14451 ^ n14450;
  assign n14458 = n14457 ^ n14452;
  assign n14461 = n14460 ^ n14458;
  assign n14466 = n14465 ^ n14461;
  assign n14487 = n14466 ^ n14396;
  assign n14467 = n14466 ^ n14415;
  assign n14495 = n14475 ^ n14467;
  assign n14496 = n14487 & n14495;
  assign n14473 = n14467 & n14472;
  assign n14497 = n14496 ^ n14473;
  assign n14509 = n14508 ^ n14497;
  assign n14512 = n14511 ^ n14509;
  assign n14478 = n14466 ^ n14328;
  assign n14479 = n14478 ^ n14467;
  assign n14477 = n14476 ^ n14328;
  assign n14485 = n14479 ^ n14477;
  assign n14480 = n14477 & n14479;
  assign n14483 = n14482 ^ n14480;
  assign n14416 = n14415 ^ n14396;
  assign n14468 = n14467 ^ n14447;
  assign n14469 = n14468 ^ n14282;
  assign n14470 = n14416 & n14469;
  assign n14474 = n14473 ^ n14470;
  assign n14484 = n14483 ^ n14474;
  assign n14486 = n14485 ^ n14484;
  assign n14526 = n14512 ^ n14486;
  assign n14494 = n14471 ^ n14468;
  assign n14498 = n14497 ^ n14494;
  assign n14490 = n14468 ^ n14327;
  assign n14362 = n14361 ^ n14328;
  assign n14491 = n14416 ^ n14362;
  assign n14492 = n14490 & n14491;
  assign n14488 = n14487 ^ n14481;
  assign n14489 = n14468 & n14488;
  assign n14493 = n14492 ^ n14489;
  assign n14499 = n14498 ^ n14493;
  assign n14513 = n14499 & n14512;
  assign n14502 = n14469 ^ n14416;
  assign n14500 = n14327 & n14478;
  assign n14501 = n14500 ^ n14489;
  assign n14503 = n14502 ^ n14501;
  assign n14504 = n14503 ^ n14474;
  assign n14532 = n14513 ^ n14504;
  assign n14533 = n14526 & n14532;
  assign n14534 = n14533 ^ n14486;
  assign n14507 = n14504 ^ n14499;
  assign n14517 = n14513 ^ n14486;
  assign n14518 = n14507 & n14517;
  assign n14519 = n14518 ^ n14504;
  assign n14535 = n14534 ^ n14519;
  assign n16585 = n14472 & n14535;
  assign n14527 = n14526 ^ n14513;
  assign n14524 = n14504 & n14512;
  assign n14525 = ~n14486 & n14524;
  assign n14528 = n14527 ^ n14525;
  assign n14514 = n14513 ^ n14507;
  assign n14505 = n14499 & ~n14504;
  assign n14506 = n14486 & n14505;
  assign n14515 = n14514 ^ n14506;
  assign n14529 = n14528 ^ n14515;
  assign n14536 = n14535 ^ n14529;
  assign n14537 = n14495 & n14536;
  assign n16696 = n16585 ^ n14537;
  assign n16561 = n14491 & n14528;
  assign n14543 = n14328 & n14515;
  assign n16562 = n16561 ^ n14543;
  assign n16726 = n16696 ^ n16562;
  assign n14522 = n14519 ^ n14515;
  assign n16631 = n14476 & n14522;
  assign n14541 = n14467 & n14535;
  assign n14540 = n14487 & n14536;
  assign n14542 = n14541 ^ n14540;
  assign n16632 = n16631 ^ n14542;
  assign n16567 = n14534 ^ n14528;
  assign n16568 = n14488 & n16567;
  assign n16725 = n16632 ^ n16568;
  assign n16727 = n16726 ^ n16725;
  assign n13526 = n13525 ^ n13519;
  assign n13514 = n13513 ^ n13507;
  assign n13527 = n13526 ^ n13514;
  assign n13470 = n13469 ^ n13465;
  assign n13462 = n13461 ^ n13457;
  assign n13471 = n13470 ^ n13462;
  assign n13536 = n13527 ^ n13471;
  assign n13424 = n13423 ^ n13417;
  assign n13412 = n13411 ^ n13400;
  assign n13425 = n13424 ^ n13412;
  assign n13384 = n13383 ^ n13372;
  assign n13344 = n13343 ^ n13335;
  assign n13362 = n13361 ^ n13344;
  assign n13385 = n13384 ^ n13362;
  assign n13392 = n13391 ^ n13385;
  assign n13426 = n13425 ^ n13392;
  assign n13541 = n13536 ^ n13426;
  assign n13499 = n13498 ^ n13490;
  assign n13483 = n13482 ^ n13474;
  assign n13500 = n13499 ^ n13483;
  assign n13501 = n13500 ^ n13471;
  assign n13444 = n13443 ^ n13438;
  assign n13434 = n13433 ^ n13428;
  assign n13445 = n13444 ^ n13434;
  assign n13502 = n13501 ^ n13445;
  assign n13325 = n13324 ^ n13317;
  assign n13301 = n13300 ^ n13285;
  assign n13311 = n13310 ^ n13301;
  assign n13326 = n13325 ^ n13311;
  assign n13546 = n13502 ^ n13326;
  assign n13277 = n13276 ^ n13174;
  assign n12258 = n12257 ^ n11318;
  assign n13278 = n13277 ^ n12258;
  assign n13327 = n13326 ^ n13278;
  assign n13565 = n13546 ^ n13327;
  assign n13538 = n13527 ^ n13500;
  assign n13556 = n13538 ^ n13426;
  assign n13564 = n13556 ^ n13502;
  assign n13569 = n13565 ^ n13564;
  assign n13566 = n13564 & ~n13565;
  assign n13532 = n13385 ^ n13278;
  assign n13560 = ~n13532 & ~n13556;
  assign n13567 = n13566 ^ n13560;
  assign n13528 = n13527 ^ n13278;
  assign n13427 = n13426 ^ n13327;
  assign n13549 = n13501 ^ n13427;
  assign n13552 = ~n13528 & ~n13549;
  assign n13542 = ~n13327 & ~n13541;
  assign n13553 = n13552 ^ n13542;
  assign n13568 = n13567 ^ n13553;
  assign n13570 = n13569 ^ n13568;
  assign n13559 = n13385 & ~n13502;
  assign n13561 = n13560 ^ n13559;
  assign n13557 = n13556 ^ n13532;
  assign n13531 = n13527 ^ n13326;
  assign n13539 = n13538 ^ n13327;
  assign n13540 = n13531 & n13539;
  assign n13543 = n13542 ^ n13540;
  assign n13558 = n13557 ^ n13543;
  assign n13562 = n13561 ^ n13558;
  assign n13574 = n13570 ^ n13562;
  assign n13537 = n13536 ^ n13427;
  assign n13544 = n13543 ^ n13537;
  assign n13533 = n13532 ^ n13531;
  assign n13534 = ~n13427 & ~n13533;
  assign n13446 = n13445 ^ n13427;
  assign n13503 = n13502 ^ n13385;
  assign n13529 = n13528 ^ n13503;
  assign n13530 = n13446 & ~n13529;
  assign n13535 = n13534 ^ n13530;
  assign n13545 = n13544 ^ n13535;
  assign n13563 = n13545 & n13562;
  assign n13550 = n13549 ^ n13528;
  assign n13547 = ~n13445 & n13546;
  assign n13548 = n13547 ^ n13534;
  assign n13551 = n13550 ^ n13548;
  assign n13554 = n13553 ^ n13551;
  assign n13575 = n13563 ^ n13554;
  assign n13576 = ~n13574 & n13575;
  assign n13577 = n13576 ^ n13570;
  assign n13555 = n13554 ^ n13545;
  assign n13571 = n13570 ^ n13563;
  assign n13572 = n13555 & ~n13571;
  assign n13573 = n13572 ^ n13554;
  assign n13578 = n13577 ^ n13573;
  assign n16575 = ~n13541 & ~n13578;
  assign n13585 = n13554 & n13562;
  assign n13586 = n13570 & n13585;
  assign n13584 = n13574 ^ n13563;
  assign n13587 = n13586 ^ n13584;
  assign n13582 = n13563 ^ n13555;
  assign n13580 = n13545 & ~n13554;
  assign n13581 = ~n13570 & n13580;
  assign n13583 = n13582 ^ n13581;
  assign n13588 = n13587 ^ n13583;
  assign n13589 = n13588 ^ n13578;
  assign n13601 = n13539 & n13589;
  assign n16692 = n16575 ^ n13601;
  assign n16550 = ~n13529 & ~n13587;
  assign n13592 = ~n13502 & n13583;
  assign n16551 = n16550 ^ n13592;
  assign n16723 = n16692 ^ n16551;
  assign n13597 = n13583 ^ n13573;
  assign n16624 = ~n13556 & n13597;
  assign n13590 = n13531 & n13589;
  assign n13579 = ~n13327 & ~n13578;
  assign n13591 = n13590 ^ n13579;
  assign n16625 = n16624 ^ n13591;
  assign n16556 = n13587 ^ n13577;
  assign n16557 = ~n13533 & n16556;
  assign n16722 = n16625 ^ n16557;
  assign n16724 = n16723 ^ n16722;
  assign n16728 = n16727 ^ n16724;
  assign n16733 = n16732 ^ n16728;
  assign n16739 = n16738 ^ n16733;
  assign n16602 = n16601 ^ n15498;
  assign n16603 = n16602 ^ n15480;
  assign n16690 = n16689 ^ n16603;
  assign n16400 = n16327 & n16375;
  assign n16395 = n16273 & n16386;
  assign n16680 = n16400 ^ n16395;
  assign n16681 = n16680 ^ n16597;
  assign n16406 = n16303 & n16372;
  assign n16408 = n16407 ^ n16406;
  assign n16679 = n16408 ^ n16391;
  assign n16682 = n16681 ^ n16679;
  assign n16412 = n16411 ^ n16408;
  assign n16376 = n16375 ^ n16372;
  assign n16377 = n16234 & n16376;
  assign n16392 = n16391 ^ n16377;
  assign n16405 = n16404 ^ n16392;
  assign n16413 = n16412 ^ n16405;
  assign n16683 = n16682 ^ n16413;
  assign n15485 = ~n15322 & n15468;
  assign n15482 = ~n15450 & ~n15458;
  assign n16511 = n15485 ^ n15482;
  assign n16514 = n16513 ^ n16511;
  assign n16510 = n15498 ^ n15478;
  assign n16515 = n16514 ^ n16510;
  assign n16678 = n16515 ^ n15500;
  assign n16684 = n16683 ^ n16678;
  assign n16587 = n14468 & n16567;
  assign n16566 = n14490 & n14528;
  assign n16569 = n16568 ^ n16566;
  assign n16674 = n16587 ^ n16569;
  assign n16675 = n16674 ^ n16562;
  assign n16676 = n16675 ^ n16632;
  assign n16577 = ~n13427 & n16556;
  assign n16555 = n13446 & ~n13587;
  assign n16558 = n16557 ^ n16555;
  assign n16671 = n16577 ^ n16558;
  assign n16672 = n16671 ^ n16551;
  assign n16673 = n16672 ^ n16625;
  assign n16677 = n16676 ^ n16673;
  assign n16685 = n16684 ^ n16677;
  assign n16691 = n16690 ^ n16685;
  assign n16740 = n16739 ^ n16691;
  assign n16564 = n14327 & n14534;
  assign n14520 = n14477 & n14519;
  assign n16565 = n16564 ^ n14520;
  assign n16570 = n16569 ^ n16565;
  assign n16563 = n16562 ^ n14542;
  assign n16571 = n16570 ^ n16563;
  assign n16553 = ~n13445 & ~n13577;
  assign n13594 = n13564 & n13573;
  assign n16554 = n16553 ^ n13594;
  assign n16559 = n16558 ^ n16554;
  assign n16552 = n16551 ^ n13591;
  assign n16560 = n16559 ^ n16552;
  assign n16572 = n16571 ^ n16560;
  assign n16544 = n16326 & n16375;
  assign n16398 = n16397 ^ n16395;
  assign n16545 = n16544 ^ n16398;
  assign n16542 = n16304 & n16386;
  assign n16543 = n16542 ^ n16408;
  assign n16546 = n16545 ^ n16543;
  assign n16538 = n16334 & n16383;
  assign n16393 = n16329 & n16376;
  assign n16539 = n16538 ^ n16393;
  assign n16540 = n16539 ^ n16409;
  assign n16541 = n16540 ^ n16392;
  assign n16547 = n16546 ^ n16541;
  assign n16548 = n16547 ^ n16413;
  assign n16533 = ~n15431 & n15468;
  assign n16534 = n16533 ^ n15498;
  assign n16531 = ~n15449 & ~n15458;
  assign n15488 = n15487 ^ n15485;
  assign n16532 = n16531 ^ n15488;
  assign n16535 = n16534 ^ n16532;
  assign n16418 = ~n15434 & n15475;
  assign n15464 = ~n15217 & n15463;
  assign n16419 = n16418 ^ n15464;
  assign n16420 = n16419 ^ n15494;
  assign n16530 = n16420 ^ n15480;
  assign n16536 = n16535 ^ n16530;
  assign n16537 = n16536 ^ n15500;
  assign n16549 = n16548 ^ n16537;
  assign n16573 = n16572 ^ n16549;
  assign n16528 = n16527 ^ n16515;
  assign n15483 = n15386 & ~n15462;
  assign n15484 = n15483 ^ n15482;
  assign n16421 = n16420 ^ n15484;
  assign n16417 = n15497 ^ n15478;
  assign n16422 = n16421 ^ n16417;
  assign n16508 = n16507 ^ n16422;
  assign n16399 = n16346 & n16372;
  assign n16401 = n16400 ^ n16399;
  assign n16402 = n16401 ^ n16398;
  assign n16394 = n16393 ^ n16392;
  assign n16403 = n16402 ^ n16394;
  assign n16414 = n16413 ^ n16403;
  assign n15489 = n15488 ^ n15484;
  assign n15481 = n15480 ^ n15464;
  assign n15490 = n15489 ^ n15481;
  assign n15501 = n15500 ^ n15490;
  assign n16415 = n16414 ^ n15501;
  assign n14544 = n14543 ^ n14542;
  assign n14530 = n14469 & n14529;
  assign n14523 = n14481 & n14522;
  assign n14531 = n14530 ^ n14523;
  assign n14538 = n14537 ^ n14531;
  assign n14516 = n14362 & n14515;
  assign n14521 = n14520 ^ n14516;
  assign n14539 = n14538 ^ n14521;
  assign n14545 = n14544 ^ n14539;
  assign n13599 = ~n13549 & ~n13588;
  assign n13598 = ~n13532 & n13597;
  assign n13600 = n13599 ^ n13598;
  assign n13602 = n13601 ^ n13600;
  assign n13595 = n13503 & n13583;
  assign n13596 = n13595 ^ n13594;
  assign n13603 = n13602 ^ n13596;
  assign n13593 = n13592 ^ n13591;
  assign n13604 = n13603 ^ n13593;
  assign n14546 = n14545 ^ n13604;
  assign n16416 = n16415 ^ n14546;
  assign n16509 = n16508 ^ n16416;
  assign n16529 = n16528 ^ n16509;
  assign n16574 = n16573 ^ n16529;
  assign n16741 = n16740 ^ n16574;
  assign n16669 = n16668 ^ n15490;
  assign n16663 = n16413 ^ n15500;
  assign n16588 = n16587 ^ n16564;
  assign n16660 = n16588 ^ n14521;
  assign n16659 = n16632 ^ n14523;
  assign n16661 = n16660 ^ n16659;
  assign n16578 = n16577 ^ n16553;
  assign n16657 = n16578 ^ n13596;
  assign n16656 = n16625 ^ n13598;
  assign n16658 = n16657 ^ n16656;
  assign n16662 = n16661 ^ n16658;
  assign n16664 = n16663 ^ n16662;
  assign n16670 = n16669 ^ n16664;
  assign n16759 = n16741 ^ n16670;
  assign n16716 = n16715 ^ n16710;
  assign n16703 = n16332 & n16383;
  assign n16704 = n16703 ^ n16539;
  assign n16701 = n16410 ^ n16390;
  assign n16702 = n16701 ^ n16545;
  assign n16705 = n16704 ^ n16702;
  assign n16608 = n15414 & n15475;
  assign n16609 = n16608 ^ n16419;
  assign n16606 = n15493 ^ n15470;
  assign n16607 = n16606 ^ n16532;
  assign n16610 = n16609 ^ n16607;
  assign n16706 = n16705 ^ n16610;
  assign n16698 = n16561 ^ n14542;
  assign n16697 = n16696 ^ n16674;
  assign n16699 = n16698 ^ n16697;
  assign n16694 = n16550 ^ n13591;
  assign n16693 = n16692 ^ n16671;
  assign n16695 = n16694 ^ n16693;
  assign n16700 = n16699 ^ n16695;
  assign n16707 = n16706 ^ n16700;
  assign n16717 = n16716 ^ n16707;
  assign n16622 = n16621 ^ n16610;
  assign n16599 = n16598 ^ n16408;
  assign n16600 = n16599 ^ n16392;
  assign n16604 = n16603 ^ n16600;
  assign n16592 = n14416 & n14529;
  assign n16593 = n16592 ^ n14531;
  assign n16589 = n14479 & n14519;
  assign n16590 = n16589 ^ n16588;
  assign n16586 = n16585 ^ n14541;
  assign n16591 = n16590 ^ n16586;
  assign n16594 = n16593 ^ n16591;
  assign n16582 = ~n13528 & ~n13588;
  assign n16583 = n16582 ^ n13600;
  assign n16579 = ~n13565 & n13573;
  assign n16580 = n16579 ^ n16578;
  assign n16576 = n16575 ^ n13579;
  assign n16581 = n16580 ^ n16576;
  assign n16584 = n16583 ^ n16581;
  assign n16595 = n16594 ^ n16584;
  assign n16605 = n16604 ^ n16595;
  assign n16623 = n16622 ^ n16605;
  assign n16718 = n16717 ^ n16623;
  assign n16719 = n16718 ^ n16670;
  assign n16652 = n16651 ^ n16536;
  assign n16640 = n16406 ^ n16391;
  assign n16639 = n16540 ^ n16401;
  assign n16641 = n16640 ^ n16639;
  assign n16642 = n16641 ^ n16422;
  assign n16634 = n14478 & n14534;
  assign n16635 = n16634 ^ n16562;
  assign n16636 = n16635 ^ n16590;
  assign n16633 = n16632 ^ n14538;
  assign n16637 = n16636 ^ n16633;
  assign n16627 = n13546 & ~n13577;
  assign n16628 = n16627 ^ n16551;
  assign n16629 = n16628 ^ n16580;
  assign n16626 = n16625 ^ n13602;
  assign n16630 = n16629 ^ n16626;
  assign n16638 = n16637 ^ n16630;
  assign n16643 = n16642 ^ n16638;
  assign n16653 = n16652 ^ n16643;
  assign n16654 = n16653 ^ n16623;
  assign n16655 = n16654 ^ n16574;
  assign n16777 = n16719 ^ n16655;
  assign n16720 = n16719 ^ n16691;
  assign n16776 = n16740 ^ n16720;
  assign n16781 = n16777 ^ n16776;
  assign n16778 = ~n16776 & ~n16777;
  assign n16743 = n16739 ^ n16509;
  assign n16772 = n16655 & ~n16743;
  assign n16779 = n16778 ^ n16772;
  assign n16747 = n16741 ^ n16718;
  assign n16748 = n16739 ^ n16653;
  assign n16754 = ~n16747 & n16748;
  assign n16751 = n16717 ^ n16653;
  assign n16752 = n16751 ^ n16574;
  assign n16753 = n16740 & n16752;
  assign n16755 = n16754 ^ n16753;
  assign n16780 = n16779 ^ n16755;
  assign n16782 = n16781 ^ n16780;
  assign n16771 = n16509 & ~n16719;
  assign n16773 = n16772 ^ n16771;
  assign n16769 = n16743 ^ n16655;
  assign n16742 = n16691 ^ n16653;
  assign n16762 = n16740 ^ n16654;
  assign n16763 = n16742 & ~n16762;
  assign n16764 = n16763 ^ n16753;
  assign n16770 = n16769 ^ n16764;
  assign n16774 = n16773 ^ n16770;
  assign n16792 = n16782 ^ n16774;
  assign n16765 = n16751 ^ n16741;
  assign n16766 = n16765 ^ n16764;
  assign n16757 = n16719 ^ n16509;
  assign n16758 = n16757 ^ n16748;
  assign n16760 = n16758 & n16759;
  assign n16744 = n16743 ^ n16742;
  assign n16745 = ~n16741 & ~n16744;
  assign n16761 = n16760 ^ n16745;
  assign n16767 = n16766 ^ n16761;
  assign n16775 = n16767 & ~n16774;
  assign n16799 = n16792 ^ n16775;
  assign n16749 = n16748 ^ n16747;
  assign n16721 = ~n16670 & ~n16720;
  assign n16746 = n16745 ^ n16721;
  assign n16750 = n16749 ^ n16746;
  assign n16756 = n16755 ^ n16750;
  assign n16797 = ~n16756 & ~n16774;
  assign n16798 = ~n16782 & n16797;
  assign n16800 = n16799 ^ n16798;
  assign n19873 = n16759 & ~n16800;
  assign n16793 = n16775 ^ n16756;
  assign n16794 = ~n16792 & ~n16793;
  assign n16795 = n16794 ^ n16782;
  assign n16807 = n16800 ^ n16795;
  assign n16808 = ~n16744 & ~n16807;
  assign n19874 = n19873 ^ n16808;
  assign n16824 = ~n16741 & ~n16807;
  assign n19875 = n19874 ^ n16824;
  assign n16811 = n16758 & ~n16800;
  assign n16787 = n16756 & n16767;
  assign n16788 = n16782 & n16787;
  assign n16768 = n16767 ^ n16756;
  assign n16786 = n16775 ^ n16768;
  assign n16789 = n16788 ^ n16786;
  assign n16810 = ~n16719 & ~n16789;
  assign n16812 = n16811 ^ n16810;
  assign n19876 = n19875 ^ n16812;
  assign n16783 = n16782 ^ n16775;
  assign n16784 = ~n16768 & n16783;
  assign n16785 = n16784 ^ n16756;
  assign n16796 = n16795 ^ n16785;
  assign n16804 = n16740 & ~n16796;
  assign n16801 = n16800 ^ n16789;
  assign n16802 = n16801 ^ n16796;
  assign n16803 = n16742 & ~n16802;
  assign n16805 = n16804 ^ n16803;
  assign n16790 = n16789 ^ n16785;
  assign n16791 = n16655 & n16790;
  assign n16806 = n16805 ^ n16791;
  assign n19877 = n19876 ^ n16806;
  assign n23305 = n19925 ^ n19877;
  assign n25582 = n25581 ^ n23305;
  assign n25584 = n25583 ^ n25582;
  assign n19649 = n17800 ^ n17782;
  assign n19645 = n17722 & n17774;
  assign n17768 = n17533 & n17767;
  assign n19646 = n19645 ^ n17768;
  assign n19647 = n19646 ^ n17797;
  assign n17786 = n17732 & n17766;
  assign n17788 = n17787 ^ n17786;
  assign n19648 = n19647 ^ n17788;
  assign n19650 = n19649 ^ n19648;
  assign n25568 = n22652 ^ n19650;
  assign n19845 = ~n19516 & n19615;
  assign n19844 = n19843 ^ n19816;
  assign n19846 = n19845 ^ n19844;
  assign n19841 = n19515 & n19611;
  assign n19842 = n19841 ^ n19814;
  assign n19847 = n19846 ^ n19842;
  assign n19630 = n19570 & n19629;
  assign n19628 = n19575 & n19625;
  assign n19631 = n19630 ^ n19628;
  assign n19632 = n19631 ^ n19627;
  assign n19840 = n19839 ^ n19632;
  assign n19848 = n19847 ^ n19840;
  assign n19641 = n19640 ^ n19637;
  assign n19633 = ~n19596 & n19624;
  assign n19635 = n19634 ^ n19633;
  assign n19636 = n19635 ^ n19632;
  assign n19642 = n19641 ^ n19636;
  assign n25566 = n19848 ^ n19642;
  assign n19834 = ~n18702 & ~n18719;
  assign n19805 = ~n18508 & n18716;
  assign n19833 = n19832 ^ n19805;
  assign n19835 = n19834 ^ n19833;
  assign n19830 = ~n18543 & n18716;
  assign n19831 = n19830 ^ n19803;
  assign n19836 = n19835 ^ n19831;
  assign n18734 = ~n18666 & n18733;
  assign n18732 = ~n18670 & n18725;
  assign n18735 = n18734 ^ n18732;
  assign n18731 = ~n18687 & ~n18726;
  assign n18736 = n18735 ^ n18731;
  assign n19829 = n19828 ^ n18736;
  assign n19837 = n19836 ^ n19829;
  assign n19788 = ~n16776 & ~n16785;
  assign n16823 = ~n16670 & n16795;
  assign n16825 = n16824 ^ n16823;
  assign n19789 = n19788 ^ n16825;
  assign n19786 = ~n16720 & n16795;
  assign n19787 = n19786 ^ n16812;
  assign n19790 = n19789 ^ n19787;
  assign n19782 = ~n16747 & n16801;
  assign n16818 = ~n16743 & n16790;
  assign n19783 = n19782 ^ n16818;
  assign n16813 = ~n16762 & ~n16802;
  assign n19784 = n19783 ^ n16813;
  assign n19785 = n19784 ^ n16806;
  assign n19791 = n19790 ^ n19785;
  assign n24242 = n19837 ^ n19791;
  assign n25567 = n25566 ^ n24242;
  assign n25569 = n25568 ^ n25567;
  assign n25606 = n25584 ^ n25569;
  assign n17791 = n17692 & n17790;
  assign n19878 = n19761 ^ n17791;
  assign n19879 = n19878 ^ n17802;
  assign n19880 = n19879 ^ n17784;
  assign n25561 = n22692 ^ n19880;
  assign n19891 = n19573 & n19625;
  assign n19892 = n19891 ^ n19631;
  assign n19889 = n19888 ^ n19639;
  assign n19890 = n19889 ^ n19846;
  assign n19893 = n19892 ^ n19890;
  assign n25559 = n19928 ^ n19893;
  assign n19997 = n16748 & n16801;
  assign n19998 = n19997 ^ n19783;
  assign n16814 = n16752 & ~n16796;
  assign n19995 = n16814 ^ n16804;
  assign n19996 = n19995 ^ n19789;
  assign n19999 = n19998 ^ n19996;
  assign n19885 = n18671 & n18725;
  assign n19886 = n19885 ^ n18735;
  assign n19882 = n18676 & ~n18720;
  assign n19883 = n19882 ^ n18728;
  assign n19884 = n19883 ^ n19835;
  assign n19887 = n19886 ^ n19884;
  assign n23327 = n19999 ^ n19887;
  assign n25560 = n25559 ^ n23327;
  assign n25562 = n25561 ^ n25560;
  assign n25593 = n25569 ^ n25562;
  assign n19796 = n17753 & n17762;
  assign n17792 = n17791 ^ n17789;
  assign n19797 = n19796 ^ n17792;
  assign n19794 = n17656 & n17777;
  assign n19795 = n19794 ^ n17802;
  assign n19798 = n19797 ^ n19795;
  assign n19793 = n19647 ^ n17784;
  assign n19799 = n19798 ^ n19793;
  assign n19800 = n19799 ^ n17804;
  assign n25578 = n22606 ^ n19800;
  assign n24260 = n19955 ^ n19848;
  assign n25577 = n24260 ^ n19823;
  assign n25579 = n25578 ^ n25577;
  assign n17793 = n17792 ^ n17788;
  assign n17785 = n17784 ^ n17768;
  assign n17794 = n17793 ^ n17785;
  assign n17805 = n17804 ^ n17794;
  assign n25550 = n22539 ^ n17805;
  assign n19981 = n19844 ^ n19635;
  assign n19980 = n19839 ^ n19630;
  assign n19982 = n19981 ^ n19980;
  assign n24252 = n19982 ^ n19955;
  assign n25548 = n24252 ^ n19642;
  assign n16821 = n16757 & ~n16789;
  assign n16820 = ~n16777 & ~n16785;
  assign n16822 = n16821 ^ n16820;
  assign n19851 = n19784 ^ n16822;
  assign n19850 = n16810 ^ n16805;
  assign n19852 = n19851 ^ n19850;
  assign n18738 = ~n18703 & ~n18719;
  assign n18737 = n18680 & ~n18711;
  assign n18739 = n18738 ^ n18737;
  assign n18740 = n18739 ^ n18736;
  assign n18730 = n18729 ^ n18712;
  assign n18741 = n18740 ^ n18730;
  assign n23299 = n19852 ^ n18741;
  assign n25549 = n25548 ^ n23299;
  assign n25551 = n25550 ^ n25549;
  assign n19917 = n16823 ^ n16820;
  assign n19918 = n19917 ^ n19874;
  assign n19916 = n16812 ^ n16805;
  assign n19919 = n19918 ^ n19916;
  assign n19806 = n19805 ^ n18738;
  assign n19811 = n19810 ^ n19806;
  assign n19804 = n19803 ^ n18729;
  assign n19812 = n19811 ^ n19804;
  assign n24258 = n19919 ^ n19812;
  assign n25576 = n25551 ^ n24258;
  assign n25580 = n25579 ^ n25576;
  assign n25594 = n25593 ^ n25580;
  assign n19898 = n17723 & n17774;
  assign n19899 = n19898 ^ n19646;
  assign n19896 = n17798 ^ n17781;
  assign n19897 = n19896 ^ n19797;
  assign n19900 = n19899 ^ n19897;
  assign n25557 = n22793 ^ n19900;
  assign n20005 = n19813 ^ n19640;
  assign n20004 = n19953 ^ n19926;
  assign n20006 = n20005 ^ n20004;
  assign n25555 = n20006 ^ n19893;
  assign n20002 = n19802 ^ n18729;
  assign n19949 = n19882 ^ n18731;
  assign n20001 = n19949 ^ n19923;
  assign n20003 = n20002 ^ n20001;
  assign n19945 = n16811 ^ n16805;
  assign n16815 = n16814 ^ n16813;
  assign n19944 = n19875 ^ n16815;
  assign n19946 = n19945 ^ n19944;
  assign n23310 = n20003 ^ n19946;
  assign n25556 = n25555 ^ n23310;
  assign n25558 = n25557 ^ n25556;
  assign n25563 = n25562 ^ n25558;
  assign n25553 = n22768 ^ n17804;
  assign n19977 = n19833 ^ n18739;
  assign n19976 = n19828 ^ n18734;
  assign n19978 = n19977 ^ n19976;
  assign n16826 = n16825 ^ n16822;
  assign n16819 = n16818 ^ n16806;
  assign n16827 = n16826 ^ n16819;
  assign n24267 = n19978 ^ n16827;
  assign n25552 = n24267 ^ n24252;
  assign n25554 = n25553 ^ n25552;
  assign n25564 = n25563 ^ n25554;
  assign n25599 = n25594 ^ n25564;
  assign n25597 = n25584 ^ n25564;
  assign n19942 = n17801 ^ n17782;
  assign n19941 = n19878 ^ n17799;
  assign n19943 = n19942 ^ n19941;
  assign n25572 = n22745 ^ n19943;
  assign n25570 = n20006 ^ n19955;
  assign n19950 = n19949 ^ n19803;
  assign n19948 = n19828 ^ n19808;
  assign n19951 = n19950 ^ n19948;
  assign n16816 = n16815 ^ n16812;
  assign n16809 = n16808 ^ n16806;
  assign n16817 = n16816 ^ n16809;
  assign n24286 = n19951 ^ n16817;
  assign n25571 = n25570 ^ n24286;
  assign n25573 = n25572 ^ n25571;
  assign n25585 = n25584 ^ n25573;
  assign n25598 = n25597 ^ n25585;
  assign n25603 = n25599 ^ n25598;
  assign n25600 = ~n25598 & ~n25599;
  assign n25595 = n25573 ^ n25551;
  assign n25596 = n25594 & ~n25595;
  assign n25601 = n25600 ^ n25596;
  assign n25589 = n25569 ^ n25558;
  assign n25590 = n25589 ^ n25580;
  assign n25591 = n25585 & n25590;
  assign n25574 = n25573 ^ n25569;
  assign n25586 = n25585 ^ n25580;
  assign n25587 = n25586 ^ n25563;
  assign n25588 = n25574 & ~n25587;
  assign n25592 = n25591 ^ n25588;
  assign n25602 = n25601 ^ n25592;
  assign n25604 = n25603 ^ n25602;
  assign n25610 = n25587 ^ n25574;
  assign n25607 = n25606 ^ n25595;
  assign n25608 = ~n25586 & ~n25607;
  assign n25605 = ~n25554 & ~n25597;
  assign n25609 = n25608 ^ n25605;
  assign n25611 = n25610 ^ n25609;
  assign n25612 = n25611 ^ n25592;
  assign n25627 = n25589 ^ n25586;
  assign n25614 = n25593 ^ n25585;
  assign n25615 = n25606 & ~n25614;
  assign n25616 = n25615 ^ n25591;
  assign n25628 = n25627 ^ n25616;
  assign n25565 = n25564 ^ n25551;
  assign n25575 = n25574 ^ n25565;
  assign n25624 = n25586 ^ n25554;
  assign n25625 = n25575 & n25624;
  assign n25626 = n25625 ^ n25608;
  assign n25629 = n25628 ^ n25626;
  assign n25636 = n25612 & n25629;
  assign n25637 = n25604 & n25636;
  assign n25634 = n25629 ^ n25612;
  assign n25618 = n25551 & ~n25564;
  assign n25619 = n25618 ^ n25596;
  assign n25613 = n25595 ^ n25594;
  assign n25617 = n25616 ^ n25613;
  assign n25620 = n25619 ^ n25617;
  assign n25630 = ~n25620 & n25629;
  assign n25635 = n25634 ^ n25630;
  assign n25638 = n25637 ^ n25635;
  assign n25623 = n25620 ^ n25604;
  assign n25631 = n25630 ^ n25623;
  assign n25621 = ~n25612 & ~n25620;
  assign n25622 = ~n25604 & n25621;
  assign n25632 = n25631 ^ n25622;
  assign n25658 = n25638 ^ n25632;
  assign n25651 = n25630 ^ n25604;
  assign n25652 = ~n25634 & n25651;
  assign n25653 = n25652 ^ n25612;
  assign n25641 = n25630 ^ n25612;
  assign n25642 = ~n25623 & ~n25641;
  assign n25643 = n25642 ^ n25604;
  assign n25656 = n25653 ^ n25643;
  assign n25659 = n25658 ^ n25656;
  assign n25660 = n25606 & ~n25659;
  assign n25657 = n25585 & ~n25656;
  assign n25661 = n25660 ^ n25657;
  assign n25633 = n25575 & ~n25632;
  assign n25895 = n25661 ^ n25633;
  assign n25858 = n25590 & ~n25656;
  assign n25806 = ~n25614 & ~n25659;
  assign n25859 = n25858 ^ n25806;
  assign n25647 = n25624 & ~n25632;
  assign n25644 = n25643 ^ n25632;
  assign n25646 = ~n25607 & ~n25644;
  assign n25648 = n25647 ^ n25646;
  assign n25645 = ~n25586 & ~n25644;
  assign n25649 = n25648 ^ n25645;
  assign n25894 = n25859 ^ n25649;
  assign n25896 = n25895 ^ n25894;
  assign n25905 = n25904 ^ n25896;
  assign n22362 = n19653 ^ n19475;
  assign n22360 = n19436 ^ n19410;
  assign n22361 = n22360 ^ n19442;
  assign n22363 = n22362 ^ n22361;
  assign n21314 = n19556 ^ n19447;
  assign n22350 = n21314 ^ n19674;
  assign n22348 = n19411 ^ n19086;
  assign n22349 = n22348 ^ n19391;
  assign n22351 = n22350 ^ n22349;
  assign n22364 = n22363 ^ n22351;
  assign n22332 = n19551 ^ n19405;
  assign n21347 = n19447 ^ n19363;
  assign n22331 = n21347 ^ n19663;
  assign n22333 = n22332 ^ n22331;
  assign n21320 = n19502 ^ n19447;
  assign n22328 = n21320 ^ n19655;
  assign n22326 = n19525 ^ n19325;
  assign n22327 = n22326 ^ n19520;
  assign n22329 = n22328 ^ n22327;
  assign n22330 = n22329 ^ n19543;
  assign n22334 = n22333 ^ n22330;
  assign n22365 = n22364 ^ n22334;
  assign n22346 = n19670 ^ n19447;
  assign n22345 = n19525 ^ n19495;
  assign n22347 = n22346 ^ n22345;
  assign n22383 = n22365 ^ n22347;
  assign n22354 = n19667 ^ n19217;
  assign n22352 = n19470 ^ n19436;
  assign n22353 = n22352 ^ n19462;
  assign n22355 = n22354 ^ n22353;
  assign n22341 = n19660 ^ n19419;
  assign n22339 = n19470 ^ n19086;
  assign n22340 = n22339 ^ n18974;
  assign n22342 = n22341 ^ n22340;
  assign n22356 = n22355 ^ n22342;
  assign n22357 = n22356 ^ n22347;
  assign n22403 = n22329 & ~n22357;
  assign n22337 = n19658 ^ n19530;
  assign n22335 = n19550 ^ n19325;
  assign n22336 = n22335 ^ n19347;
  assign n22338 = n22337 ^ n22336;
  assign n22343 = n22342 ^ n22338;
  assign n22344 = n22343 ^ n22334;
  assign n22367 = n22363 ^ n22329;
  assign n22396 = n22344 & ~n22367;
  assign n22404 = n22403 ^ n22396;
  assign n22401 = n22367 ^ n22344;
  assign n22366 = n22351 ^ n22338;
  assign n22387 = n22364 ^ n22343;
  assign n22388 = n22366 & ~n22387;
  assign n22376 = n22355 ^ n22338;
  assign n22377 = n22376 ^ n22334;
  assign n22378 = n22364 & n22377;
  assign n22389 = n22388 ^ n22378;
  assign n22402 = n22401 ^ n22389;
  assign n22405 = n22404 ^ n22402;
  assign n22394 = n22357 ^ n22344;
  assign n22358 = n22357 ^ n22351;
  assign n22393 = n22364 ^ n22358;
  assign n22399 = n22394 ^ n22393;
  assign n22395 = ~n22393 & ~n22394;
  assign n22397 = n22396 ^ n22395;
  assign n22371 = n22365 ^ n22356;
  assign n22372 = n22363 ^ n22338;
  assign n22375 = ~n22371 & n22372;
  assign n22379 = n22378 ^ n22375;
  assign n22398 = n22397 ^ n22379;
  assign n22400 = n22399 ^ n22398;
  assign n22416 = n22405 ^ n22400;
  assign n22386 = n22376 ^ n22365;
  assign n22390 = n22389 ^ n22386;
  assign n22381 = n22357 ^ n22329;
  assign n22382 = n22381 ^ n22372;
  assign n22384 = n22382 & n22383;
  assign n22368 = n22367 ^ n22366;
  assign n22369 = ~n22365 & ~n22368;
  assign n22385 = n22384 ^ n22369;
  assign n22391 = n22390 ^ n22385;
  assign n22406 = n22391 & ~n22405;
  assign n22424 = n22416 ^ n22406;
  assign n22373 = n22372 ^ n22371;
  assign n22359 = ~n22347 & ~n22358;
  assign n22370 = n22369 ^ n22359;
  assign n22374 = n22373 ^ n22370;
  assign n22380 = n22379 ^ n22374;
  assign n22422 = ~n22380 & ~n22405;
  assign n22423 = ~n22400 & n22422;
  assign n22425 = n22424 ^ n22423;
  assign n22679 = n22383 & ~n22425;
  assign n22417 = n22406 ^ n22380;
  assign n22418 = ~n22416 & ~n22417;
  assign n22419 = n22418 ^ n22400;
  assign n22431 = n22425 ^ n22419;
  assign n22432 = ~n22368 & ~n22431;
  assign n22680 = n22679 ^ n22432;
  assign n22448 = ~n22365 & ~n22431;
  assign n22681 = n22680 ^ n22448;
  assign n22435 = n22382 & ~n22425;
  assign n22411 = n22380 & n22391;
  assign n22412 = n22400 & n22411;
  assign n22392 = n22391 ^ n22380;
  assign n22410 = n22406 ^ n22392;
  assign n22413 = n22412 ^ n22410;
  assign n22434 = ~n22357 & ~n22413;
  assign n22436 = n22435 ^ n22434;
  assign n22682 = n22681 ^ n22436;
  assign n22426 = n22425 ^ n22413;
  assign n22407 = n22406 ^ n22400;
  assign n22408 = ~n22392 & n22407;
  assign n22409 = n22408 ^ n22380;
  assign n22420 = n22419 ^ n22409;
  assign n22427 = n22426 ^ n22420;
  assign n22428 = n22366 & ~n22427;
  assign n22421 = n22364 & ~n22420;
  assign n22429 = n22428 ^ n22421;
  assign n22414 = n22413 ^ n22409;
  assign n22415 = n22344 & n22414;
  assign n22430 = n22429 ^ n22415;
  assign n22683 = n22682 ^ n22430;
  assign n25441 = n25440 ^ n22683;
  assign n20491 = n16641 ^ n14545;
  assign n22243 = n20491 ^ n16536;
  assign n22244 = n22243 ^ n16547;
  assign n22245 = n22244 ^ n16630;
  assign n22246 = n22245 ^ n18659;
  assign n22213 = n18385 ^ n16710;
  assign n20503 = n16705 ^ n16594;
  assign n22211 = n20503 ^ n16695;
  assign n22212 = n22211 ^ n16731;
  assign n22214 = n22213 ^ n22212;
  assign n22257 = n22246 ^ n22214;
  assign n21077 = n16727 ^ n16637;
  assign n22235 = n21077 ^ n16560;
  assign n22234 = n16682 ^ n16548;
  assign n22236 = n22235 ^ n22234;
  assign n22231 = n18570 ^ n16422;
  assign n21046 = n16727 ^ n16661;
  assign n22229 = n21046 ^ n13604;
  assign n22228 = n16641 ^ n16414;
  assign n22230 = n22229 ^ n22228;
  assign n22232 = n22231 ^ n22230;
  assign n22227 = n18585 ^ n16515;
  assign n22233 = n22232 ^ n22227;
  assign n22237 = n22236 ^ n22233;
  assign n22258 = n22257 ^ n22237;
  assign n22221 = n16683 ^ n16604;
  assign n21052 = n16727 ^ n16571;
  assign n22222 = n22221 ^ n21052;
  assign n22223 = n22222 ^ n16673;
  assign n22224 = n22223 ^ n18537;
  assign n22247 = n22246 ^ n22224;
  assign n22208 = n16706 ^ n16584;
  assign n22209 = n22208 ^ n18454;
  assign n20520 = n16676 ^ n16600;
  assign n22210 = n22209 ^ n20520;
  assign n22268 = n22246 ^ n22210;
  assign n20525 = n16731 ^ n16699;
  assign n22238 = n20525 ^ n16724;
  assign n22239 = n22238 ^ n16663;
  assign n22240 = n22239 ^ n18628;
  assign n22241 = n22240 ^ n22224;
  assign n22269 = n22268 ^ n22241;
  assign n22270 = n22247 & ~n22269;
  assign n22259 = n22241 & n22258;
  assign n22271 = n22270 ^ n22259;
  assign n22242 = n22241 ^ n22237;
  assign n22267 = n22257 ^ n22242;
  assign n22272 = n22271 ^ n22267;
  assign n22218 = n18502 ^ n15490;
  assign n22216 = n16727 ^ n16658;
  assign n22217 = n22216 ^ n16414;
  assign n22219 = n22218 ^ n22217;
  assign n22215 = n22214 ^ n22210;
  assign n22220 = n22219 ^ n22215;
  assign n22262 = n22232 ^ n22220;
  assign n22253 = n22246 ^ n22240;
  assign n22263 = n22262 ^ n22253;
  assign n22264 = n22242 ^ n22219;
  assign n22265 = n22263 & n22264;
  assign n22248 = n22240 ^ n22232;
  assign n22249 = n22248 ^ n22247;
  assign n22250 = ~n22242 & ~n22249;
  assign n22266 = n22265 ^ n22250;
  assign n22273 = n22272 ^ n22266;
  assign n22252 = n22242 ^ n22215;
  assign n22256 = ~n22252 & n22253;
  assign n22260 = n22259 ^ n22256;
  assign n22254 = n22253 ^ n22252;
  assign n22225 = n22224 ^ n22220;
  assign n22226 = ~n22219 & ~n22225;
  assign n22251 = n22250 ^ n22226;
  assign n22255 = n22254 ^ n22251;
  assign n22261 = n22260 ^ n22255;
  assign n22274 = n22273 ^ n22261;
  assign n22275 = n22268 ^ n22237;
  assign n22285 = n22275 ^ n22220;
  assign n22284 = n22241 ^ n22225;
  assign n22289 = n22285 ^ n22284;
  assign n22286 = ~n22284 & ~n22285;
  assign n22279 = ~n22248 & n22275;
  assign n22287 = n22286 ^ n22279;
  assign n22288 = n22287 ^ n22260;
  assign n22290 = n22289 ^ n22288;
  assign n22278 = ~n22220 & n22232;
  assign n22280 = n22279 ^ n22278;
  assign n22276 = n22275 ^ n22248;
  assign n22277 = n22276 ^ n22271;
  assign n22281 = n22280 ^ n22277;
  assign n22282 = n22273 & ~n22281;
  assign n22299 = n22290 ^ n22282;
  assign n22300 = ~n22274 & n22299;
  assign n22301 = n22300 ^ n22261;
  assign n22295 = n22290 ^ n22281;
  assign n22296 = n22282 ^ n22261;
  assign n22297 = ~n22295 & ~n22296;
  assign n22298 = n22297 ^ n22290;
  assign n22302 = n22301 ^ n22298;
  assign n22671 = n22258 & ~n22302;
  assign n22305 = n22295 ^ n22282;
  assign n22303 = ~n22261 & ~n22281;
  assign n22304 = ~n22290 & n22303;
  assign n22306 = n22305 ^ n22304;
  assign n22291 = n22261 & n22273;
  assign n22292 = n22290 & n22291;
  assign n22283 = n22282 ^ n22274;
  assign n22293 = n22292 ^ n22283;
  assign n22307 = n22306 ^ n22293;
  assign n22308 = n22307 ^ n22302;
  assign n22313 = ~n22269 & ~n22308;
  assign n22731 = n22671 ^ n22313;
  assign n22554 = n22263 & ~n22306;
  assign n22294 = ~n22220 & ~n22293;
  assign n22555 = n22554 ^ n22294;
  assign n22732 = n22731 ^ n22555;
  assign n22314 = n22301 ^ n22293;
  assign n22623 = n22275 & n22314;
  assign n22310 = n22241 & ~n22302;
  assign n22309 = n22247 & ~n22308;
  assign n22311 = n22310 ^ n22309;
  assign n22624 = n22623 ^ n22311;
  assign n22559 = n22306 ^ n22298;
  assign n22560 = ~n22249 & ~n22559;
  assign n22730 = n22624 ^ n22560;
  assign n22733 = n22732 ^ n22730;
  assign n22561 = n22264 & ~n22306;
  assign n22562 = n22561 ^ n22560;
  assign n22557 = ~n22219 & n22298;
  assign n22320 = ~n22285 & ~n22301;
  assign n22558 = n22557 ^ n22320;
  assign n22563 = n22562 ^ n22558;
  assign n22556 = n22555 ^ n22311;
  assign n22564 = n22563 ^ n22556;
  assign n24395 = n22733 ^ n22564;
  assign n21996 = n21995 ^ n18523;
  assign n21446 = n18615 ^ n18595;
  assign n21993 = n21446 ^ n18519;
  assign n21994 = n21993 ^ n18411;
  assign n21997 = n21996 ^ n21994;
  assign n21989 = n21988 ^ n18624;
  assign n21466 = n18483 ^ n18469;
  assign n20378 = n18618 ^ n17920;
  assign n21987 = n21466 ^ n20378;
  assign n21990 = n21989 ^ n21987;
  assign n21998 = n21997 ^ n21990;
  assign n21978 = n21977 ^ n18580;
  assign n21459 = n18641 ^ n18615;
  assign n21976 = n21459 ^ n18602;
  assign n21979 = n21978 ^ n21976;
  assign n21958 = n21957 ^ n18565;
  assign n21441 = n18615 ^ n18478;
  assign n21955 = n21441 ^ n18554;
  assign n21956 = n21955 ^ n18650;
  assign n21959 = n21958 ^ n21956;
  assign n21457 = n18528 ^ n18518;
  assign n21975 = n21959 ^ n21457;
  assign n21980 = n21979 ^ n21975;
  assign n22008 = n21998 ^ n21980;
  assign n21442 = n18553 ^ n18466;
  assign n20394 = n18615 ^ n18483;
  assign n21971 = n21442 ^ n20394;
  assign n21970 = n21969 ^ n18493;
  assign n21972 = n21971 ^ n21970;
  assign n22029 = n22008 ^ n21972;
  assign n21983 = n21982 ^ n18646;
  assign n21473 = n18608 ^ n18601;
  assign n20349 = n18649 ^ n18548;
  assign n21981 = n21473 ^ n20349;
  assign n21984 = n21983 ^ n21981;
  assign n21966 = n21965 ^ n18437;
  assign n20387 = n18513 ^ n18404;
  assign n21964 = n20387 ^ n18298;
  assign n21967 = n21966 ^ n21964;
  assign n21985 = n21984 ^ n21967;
  assign n21986 = n21985 ^ n21980;
  assign n21962 = n21961 ^ n18043;
  assign n20360 = n18424 ^ n18284;
  assign n21960 = n20360 ^ n18619;
  assign n21963 = n21962 ^ n21960;
  assign n21968 = n21967 ^ n21963;
  assign n21973 = n21972 ^ n21968;
  assign n22001 = n21986 ^ n21973;
  assign n21999 = n21997 ^ n21973;
  assign n22000 = n21999 ^ n21998;
  assign n22013 = n22001 ^ n22000;
  assign n22007 = n21990 ^ n21984;
  assign n22009 = n22008 ^ n21968;
  assign n22010 = n22007 & ~n22009;
  assign n22004 = n21984 ^ n21963;
  assign n22005 = n22004 ^ n21980;
  assign n22006 = n21998 & ~n22005;
  assign n22011 = n22010 ^ n22006;
  assign n22002 = n22000 & n22001;
  assign n21991 = n21990 ^ n21959;
  assign n21992 = n21986 & n21991;
  assign n22003 = n22002 ^ n21992;
  assign n22012 = n22011 ^ n22003;
  assign n22014 = n22013 ^ n22012;
  assign n22020 = n22009 ^ n22007;
  assign n22018 = ~n21972 & n21999;
  assign n22015 = n21997 ^ n21984;
  assign n22016 = n22015 ^ n21991;
  assign n22017 = n22008 & n22016;
  assign n22019 = n22018 ^ n22017;
  assign n22021 = n22020 ^ n22019;
  assign n22022 = n22021 ^ n22011;
  assign n22038 = ~n21959 & n21973;
  assign n22039 = n22038 ^ n21992;
  assign n22036 = n21991 ^ n21986;
  assign n22024 = n21998 ^ n21985;
  assign n22025 = n22015 & n22024;
  assign n22026 = n22025 ^ n22006;
  assign n22037 = n22036 ^ n22026;
  assign n22040 = n22039 ^ n22037;
  assign n22056 = ~n22022 & n22040;
  assign n22057 = ~n22014 & n22056;
  assign n22050 = n22040 ^ n22014;
  assign n21974 = n21973 ^ n21959;
  assign n22028 = n22007 ^ n21974;
  assign n22030 = n22028 & ~n22029;
  assign n22031 = n22030 ^ n22017;
  assign n22023 = n22008 ^ n22004;
  assign n22027 = n22026 ^ n22023;
  assign n22032 = n22031 ^ n22027;
  assign n22041 = ~n22032 & n22040;
  assign n22055 = n22050 ^ n22041;
  assign n22058 = n22057 ^ n22055;
  assign n22577 = ~n22029 & n22058;
  assign n22051 = n22041 ^ n22022;
  assign n22052 = n22050 & ~n22051;
  assign n22053 = n22052 ^ n22014;
  assign n22078 = n22058 ^ n22053;
  assign n22083 = n22016 & n22078;
  assign n22578 = n22577 ^ n22083;
  assign n22077 = ~n21972 & n22053;
  assign n22035 = n22032 ^ n22022;
  assign n22045 = n22041 ^ n22014;
  assign n22046 = n22035 & n22045;
  assign n22047 = n22046 ^ n22022;
  assign n22048 = n22001 & ~n22047;
  assign n22576 = n22077 ^ n22048;
  assign n22579 = n22578 ^ n22576;
  assign n22087 = n22028 & n22058;
  assign n22042 = n22041 ^ n22035;
  assign n22033 = n22022 & ~n22032;
  assign n22034 = n22014 & n22033;
  assign n22043 = n22042 ^ n22034;
  assign n22071 = n21973 & n22043;
  assign n22088 = n22087 ^ n22071;
  assign n22054 = n22053 ^ n22047;
  assign n22069 = n21998 & ~n22054;
  assign n22059 = n22058 ^ n22043;
  assign n22060 = n22059 ^ n22054;
  assign n22068 = n22015 & ~n22060;
  assign n22070 = n22069 ^ n22068;
  assign n22575 = n22088 ^ n22070;
  assign n22580 = n22579 ^ n22575;
  assign n22085 = ~n22005 & ~n22054;
  assign n22061 = n22024 & ~n22060;
  assign n22086 = n22085 ^ n22061;
  assign n22089 = n22088 ^ n22086;
  assign n22062 = n22047 ^ n22043;
  assign n22074 = n21986 & ~n22062;
  assign n22075 = n22074 ^ n22070;
  assign n22084 = n22083 ^ n22075;
  assign n22090 = n22089 ^ n22084;
  assign n22698 = n22580 ^ n22090;
  assign n25438 = n24395 ^ n22698;
  assign n22628 = ~n22242 & ~n22559;
  assign n22703 = n22628 ^ n22562;
  assign n22704 = n22703 ^ n22555;
  assign n22705 = n22704 ^ n22624;
  assign n22129 = n17662 ^ n17641;
  assign n21195 = n17697 ^ n17095;
  assign n22128 = n21195 ^ n17682;
  assign n22130 = n22129 ^ n22128;
  assign n22126 = n19764 ^ n17648;
  assign n22095 = n19651 ^ n17708;
  assign n21174 = n17539 ^ n17095;
  assign n22093 = n21174 ^ n17518;
  assign n20112 = n17492 ^ n17471;
  assign n22094 = n22093 ^ n20112;
  assign n22096 = n22095 ^ n22094;
  assign n22127 = n22126 ^ n22096;
  assign n22131 = n22130 ^ n22127;
  assign n22115 = n19931 ^ n17619;
  assign n21186 = n17666 ^ n17095;
  assign n22113 = n21186 ^ n17649;
  assign n20116 = n17636 ^ n17615;
  assign n22114 = n22113 ^ n20116;
  assign n22116 = n22115 ^ n22114;
  assign n22098 = n19958 ^ n17517;
  assign n21205 = n17563 ^ n17356;
  assign n20147 = n17236 ^ n16960;
  assign n22097 = n21205 ^ n20147;
  assign n22099 = n22098 ^ n22097;
  assign n22118 = n22116 ^ n22099;
  assign n22138 = n22131 ^ n22118;
  assign n22108 = n17518 ^ n17095;
  assign n22109 = n22108 ^ n17545;
  assign n22110 = n22109 ^ n17497;
  assign n22111 = n22110 ^ n19984;
  assign n22105 = n20009 ^ n17356;
  assign n21201 = n17612 ^ n17588;
  assign n20127 = n17569 ^ n17228;
  assign n22104 = n21201 ^ n20127;
  assign n22106 = n22105 ^ n22104;
  assign n22102 = n19901 ^ n17588;
  assign n21187 = n17634 ^ n17619;
  assign n20132 = n17605 ^ n17577;
  assign n22101 = n21187 ^ n20132;
  assign n22103 = n22102 ^ n22101;
  assign n22107 = n22106 ^ n22103;
  assign n22112 = n22111 ^ n22107;
  assign n22171 = ~n22096 & n22112;
  assign n22100 = n22099 ^ n22096;
  assign n22123 = n19855 ^ n17681;
  assign n22121 = n17702 ^ n17673;
  assign n22120 = n17708 ^ n17481;
  assign n22122 = n22121 ^ n22120;
  assign n22124 = n22123 ^ n22122;
  assign n22125 = n22124 ^ n22103;
  assign n22132 = n22131 ^ n22125;
  assign n22135 = n22100 & n22132;
  assign n22172 = n22171 ^ n22135;
  assign n22169 = n22132 ^ n22100;
  assign n22148 = n22124 ^ n22116;
  assign n22156 = n22125 ^ n22118;
  assign n22157 = n22148 & n22156;
  assign n22141 = n22124 ^ n22106;
  assign n22142 = n22141 ^ n22131;
  assign n22143 = n22118 & n22142;
  assign n22158 = n22157 ^ n22143;
  assign n22170 = n22169 ^ n22158;
  assign n22173 = n22172 ^ n22170;
  assign n22133 = n22132 ^ n22112;
  assign n22117 = n22116 ^ n22112;
  assign n22119 = n22118 ^ n22117;
  assign n22146 = n22133 ^ n22119;
  assign n22137 = n22124 ^ n22099;
  assign n22139 = n22138 ^ n22107;
  assign n22140 = n22137 & n22139;
  assign n22144 = n22143 ^ n22140;
  assign n22134 = n22119 & n22133;
  assign n22136 = n22135 ^ n22134;
  assign n22145 = n22144 ^ n22136;
  assign n22147 = n22146 ^ n22145;
  assign n22185 = n22173 ^ n22147;
  assign n22159 = n22141 ^ n22138;
  assign n22160 = n22159 ^ n22158;
  assign n22151 = n22138 ^ n22111;
  assign n22152 = n22112 ^ n22096;
  assign n22153 = n22152 ^ n22137;
  assign n22154 = n22151 & n22153;
  assign n22149 = n22148 ^ n22100;
  assign n22150 = n22138 & n22149;
  assign n22155 = n22154 ^ n22150;
  assign n22161 = n22160 ^ n22155;
  assign n22174 = n22161 & n22173;
  assign n22164 = n22139 ^ n22137;
  assign n22162 = n22111 & n22117;
  assign n22163 = n22162 ^ n22150;
  assign n22165 = n22164 ^ n22163;
  assign n22166 = n22165 ^ n22144;
  assign n22191 = n22174 ^ n22166;
  assign n22192 = n22185 & n22191;
  assign n22193 = n22192 ^ n22147;
  assign n22186 = n22185 ^ n22174;
  assign n22183 = n22166 & n22173;
  assign n22184 = ~n22147 & n22183;
  assign n22187 = n22186 ^ n22184;
  assign n22549 = n22193 ^ n22187;
  assign n22617 = n22138 & n22549;
  assign n22550 = n22149 & n22549;
  assign n22548 = n22151 & n22187;
  assign n22551 = n22550 ^ n22548;
  assign n22700 = n22617 ^ n22551;
  assign n22543 = n22153 & n22187;
  assign n22175 = n22166 ^ n22161;
  assign n22176 = n22175 ^ n22174;
  assign n22167 = n22161 & ~n22166;
  assign n22168 = n22147 & n22167;
  assign n22177 = n22176 ^ n22168;
  assign n22202 = n22112 & n22177;
  assign n22544 = n22543 ^ n22202;
  assign n22701 = n22700 ^ n22544;
  assign n22178 = n22174 ^ n22147;
  assign n22179 = n22175 & n22178;
  assign n22180 = n22179 ^ n22166;
  assign n22181 = n22180 ^ n22177;
  assign n22612 = n22132 & n22181;
  assign n22194 = n22193 ^ n22180;
  assign n22204 = n22118 & n22194;
  assign n22188 = n22187 ^ n22177;
  assign n22195 = n22194 ^ n22188;
  assign n22203 = n22148 & n22195;
  assign n22205 = n22204 ^ n22203;
  assign n22613 = n22612 ^ n22205;
  assign n22702 = n22701 ^ n22613;
  assign n22706 = n22705 ^ n22702;
  assign n25439 = n25438 ^ n22706;
  assign n25442 = n25441 ^ n25439;
  assign n22588 = ~n22393 & ~n22409;
  assign n22447 = ~n22347 & n22419;
  assign n22449 = n22448 ^ n22447;
  assign n22589 = n22588 ^ n22449;
  assign n22586 = ~n22358 & n22419;
  assign n22587 = n22586 ^ n22436;
  assign n22590 = n22589 ^ n22587;
  assign n22582 = ~n22371 & n22426;
  assign n22442 = ~n22367 & n22414;
  assign n22583 = n22582 ^ n22442;
  assign n22438 = ~n22387 & ~n22427;
  assign n22584 = n22583 ^ n22438;
  assign n22585 = n22584 ^ n22430;
  assign n22591 = n22590 ^ n22585;
  assign n25415 = n25414 ^ n22591;
  assign n22319 = n22262 & ~n22293;
  assign n22321 = n22320 ^ n22319;
  assign n22316 = ~n22252 & n22307;
  assign n22315 = ~n22248 & n22314;
  assign n22317 = n22316 ^ n22315;
  assign n22318 = n22317 ^ n22313;
  assign n22322 = n22321 ^ n22318;
  assign n22312 = n22311 ^ n22294;
  assign n22323 = n22322 ^ n22312;
  assign n22072 = n22071 ^ n22070;
  assign n22064 = ~n22009 & n22059;
  assign n22063 = n21991 & ~n22062;
  assign n22065 = n22064 ^ n22063;
  assign n22066 = n22065 ^ n22061;
  assign n22044 = n21974 & n22043;
  assign n22049 = n22048 ^ n22044;
  assign n22067 = n22066 ^ n22049;
  assign n22073 = n22072 ^ n22067;
  assign n23421 = n22323 ^ n22073;
  assign n22630 = ~n22284 & ~n22301;
  assign n22629 = n22628 ^ n22557;
  assign n22631 = n22630 ^ n22629;
  assign n22626 = ~n22225 & n22298;
  assign n22627 = n22626 ^ n22555;
  assign n22632 = n22631 ^ n22627;
  assign n22625 = n22624 ^ n22318;
  assign n22633 = n22632 ^ n22625;
  assign n22619 = n22119 & n22180;
  assign n22546 = n22111 & n22193;
  assign n22618 = n22617 ^ n22546;
  assign n22620 = n22619 ^ n22618;
  assign n22615 = n22117 & n22193;
  assign n22616 = n22615 ^ n22544;
  assign n22621 = n22620 ^ n22616;
  assign n22196 = n22156 & n22195;
  assign n22189 = n22139 & n22188;
  assign n22182 = n22100 & n22181;
  assign n22190 = n22189 ^ n22182;
  assign n22197 = n22196 ^ n22190;
  assign n22614 = n22613 ^ n22197;
  assign n22622 = n22621 ^ n22614;
  assign n22634 = n22633 ^ n22622;
  assign n25413 = n23421 ^ n22634;
  assign n25416 = n25415 ^ n25413;
  assign n25457 = n25442 ^ n25416;
  assign n22785 = n22372 & n22426;
  assign n22786 = n22785 ^ n22583;
  assign n22437 = n22377 & ~n22420;
  assign n22783 = n22437 ^ n22421;
  assign n22784 = n22783 ^ n22589;
  assign n22787 = n22786 ^ n22784;
  assign n25445 = n25444 ^ n22787;
  assign n22079 = n22008 & n22078;
  assign n22656 = n22578 ^ n22079;
  assign n22657 = n22656 ^ n22088;
  assign n22658 = n22657 ^ n22075;
  assign n23462 = n22705 ^ n22658;
  assign n22674 = n22253 & n22307;
  assign n22675 = n22674 ^ n22317;
  assign n22672 = n22671 ^ n22310;
  assign n22673 = n22672 ^ n22631;
  assign n22676 = n22675 ^ n22673;
  assign n22668 = n22137 & n22188;
  assign n22669 = n22668 ^ n22190;
  assign n22665 = n22142 & n22194;
  assign n22666 = n22665 ^ n22204;
  assign n22667 = n22666 ^ n22620;
  assign n22670 = n22669 ^ n22667;
  assign n22677 = n22676 ^ n22670;
  assign n25443 = n23462 ^ n22677;
  assign n25446 = n25445 ^ n25443;
  assign n25476 = n25446 ^ n25416;
  assign n22439 = n22438 ^ n22437;
  assign n22440 = n22439 ^ n22436;
  assign n22433 = n22432 ^ n22430;
  assign n22441 = n22440 ^ n22433;
  assign n25453 = n25452 ^ n22441;
  assign n22779 = n22554 ^ n22311;
  assign n22778 = n22731 ^ n22703;
  assign n22780 = n22779 ^ n22778;
  assign n22723 = n22087 ^ n22070;
  assign n22722 = n22656 ^ n22086;
  assign n22724 = n22723 ^ n22722;
  assign n23427 = n22780 ^ n22724;
  assign n22727 = n22665 ^ n22196;
  assign n22728 = n22727 ^ n22544;
  assign n22726 = n22613 ^ n22550;
  assign n22729 = n22728 ^ n22726;
  assign n22734 = n22733 ^ n22729;
  assign n25451 = n23427 ^ n22734;
  assign n25454 = n25453 ^ n25451;
  assign n25455 = n25454 ^ n25442;
  assign n25477 = n25476 ^ n25455;
  assign n25478 = ~n25457 & n25477;
  assign n22444 = ~n22394 & ~n22409;
  assign n22709 = n22447 ^ n22444;
  assign n22710 = n22709 ^ n22680;
  assign n22708 = n22436 ^ n22429;
  assign n22711 = n22710 ^ n22708;
  assign n25430 = n25429 ^ n22711;
  assign n24384 = n22733 ^ n22633;
  assign n22570 = n22000 & ~n22047;
  assign n22080 = n22079 ^ n22077;
  assign n22571 = n22570 ^ n22080;
  assign n22568 = n21999 & n22053;
  assign n22569 = n22568 ^ n22088;
  assign n22572 = n22571 ^ n22569;
  assign n22567 = n22075 ^ n22066;
  assign n22573 = n22572 ^ n22567;
  assign n22574 = n22573 ^ n22090;
  assign n25428 = n24384 ^ n22574;
  assign n25431 = n25430 ^ n25428;
  assign n22445 = n22381 & ~n22413;
  assign n22446 = n22445 ^ n22444;
  assign n22637 = n22584 ^ n22446;
  assign n22636 = n22434 ^ n22429;
  assign n22638 = n22637 ^ n22636;
  assign n25425 = n25424 ^ n22638;
  assign n22759 = n22629 ^ n22321;
  assign n22758 = n22624 ^ n22315;
  assign n22760 = n22759 ^ n22758;
  assign n24377 = n22760 ^ n22733;
  assign n22081 = n22080 ^ n22049;
  assign n22076 = n22075 ^ n22063;
  assign n22082 = n22081 ^ n22076;
  assign n22091 = n22090 ^ n22082;
  assign n25422 = n24377 ^ n22091;
  assign n22206 = n22205 ^ n22202;
  assign n22199 = n22133 & n22180;
  assign n22198 = n22152 & n22177;
  assign n22200 = n22199 ^ n22198;
  assign n22201 = n22200 ^ n22197;
  assign n22207 = n22206 ^ n22201;
  assign n22324 = n22323 ^ n22207;
  assign n25423 = n25422 ^ n22324;
  assign n25426 = n25425 ^ n25423;
  assign n22547 = n22546 ^ n22199;
  assign n22552 = n22551 ^ n22547;
  assign n22545 = n22544 ^ n22205;
  assign n22553 = n22552 ^ n22545;
  assign n22565 = n22564 ^ n22553;
  assign n25427 = n25426 ^ n22565;
  assign n25432 = n25431 ^ n25427;
  assign n22737 = n22435 ^ n22429;
  assign n22736 = n22681 ^ n22439;
  assign n22738 = n22737 ^ n22736;
  assign n25419 = n25418 ^ n22738;
  assign n22661 = n22007 & n22059;
  assign n22662 = n22661 ^ n22065;
  assign n22659 = n22085 ^ n22069;
  assign n22660 = n22659 ^ n22571;
  assign n22663 = n22662 ^ n22660;
  assign n23433 = n22676 ^ n22663;
  assign n22776 = n22543 ^ n22205;
  assign n22775 = n22727 ^ n22700;
  assign n22777 = n22776 ^ n22775;
  assign n22781 = n22780 ^ n22777;
  assign n25417 = n23433 ^ n22781;
  assign n25420 = n25419 ^ n25417;
  assign n25421 = n25420 ^ n25416;
  assign n25433 = n25432 ^ n25421;
  assign n25466 = n25433 & n25455;
  assign n25479 = n25478 ^ n25466;
  assign n25456 = n25455 ^ n25432;
  assign n25475 = n25456 ^ n25421;
  assign n25480 = n25479 ^ n25475;
  assign n25447 = n25446 ^ n25420;
  assign n22450 = n22449 ^ n22446;
  assign n22443 = n22442 ^ n22430;
  assign n22451 = n22450 ^ n22443;
  assign n25436 = n25435 ^ n22451;
  assign n23447 = n22733 ^ n22090;
  assign n22756 = n22618 ^ n22200;
  assign n22755 = n22613 ^ n22182;
  assign n22757 = n22756 ^ n22755;
  assign n22761 = n22760 ^ n22757;
  assign n25434 = n23447 ^ n22761;
  assign n25437 = n25436 ^ n25434;
  assign n25448 = n25447 ^ n25437;
  assign n25470 = n25448 ^ n25426;
  assign n25463 = n25454 ^ n25416;
  assign n25471 = n25470 ^ n25463;
  assign n25472 = n25456 ^ n25437;
  assign n25473 = n25471 & n25472;
  assign n25458 = n25454 ^ n25426;
  assign n25459 = n25458 ^ n25457;
  assign n25460 = ~n25456 & n25459;
  assign n25474 = n25473 ^ n25460;
  assign n25481 = n25480 ^ n25474;
  assign n25483 = n25476 ^ n25432;
  assign n25487 = ~n25458 & ~n25483;
  assign n25486 = n25426 & n25448;
  assign n25488 = n25487 ^ n25486;
  assign n25484 = n25483 ^ n25458;
  assign n25485 = n25484 ^ n25479;
  assign n25489 = n25488 ^ n25485;
  assign n25490 = n25481 & n25489;
  assign n25462 = n25456 ^ n25447;
  assign n25467 = n25462 & ~n25463;
  assign n25468 = n25467 ^ n25466;
  assign n25464 = n25463 ^ n25462;
  assign n25449 = n25448 ^ n25442;
  assign n25450 = ~n25437 & n25449;
  assign n25461 = n25460 ^ n25450;
  assign n25465 = n25464 ^ n25461;
  assign n25469 = n25468 ^ n25465;
  assign n25482 = n25481 ^ n25469;
  assign n25522 = n25490 ^ n25482;
  assign n25492 = n25483 ^ n25448;
  assign n25491 = n25455 ^ n25449;
  assign n25496 = n25492 ^ n25491;
  assign n25493 = n25491 & ~n25492;
  assign n25494 = n25493 ^ n25487;
  assign n25495 = n25494 ^ n25468;
  assign n25497 = n25496 ^ n25495;
  assign n25520 = n25469 & n25481;
  assign n25521 = ~n25497 & n25520;
  assign n25523 = n25522 ^ n25521;
  assign n25501 = n25497 ^ n25489;
  assign n25511 = n25501 ^ n25490;
  assign n25509 = ~n25469 & n25489;
  assign n25510 = n25497 & n25509;
  assign n25512 = n25511 ^ n25510;
  assign n25524 = n25523 ^ n25512;
  assign n25502 = n25490 ^ n25469;
  assign n25503 = ~n25501 & ~n25502;
  assign n25504 = n25503 ^ n25497;
  assign n25498 = n25497 ^ n25490;
  assign n25499 = ~n25482 & ~n25498;
  assign n25500 = n25499 ^ n25469;
  assign n25505 = n25504 ^ n25500;
  assign n25540 = n25524 ^ n25505;
  assign n25541 = ~n25457 & n25540;
  assign n25507 = n25455 & n25505;
  assign n25542 = n25541 ^ n25507;
  assign n25536 = n25471 & ~n25512;
  assign n25890 = n25542 ^ n25536;
  assign n25757 = n25477 & n25540;
  assign n25506 = n25433 & n25505;
  assign n25838 = n25757 ^ n25506;
  assign n25513 = n25512 ^ n25504;
  assign n25533 = n25459 & n25513;
  assign n25532 = n25472 & ~n25512;
  assign n25534 = n25533 ^ n25532;
  assign n25514 = ~n25456 & n25513;
  assign n25535 = n25534 ^ n25514;
  assign n25889 = n25838 ^ n25535;
  assign n25891 = n25890 ^ n25889;
  assign n25537 = n25448 & ~n25523;
  assign n25538 = n25537 ^ n25536;
  assign n25839 = n25838 ^ n25538;
  assign n25526 = n25523 ^ n25500;
  assign n25543 = ~n25483 & n25526;
  assign n25544 = n25543 ^ n25542;
  assign n25837 = n25544 ^ n25533;
  assign n25840 = n25839 ^ n25837;
  assign n25892 = n25891 ^ n25840;
  assign n21472 = n18641 ^ n18548;
  assign n21474 = n21473 ^ n21472;
  assign n21471 = n19659 ^ n18565;
  assign n21475 = n21474 ^ n21471;
  assign n21465 = n18615 ^ n17920;
  assign n21467 = n21466 ^ n21465;
  assign n21464 = n19654 ^ n18043;
  assign n21468 = n21467 ^ n21464;
  assign n21481 = n21475 ^ n21468;
  assign n21432 = n18513 ^ n18424;
  assign n21433 = n21432 ^ n18298;
  assign n21431 = n19661 ^ n18523;
  assign n21434 = n21433 ^ n21431;
  assign n21497 = n21475 ^ n21434;
  assign n20356 = n18646 ^ n18624;
  assign n21461 = n20356 ^ n19664;
  assign n21460 = n21459 ^ n18595;
  assign n21462 = n21461 ^ n21460;
  assign n20347 = n18624 ^ n18493;
  assign n21455 = n20347 ^ n19656;
  assign n21453 = n21441 ^ n18548;
  assign n21454 = n21453 ^ n18650;
  assign n21456 = n21455 ^ n21454;
  assign n21458 = n21457 ^ n21456;
  assign n21463 = n21462 ^ n21458;
  assign n21504 = n21497 ^ n21463;
  assign n21443 = n21442 ^ n21441;
  assign n21440 = n19671 ^ n18624;
  assign n21444 = n21443 ^ n21440;
  assign n21436 = n18424 ^ n17920;
  assign n21437 = n21436 ^ n18619;
  assign n21435 = n19668 ^ n18437;
  assign n21438 = n21437 ^ n21435;
  assign n21439 = n21438 ^ n21434;
  assign n21445 = n21444 ^ n21439;
  assign n21514 = n21504 ^ n21445;
  assign n20385 = n18624 ^ n18580;
  assign n21449 = n20385 ^ n19675;
  assign n21447 = n21446 ^ n18513;
  assign n21448 = n21447 ^ n18411;
  assign n21450 = n21449 ^ n21448;
  assign n21469 = n21468 ^ n21450;
  assign n21451 = n21450 ^ n21445;
  assign n21513 = n21469 ^ n21451;
  assign n21518 = n21514 ^ n21513;
  assign n21515 = ~n21513 & ~n21514;
  assign n21477 = n21468 ^ n21456;
  assign n21508 = ~n21477 & n21504;
  assign n21516 = n21515 ^ n21508;
  assign n21486 = n21475 ^ n21438;
  assign n21487 = n21486 ^ n21463;
  assign n21488 = n21469 & n21487;
  assign n21470 = n21469 ^ n21463;
  assign n21482 = n21470 ^ n21439;
  assign n21485 = n21481 & ~n21482;
  assign n21489 = n21488 ^ n21485;
  assign n21517 = n21516 ^ n21489;
  assign n21519 = n21518 ^ n21517;
  assign n21507 = ~n21445 & n21456;
  assign n21509 = n21508 ^ n21507;
  assign n21505 = n21504 ^ n21477;
  assign n21476 = n21475 ^ n21450;
  assign n21498 = n21497 ^ n21469;
  assign n21499 = n21476 & ~n21498;
  assign n21500 = n21499 ^ n21488;
  assign n21506 = n21505 ^ n21500;
  assign n21510 = n21509 ^ n21506;
  assign n21527 = n21519 ^ n21510;
  assign n21496 = n21486 ^ n21470;
  assign n21501 = n21500 ^ n21496;
  assign n21491 = n21456 ^ n21445;
  assign n21492 = n21491 ^ n21481;
  assign n21493 = n21470 ^ n21444;
  assign n21494 = n21492 & n21493;
  assign n21478 = n21477 ^ n21476;
  assign n21479 = ~n21470 & ~n21478;
  assign n21495 = n21494 ^ n21479;
  assign n21502 = n21501 ^ n21495;
  assign n21511 = n21502 & ~n21510;
  assign n21535 = n21527 ^ n21511;
  assign n21483 = n21482 ^ n21481;
  assign n21452 = ~n21444 & ~n21451;
  assign n21480 = n21479 ^ n21452;
  assign n21484 = n21483 ^ n21480;
  assign n21490 = n21489 ^ n21484;
  assign n21533 = ~n21490 & ~n21510;
  assign n21534 = ~n21519 & n21533;
  assign n21536 = n21535 ^ n21534;
  assign n21520 = n21490 & n21502;
  assign n21521 = n21519 & n21520;
  assign n21503 = n21502 ^ n21490;
  assign n21512 = n21511 ^ n21503;
  assign n21522 = n21521 ^ n21512;
  assign n21537 = n21536 ^ n21522;
  assign n21772 = n21481 & n21537;
  assign n21524 = n21519 ^ n21511;
  assign n21525 = ~n21503 & n21524;
  assign n21526 = n21525 ^ n21490;
  assign n21543 = n21526 ^ n21522;
  assign n21544 = ~n21477 & n21543;
  assign n21542 = ~n21482 & n21537;
  assign n21545 = n21544 ^ n21542;
  assign n21773 = n21772 ^ n21545;
  assign n21528 = n21511 ^ n21490;
  assign n21529 = ~n21527 & ~n21528;
  assign n21530 = n21529 ^ n21519;
  assign n21531 = n21530 ^ n21526;
  assign n21769 = n21487 & ~n21531;
  assign n21532 = n21469 & ~n21531;
  assign n21770 = n21769 ^ n21532;
  assign n21685 = n21536 ^ n21530;
  assign n21711 = ~n21470 & ~n21685;
  assign n21682 = ~n21444 & n21530;
  assign n21712 = n21711 ^ n21682;
  assign n21710 = ~n21513 & ~n21526;
  assign n21713 = n21712 ^ n21710;
  assign n21771 = n21770 ^ n21713;
  assign n21774 = n21773 ^ n21771;
  assign n21341 = n19856 ^ n19363;
  assign n21339 = n19530 ^ n19519;
  assign n21338 = n19550 ^ n19346;
  assign n21340 = n21339 ^ n21338;
  assign n21342 = n21341 ^ n21340;
  assign n21312 = n19959 ^ n19447;
  assign n20254 = n19475 ^ n19461;
  assign n21311 = n20254 ^ n19485;
  assign n21313 = n21312 ^ n21311;
  assign n21343 = n21342 ^ n21313;
  assign n21333 = n19902 ^ n19217;
  assign n20249 = n19419 ^ n19390;
  assign n21332 = n20249 ^ n19471;
  assign n21334 = n21333 ^ n21332;
  assign n21362 = n21342 ^ n21334;
  assign n21349 = n19405 ^ n19395;
  assign n20239 = n19441 ^ n19341;
  assign n21348 = n21347 ^ n20239;
  assign n21350 = n21349 ^ n21348;
  assign n21345 = n19765 ^ n19556;
  assign n21323 = n19652 ^ n19530;
  assign n20232 = n19491 ^ n19441;
  assign n21321 = n21320 ^ n20232;
  assign n21322 = n21321 ^ n19326;
  assign n21324 = n21323 ^ n21322;
  assign n21346 = n21345 ^ n21324;
  assign n21351 = n21350 ^ n21346;
  assign n21380 = n21362 ^ n21351;
  assign n21330 = n20010 ^ n19475;
  assign n20225 = n19217 ^ n18857;
  assign n21329 = n20225 ^ n19437;
  assign n21331 = n21330 ^ n21329;
  assign n21335 = n21334 ^ n21331;
  assign n21325 = n21320 ^ n19441;
  assign n21326 = n21325 ^ n19494;
  assign n21327 = n21326 ^ n19524;
  assign n21328 = n21327 ^ n19985;
  assign n21336 = n21335 ^ n21328;
  assign n21389 = n21380 ^ n21336;
  assign n21317 = n19932 ^ n19419;
  assign n20248 = n19542 ^ n19441;
  assign n21315 = n21314 ^ n20248;
  assign n21316 = n21315 ^ n19101;
  assign n21318 = n21317 ^ n21316;
  assign n21370 = n21336 ^ n21318;
  assign n21319 = n21318 ^ n21313;
  assign n21388 = n21370 ^ n21319;
  assign n21393 = n21389 ^ n21388;
  assign n21390 = ~n21388 & ~n21389;
  assign n21356 = n21324 ^ n21313;
  assign n21384 = ~n21356 & n21380;
  assign n21391 = n21390 ^ n21384;
  assign n21352 = n21351 ^ n21319;
  assign n21373 = n21352 ^ n21335;
  assign n21376 = n21343 & ~n21373;
  assign n21360 = n21342 ^ n21331;
  assign n21365 = n21360 ^ n21351;
  assign n21366 = n21319 & n21365;
  assign n21377 = n21376 ^ n21366;
  assign n21392 = n21391 ^ n21377;
  assign n21394 = n21393 ^ n21392;
  assign n21355 = n21342 ^ n21318;
  assign n21363 = n21362 ^ n21319;
  assign n21364 = n21355 & ~n21363;
  assign n21367 = n21366 ^ n21364;
  assign n21361 = n21360 ^ n21352;
  assign n21368 = n21367 ^ n21361;
  assign n21357 = n21356 ^ n21355;
  assign n21358 = ~n21352 & ~n21357;
  assign n21337 = n21336 ^ n21324;
  assign n21344 = n21343 ^ n21337;
  assign n21353 = n21352 ^ n21328;
  assign n21354 = n21344 & n21353;
  assign n21359 = n21358 ^ n21354;
  assign n21369 = n21368 ^ n21359;
  assign n21374 = n21373 ^ n21343;
  assign n21371 = ~n21328 & ~n21370;
  assign n21372 = n21371 ^ n21358;
  assign n21375 = n21374 ^ n21372;
  assign n21378 = n21377 ^ n21375;
  assign n21409 = n21369 & n21378;
  assign n21410 = n21394 & n21409;
  assign n21383 = n21324 & ~n21336;
  assign n21385 = n21384 ^ n21383;
  assign n21381 = n21380 ^ n21356;
  assign n21382 = n21381 ^ n21367;
  assign n21386 = n21385 ^ n21382;
  assign n21387 = n21369 & ~n21386;
  assign n21379 = n21378 ^ n21369;
  assign n21408 = n21387 ^ n21379;
  assign n21411 = n21410 ^ n21408;
  assign n21398 = n21394 ^ n21386;
  assign n21406 = n21398 ^ n21387;
  assign n21404 = ~n21378 & ~n21386;
  assign n21405 = ~n21394 & n21404;
  assign n21407 = n21406 ^ n21405;
  assign n21412 = n21411 ^ n21407;
  assign n21764 = n21343 & n21412;
  assign n21395 = n21394 ^ n21387;
  assign n21396 = ~n21379 & n21395;
  assign n21397 = n21396 ^ n21378;
  assign n21419 = n21411 ^ n21397;
  assign n21420 = ~n21356 & n21419;
  assign n21418 = ~n21373 & n21412;
  assign n21421 = n21420 ^ n21418;
  assign n21765 = n21764 ^ n21421;
  assign n21399 = n21387 ^ n21378;
  assign n21400 = ~n21398 & ~n21399;
  assign n21401 = n21400 ^ n21394;
  assign n21402 = n21401 ^ n21397;
  assign n21761 = n21365 & ~n21402;
  assign n21403 = n21319 & ~n21402;
  assign n21762 = n21761 ^ n21403;
  assign n21652 = n21407 ^ n21401;
  assign n21735 = ~n21352 & ~n21652;
  assign n21649 = ~n21328 & n21401;
  assign n21736 = n21735 ^ n21649;
  assign n21734 = ~n21388 & ~n21397;
  assign n21737 = n21736 ^ n21734;
  assign n21763 = n21762 ^ n21737;
  assign n21766 = n21765 ^ n21763;
  assign n24505 = n21774 ^ n21766;
  assign n20508 = n16637 ^ n16547;
  assign n21058 = n20508 ^ n14546;
  assign n21057 = n19379 ^ n16536;
  assign n21059 = n21058 ^ n21057;
  assign n20534 = n16727 ^ n16413;
  assign n21044 = n20534 ^ n16700;
  assign n21043 = n19452 ^ n15500;
  assign n21045 = n21044 ^ n21043;
  assign n21088 = n21059 ^ n21045;
  assign n21069 = n20525 ^ n16595;
  assign n21068 = n19479 ^ n16710;
  assign n21070 = n21069 ^ n21068;
  assign n21092 = n21070 ^ n21059;
  assign n21079 = n19561 ^ n16515;
  assign n20498 = n16724 ^ n16630;
  assign n21078 = n21077 ^ n20498;
  assign n21080 = n21079 ^ n21078;
  assign n21049 = n19534 ^ n16422;
  assign n20489 = n16724 ^ n16658;
  assign n21047 = n21046 ^ n20489;
  assign n21048 = n21047 ^ n20491;
  assign n21050 = n21049 ^ n21048;
  assign n20495 = n16682 ^ n16571;
  assign n21076 = n21050 ^ n20495;
  assign n21081 = n21080 ^ n21076;
  assign n21055 = n19426 ^ n16603;
  assign n20518 = n16724 ^ n16560;
  assign n21053 = n21052 ^ n20518;
  assign n21054 = n21053 ^ n20520;
  assign n21056 = n21055 ^ n21054;
  assign n21074 = n21056 ^ n21045;
  assign n21089 = n21081 ^ n21074;
  assign n21121 = n21092 ^ n21089;
  assign n21060 = n21059 ^ n21056;
  assign n21066 = n20503 ^ n16677;
  assign n21065 = n19302 ^ n16610;
  assign n21067 = n21066 ^ n21065;
  assign n21082 = n21067 ^ n21059;
  assign n21100 = n21082 ^ n21074;
  assign n21101 = n21060 & n21100;
  assign n21093 = n21092 ^ n21081;
  assign n21094 = ~n21074 & ~n21093;
  assign n21102 = n21101 ^ n21094;
  assign n21122 = n21121 ^ n21102;
  assign n21071 = n21070 ^ n21067;
  assign n20514 = n16661 ^ n16403;
  assign n21063 = n20514 ^ n16728;
  assign n21062 = n19509 ^ n15490;
  assign n21064 = n21063 ^ n21062;
  assign n21072 = n21071 ^ n21064;
  assign n21116 = n21072 ^ n21050;
  assign n21117 = n21116 ^ n21088;
  assign n21118 = n21089 ^ n21064;
  assign n21119 = n21117 & n21118;
  assign n21051 = n21050 ^ n21045;
  assign n21061 = n21060 ^ n21051;
  assign n21108 = n21061 & n21089;
  assign n21120 = n21119 ^ n21108;
  assign n21123 = n21122 ^ n21120;
  assign n21090 = n21089 ^ n21071;
  assign n21110 = n21090 ^ n21088;
  assign n21073 = n21072 ^ n21056;
  assign n21107 = n21064 & n21073;
  assign n21109 = n21108 ^ n21107;
  assign n21111 = n21110 ^ n21109;
  assign n21091 = ~n21088 & ~n21090;
  assign n21095 = n21094 ^ n21091;
  assign n21112 = n21111 ^ n21095;
  assign n21134 = n21123 ^ n21112;
  assign n21104 = ~n21050 & ~n21072;
  assign n21083 = n21082 ^ n21081;
  assign n21086 = n21051 & n21083;
  assign n21105 = n21104 ^ n21086;
  assign n21099 = n21083 ^ n21051;
  assign n21103 = n21102 ^ n21099;
  assign n21106 = n21105 ^ n21103;
  assign n21124 = n21106 & n21123;
  assign n21135 = n21134 ^ n21124;
  assign n21084 = n21083 ^ n21072;
  assign n21075 = n21074 ^ n21073;
  assign n21097 = n21084 ^ n21075;
  assign n21085 = ~n21075 & ~n21084;
  assign n21087 = n21086 ^ n21085;
  assign n21096 = n21095 ^ n21087;
  assign n21098 = n21097 ^ n21096;
  assign n21132 = ~n21112 & n21123;
  assign n21133 = n21098 & n21132;
  assign n21136 = n21135 ^ n21133;
  assign n21115 = n21106 ^ n21098;
  assign n21125 = n21124 ^ n21115;
  assign n21113 = n21106 & n21112;
  assign n21114 = ~n21098 & n21113;
  assign n21126 = n21125 ^ n21114;
  assign n21137 = n21136 ^ n21126;
  assign n21815 = ~n21088 & n21137;
  assign n21659 = ~n21090 & n21137;
  assign n21138 = n21124 ^ n21098;
  assign n21139 = n21134 & n21138;
  assign n21140 = n21139 ^ n21112;
  assign n21146 = n21140 ^ n21136;
  assign n21158 = n21051 & n21146;
  assign n21660 = n21659 ^ n21158;
  assign n21816 = n21815 ^ n21660;
  assign n21127 = n21124 ^ n21112;
  assign n21128 = n21115 & n21127;
  assign n21129 = n21128 ^ n21098;
  assign n21141 = n21140 ^ n21129;
  assign n21154 = ~n21093 & n21141;
  assign n21144 = ~n21074 & n21141;
  assign n21813 = n21154 ^ n21144;
  assign n21665 = ~n21075 & n21140;
  assign n21130 = n21129 ^ n21126;
  assign n21161 = n21089 & n21130;
  assign n21160 = n21064 & n21129;
  assign n21162 = n21161 ^ n21160;
  assign n21666 = n21665 ^ n21162;
  assign n21814 = n21813 ^ n21666;
  assign n21817 = n21816 ^ n21814;
  assign n25325 = n24505 ^ n21817;
  assign n25326 = n25325 ^ n20866;
  assign n21653 = ~n21357 & ~n21652;
  assign n21651 = n21353 & ~n21407;
  assign n21654 = n21653 ^ n21651;
  assign n21822 = n21735 ^ n21654;
  assign n21646 = n21344 & ~n21407;
  assign n21416 = ~n21336 & ~n21411;
  assign n21647 = n21646 ^ n21416;
  assign n21840 = n21822 ^ n21647;
  assign n21729 = n21380 & n21419;
  assign n21413 = n21412 ^ n21402;
  assign n21414 = n21355 & ~n21413;
  assign n21415 = n21414 ^ n21403;
  assign n21730 = n21729 ^ n21415;
  assign n21841 = n21840 ^ n21730;
  assign n21218 = n18503 ^ n17512;
  assign n21216 = n17497 ^ n16960;
  assign n21217 = n21216 ^ n21174;
  assign n21219 = n21218 ^ n21217;
  assign n20107 = n17702 ^ n16960;
  assign n21197 = n20107 ^ n17641;
  assign n21196 = n21195 ^ n17666;
  assign n21198 = n21197 ^ n21196;
  assign n21193 = n18586 ^ n17648;
  assign n21178 = n18571 ^ n17708;
  assign n20101 = n17545 ^ n16960;
  assign n21176 = n20101 ^ n17492;
  assign n21175 = n21174 ^ n17481;
  assign n21177 = n21176 ^ n21175;
  assign n21179 = n21178 ^ n21177;
  assign n21194 = n21193 ^ n21179;
  assign n21199 = n21198 ^ n21194;
  assign n21188 = n21187 ^ n21186;
  assign n20122 = n17662 ^ n16960;
  assign n21189 = n21188 ^ n20122;
  assign n21190 = n21189 ^ n17615;
  assign n21191 = n21190 ^ n18538;
  assign n21172 = n18629 ^ n17517;
  assign n21170 = n17569 ^ n17236;
  assign n21169 = n17563 ^ n17095;
  assign n21171 = n21170 ^ n21169;
  assign n21173 = n21172 ^ n21171;
  assign n21192 = n21191 ^ n21173;
  assign n21200 = n21199 ^ n21192;
  assign n21234 = n21219 ^ n21200;
  assign n21206 = n21205 ^ n17613;
  assign n21207 = n21206 ^ n17228;
  assign n21208 = n21207 ^ n18386;
  assign n21202 = n21201 ^ n17577;
  assign n21203 = n21202 ^ n17637;
  assign n21204 = n21203 ^ n18455;
  assign n21209 = n21208 ^ n21204;
  assign n21220 = n21219 ^ n21209;
  assign n21256 = ~n21179 & n21220;
  assign n21180 = n21179 ^ n21173;
  assign n21181 = n17681 ^ n17482;
  assign n21182 = n21181 ^ n17697;
  assign n21183 = n21182 ^ n17673;
  assign n21184 = n21183 ^ n18660;
  assign n21223 = n21204 ^ n21184;
  assign n21224 = n21223 ^ n21199;
  assign n21227 = n21180 & n21224;
  assign n21257 = n21256 ^ n21227;
  assign n21254 = n21224 ^ n21180;
  assign n21236 = n21191 ^ n21184;
  assign n21241 = n21223 ^ n21192;
  assign n21242 = n21236 & n21241;
  assign n21212 = n21208 ^ n21184;
  assign n21213 = n21212 ^ n21199;
  assign n21214 = n21192 & n21213;
  assign n21243 = n21242 ^ n21214;
  assign n21255 = n21254 ^ n21243;
  assign n21258 = n21257 ^ n21255;
  assign n21225 = n21224 ^ n21220;
  assign n21221 = n21220 ^ n21191;
  assign n21222 = n21221 ^ n21192;
  assign n21230 = n21225 ^ n21222;
  assign n21226 = n21222 & n21225;
  assign n21228 = n21227 ^ n21226;
  assign n21185 = n21184 ^ n21173;
  assign n21210 = n21209 ^ n21200;
  assign n21211 = n21185 & n21210;
  assign n21215 = n21214 ^ n21211;
  assign n21229 = n21228 ^ n21215;
  assign n21231 = n21230 ^ n21229;
  assign n21270 = n21258 ^ n21231;
  assign n21240 = n21212 ^ n21200;
  assign n21244 = n21243 ^ n21240;
  assign n21237 = n21236 ^ n21180;
  assign n21238 = n21200 & n21237;
  assign n21232 = n21220 ^ n21179;
  assign n21233 = n21232 ^ n21185;
  assign n21235 = n21233 & n21234;
  assign n21239 = n21238 ^ n21235;
  assign n21245 = n21244 ^ n21239;
  assign n21259 = n21245 & n21258;
  assign n21271 = n21270 ^ n21259;
  assign n21248 = n21210 ^ n21185;
  assign n21246 = n21219 & n21221;
  assign n21247 = n21246 ^ n21238;
  assign n21249 = n21248 ^ n21247;
  assign n21250 = n21249 ^ n21215;
  assign n21268 = n21250 & n21258;
  assign n21269 = ~n21231 & n21268;
  assign n21272 = n21271 ^ n21269;
  assign n21642 = n21234 & n21272;
  assign n21274 = n21259 ^ n21250;
  assign n21275 = n21270 & n21274;
  assign n21276 = n21275 ^ n21231;
  assign n21288 = n21276 ^ n21272;
  assign n21293 = n21237 & n21288;
  assign n21643 = n21642 ^ n21293;
  assign n21289 = n21200 & n21288;
  assign n21752 = n21643 ^ n21289;
  assign n21296 = n21233 & n21272;
  assign n21253 = n21250 ^ n21245;
  assign n21260 = n21259 ^ n21253;
  assign n21251 = n21245 & ~n21250;
  assign n21252 = n21231 & n21251;
  assign n21261 = n21260 ^ n21252;
  assign n21295 = n21220 & n21261;
  assign n21297 = n21296 ^ n21295;
  assign n21753 = n21752 ^ n21297;
  assign n21262 = n21259 ^ n21231;
  assign n21263 = n21253 & n21262;
  assign n21264 = n21263 ^ n21250;
  assign n21277 = n21276 ^ n21264;
  assign n21280 = n21192 & n21277;
  assign n21273 = n21272 ^ n21261;
  assign n21278 = n21277 ^ n21273;
  assign n21279 = n21236 & n21278;
  assign n21281 = n21280 ^ n21279;
  assign n21265 = n21264 ^ n21261;
  assign n21267 = n21224 & n21265;
  assign n21282 = n21281 ^ n21267;
  assign n21754 = n21753 ^ n21282;
  assign n21842 = n21841 ^ n21754;
  assign n25327 = n25326 ^ n21842;
  assign n21708 = ~n21451 & n21530;
  assign n21679 = n21492 & ~n21536;
  assign n21523 = ~n21445 & ~n21522;
  assign n21680 = n21679 ^ n21523;
  assign n21709 = n21708 ^ n21680;
  assign n21714 = n21713 ^ n21709;
  assign n21705 = n21504 & n21543;
  assign n21538 = n21537 ^ n21531;
  assign n21539 = n21476 & ~n21538;
  assign n21540 = n21539 ^ n21532;
  assign n21706 = n21705 ^ n21540;
  assign n21546 = ~n21498 & ~n21538;
  assign n21547 = n21546 ^ n21545;
  assign n21707 = n21706 ^ n21547;
  assign n21715 = n21714 ^ n21707;
  assign n21425 = ~n21389 & ~n21397;
  assign n21424 = n21337 & ~n21411;
  assign n21426 = n21425 ^ n21424;
  assign n21422 = ~n21363 & ~n21413;
  assign n21423 = n21422 ^ n21421;
  assign n21427 = n21426 ^ n21423;
  assign n21417 = n21416 ^ n21415;
  assign n21428 = n21427 ^ n21417;
  assign n21309 = n21295 ^ n21281;
  assign n21305 = n21210 & n21273;
  assign n21266 = n21180 & n21265;
  assign n21306 = n21305 ^ n21266;
  assign n21298 = n21241 & n21278;
  assign n21307 = n21306 ^ n21298;
  assign n21285 = n21225 & n21264;
  assign n21284 = n21232 & n21261;
  assign n21286 = n21285 ^ n21284;
  assign n21308 = n21307 ^ n21286;
  assign n21310 = n21309 ^ n21308;
  assign n21429 = n21428 ^ n21310;
  assign n25296 = n21715 ^ n21429;
  assign n21732 = ~n21370 & n21401;
  assign n21733 = n21732 ^ n21647;
  assign n21738 = n21737 ^ n21733;
  assign n21731 = n21730 ^ n21423;
  assign n21739 = n21738 ^ n21731;
  assign n25297 = n25296 ^ n21739;
  assign n21663 = n21073 & n21129;
  assign n21151 = n21117 & n21126;
  assign n21150 = ~n21072 & n21136;
  assign n21152 = n21151 ^ n21150;
  assign n21664 = n21663 ^ n21152;
  assign n21667 = n21666 ^ n21664;
  assign n21142 = n21141 ^ n21137;
  assign n21153 = n21100 & n21142;
  assign n21661 = n21660 ^ n21153;
  assign n21147 = n21083 & n21146;
  assign n21143 = n21060 & n21142;
  assign n21145 = n21144 ^ n21143;
  assign n21148 = n21147 ^ n21145;
  assign n21662 = n21661 ^ n21148;
  assign n21668 = n21667 ^ n21662;
  assign n25298 = n25297 ^ n21668;
  assign n25299 = n25298 ^ n20835;
  assign n25356 = n25327 ^ n25299;
  assign n21825 = n21646 ^ n21415;
  assign n21823 = n21761 ^ n21422;
  assign n21824 = n21823 ^ n21822;
  assign n21826 = n21825 ^ n21824;
  assign n21820 = n21296 ^ n21281;
  assign n21299 = n21213 & n21277;
  assign n21300 = n21299 ^ n21298;
  assign n21819 = n21752 ^ n21300;
  assign n21821 = n21820 ^ n21819;
  assign n21827 = n21826 ^ n21821;
  assign n21155 = n21154 ^ n21153;
  assign n21156 = n21155 ^ n21152;
  assign n21131 = n21061 & n21130;
  assign n21149 = n21148 ^ n21131;
  assign n21157 = n21156 ^ n21149;
  assign n25332 = n21827 ^ n21157;
  assign n21862 = n21823 ^ n21647;
  assign n21861 = n21730 ^ n21653;
  assign n21863 = n21862 ^ n21861;
  assign n21802 = n21769 ^ n21546;
  assign n21854 = n21802 ^ n21680;
  assign n21686 = ~n21478 & ~n21685;
  assign n21853 = n21706 ^ n21686;
  assign n21855 = n21854 ^ n21853;
  assign n24515 = n21863 ^ n21855;
  assign n25333 = n25332 ^ n24515;
  assign n25334 = n25333 ^ n20792;
  assign n21650 = n21649 ^ n21425;
  assign n21655 = n21654 ^ n21650;
  assign n21648 = n21647 ^ n21415;
  assign n21656 = n21655 ^ n21648;
  assign n24521 = n21863 ^ n21656;
  assign n21684 = n21493 & ~n21536;
  assign n21687 = n21686 ^ n21684;
  assign n21801 = n21711 ^ n21687;
  assign n21844 = n21801 ^ n21680;
  assign n21845 = n21844 ^ n21706;
  assign n24509 = n21845 ^ n21841;
  assign n25321 = n24521 ^ n24509;
  assign n21287 = n21219 & n21276;
  assign n21641 = n21287 ^ n21285;
  assign n21644 = n21643 ^ n21641;
  assign n21640 = n21297 ^ n21281;
  assign n21645 = n21644 ^ n21640;
  assign n21301 = n21300 ^ n21297;
  assign n21294 = n21293 ^ n21282;
  assign n21302 = n21301 ^ n21294;
  assign n21838 = n21645 ^ n21302;
  assign n25322 = n25321 ^ n21838;
  assign n21747 = n21118 & n21126;
  assign n21748 = n21747 ^ n21131;
  assign n21749 = n21748 ^ n21161;
  assign n21750 = n21749 ^ n21152;
  assign n21751 = n21750 ^ n21148;
  assign n25323 = n25322 ^ n21751;
  assign n25324 = n25323 ^ n20930;
  assign n25335 = n25334 ^ n25324;
  assign n25357 = n25356 ^ n25335;
  assign n25337 = n25324 ^ n25299;
  assign n25358 = n25337 & n25357;
  assign n21163 = ~n21084 & n21140;
  assign n21834 = n21163 ^ n21160;
  assign n21835 = n21834 ^ n21748;
  assign n21833 = n21152 ^ n21145;
  assign n21836 = n21835 ^ n21833;
  assign n21673 = n21222 & n21264;
  assign n21290 = n21289 ^ n21287;
  assign n21674 = n21673 ^ n21290;
  assign n21671 = n21221 & n21276;
  assign n21672 = n21671 ^ n21297;
  assign n21675 = n21674 ^ n21672;
  assign n21670 = n21307 ^ n21282;
  assign n21676 = n21675 ^ n21670;
  assign n21677 = n21676 ^ n21302;
  assign n25313 = n21836 ^ n21677;
  assign n24532 = n21863 ^ n21739;
  assign n25312 = n24532 ^ n21656;
  assign n25314 = n25313 ^ n25312;
  assign n21549 = ~n21514 & ~n21526;
  assign n21683 = n21682 ^ n21549;
  assign n21688 = n21687 ^ n21683;
  assign n21681 = n21680 ^ n21540;
  assign n21689 = n21688 ^ n21681;
  assign n25310 = n21689 ^ n20882;
  assign n21548 = n21491 & ~n21522;
  assign n21550 = n21549 ^ n21548;
  assign n21551 = n21550 ^ n21547;
  assign n21541 = n21540 ^ n21523;
  assign n21552 = n21551 ^ n21541;
  assign n25308 = n21552 ^ n20749;
  assign n21742 = n21150 ^ n21145;
  assign n21164 = ~n21116 & n21136;
  assign n21165 = n21164 ^ n21163;
  assign n21741 = n21661 ^ n21165;
  assign n21743 = n21742 ^ n21741;
  assign n21291 = n21290 ^ n21286;
  assign n21283 = n21282 ^ n21266;
  assign n21292 = n21291 ^ n21283;
  assign n21303 = n21302 ^ n21292;
  assign n25306 = n21743 ^ n21303;
  assign n21787 = n21736 ^ n21426;
  assign n21786 = n21730 ^ n21420;
  assign n21788 = n21787 ^ n21786;
  assign n24499 = n21863 ^ n21788;
  assign n25305 = n24499 ^ n21428;
  assign n25307 = n25306 ^ n25305;
  assign n25309 = n25308 ^ n25307;
  assign n25311 = n25310 ^ n25309;
  assign n25315 = n25314 ^ n25311;
  assign n21804 = n21679 ^ n21540;
  assign n21803 = n21802 ^ n21801;
  assign n21805 = n21804 ^ n21803;
  assign n25302 = n21805 ^ n20955;
  assign n21866 = n21151 ^ n21145;
  assign n21865 = n21749 ^ n21155;
  assign n21867 = n21866 ^ n21865;
  assign n21758 = n21185 & n21273;
  assign n21759 = n21758 ^ n21306;
  assign n21756 = n21299 ^ n21280;
  assign n21757 = n21756 ^ n21674;
  assign n21760 = n21759 ^ n21757;
  assign n21767 = n21766 ^ n21760;
  assign n25300 = n21867 ^ n21767;
  assign n25301 = n25300 ^ n21826;
  assign n25303 = n25302 ^ n25301;
  assign n25304 = n25303 ^ n25299;
  assign n25316 = n25315 ^ n25304;
  assign n25346 = n25316 & n25335;
  assign n25359 = n25358 ^ n25346;
  assign n25336 = n25335 ^ n25315;
  assign n25355 = n25336 ^ n25304;
  assign n25360 = n25359 ^ n25355;
  assign n25328 = n25327 ^ n25303;
  assign n21166 = n21165 ^ n21162;
  assign n21159 = n21158 ^ n21148;
  assign n21167 = n21166 ^ n21159;
  assign n25318 = n21302 ^ n21167;
  assign n25319 = n25318 ^ n24499;
  assign n21793 = n21712 ^ n21550;
  assign n21792 = n21706 ^ n21544;
  assign n21794 = n21793 ^ n21792;
  assign n25317 = n21794 ^ n20701;
  assign n25320 = n25319 ^ n25317;
  assign n25329 = n25328 ^ n25320;
  assign n25350 = n25329 ^ n25309;
  assign n25343 = n25334 ^ n25299;
  assign n25351 = n25350 ^ n25343;
  assign n25352 = n25336 ^ n25320;
  assign n25353 = n25351 & n25352;
  assign n25338 = n25334 ^ n25309;
  assign n25339 = n25338 ^ n25337;
  assign n25340 = n25336 & n25339;
  assign n25354 = n25353 ^ n25340;
  assign n25361 = n25360 ^ n25354;
  assign n25363 = n25356 ^ n25315;
  assign n25367 = n25338 & n25363;
  assign n25366 = ~n25309 & n25329;
  assign n25368 = n25367 ^ n25366;
  assign n25364 = n25363 ^ n25338;
  assign n25365 = n25364 ^ n25359;
  assign n25369 = n25368 ^ n25365;
  assign n25370 = n25361 & n25369;
  assign n25342 = n25336 ^ n25328;
  assign n25347 = n25342 & n25343;
  assign n25348 = n25347 ^ n25346;
  assign n25344 = n25343 ^ n25342;
  assign n25330 = n25329 ^ n25324;
  assign n25331 = n25320 & n25330;
  assign n25341 = n25340 ^ n25331;
  assign n25345 = n25344 ^ n25341;
  assign n25349 = n25348 ^ n25345;
  assign n25362 = n25361 ^ n25349;
  assign n25402 = n25370 ^ n25362;
  assign n25372 = n25363 ^ n25329;
  assign n25371 = n25335 ^ n25330;
  assign n25376 = n25372 ^ n25371;
  assign n25373 = n25371 & n25372;
  assign n25374 = n25373 ^ n25367;
  assign n25375 = n25374 ^ n25348;
  assign n25377 = n25376 ^ n25375;
  assign n25400 = ~n25349 & n25361;
  assign n25401 = n25377 & n25400;
  assign n25403 = n25402 ^ n25401;
  assign n25381 = n25377 ^ n25369;
  assign n25391 = n25381 ^ n25370;
  assign n25389 = n25349 & n25369;
  assign n25390 = ~n25377 & n25389;
  assign n25392 = n25391 ^ n25390;
  assign n25404 = n25403 ^ n25392;
  assign n25382 = n25370 ^ n25349;
  assign n25383 = n25381 & n25382;
  assign n25384 = n25383 ^ n25377;
  assign n25378 = n25377 ^ n25370;
  assign n25379 = n25362 & n25378;
  assign n25380 = n25379 ^ n25349;
  assign n25385 = n25384 ^ n25380;
  assign n25783 = n25404 ^ n25385;
  assign n25788 = n25357 & n25783;
  assign n25386 = n25316 & n25385;
  assign n25885 = n25788 ^ n25386;
  assign n25792 = n25329 & n25403;
  assign n25791 = n25351 & n25392;
  assign n25793 = n25792 ^ n25791;
  assign n25886 = n25885 ^ n25793;
  assign n25393 = n25392 ^ n25384;
  assign n25850 = n25339 & n25393;
  assign n25406 = n25403 ^ n25380;
  assign n25786 = n25363 & n25406;
  assign n25784 = n25337 & n25783;
  assign n25387 = n25335 & n25385;
  assign n25785 = n25784 ^ n25387;
  assign n25787 = n25786 ^ n25785;
  assign n25884 = n25850 ^ n25787;
  assign n25887 = n25886 ^ n25884;
  assign n20536 = n17458 ^ n16710;
  assign n20533 = n16724 ^ n16695;
  assign n20535 = n20534 ^ n20533;
  assign n20537 = n20536 ^ n20535;
  assign n20510 = n17714 ^ n16422;
  assign n20507 = n16630 ^ n13604;
  assign n20509 = n20508 ^ n20507;
  assign n20511 = n20510 ^ n20509;
  assign n20546 = n20537 ^ n20511;
  assign n20527 = n17595 ^ n16610;
  assign n20524 = n16695 ^ n16584;
  assign n20526 = n20525 ^ n20524;
  assign n20528 = n20527 ^ n20526;
  assign n20505 = n17627 ^ n16603;
  assign n20502 = n16673 ^ n16584;
  assign n20504 = n20503 ^ n20502;
  assign n20506 = n20505 ^ n20504;
  assign n20529 = n20528 ^ n20506;
  assign n20516 = n17554 ^ n15500;
  assign n20515 = n20514 ^ n20489;
  assign n20517 = n20516 ^ n20515;
  assign n20530 = n20529 ^ n20517;
  assign n20512 = n20511 ^ n20506;
  assign n20499 = n20498 ^ n16560;
  assign n20497 = n17687 ^ n16537;
  assign n20500 = n20499 ^ n20497;
  assign n20493 = n17529 ^ n15501;
  assign n20490 = n20489 ^ n13604;
  assign n20492 = n20491 ^ n20490;
  assign n20494 = n20493 ^ n20492;
  assign n20496 = n20495 ^ n20494;
  assign n20501 = n20500 ^ n20496;
  assign n20513 = n20512 ^ n20501;
  assign n20575 = n20530 ^ n20513;
  assign n20522 = n17652 ^ n16678;
  assign n20519 = n20518 ^ n16673;
  assign n20521 = n20520 ^ n20519;
  assign n20523 = n20522 ^ n20521;
  assign n20538 = n20537 ^ n20523;
  assign n20531 = n20530 ^ n20523;
  assign n20574 = n20538 ^ n20531;
  assign n20579 = n20575 ^ n20574;
  assign n20576 = ~n20574 & ~n20575;
  assign n20541 = n20537 ^ n20494;
  assign n20570 = n20513 & ~n20541;
  assign n20577 = n20576 ^ n20570;
  assign n20539 = n20538 ^ n20501;
  assign n20545 = n20539 ^ n20529;
  assign n20552 = ~n20545 & n20546;
  assign n20549 = n20528 ^ n20511;
  assign n20550 = n20549 ^ n20501;
  assign n20551 = n20538 & n20550;
  assign n20553 = n20552 ^ n20551;
  assign n20578 = n20577 ^ n20553;
  assign n20580 = n20579 ^ n20578;
  assign n20569 = n20494 & ~n20530;
  assign n20571 = n20570 ^ n20569;
  assign n20567 = n20541 ^ n20513;
  assign n20540 = n20523 ^ n20511;
  assign n20561 = n20538 ^ n20512;
  assign n20562 = n20540 & ~n20561;
  assign n20563 = n20562 ^ n20551;
  assign n20568 = n20567 ^ n20563;
  assign n20572 = n20571 ^ n20568;
  assign n20590 = n20580 ^ n20572;
  assign n20560 = n20549 ^ n20539;
  assign n20564 = n20563 ^ n20560;
  assign n20555 = n20530 ^ n20494;
  assign n20556 = n20555 ^ n20546;
  assign n20557 = n20539 ^ n20517;
  assign n20558 = n20556 & n20557;
  assign n20542 = n20541 ^ n20540;
  assign n20543 = ~n20539 & ~n20542;
  assign n20559 = n20558 ^ n20543;
  assign n20565 = n20564 ^ n20559;
  assign n20573 = n20565 & ~n20572;
  assign n20598 = n20590 ^ n20573;
  assign n20547 = n20546 ^ n20545;
  assign n20532 = ~n20517 & ~n20531;
  assign n20544 = n20543 ^ n20532;
  assign n20548 = n20547 ^ n20544;
  assign n20554 = n20553 ^ n20548;
  assign n20596 = ~n20554 & ~n20572;
  assign n20597 = ~n20580 & n20596;
  assign n20599 = n20598 ^ n20597;
  assign n20585 = n20554 & n20565;
  assign n20586 = n20580 & n20585;
  assign n20566 = n20565 ^ n20554;
  assign n20584 = n20573 ^ n20566;
  assign n20587 = n20586 ^ n20584;
  assign n20600 = n20599 ^ n20587;
  assign n20850 = n20546 & n20600;
  assign n20735 = ~n20545 & n20600;
  assign n20581 = n20580 ^ n20573;
  assign n20582 = ~n20566 & n20581;
  assign n20583 = n20582 ^ n20554;
  assign n20588 = n20587 ^ n20583;
  assign n20605 = ~n20541 & n20588;
  assign n20736 = n20735 ^ n20605;
  assign n20851 = n20850 ^ n20736;
  assign n20591 = n20573 ^ n20554;
  assign n20592 = ~n20590 & ~n20591;
  assign n20593 = n20592 ^ n20580;
  assign n20594 = n20593 ^ n20583;
  assign n20780 = n20550 & ~n20594;
  assign n20595 = n20538 & ~n20594;
  assign n20848 = n20780 ^ n20595;
  assign n20807 = ~n20574 & ~n20583;
  assign n20611 = n20599 ^ n20593;
  assign n20612 = ~n20539 & ~n20611;
  assign n20610 = ~n20517 & n20593;
  assign n20613 = n20612 ^ n20610;
  assign n20808 = n20807 ^ n20613;
  assign n20849 = n20848 ^ n20808;
  assign n20852 = n20851 ^ n20849;
  assign n25211 = n20852 ^ n19910;
  assign n20264 = n19447 ^ n18630;
  assign n20262 = n19462 ^ n19410;
  assign n20263 = n20262 ^ n19441;
  assign n20265 = n20264 ^ n20263;
  assign n20221 = n19520 ^ n19363;
  assign n20222 = n20221 ^ n19341;
  assign n20223 = n20222 ^ n19550;
  assign n20224 = n20223 ^ n18661;
  assign n20274 = n20265 ^ n20224;
  assign n20235 = n19530 ^ n18572;
  assign n20233 = n20232 ^ n19519;
  assign n20231 = n19521 ^ n19325;
  assign n20234 = n20233 ^ n20231;
  assign n20236 = n20235 ^ n20234;
  assign n20255 = n20254 ^ n18974;
  assign n20256 = n20255 ^ n19436;
  assign n20257 = n20256 ^ n18387;
  assign n20226 = n20225 ^ n19470;
  assign n20227 = n20226 ^ n19391;
  assign n20228 = n20227 ^ n18456;
  assign n20258 = n20257 ^ n20228;
  assign n20246 = n19502 ^ n18504;
  assign n20244 = n19524 ^ n19399;
  assign n20245 = n20244 ^ n20232;
  assign n20247 = n20246 ^ n20245;
  assign n20259 = n20258 ^ n20247;
  assign n20305 = n20236 & ~n20259;
  assign n20240 = n20239 ^ n19542;
  assign n20238 = n19545 ^ n19405;
  assign n20241 = n20240 ^ n20238;
  assign n20230 = n19556 ^ n18587;
  assign n20237 = n20236 ^ n20230;
  assign n20242 = n20241 ^ n20237;
  assign n20229 = n20228 ^ n20224;
  assign n20243 = n20242 ^ n20229;
  assign n20269 = n20265 ^ n20236;
  assign n20298 = n20243 & ~n20269;
  assign n20306 = n20305 ^ n20298;
  assign n20303 = n20269 ^ n20243;
  assign n20250 = n20249 ^ n20248;
  assign n20251 = n20250 ^ n19400;
  assign n20252 = n20251 ^ n19086;
  assign n20253 = n20252 ^ n18539;
  assign n20268 = n20253 ^ n20224;
  assign n20266 = n20265 ^ n20253;
  assign n20289 = n20266 ^ n20229;
  assign n20290 = n20268 & ~n20289;
  assign n20278 = n20257 ^ n20224;
  assign n20279 = n20278 ^ n20242;
  assign n20280 = n20266 & n20279;
  assign n20291 = n20290 ^ n20280;
  assign n20304 = n20303 ^ n20291;
  assign n20307 = n20306 ^ n20304;
  assign n20296 = n20259 ^ n20243;
  assign n20260 = n20259 ^ n20253;
  assign n20295 = n20266 ^ n20260;
  assign n20301 = n20296 ^ n20295;
  assign n20297 = ~n20295 & ~n20296;
  assign n20299 = n20298 ^ n20297;
  assign n20267 = n20266 ^ n20242;
  assign n20273 = n20267 ^ n20258;
  assign n20277 = ~n20273 & n20274;
  assign n20281 = n20280 ^ n20277;
  assign n20300 = n20299 ^ n20281;
  assign n20302 = n20301 ^ n20300;
  assign n20318 = n20307 ^ n20302;
  assign n20288 = n20278 ^ n20267;
  assign n20292 = n20291 ^ n20288;
  assign n20283 = n20259 ^ n20236;
  assign n20284 = n20283 ^ n20274;
  assign n20285 = n20267 ^ n20247;
  assign n20286 = n20284 & n20285;
  assign n20270 = n20269 ^ n20268;
  assign n20271 = ~n20267 & ~n20270;
  assign n20287 = n20286 ^ n20271;
  assign n20293 = n20292 ^ n20287;
  assign n20308 = n20293 & ~n20307;
  assign n20326 = n20318 ^ n20308;
  assign n20275 = n20274 ^ n20273;
  assign n20261 = ~n20247 & ~n20260;
  assign n20272 = n20271 ^ n20261;
  assign n20276 = n20275 ^ n20272;
  assign n20282 = n20281 ^ n20276;
  assign n20324 = ~n20282 & ~n20307;
  assign n20325 = ~n20302 & n20324;
  assign n20327 = n20326 ^ n20325;
  assign n20313 = n20282 & n20293;
  assign n20314 = n20302 & n20313;
  assign n20294 = n20293 ^ n20282;
  assign n20312 = n20308 ^ n20294;
  assign n20315 = n20314 ^ n20312;
  assign n20328 = n20327 ^ n20315;
  assign n20939 = n20274 & n20328;
  assign n20797 = ~n20273 & n20328;
  assign n20309 = n20308 ^ n20302;
  assign n20310 = ~n20294 & n20309;
  assign n20311 = n20310 ^ n20282;
  assign n20316 = n20315 ^ n20311;
  assign n20705 = ~n20269 & n20316;
  assign n20798 = n20797 ^ n20705;
  assign n20940 = n20939 ^ n20798;
  assign n20319 = n20308 ^ n20282;
  assign n20320 = ~n20318 & ~n20319;
  assign n20321 = n20320 ^ n20302;
  assign n20322 = n20321 ^ n20311;
  assign n20339 = n20279 & ~n20322;
  assign n20323 = n20266 & ~n20322;
  assign n20937 = n20339 ^ n20323;
  assign n20888 = ~n20295 & ~n20311;
  assign n20333 = n20327 ^ n20321;
  assign n20711 = ~n20267 & ~n20333;
  assign n20710 = ~n20247 & n20321;
  assign n20712 = n20711 ^ n20710;
  assign n20889 = n20888 ^ n20712;
  assign n20938 = n20937 ^ n20889;
  assign n20941 = n20940 ^ n20938;
  assign n20129 = n19453 ^ n17517;
  assign n20128 = n20127 ^ n17096;
  assign n20130 = n20129 ^ n20128;
  assign n20114 = n19380 ^ n17681;
  assign n20113 = n20112 ^ n17703;
  assign n20115 = n20114 ^ n20113;
  assign n20139 = n20130 ^ n20115;
  assign n20104 = n19535 ^ n17708;
  assign n20102 = n20101 ^ n17498;
  assign n20103 = n20102 ^ n17482;
  assign n20105 = n20104 ^ n20103;
  assign n20149 = n19510 ^ n17512;
  assign n20148 = n20147 ^ n17546;
  assign n20150 = n20149 ^ n20148;
  assign n20134 = n19480 ^ n17356;
  assign n20133 = n20132 ^ n17570;
  assign n20135 = n20134 ^ n20133;
  assign n20118 = n19303 ^ n17588;
  assign n20117 = n20116 ^ n17613;
  assign n20119 = n20118 ^ n20117;
  assign n20141 = n20135 ^ n20119;
  assign n20151 = n20150 ^ n20141;
  assign n20184 = n20105 & ~n20151;
  assign n20120 = n20119 ^ n20115;
  assign n20109 = n19562 ^ n17648;
  assign n20108 = n20107 ^ n17674;
  assign n20110 = n20109 ^ n20108;
  assign n20106 = n20105 ^ n17667;
  assign n20111 = n20110 ^ n20106;
  assign n20121 = n20120 ^ n20111;
  assign n20145 = n20130 ^ n20105;
  assign n20146 = ~n20121 & ~n20145;
  assign n20185 = n20184 ^ n20146;
  assign n20182 = n20145 ^ n20121;
  assign n20125 = n19427 ^ n17619;
  assign n20123 = n20122 ^ n17642;
  assign n20124 = n20123 ^ n17637;
  assign n20126 = n20125 ^ n20124;
  assign n20160 = n20126 ^ n20115;
  assign n20131 = n20130 ^ n20126;
  assign n20169 = n20131 ^ n20120;
  assign n20170 = n20160 & ~n20169;
  assign n20136 = n20135 ^ n20115;
  assign n20137 = n20136 ^ n20111;
  assign n20138 = n20131 & n20137;
  assign n20171 = n20170 ^ n20138;
  assign n20183 = n20182 ^ n20171;
  assign n20186 = n20185 ^ n20183;
  assign n20154 = n20151 ^ n20121;
  assign n20152 = n20151 ^ n20126;
  assign n20153 = n20152 ^ n20131;
  assign n20158 = n20154 ^ n20153;
  assign n20155 = ~n20153 & n20154;
  assign n20156 = n20155 ^ n20146;
  assign n20140 = n20131 ^ n20111;
  assign n20142 = n20141 ^ n20140;
  assign n20143 = n20139 & ~n20142;
  assign n20144 = n20143 ^ n20138;
  assign n20157 = n20156 ^ n20144;
  assign n20159 = n20158 ^ n20157;
  assign n20197 = n20186 ^ n20159;
  assign n20168 = n20140 ^ n20136;
  assign n20172 = n20171 ^ n20168;
  assign n20163 = n20151 ^ n20105;
  assign n20164 = n20163 ^ n20139;
  assign n20165 = n20150 ^ n20140;
  assign n20166 = n20164 & n20165;
  assign n20161 = n20160 ^ n20145;
  assign n20162 = n20140 & ~n20161;
  assign n20167 = n20166 ^ n20162;
  assign n20173 = n20172 ^ n20167;
  assign n20187 = n20173 & n20186;
  assign n20198 = n20197 ^ n20187;
  assign n20176 = n20142 ^ n20139;
  assign n20174 = n20150 & ~n20152;
  assign n20175 = n20174 ^ n20162;
  assign n20177 = n20176 ^ n20175;
  assign n20178 = n20177 ^ n20144;
  assign n20195 = ~n20178 & n20186;
  assign n20196 = n20159 & n20195;
  assign n20199 = n20198 ^ n20196;
  assign n20181 = n20178 ^ n20173;
  assign n20188 = n20187 ^ n20181;
  assign n20179 = n20173 & n20178;
  assign n20180 = ~n20159 & n20179;
  assign n20189 = n20188 ^ n20180;
  assign n20200 = n20199 ^ n20189;
  assign n20840 = n20139 & n20200;
  assign n20716 = ~n20142 & n20200;
  assign n20190 = n20187 ^ n20159;
  assign n20191 = ~n20181 & ~n20190;
  assign n20192 = n20191 ^ n20178;
  assign n20193 = n20192 ^ n20189;
  assign n20210 = ~n20145 & n20193;
  assign n20717 = n20716 ^ n20210;
  assign n20841 = n20840 ^ n20717;
  assign n20201 = n20187 ^ n20178;
  assign n20202 = ~n20197 & ~n20201;
  assign n20203 = n20202 ^ n20159;
  assign n20204 = n20203 ^ n20192;
  assign n20770 = n20137 & n20204;
  assign n20207 = n20131 & n20204;
  assign n20838 = n20770 ^ n20207;
  assign n20823 = ~n20153 & ~n20192;
  assign n20216 = n20203 ^ n20199;
  assign n20217 = n20140 & n20216;
  assign n20215 = n20150 & ~n20203;
  assign n20218 = n20217 ^ n20215;
  assign n20824 = n20823 ^ n20218;
  assign n20839 = n20838 ^ n20824;
  assign n20842 = n20841 ^ n20839;
  assign n23730 = n20941 ^ n20842;
  assign n20872 = n20557 & ~n20599;
  assign n20776 = ~n20542 & ~n20611;
  assign n20873 = n20872 ^ n20776;
  assign n20912 = n20873 ^ n20612;
  assign n20778 = n20556 & ~n20599;
  assign n20733 = ~n20530 & ~n20587;
  assign n20779 = n20778 ^ n20733;
  assign n20913 = n20912 ^ n20779;
  assign n20601 = n20600 ^ n20594;
  assign n20602 = n20540 & ~n20601;
  assign n20603 = n20602 ^ n20595;
  assign n20589 = n20513 & n20588;
  assign n20604 = n20603 ^ n20589;
  assign n20914 = n20913 ^ n20604;
  assign n20397 = n20396 ^ n18624;
  assign n20395 = n20394 ^ n18162;
  assign n20398 = n20397 ^ n20395;
  assign n20390 = n20389 ^ n18523;
  assign n20386 = n20385 ^ n18529;
  assign n20388 = n20387 ^ n20386;
  assign n20391 = n20390 ^ n20388;
  assign n20399 = n20398 ^ n20391;
  assign n20357 = n20356 ^ n18609;
  assign n20355 = n18595 ^ n18518;
  assign n20358 = n20357 ^ n20355;
  assign n20352 = n20351 ^ n18565;
  assign n20348 = n20347 ^ n18470;
  assign n20350 = n20349 ^ n20348;
  assign n20353 = n20352 ^ n20350;
  assign n20346 = n20345 ^ n18580;
  assign n20354 = n20353 ^ n20346;
  assign n20359 = n20358 ^ n20354;
  assign n20400 = n20399 ^ n20359;
  assign n20373 = n20347 ^ n18469;
  assign n20374 = n20373 ^ n18553;
  assign n20375 = n20374 ^ n18478;
  assign n20377 = n20376 ^ n20375;
  assign n20418 = n20400 ^ n20377;
  assign n20381 = n20380 ^ n18043;
  assign n20379 = n20378 ^ n18438;
  assign n20382 = n20381 ^ n20379;
  assign n20363 = n20362 ^ n18437;
  assign n20361 = n20360 ^ n18524;
  assign n20364 = n20363 ^ n20361;
  assign n20383 = n20382 ^ n20364;
  assign n20384 = n20383 ^ n20377;
  assign n20369 = n20368 ^ n18646;
  assign n20366 = n18565 ^ n18559;
  assign n20365 = n18641 ^ n18601;
  assign n20367 = n20366 ^ n20365;
  assign n20370 = n20369 ^ n20367;
  assign n20371 = n20370 ^ n20364;
  assign n20372 = n20371 ^ n20359;
  assign n20436 = n20384 ^ n20372;
  assign n20392 = n20391 ^ n20384;
  assign n20435 = n20399 ^ n20392;
  assign n20440 = n20436 ^ n20435;
  assign n20437 = ~n20435 & ~n20436;
  assign n20402 = n20398 ^ n20353;
  assign n20431 = n20372 & ~n20402;
  assign n20438 = n20437 ^ n20431;
  assign n20411 = n20382 ^ n20370;
  assign n20412 = n20411 ^ n20359;
  assign n20413 = n20399 & n20412;
  assign n20406 = n20400 ^ n20383;
  assign n20407 = n20398 ^ n20370;
  assign n20410 = ~n20406 & n20407;
  assign n20414 = n20413 ^ n20410;
  assign n20439 = n20438 ^ n20414;
  assign n20441 = n20440 ^ n20439;
  assign n20430 = n20353 & ~n20384;
  assign n20432 = n20431 ^ n20430;
  assign n20428 = n20402 ^ n20372;
  assign n20401 = n20391 ^ n20370;
  assign n20422 = n20399 ^ n20371;
  assign n20423 = n20401 & ~n20422;
  assign n20424 = n20423 ^ n20413;
  assign n20429 = n20428 ^ n20424;
  assign n20433 = n20432 ^ n20429;
  assign n20451 = n20441 ^ n20433;
  assign n20421 = n20411 ^ n20400;
  assign n20425 = n20424 ^ n20421;
  assign n20416 = n20384 ^ n20353;
  assign n20417 = n20416 ^ n20407;
  assign n20419 = n20417 & n20418;
  assign n20403 = n20402 ^ n20401;
  assign n20404 = ~n20400 & ~n20403;
  assign n20420 = n20419 ^ n20404;
  assign n20426 = n20425 ^ n20420;
  assign n20434 = n20426 & ~n20433;
  assign n20458 = n20451 ^ n20434;
  assign n20408 = n20407 ^ n20406;
  assign n20393 = ~n20377 & ~n20392;
  assign n20405 = n20404 ^ n20393;
  assign n20409 = n20408 ^ n20405;
  assign n20415 = n20414 ^ n20409;
  assign n20456 = ~n20415 & ~n20433;
  assign n20457 = ~n20441 & n20456;
  assign n20459 = n20458 ^ n20457;
  assign n20753 = n20418 & ~n20459;
  assign n20452 = n20434 ^ n20415;
  assign n20453 = ~n20451 & ~n20452;
  assign n20454 = n20453 ^ n20441;
  assign n20472 = n20459 ^ n20454;
  assign n20477 = ~n20403 & ~n20472;
  assign n20754 = n20753 ^ n20477;
  assign n20473 = ~n20400 & ~n20472;
  assign n20755 = n20754 ^ n20473;
  assign n20446 = n20415 & n20426;
  assign n20447 = n20441 & n20446;
  assign n20427 = n20426 ^ n20415;
  assign n20445 = n20434 ^ n20427;
  assign n20448 = n20447 ^ n20445;
  assign n20483 = ~n20384 & ~n20448;
  assign n20482 = n20417 & ~n20459;
  assign n20484 = n20483 ^ n20482;
  assign n20857 = n20755 ^ n20484;
  assign n20442 = n20441 ^ n20434;
  assign n20443 = ~n20427 & n20442;
  assign n20444 = n20443 ^ n20415;
  assign n20455 = n20454 ^ n20444;
  assign n20463 = n20399 & ~n20455;
  assign n20460 = n20459 ^ n20448;
  assign n20461 = n20460 ^ n20455;
  assign n20462 = n20401 & ~n20461;
  assign n20464 = n20463 ^ n20462;
  assign n20449 = n20448 ^ n20444;
  assign n20450 = n20372 & n20449;
  assign n20465 = n20464 ^ n20450;
  assign n20858 = n20857 ^ n20465;
  assign n20915 = n20914 ^ n20858;
  assign n25210 = n23730 ^ n20915;
  assign n25212 = n25211 ^ n25210;
  assign n20805 = ~n20531 & n20593;
  assign n20806 = n20805 ^ n20779;
  assign n20809 = n20808 ^ n20806;
  assign n20737 = ~n20561 & ~n20601;
  assign n20738 = n20737 ^ n20736;
  assign n20804 = n20738 ^ n20604;
  assign n20810 = n20809 ^ n20804;
  assign n25184 = n20810 ^ n19869;
  assign n20608 = ~n20575 & ~n20583;
  assign n20607 = n20555 & ~n20587;
  assign n20609 = n20608 ^ n20607;
  assign n20739 = n20738 ^ n20609;
  assign n20734 = n20733 ^ n20603;
  assign n20740 = n20739 ^ n20734;
  assign n20726 = ~n20406 & n20460;
  assign n20466 = ~n20402 & n20449;
  assign n20727 = n20726 ^ n20466;
  assign n20479 = ~n20422 & ~n20461;
  assign n20728 = n20727 ^ n20479;
  assign n20469 = n20416 & ~n20448;
  assign n20468 = ~n20436 & ~n20444;
  assign n20470 = n20469 ^ n20468;
  assign n20729 = n20728 ^ n20470;
  assign n20725 = n20483 ^ n20464;
  assign n20730 = n20729 ^ n20725;
  assign n25182 = n20740 ^ n20730;
  assign n20329 = n20328 ^ n20322;
  assign n20340 = ~n20289 & ~n20329;
  assign n20799 = n20798 ^ n20340;
  assign n20330 = n20268 & ~n20329;
  assign n20331 = n20330 ^ n20323;
  assign n20317 = n20243 & n20316;
  assign n20332 = n20331 ^ n20317;
  assign n20891 = n20799 ^ n20332;
  assign n20886 = ~n20260 & n20321;
  assign n20337 = n20284 & ~n20327;
  assign n20336 = ~n20259 & ~n20315;
  assign n20338 = n20337 ^ n20336;
  assign n20887 = n20886 ^ n20338;
  assign n20890 = n20889 ^ n20887;
  assign n20892 = n20891 ^ n20890;
  assign n20821 = ~n20152 & ~n20203;
  assign n20768 = n20164 & ~n20199;
  assign n20721 = ~n20151 & ~n20189;
  assign n20769 = n20768 ^ n20721;
  assign n20822 = n20821 ^ n20769;
  assign n20825 = n20824 ^ n20822;
  assign n20205 = n20204 ^ n20200;
  assign n20718 = ~n20169 & n20205;
  assign n20719 = n20718 ^ n20717;
  assign n20206 = n20160 & n20205;
  assign n20208 = n20207 ^ n20206;
  assign n20194 = ~n20121 & n20193;
  assign n20209 = n20208 ^ n20194;
  assign n20820 = n20719 ^ n20209;
  assign n20826 = n20825 ^ n20820;
  assign n25181 = n20892 ^ n20826;
  assign n25183 = n25182 ^ n25181;
  assign n25185 = n25184 ^ n25183;
  assign n25219 = n25212 ^ n25185;
  assign n20781 = n20780 ^ n20737;
  assign n20782 = n20781 ^ n20779;
  assign n20777 = n20776 ^ n20604;
  assign n20783 = n20782 ^ n20777;
  assign n25206 = n20783 ^ n19965;
  assign n20771 = n20770 ^ n20718;
  assign n20772 = n20771 ^ n20769;
  assign n20766 = ~n20161 & n20216;
  assign n20767 = n20766 ^ n20209;
  assign n20773 = n20772 ^ n20767;
  assign n20341 = n20340 ^ n20339;
  assign n20342 = n20341 ^ n20338;
  assign n20334 = ~n20270 & ~n20333;
  assign n20335 = n20334 ^ n20332;
  assign n20343 = n20342 ^ n20335;
  assign n23718 = n20773 ^ n20343;
  assign n20944 = n20778 ^ n20603;
  assign n20943 = n20912 ^ n20781;
  assign n20945 = n20944 ^ n20943;
  assign n20757 = n20482 ^ n20464;
  assign n20480 = n20412 & ~n20455;
  assign n20481 = n20480 ^ n20479;
  assign n20756 = n20755 ^ n20481;
  assign n20758 = n20757 ^ n20756;
  assign n20946 = n20945 ^ n20758;
  assign n25205 = n23718 ^ n20946;
  assign n25207 = n25206 ^ n25205;
  assign n25203 = n20914 ^ n19937;
  assign n20871 = n20610 ^ n20608;
  assign n20874 = n20873 ^ n20871;
  assign n20870 = n20779 ^ n20603;
  assign n20875 = n20874 ^ n20870;
  assign n24618 = n20875 ^ n20783;
  assign n20471 = ~n20377 & n20454;
  assign n20902 = n20471 ^ n20468;
  assign n20903 = n20902 ^ n20754;
  assign n20901 = n20484 ^ n20464;
  assign n20904 = n20903 ^ n20901;
  assign n20485 = n20484 ^ n20481;
  assign n20478 = n20477 ^ n20465;
  assign n20486 = n20485 ^ n20478;
  assign n20911 = n20904 ^ n20486;
  assign n25201 = n24618 ^ n20911;
  assign n20896 = n20165 & ~n20199;
  assign n20897 = n20896 ^ n20766;
  assign n20923 = n20897 ^ n20217;
  assign n20924 = n20923 ^ n20769;
  assign n20925 = n20924 ^ n20209;
  assign n20759 = n20285 & ~n20327;
  assign n20760 = n20759 ^ n20334;
  assign n20761 = n20760 ^ n20711;
  assign n20855 = n20761 ^ n20338;
  assign n20856 = n20855 ^ n20332;
  assign n23739 = n20925 ^ n20856;
  assign n25202 = n25201 ^ n23739;
  assign n25204 = n25203 ^ n25202;
  assign n25208 = n25207 ^ n25204;
  assign n25236 = n25219 ^ n25208;
  assign n20614 = n20613 ^ n20609;
  assign n20606 = n20605 ^ n20604;
  assign n20615 = n20614 ^ n20606;
  assign n24624 = n20783 ^ n20615;
  assign n25221 = n24624 ^ n20486;
  assign n20708 = ~n20296 & ~n20311;
  assign n20707 = n20283 & ~n20315;
  assign n20709 = n20708 ^ n20707;
  assign n20713 = n20712 ^ n20709;
  assign n20706 = n20705 ^ n20332;
  assign n20714 = n20713 ^ n20706;
  assign n25222 = n25221 ^ n20714;
  assign n20213 = n20154 & ~n20192;
  assign n20212 = n20163 & ~n20189;
  assign n20214 = n20213 ^ n20212;
  assign n20219 = n20218 ^ n20214;
  assign n20211 = n20210 ^ n20209;
  assign n20220 = n20219 ^ n20211;
  assign n25223 = n25222 ^ n20220;
  assign n25224 = n25223 ^ n19990;
  assign n25187 = n20945 ^ n20015;
  assign n20949 = n20768 ^ n20208;
  assign n20948 = n20923 ^ n20771;
  assign n20950 = n20949 ^ n20948;
  assign n20763 = n20337 ^ n20331;
  assign n20762 = n20761 ^ n20341;
  assign n20764 = n20763 ^ n20762;
  assign n23690 = n20950 ^ n20764;
  assign n20845 = n20407 & n20460;
  assign n20846 = n20845 ^ n20727;
  assign n20843 = n20480 ^ n20463;
  assign n20815 = ~n20435 & ~n20444;
  assign n20474 = n20473 ^ n20471;
  assign n20816 = n20815 ^ n20474;
  assign n20844 = n20843 ^ n20816;
  assign n20847 = n20846 ^ n20844;
  assign n20853 = n20852 ^ n20847;
  assign n25186 = n23690 ^ n20853;
  assign n25188 = n25187 ^ n25186;
  assign n25213 = n25212 ^ n25188;
  assign n25225 = n25224 ^ n25213;
  assign n25227 = n25225 ^ n25204;
  assign n25228 = n25227 ^ n25208;
  assign n24628 = n20810 ^ n20783;
  assign n20813 = ~n20392 & n20454;
  assign n20814 = n20813 ^ n20484;
  assign n20817 = n20816 ^ n20814;
  assign n20812 = n20728 ^ n20465;
  assign n20818 = n20817 ^ n20812;
  assign n20905 = n20818 ^ n20486;
  assign n25197 = n24628 ^ n20905;
  assign n20919 = n20338 ^ n20331;
  assign n20917 = n20710 ^ n20708;
  assign n20918 = n20917 ^ n20760;
  assign n20920 = n20919 ^ n20918;
  assign n20895 = n20215 ^ n20213;
  assign n20898 = n20897 ^ n20895;
  assign n20894 = n20769 ^ n20208;
  assign n20899 = n20898 ^ n20894;
  assign n25196 = n20920 ^ n20899;
  assign n25198 = n25197 ^ n25196;
  assign n25193 = n20740 ^ n19754;
  assign n20475 = n20474 ^ n20470;
  assign n20467 = n20466 ^ n20465;
  assign n20476 = n20475 ^ n20467;
  assign n20487 = n20486 ^ n20476;
  assign n25191 = n24624 ^ n20487;
  assign n20801 = n20336 ^ n20331;
  assign n20800 = n20799 ^ n20709;
  assign n20802 = n20801 ^ n20800;
  assign n20722 = n20721 ^ n20208;
  assign n20720 = n20719 ^ n20214;
  assign n20723 = n20722 ^ n20720;
  assign n23725 = n20802 ^ n20723;
  assign n25192 = n25191 ^ n23725;
  assign n25194 = n25193 ^ n25192;
  assign n25190 = n20875 ^ n19778;
  assign n25195 = n25194 ^ n25190;
  assign n25199 = n25198 ^ n25195;
  assign n25220 = n25219 ^ n25199;
  assign n25226 = n25225 ^ n25220;
  assign n25234 = n25228 ^ n25226;
  assign n25230 = n25207 ^ n25194;
  assign n25231 = n25220 & ~n25230;
  assign n25229 = ~n25226 & ~n25228;
  assign n25232 = n25231 ^ n25229;
  assign n25189 = n25188 ^ n25185;
  assign n25200 = n25199 ^ n25189;
  assign n25217 = n25200 & n25208;
  assign n25209 = n25208 ^ n25199;
  assign n25214 = n25213 ^ n25209;
  assign n25215 = n25207 ^ n25185;
  assign n25216 = ~n25214 & n25215;
  assign n25218 = n25217 ^ n25216;
  assign n25233 = n25232 ^ n25218;
  assign n25235 = n25234 ^ n25233;
  assign n25250 = n25215 ^ n25214;
  assign n25237 = n25204 ^ n25185;
  assign n25247 = n25237 ^ n25230;
  assign n25248 = ~n25209 & ~n25247;
  assign n25246 = ~n25224 & ~n25227;
  assign n25249 = n25248 ^ n25246;
  assign n25251 = n25250 ^ n25249;
  assign n25252 = n25251 ^ n25218;
  assign n25258 = n25209 ^ n25189;
  assign n25238 = ~n25236 & n25237;
  assign n25239 = n25238 ^ n25217;
  assign n25259 = n25258 ^ n25239;
  assign n25253 = n25224 ^ n25209;
  assign n25254 = n25225 ^ n25194;
  assign n25255 = n25254 ^ n25215;
  assign n25256 = n25253 & n25255;
  assign n25257 = n25256 ^ n25248;
  assign n25260 = n25259 ^ n25257;
  assign n25285 = n25252 & n25260;
  assign n25286 = n25235 & n25285;
  assign n25265 = n25260 ^ n25252;
  assign n25242 = n25194 & ~n25225;
  assign n25243 = n25242 ^ n25231;
  assign n25240 = n25230 ^ n25220;
  assign n25241 = n25240 ^ n25239;
  assign n25244 = n25243 ^ n25241;
  assign n25261 = ~n25244 & n25260;
  assign n25284 = n25265 ^ n25261;
  assign n25287 = n25286 ^ n25284;
  assign n25245 = n25244 ^ n25235;
  assign n25275 = n25261 ^ n25245;
  assign n25273 = ~n25244 & ~n25252;
  assign n25274 = ~n25235 & n25273;
  assign n25276 = n25275 ^ n25274;
  assign n25288 = n25287 ^ n25276;
  assign n25266 = n25261 ^ n25235;
  assign n25267 = ~n25265 & n25266;
  assign n25268 = n25267 ^ n25252;
  assign n25262 = n25261 ^ n25252;
  assign n25263 = ~n25245 & ~n25262;
  assign n25264 = n25263 ^ n25235;
  assign n25269 = n25268 ^ n25264;
  assign n25774 = n25288 ^ n25269;
  assign n25779 = ~n25236 & ~n25774;
  assign n25270 = n25200 & ~n25269;
  assign n25881 = n25779 ^ n25270;
  assign n25769 = ~n25225 & ~n25287;
  assign n25768 = n25255 & ~n25276;
  assign n25770 = n25769 ^ n25768;
  assign n25882 = n25881 ^ n25770;
  assign n25277 = n25276 ^ n25264;
  assign n25844 = ~n25247 & ~n25277;
  assign n25290 = n25287 ^ n25268;
  assign n25777 = n25220 & n25290;
  assign n25775 = n25237 & ~n25774;
  assign n25271 = n25208 & ~n25269;
  assign n25776 = n25775 ^ n25271;
  assign n25778 = n25777 ^ n25776;
  assign n25880 = n25844 ^ n25778;
  assign n25883 = n25882 ^ n25880;
  assign n25888 = n25887 ^ n25883;
  assign n25893 = n25892 ^ n25888;
  assign n25906 = n25905 ^ n25893;
  assign n25824 = ~n25698 & ~n25720;
  assign n25825 = n25824 ^ n25823;
  assign n25819 = n25818 ^ n22650;
  assign n25738 = ~n25702 & n25737;
  assign n25736 = n25667 & n25735;
  assign n25739 = n25738 ^ n25736;
  assign n25813 = n25812 ^ n25739;
  assign n25729 = ~n25699 & n25728;
  assign n25723 = n25435 & ~n25720;
  assign n25722 = n25666 & ~n25721;
  assign n25724 = n25723 ^ n25722;
  assign n25730 = n25729 ^ n25724;
  assign n25814 = n25813 ^ n25730;
  assign n25820 = n25819 ^ n25814;
  assign n25826 = n25825 ^ n25820;
  assign n25827 = n25826 ^ n22651;
  assign n25828 = n25827 ^ n22652;
  assign n25829 = n25828 ^ n22653;
  assign n25639 = ~n25564 & ~n25638;
  assign n25809 = n25661 ^ n25639;
  assign n25804 = ~n25587 & n25658;
  assign n25654 = n25653 ^ n25638;
  assign n25803 = ~n25595 & n25654;
  assign n25805 = n25804 ^ n25803;
  assign n25807 = n25806 ^ n25805;
  assign n25801 = n25565 & ~n25638;
  assign n25800 = ~n25599 & ~n25653;
  assign n25802 = n25801 ^ n25800;
  assign n25808 = n25807 ^ n25802;
  assign n25810 = n25809 ^ n25808;
  assign n25830 = n25829 ^ n25810;
  assign n25794 = n25330 & n25384;
  assign n25795 = n25794 ^ n25793;
  assign n25397 = n25371 & n25380;
  assign n25395 = n25320 & n25384;
  assign n25394 = n25336 & n25393;
  assign n25396 = n25395 ^ n25394;
  assign n25398 = n25397 ^ n25396;
  assign n25796 = n25795 ^ n25398;
  assign n25408 = n25342 & n25404;
  assign n25407 = n25338 & n25406;
  assign n25409 = n25408 ^ n25407;
  assign n25789 = n25788 ^ n25409;
  assign n25790 = n25789 ^ n25787;
  assign n25797 = n25796 ^ n25790;
  assign n25292 = ~n25214 & n25288;
  assign n25291 = ~n25230 & n25290;
  assign n25293 = n25292 ^ n25291;
  assign n25780 = n25779 ^ n25293;
  assign n25781 = n25780 ^ n25778;
  assign n25771 = ~n25227 & n25264;
  assign n25772 = n25771 ^ n25770;
  assign n25281 = ~n25228 & ~n25268;
  assign n25279 = ~n25224 & n25264;
  assign n25278 = ~n25209 & ~n25277;
  assign n25280 = n25279 ^ n25278;
  assign n25282 = n25281 ^ n25280;
  assign n25773 = n25772 ^ n25282;
  assign n25782 = n25781 ^ n25773;
  assign n25798 = n25797 ^ n25782;
  assign n25763 = n25449 & ~n25504;
  assign n25764 = n25763 ^ n25538;
  assign n25517 = n25491 & ~n25500;
  assign n25515 = ~n25437 & ~n25504;
  assign n25516 = n25515 ^ n25514;
  assign n25518 = n25517 ^ n25516;
  assign n25765 = n25764 ^ n25518;
  assign n25528 = n25462 & n25524;
  assign n25527 = ~n25458 & n25526;
  assign n25529 = n25528 ^ n25527;
  assign n25758 = n25757 ^ n25529;
  assign n25762 = n25758 ^ n25544;
  assign n25766 = n25765 ^ n25762;
  assign n25760 = n25542 ^ n25537;
  assign n25755 = ~n25470 & ~n25523;
  assign n25754 = ~n25492 & ~n25500;
  assign n25756 = n25755 ^ n25754;
  assign n25759 = n25758 ^ n25756;
  assign n25761 = n25760 ^ n25759;
  assign n25767 = n25766 ^ n25761;
  assign n25799 = n25798 ^ n25767;
  assign n25831 = n25830 ^ n25799;
  assign n26032 = n25906 ^ n25831;
  assign n25965 = n25822 ^ n25816;
  assign n25962 = n25697 & n25728;
  assign n25961 = ~n25686 & n25734;
  assign n25963 = n25962 ^ n25961;
  assign n25964 = n25963 ^ n25813;
  assign n25966 = n25965 ^ n25964;
  assign n25967 = n25966 ^ n22537;
  assign n25968 = n25967 ^ n22538;
  assign n25969 = n25968 ^ n22539;
  assign n25970 = n25969 ^ n22540;
  assign n25862 = ~n25554 & n25643;
  assign n25921 = n25862 ^ n25645;
  assign n25958 = n25921 ^ n25802;
  assign n25655 = n25594 & n25654;
  assign n25662 = n25661 ^ n25655;
  assign n25957 = n25803 ^ n25662;
  assign n25959 = n25958 ^ n25957;
  assign n25640 = n25639 ^ n25633;
  assign n25860 = n25859 ^ n25640;
  assign n25857 = n25662 ^ n25646;
  assign n25861 = n25860 ^ n25857;
  assign n25960 = n25959 ^ n25861;
  assign n25971 = n25970 ^ n25960;
  assign n25953 = n25792 ^ n25785;
  assign n25950 = n25372 & n25380;
  assign n25949 = n25350 & n25403;
  assign n25951 = n25950 ^ n25949;
  assign n25952 = n25951 ^ n25789;
  assign n25954 = n25953 ^ n25952;
  assign n25947 = n25776 ^ n25769;
  assign n25944 = ~n25226 & ~n25268;
  assign n25943 = n25254 & ~n25287;
  assign n25945 = n25944 ^ n25943;
  assign n25946 = n25945 ^ n25780;
  assign n25948 = n25947 ^ n25946;
  assign n25955 = n25954 ^ n25948;
  assign n25939 = n25756 ^ n25516;
  assign n25938 = n25544 ^ n25527;
  assign n25940 = n25939 ^ n25938;
  assign n25941 = n25940 ^ n25840;
  assign n25942 = n25941 ^ n25761;
  assign n25956 = n25955 ^ n25942;
  assign n25972 = n25971 ^ n25956;
  assign n26005 = n25972 ^ n25906;
  assign n25994 = n25962 ^ n25723;
  assign n25992 = n25816 ^ n22604;
  assign n25868 = n25685 & n25717;
  assign n25870 = n25869 ^ n25868;
  assign n25991 = n25870 ^ n25823;
  assign n25993 = n25992 ^ n25991;
  assign n25995 = n25994 ^ n25993;
  assign n25996 = n25995 ^ n22605;
  assign n25997 = n25996 ^ n22606;
  assign n25998 = n25997 ^ n22607;
  assign n25988 = n25807 ^ n25662;
  assign n25985 = ~n25597 & n25643;
  assign n25986 = n25985 ^ n25640;
  assign n25922 = ~n25598 & ~n25653;
  assign n25923 = n25922 ^ n25921;
  assign n25987 = n25986 ^ n25923;
  assign n25989 = n25988 ^ n25987;
  assign n25990 = n25989 ^ n25861;
  assign n25999 = n25998 ^ n25990;
  assign n25983 = n25840 ^ n25766;
  assign n25834 = n25754 ^ n25515;
  assign n25835 = n25834 ^ n25534;
  assign n25833 = n25542 ^ n25538;
  assign n25836 = n25835 ^ n25833;
  assign n25984 = n25983 ^ n25836;
  assign n26000 = n25999 ^ n25984;
  assign n25978 = n25950 ^ n25395;
  assign n25849 = n25352 & n25392;
  assign n25851 = n25850 ^ n25849;
  assign n25979 = n25978 ^ n25851;
  assign n25977 = n25793 ^ n25785;
  assign n25980 = n25979 ^ n25977;
  assign n25975 = n25776 ^ n25770;
  assign n25973 = n25944 ^ n25279;
  assign n25843 = n25253 & ~n25276;
  assign n25845 = n25844 ^ n25843;
  assign n25974 = n25973 ^ n25845;
  assign n25976 = n25975 ^ n25974;
  assign n25981 = n25980 ^ n25976;
  assign n25982 = n25981 ^ n25972;
  assign n26001 = n26000 ^ n25982;
  assign n25747 = n25746 ^ n25745;
  assign n25741 = ~n25687 & n25737;
  assign n25742 = n25741 ^ n22690;
  assign n25740 = n25739 ^ n25730;
  assign n25743 = n25742 ^ n25740;
  assign n25748 = n25747 ^ n25743;
  assign n25749 = n25748 ^ n22691;
  assign n25750 = n25749 ^ n22692;
  assign n25751 = n25750 ^ n22693;
  assign n25650 = n25649 ^ n25640;
  assign n25663 = n25662 ^ n25650;
  assign n25752 = n25751 ^ n25663;
  assign n25539 = n25538 ^ n25535;
  assign n25545 = n25544 ^ n25539;
  assign n25525 = ~n25463 & n25524;
  assign n25530 = n25529 ^ n25525;
  assign n25508 = n25507 ^ n25506;
  assign n25519 = n25518 ^ n25508;
  assign n25531 = n25530 ^ n25519;
  assign n25546 = n25545 ^ n25531;
  assign n25405 = n25343 & n25404;
  assign n25410 = n25409 ^ n25405;
  assign n25388 = n25387 ^ n25386;
  assign n25399 = n25398 ^ n25388;
  assign n25411 = n25410 ^ n25399;
  assign n25289 = n25215 & n25288;
  assign n25294 = n25293 ^ n25289;
  assign n25272 = n25271 ^ n25270;
  assign n25283 = n25282 ^ n25272;
  assign n25295 = n25294 ^ n25283;
  assign n25412 = n25411 ^ n25295;
  assign n25547 = n25546 ^ n25412;
  assign n25753 = n25752 ^ n25547;
  assign n25832 = n25831 ^ n25753;
  assign n26006 = n26001 ^ n25832;
  assign n26029 = ~n26005 & n26006;
  assign n26019 = n25963 ^ n25724;
  assign n26018 = n25818 ^ n25736;
  assign n26020 = n26019 ^ n26018;
  assign n26021 = n26020 ^ n22766;
  assign n26022 = n26021 ^ n22767;
  assign n26023 = n26022 ^ n22768;
  assign n26024 = n26023 ^ n22769;
  assign n26025 = n26024 ^ n25861;
  assign n26014 = n25951 ^ n25396;
  assign n26013 = n25787 ^ n25407;
  assign n26015 = n26014 ^ n26013;
  assign n26011 = n25945 ^ n25280;
  assign n26010 = n25778 ^ n25291;
  assign n26012 = n26011 ^ n26010;
  assign n26016 = n26015 ^ n26012;
  assign n26017 = n26016 ^ n25941;
  assign n26026 = n26025 ^ n26017;
  assign n25929 = n25821 ^ n25816;
  assign n25871 = n25870 ^ n25722;
  assign n25928 = n25898 ^ n25871;
  assign n25930 = n25929 ^ n25928;
  assign n25931 = n25930 ^ n22791;
  assign n25932 = n25931 ^ n22792;
  assign n25933 = n25932 ^ n22793;
  assign n25934 = n25933 ^ n22794;
  assign n25925 = n25574 & n25658;
  assign n25926 = n25925 ^ n25805;
  assign n25920 = n25858 ^ n25657;
  assign n25924 = n25923 ^ n25920;
  assign n25927 = n25926 ^ n25924;
  assign n25935 = n25934 ^ n25927;
  assign n25918 = n25891 ^ n25531;
  assign n25915 = n25791 ^ n25785;
  assign n25852 = n25851 ^ n25394;
  assign n25914 = n25885 ^ n25852;
  assign n25916 = n25915 ^ n25914;
  assign n25912 = n25776 ^ n25768;
  assign n25846 = n25845 ^ n25278;
  assign n25911 = n25881 ^ n25846;
  assign n25913 = n25912 ^ n25911;
  assign n25917 = n25916 ^ n25913;
  assign n25919 = n25918 ^ n25917;
  assign n25936 = n25935 ^ n25919;
  assign n26009 = n25936 ^ n25753;
  assign n26027 = n26026 ^ n26009;
  assign n26028 = n25972 & ~n26027;
  assign n26030 = n26029 ^ n26028;
  assign n26007 = n26006 ^ n26005;
  assign n25873 = n25818 ^ n22716;
  assign n25872 = n25871 ^ n25823;
  assign n25874 = n25873 ^ n25872;
  assign n25875 = n25874 ^ n22717;
  assign n25876 = n25875 ^ n22718;
  assign n25877 = n25876 ^ n22719;
  assign n25865 = n25661 ^ n25640;
  assign n25863 = n25862 ^ n25800;
  assign n25864 = n25863 ^ n25648;
  assign n25866 = n25865 ^ n25864;
  assign n25867 = n25866 ^ n25861;
  assign n25878 = n25877 ^ n25867;
  assign n25853 = n25852 ^ n25793;
  assign n25854 = n25853 ^ n25787;
  assign n25847 = n25846 ^ n25770;
  assign n25848 = n25847 ^ n25778;
  assign n25855 = n25854 ^ n25848;
  assign n25841 = n25840 ^ n25836;
  assign n25842 = n25841 ^ n25545;
  assign n25856 = n25855 ^ n25842;
  assign n25879 = n25878 ^ n25856;
  assign n25907 = n25906 ^ n25879;
  assign n25937 = n25936 ^ n25831;
  assign n26002 = n26001 ^ n25937;
  assign n26003 = n25907 & n26002;
  assign n25908 = n25907 ^ n25832;
  assign n25909 = n25879 ^ n25831;
  assign n25910 = ~n25908 & n25909;
  assign n26004 = n26003 ^ n25910;
  assign n26008 = n26007 ^ n26004;
  assign n26031 = n26030 ^ n26008;
  assign n26033 = n26001 ^ n25907;
  assign n26058 = n26033 ^ n25937;
  assign n26059 = n26058 ^ n26004;
  assign n26053 = n26027 ^ n25972;
  assign n26054 = n26053 ^ n26032;
  assign n26055 = n26033 ^ n26026;
  assign n26056 = n26054 & n26055;
  assign n26047 = n26005 ^ n25909;
  assign n26048 = ~n26033 & ~n26047;
  assign n26057 = n26056 ^ n26048;
  assign n26060 = n26059 ^ n26057;
  assign n26061 = ~n26031 & n26060;
  assign n26039 = n26027 ^ n26006;
  assign n26037 = n26027 ^ n25879;
  assign n26038 = n26037 ^ n25907;
  assign n26043 = n26039 ^ n26038;
  assign n26040 = ~n26038 & ~n26039;
  assign n26041 = n26040 ^ n26029;
  assign n26034 = n26033 ^ n26009;
  assign n26035 = n26032 & ~n26034;
  assign n26036 = n26035 ^ n26003;
  assign n26042 = n26041 ^ n26036;
  assign n26044 = n26043 ^ n26042;
  assign n26045 = n26044 ^ n26031;
  assign n26076 = n26061 ^ n26045;
  assign n26050 = n26034 ^ n26032;
  assign n26046 = ~n26026 & ~n26037;
  assign n26049 = n26048 ^ n26046;
  assign n26051 = n26050 ^ n26049;
  assign n26052 = n26051 ^ n26036;
  assign n26074 = ~n26031 & ~n26052;
  assign n26075 = ~n26044 & n26074;
  assign n26077 = n26076 ^ n26075;
  assign n26071 = n26052 & n26060;
  assign n26072 = n26044 & n26071;
  assign n26065 = n26060 ^ n26052;
  assign n26070 = n26065 ^ n26061;
  assign n26073 = n26072 ^ n26070;
  assign n26078 = n26077 ^ n26073;
  assign n26424 = n26032 & n26078;
  assign n26066 = n26061 ^ n26044;
  assign n26067 = ~n26065 & n26066;
  assign n26068 = n26067 ^ n26052;
  assign n26082 = n26073 ^ n26068;
  assign n26083 = ~n26005 & n26082;
  assign n26081 = ~n26034 & n26078;
  assign n26084 = n26083 ^ n26081;
  assign n26425 = n26424 ^ n26084;
  assign n26062 = n26061 ^ n26052;
  assign n26063 = ~n26045 & ~n26062;
  assign n26064 = n26063 ^ n26044;
  assign n26069 = n26068 ^ n26064;
  assign n26355 = n26002 & ~n26069;
  assign n26088 = n25907 & ~n26069;
  assign n26422 = n26355 ^ n26088;
  assign n26100 = ~n26026 & n26064;
  assign n26098 = n26077 ^ n26064;
  assign n26099 = ~n26033 & ~n26098;
  assign n26101 = n26100 ^ n26099;
  assign n26097 = ~n26038 & ~n26068;
  assign n26102 = n26101 ^ n26097;
  assign n26423 = n26422 ^ n26102;
  assign n26426 = n26425 ^ n26423;
  assign n26433 = n26432 ^ n26426;
  assign n24649 = n22691 ^ n20914;
  assign n24647 = n20925 ^ n20842;
  assign n20942 = n20941 ^ n20847;
  assign n24648 = n24647 ^ n20942;
  assign n24650 = n24649 ^ n24648;
  assign n24640 = n22651 ^ n20740;
  assign n24638 = n20826 ^ n20723;
  assign n23724 = n20892 ^ n20818;
  assign n24639 = n24638 ^ n23724;
  assign n24641 = n24640 ^ n24639;
  assign n24658 = n24650 ^ n24641;
  assign n24619 = n24618 ^ n22717;
  assign n23695 = n20899 ^ n20773;
  assign n24616 = n23695 ^ n20925;
  assign n20859 = n20858 ^ n20856;
  assign n24617 = n24616 ^ n20859;
  assign n24620 = n24619 ^ n24617;
  assign n24614 = n22744 ^ n20945;
  assign n24612 = n20950 ^ n20773;
  assign n23689 = n20486 ^ n20343;
  assign n24613 = n24612 ^ n23689;
  assign n24615 = n24614 ^ n24613;
  assign n24621 = n24620 ^ n24615;
  assign n24672 = n24658 ^ n24621;
  assign n24645 = n22792 ^ n20852;
  assign n24643 = n20950 ^ n20842;
  assign n20765 = n20764 ^ n20758;
  assign n24644 = n24643 ^ n20765;
  assign n24646 = n24645 ^ n24644;
  assign n24651 = n24650 ^ n24646;
  assign n24635 = n22767 ^ n20783;
  assign n23717 = n20714 ^ n20476;
  assign n23702 = n20773 ^ n20220;
  assign n24634 = n23717 ^ n23702;
  assign n24636 = n24635 ^ n24634;
  assign n24660 = n24651 ^ n24636;
  assign n24662 = n24660 ^ n24620;
  assign n24663 = n24662 ^ n24621;
  assign n23710 = n20826 ^ n20773;
  assign n24630 = n23710 ^ n20899;
  assign n24629 = n24628 ^ n22605;
  assign n24631 = n24630 ^ n24629;
  assign n24625 = n24624 ^ n22538;
  assign n24622 = n23702 ^ n20723;
  assign n20803 = n20802 ^ n20730;
  assign n24623 = n24622 ^ n20803;
  assign n24626 = n24625 ^ n24623;
  assign n23708 = n20920 ^ n20904;
  assign n24627 = n24626 ^ n23708;
  assign n24632 = n24631 ^ n24627;
  assign n24659 = n24658 ^ n24632;
  assign n24661 = n24660 ^ n24659;
  assign n24669 = n24663 ^ n24661;
  assign n24665 = n24626 ^ n24615;
  assign n24666 = n24659 & ~n24665;
  assign n24664 = ~n24661 & ~n24663;
  assign n24667 = n24666 ^ n24664;
  assign n24654 = n24646 ^ n24641;
  assign n24655 = n24654 ^ n24632;
  assign n24656 = n24621 & n24655;
  assign n24642 = n24641 ^ n24615;
  assign n24633 = n24632 ^ n24621;
  assign n24652 = n24651 ^ n24633;
  assign n24653 = n24642 & ~n24652;
  assign n24657 = n24656 ^ n24653;
  assign n24668 = n24667 ^ n24657;
  assign n24670 = n24669 ^ n24668;
  assign n24684 = n24652 ^ n24642;
  assign n24671 = n24641 ^ n24620;
  assign n24681 = n24671 ^ n24665;
  assign n24682 = ~n24633 & ~n24681;
  assign n24680 = ~n24636 & ~n24662;
  assign n24683 = n24682 ^ n24680;
  assign n24685 = n24684 ^ n24683;
  assign n24686 = n24685 ^ n24657;
  assign n24693 = n24654 ^ n24633;
  assign n24673 = n24671 & ~n24672;
  assign n24674 = n24673 ^ n24656;
  assign n24694 = n24693 ^ n24674;
  assign n24637 = n24636 ^ n24633;
  assign n24689 = n24660 ^ n24626;
  assign n24690 = n24689 ^ n24642;
  assign n24691 = n24637 & n24690;
  assign n24692 = n24691 ^ n24682;
  assign n24695 = n24694 ^ n24692;
  assign n24712 = n24686 & n24695;
  assign n24713 = n24670 & n24712;
  assign n24710 = n24695 ^ n24686;
  assign n24677 = n24626 & ~n24660;
  assign n24678 = n24677 ^ n24666;
  assign n24675 = n24665 ^ n24659;
  assign n24676 = n24675 ^ n24674;
  assign n24679 = n24678 ^ n24676;
  assign n24696 = ~n24679 & n24695;
  assign n24711 = n24710 ^ n24696;
  assign n24714 = n24713 ^ n24711;
  assign n24697 = n24679 ^ n24670;
  assign n24698 = n24697 ^ n24696;
  assign n24687 = ~n24679 & ~n24686;
  assign n24688 = ~n24670 & n24687;
  assign n24699 = n24698 ^ n24688;
  assign n24723 = n24714 ^ n24699;
  assign n24718 = n24696 ^ n24670;
  assign n24719 = ~n24710 & n24718;
  assign n24720 = n24719 ^ n24686;
  assign n24701 = n24696 ^ n24686;
  assign n24702 = ~n24697 & ~n24701;
  assign n24703 = n24702 ^ n24670;
  assign n24721 = n24720 ^ n24703;
  assign n24724 = n24723 ^ n24721;
  assign n24870 = ~n24672 & ~n24724;
  assign n24733 = n24655 & ~n24721;
  assign n24918 = n24870 ^ n24733;
  assign n24715 = ~n24660 & ~n24714;
  assign n24709 = n24690 & ~n24699;
  assign n24716 = n24715 ^ n24709;
  assign n24919 = n24918 ^ n24716;
  assign n24727 = n24720 ^ n24714;
  assign n24728 = n24659 & n24727;
  assign n24725 = n24671 & ~n24724;
  assign n24722 = n24621 & ~n24721;
  assign n24726 = n24725 ^ n24722;
  assign n24729 = n24728 ^ n24726;
  assign n24704 = n24703 ^ n24699;
  assign n24705 = ~n24681 & ~n24704;
  assign n24917 = n24729 ^ n24705;
  assign n24920 = n24919 ^ n24917;
  assign n24983 = n24982 ^ n24920;
  assign n24524 = n21845 ^ n19936;
  assign n23571 = n21855 ^ n21689;
  assign n24522 = n24521 ^ n23571;
  assign n21755 = n21754 ^ n21751;
  assign n24523 = n24522 ^ n21755;
  assign n24525 = n24524 ^ n24523;
  assign n24491 = n21676 ^ n21668;
  assign n24490 = n21552 ^ n21428;
  assign n24492 = n24491 ^ n24490;
  assign n24489 = n21715 ^ n19868;
  assign n24493 = n24492 ^ n24489;
  assign n24554 = n24525 ^ n24493;
  assign n21868 = n21867 ^ n21821;
  assign n24506 = n24505 ^ n21868;
  assign n24504 = n21805 ^ n20014;
  assign n24507 = n24506 ^ n24504;
  assign n24546 = n24507 ^ n24493;
  assign n24534 = n21836 ^ n21645;
  assign n23583 = n21855 ^ n21715;
  assign n24533 = n24532 ^ n23583;
  assign n24535 = n24534 ^ n24533;
  assign n24530 = n21689 ^ n19777;
  assign n24502 = n21552 ^ n19753;
  assign n23577 = n21855 ^ n21794;
  assign n24500 = n24499 ^ n23577;
  assign n21744 = n21743 ^ n21310;
  assign n24501 = n24500 ^ n21744;
  assign n24503 = n24502 ^ n24501;
  assign n24531 = n24530 ^ n24503;
  assign n24536 = n24535 ^ n24531;
  assign n24495 = n21826 ^ n21805;
  assign n21790 = n21302 ^ n21157;
  assign n24496 = n24495 ^ n21790;
  assign n24494 = n21855 ^ n19964;
  assign n24497 = n24496 ^ n24494;
  assign n24527 = n24525 ^ n24497;
  assign n24543 = n24536 ^ n24527;
  assign n24575 = n24546 ^ n24543;
  assign n21818 = n21817 ^ n21760;
  assign n24510 = n24509 ^ n21818;
  assign n24508 = n21774 ^ n19909;
  assign n24511 = n24510 ^ n24508;
  assign n24529 = n24511 ^ n24493;
  assign n24555 = n24529 ^ n24527;
  assign n24556 = n24554 & n24555;
  assign n24547 = n24546 ^ n24536;
  assign n24548 = n24527 & n24547;
  assign n24557 = n24556 ^ n24548;
  assign n24576 = n24575 ^ n24557;
  assign n24514 = n21292 ^ n21167;
  assign n24516 = n24515 ^ n24514;
  assign n24513 = n21794 ^ n19989;
  assign n24517 = n24516 ^ n24513;
  assign n24512 = n24511 ^ n24507;
  assign n24518 = n24517 ^ n24512;
  assign n24519 = n24518 ^ n24503;
  assign n24498 = n24497 ^ n24493;
  assign n24520 = n24519 ^ n24498;
  assign n24572 = n24543 ^ n24517;
  assign n24573 = n24520 & n24572;
  assign n24540 = n24503 ^ n24497;
  assign n24563 = n24554 ^ n24540;
  assign n24564 = n24543 & n24563;
  assign n24574 = n24573 ^ n24564;
  assign n24577 = n24576 ^ n24574;
  assign n24544 = n24543 ^ n24512;
  assign n24566 = n24544 ^ n24498;
  assign n24526 = n24525 ^ n24518;
  assign n24562 = n24517 & n24526;
  assign n24565 = n24564 ^ n24562;
  assign n24567 = n24566 ^ n24565;
  assign n24545 = n24498 & n24544;
  assign n24549 = n24548 ^ n24545;
  assign n24568 = n24567 ^ n24549;
  assign n24584 = n24577 ^ n24568;
  assign n24559 = ~n24503 & n24518;
  assign n24537 = n24536 ^ n24529;
  assign n24541 = n24537 & n24540;
  assign n24560 = n24559 ^ n24541;
  assign n24553 = n24540 ^ n24537;
  assign n24558 = n24557 ^ n24553;
  assign n24561 = n24560 ^ n24558;
  assign n24578 = n24561 & n24577;
  assign n24585 = n24584 ^ n24578;
  assign n24538 = n24537 ^ n24518;
  assign n24528 = n24527 ^ n24526;
  assign n24551 = n24538 ^ n24528;
  assign n24539 = n24528 & n24538;
  assign n24542 = n24541 ^ n24539;
  assign n24550 = n24549 ^ n24542;
  assign n24552 = n24551 ^ n24550;
  assign n24582 = ~n24568 & n24577;
  assign n24583 = n24552 & n24582;
  assign n24586 = n24585 ^ n24583;
  assign n24571 = n24561 ^ n24552;
  assign n24579 = n24578 ^ n24571;
  assign n24569 = n24561 & n24568;
  assign n24570 = ~n24552 & n24569;
  assign n24580 = n24579 ^ n24570;
  assign n24606 = n24586 ^ n24580;
  assign n24599 = n24578 ^ n24552;
  assign n24600 = n24584 & n24599;
  assign n24601 = n24600 ^ n24568;
  assign n24589 = n24578 ^ n24568;
  assign n24590 = n24571 & n24589;
  assign n24591 = n24590 ^ n24552;
  assign n24604 = n24601 ^ n24591;
  assign n24607 = n24606 ^ n24604;
  assign n24608 = n24554 & n24607;
  assign n24605 = n24527 & n24604;
  assign n24609 = n24608 ^ n24605;
  assign n24581 = n24520 & n24580;
  assign n24972 = n24609 ^ n24581;
  assign n24923 = n24547 & n24604;
  assign n24880 = n24555 & n24607;
  assign n24924 = n24923 ^ n24880;
  assign n24595 = n24572 & n24580;
  assign n24592 = n24591 ^ n24580;
  assign n24594 = n24563 & n24592;
  assign n24596 = n24595 ^ n24594;
  assign n24593 = n24543 & n24592;
  assign n24597 = n24596 ^ n24593;
  assign n24971 = n24924 ^ n24597;
  assign n24973 = n24972 ^ n24971;
  assign n24969 = n24726 ^ n24709;
  assign n24707 = ~n24633 & ~n24704;
  assign n24700 = n24637 & ~n24699;
  assign n24706 = n24705 ^ n24700;
  assign n24708 = n24707 ^ n24706;
  assign n24968 = n24918 ^ n24708;
  assign n24970 = n24969 ^ n24968;
  assign n24974 = n24973 ^ n24970;
  assign n23426 = n22787 ^ n22670;
  assign n24399 = n23426 ^ n22663;
  assign n24400 = n24399 ^ n22706;
  assign n24401 = n24400 ^ n22885;
  assign n24368 = n22591 ^ n22324;
  assign n24369 = n24368 ^ n22622;
  assign n24370 = n24369 ^ n22573;
  assign n24371 = n24370 ^ n22882;
  assign n24432 = n24401 ^ n24371;
  assign n24409 = n22902 ^ n22441;
  assign n24407 = n22777 ^ n22729;
  assign n24406 = n22780 ^ n22090;
  assign n24408 = n24407 ^ n24406;
  assign n24410 = n24409 ^ n24408;
  assign n23460 = n22729 ^ n22553;
  assign n23432 = n22702 ^ n22683;
  assign n24394 = n23460 ^ n23432;
  assign n24396 = n24395 ^ n24394;
  assign n24397 = n24396 ^ n22658;
  assign n24398 = n24397 ^ n22880;
  assign n24411 = n24410 ^ n24398;
  assign n24433 = n24432 ^ n24411;
  assign n23473 = n22729 ^ n22622;
  assign n24386 = n23473 ^ n22553;
  assign n24385 = n24384 ^ n22580;
  assign n24387 = n24386 ^ n24385;
  assign n24381 = n22890 ^ n22638;
  assign n23419 = n22757 ^ n22729;
  assign n24379 = n23419 ^ n22207;
  assign n24378 = n24377 ^ n22073;
  assign n24380 = n24379 ^ n24378;
  assign n24382 = n24381 ^ n24380;
  assign n24376 = n22888 ^ n22711;
  assign n24383 = n24382 ^ n24376;
  assign n24388 = n24387 ^ n24383;
  assign n24439 = n24432 ^ n24388;
  assign n23446 = n22777 ^ n22738;
  assign n24372 = n23446 ^ n22677;
  assign n24373 = n24372 ^ n22724;
  assign n24374 = n24373 ^ n22894;
  assign n24402 = n24401 ^ n24374;
  assign n24392 = n22897 ^ n22451;
  assign n24390 = n22733 ^ n22082;
  assign n24391 = n24390 ^ n23419;
  assign n24393 = n24392 ^ n24391;
  assign n24403 = n24402 ^ n24393;
  assign n24448 = n24439 ^ n24403;
  assign n24404 = n24403 ^ n24398;
  assign n24447 = n24411 ^ n24404;
  assign n24452 = n24448 ^ n24447;
  assign n24449 = ~n24447 & ~n24448;
  assign n24414 = n24410 ^ n24382;
  assign n24442 = ~n24414 & n24439;
  assign n24450 = n24449 ^ n24442;
  assign n24375 = n24374 ^ n24371;
  assign n24389 = n24388 ^ n24375;
  assign n24423 = n24389 & n24411;
  assign n24412 = n24411 ^ n24388;
  assign n24418 = n24412 ^ n24402;
  assign n24419 = n24410 ^ n24371;
  assign n24422 = ~n24418 & n24419;
  assign n24424 = n24423 ^ n24422;
  assign n24451 = n24450 ^ n24424;
  assign n24453 = n24452 ^ n24451;
  assign n24420 = n24419 ^ n24418;
  assign n24413 = n24398 ^ n24371;
  assign n24415 = n24414 ^ n24413;
  assign n24416 = ~n24412 & ~n24415;
  assign n24405 = ~n24393 & ~n24404;
  assign n24417 = n24416 ^ n24405;
  assign n24421 = n24420 ^ n24417;
  assign n24425 = n24424 ^ n24421;
  assign n24434 = n24413 & ~n24433;
  assign n24435 = n24434 ^ n24423;
  assign n24431 = n24412 ^ n24375;
  assign n24436 = n24435 ^ n24431;
  assign n24426 = n24403 ^ n24382;
  assign n24427 = n24426 ^ n24419;
  assign n24428 = n24412 ^ n24393;
  assign n24429 = n24427 & n24428;
  assign n24430 = n24429 ^ n24416;
  assign n24437 = n24436 ^ n24430;
  assign n24477 = n24425 & n24437;
  assign n24478 = n24453 & n24477;
  assign n24443 = n24382 & ~n24403;
  assign n24444 = n24443 ^ n24442;
  assign n24440 = n24439 ^ n24414;
  assign n24441 = n24440 ^ n24435;
  assign n24445 = n24444 ^ n24441;
  assign n24446 = n24437 & ~n24445;
  assign n24438 = n24437 ^ n24425;
  assign n24476 = n24446 ^ n24438;
  assign n24479 = n24478 ^ n24476;
  assign n24457 = n24453 ^ n24445;
  assign n24467 = n24457 ^ n24446;
  assign n24465 = ~n24425 & ~n24445;
  assign n24466 = ~n24453 & n24465;
  assign n24468 = n24467 ^ n24466;
  assign n24480 = n24479 ^ n24468;
  assign n24458 = n24446 ^ n24425;
  assign n24459 = ~n24457 & ~n24458;
  assign n24460 = n24459 ^ n24453;
  assign n24454 = n24453 ^ n24446;
  assign n24455 = ~n24438 & n24454;
  assign n24456 = n24455 ^ n24425;
  assign n24461 = n24460 ^ n24456;
  assign n24850 = n24480 ^ n24461;
  assign n24855 = ~n24433 & ~n24850;
  assign n24462 = n24389 & ~n24461;
  assign n24964 = n24855 ^ n24462;
  assign n24859 = ~n24403 & ~n24479;
  assign n24858 = n24427 & ~n24468;
  assign n24860 = n24859 ^ n24858;
  assign n24965 = n24964 ^ n24860;
  assign n24469 = n24468 ^ n24460;
  assign n24941 = ~n24415 & ~n24469;
  assign n24483 = n24479 ^ n24456;
  assign n24853 = n24439 & n24483;
  assign n24851 = n24413 & ~n24850;
  assign n24463 = n24411 & ~n24461;
  assign n24852 = n24851 ^ n24463;
  assign n24854 = n24853 ^ n24852;
  assign n24963 = n24941 ^ n24854;
  assign n24966 = n24965 ^ n24963;
  assign n24280 = n24279 ^ n19900;
  assign n19929 = n19928 ^ n19925;
  assign n24278 = n23327 ^ n19929;
  assign n24281 = n24280 ^ n24278;
  assign n24245 = n24244 ^ n19799;
  assign n19643 = n19642 ^ n18741;
  assign n24243 = n24242 ^ n19643;
  assign n24246 = n24245 ^ n24243;
  assign n24307 = n24281 ^ n24246;
  assign n24289 = n24288 ^ n17804;
  assign n20007 = n20006 ^ n20003;
  assign n24287 = n24286 ^ n20007;
  assign n24290 = n24289 ^ n24287;
  assign n24276 = n24275 ^ n19880;
  assign n23316 = n19951 ^ n19812;
  assign n24273 = n24272 ^ n23316;
  assign n24274 = n24273 ^ n23305;
  assign n24277 = n24276 ^ n24274;
  assign n24291 = n24290 ^ n24277;
  assign n24308 = n24307 ^ n24291;
  assign n24249 = n24248 ^ n19943;
  assign n19894 = n19893 ^ n19887;
  assign n24247 = n23310 ^ n19894;
  assign n24250 = n24249 ^ n24247;
  assign n24282 = n24281 ^ n24250;
  assign n24270 = n24269 ^ n17794;
  assign n19956 = n19955 ^ n19951;
  assign n24268 = n24267 ^ n19956;
  assign n24271 = n24270 ^ n24268;
  assign n24283 = n24282 ^ n24271;
  assign n24256 = n24255 ^ n19650;
  assign n23288 = n19978 ^ n19951;
  assign n24253 = n24252 ^ n23288;
  assign n24254 = n24253 ^ n23299;
  assign n24257 = n24256 ^ n24254;
  assign n24312 = n24283 ^ n24257;
  assign n24299 = n24290 ^ n24246;
  assign n24313 = n24312 ^ n24299;
  assign n24263 = n24262 ^ n19763;
  assign n23295 = n19951 ^ n19837;
  assign n24261 = n24260 ^ n23295;
  assign n24264 = n24263 ^ n24261;
  assign n24259 = n24258 ^ n24257;
  assign n24265 = n24264 ^ n24259;
  assign n24292 = n24291 ^ n24265;
  assign n24314 = n24292 ^ n24271;
  assign n24315 = n24313 & ~n24314;
  assign n24294 = n24290 ^ n24257;
  assign n24293 = n24277 ^ n24246;
  assign n24295 = n24294 ^ n24293;
  assign n24296 = n24292 & ~n24295;
  assign n24316 = n24315 ^ n24296;
  assign n24309 = ~n24293 & ~n24308;
  assign n24251 = n24250 ^ n24246;
  assign n24266 = n24265 ^ n24251;
  assign n24303 = ~n24266 & n24291;
  assign n24310 = n24309 ^ n24303;
  assign n24306 = n24292 ^ n24251;
  assign n24311 = n24310 ^ n24306;
  assign n24317 = n24316 ^ n24311;
  assign n24323 = ~n24257 & ~n24283;
  assign n24319 = n24307 ^ n24265;
  assign n24322 = n24294 & ~n24319;
  assign n24324 = n24323 ^ n24322;
  assign n24320 = n24319 ^ n24294;
  assign n24321 = n24320 ^ n24310;
  assign n24325 = n24324 ^ n24321;
  assign n24326 = ~n24317 & ~n24325;
  assign n24298 = n24292 ^ n24282;
  assign n24302 = n24298 & ~n24299;
  assign n24304 = n24303 ^ n24302;
  assign n24300 = n24299 ^ n24298;
  assign n24284 = n24283 ^ n24277;
  assign n24285 = ~n24271 & ~n24284;
  assign n24297 = n24296 ^ n24285;
  assign n24301 = n24300 ^ n24297;
  assign n24305 = n24304 ^ n24301;
  assign n24318 = n24317 ^ n24305;
  assign n24358 = n24326 ^ n24318;
  assign n24328 = n24319 ^ n24283;
  assign n24327 = n24291 ^ n24284;
  assign n24332 = n24328 ^ n24327;
  assign n24329 = ~n24327 & n24328;
  assign n24330 = n24329 ^ n24322;
  assign n24331 = n24330 ^ n24304;
  assign n24333 = n24332 ^ n24331;
  assign n24356 = n24305 & ~n24317;
  assign n24357 = ~n24333 & n24356;
  assign n24359 = n24358 ^ n24357;
  assign n24337 = n24333 ^ n24325;
  assign n24347 = n24337 ^ n24326;
  assign n24345 = ~n24305 & ~n24325;
  assign n24346 = n24333 & n24345;
  assign n24348 = n24347 ^ n24346;
  assign n24360 = n24359 ^ n24348;
  assign n24338 = n24326 ^ n24305;
  assign n24339 = n24337 & ~n24338;
  assign n24340 = n24339 ^ n24333;
  assign n24334 = n24333 ^ n24326;
  assign n24335 = n24318 & ~n24334;
  assign n24336 = n24335 ^ n24305;
  assign n24341 = n24340 ^ n24336;
  assign n24835 = n24360 ^ n24341;
  assign n24840 = ~n24308 & n24835;
  assign n24342 = ~n24266 & n24341;
  assign n24960 = n24840 ^ n24342;
  assign n24844 = ~n24283 & n24359;
  assign n24843 = n24313 & n24348;
  assign n24845 = n24844 ^ n24843;
  assign n24961 = n24960 ^ n24845;
  assign n24349 = n24348 ^ n24340;
  assign n24935 = ~n24295 & ~n24349;
  assign n24362 = n24359 ^ n24336;
  assign n24838 = ~n24319 & ~n24362;
  assign n24836 = ~n24293 & n24835;
  assign n24343 = n24291 & n24341;
  assign n24837 = n24836 ^ n24343;
  assign n24839 = n24838 ^ n24837;
  assign n24959 = n24935 ^ n24839;
  assign n24962 = n24961 ^ n24959;
  assign n24967 = n24966 ^ n24962;
  assign n24975 = n24974 ^ n24967;
  assign n24984 = n24983 ^ n24975;
  assign n24888 = ~n24662 & n24703;
  assign n24889 = n24888 ^ n24716;
  assign n24737 = ~n24663 & ~n24720;
  assign n24735 = ~n24636 & n24703;
  assign n24736 = n24735 ^ n24707;
  assign n24738 = n24737 ^ n24736;
  assign n24890 = n24889 ^ n24738;
  assign n24742 = ~n24665 & n24727;
  assign n24741 = ~n24652 & n24723;
  assign n24743 = n24742 ^ n24741;
  assign n24871 = n24870 ^ n24743;
  assign n24887 = n24871 ^ n24729;
  assign n24891 = n24890 ^ n24887;
  assign n24910 = n24909 ^ n24891;
  assign n24587 = n24518 & n24586;
  assign n24883 = n24609 ^ n24587;
  assign n24878 = n24544 & n24606;
  assign n24602 = n24601 ^ n24586;
  assign n24877 = n24540 & n24602;
  assign n24879 = n24878 ^ n24877;
  assign n24881 = n24880 ^ n24879;
  assign n24875 = n24519 & n24586;
  assign n24874 = n24538 & n24601;
  assign n24876 = n24875 ^ n24874;
  assign n24882 = n24881 ^ n24876;
  assign n24884 = n24883 ^ n24882;
  assign n24868 = n24689 & ~n24714;
  assign n24867 = ~n24661 & ~n24720;
  assign n24869 = n24868 ^ n24867;
  assign n24872 = n24871 ^ n24869;
  assign n24866 = n24726 ^ n24715;
  assign n24873 = n24872 ^ n24866;
  assign n24885 = n24884 ^ n24873;
  assign n24861 = ~n24404 & n24460;
  assign n24862 = n24861 ^ n24860;
  assign n24473 = ~n24447 & ~n24456;
  assign n24471 = ~n24393 & n24460;
  assign n24470 = ~n24412 & ~n24469;
  assign n24472 = n24471 ^ n24470;
  assign n24474 = n24473 ^ n24472;
  assign n24863 = n24862 ^ n24474;
  assign n24484 = ~n24414 & n24483;
  assign n24482 = ~n24418 & n24480;
  assign n24485 = n24484 ^ n24482;
  assign n24856 = n24855 ^ n24485;
  assign n24857 = n24856 ^ n24854;
  assign n24864 = n24863 ^ n24857;
  assign n24846 = ~n24284 & ~n24340;
  assign n24847 = n24846 ^ n24845;
  assign n24353 = ~n24327 & ~n24336;
  assign n24351 = ~n24271 & ~n24340;
  assign n24350 = n24292 & ~n24349;
  assign n24352 = n24351 ^ n24350;
  assign n24354 = n24353 ^ n24352;
  assign n24848 = n24847 ^ n24354;
  assign n24364 = n24298 & n24360;
  assign n24363 = n24294 & ~n24362;
  assign n24365 = n24364 ^ n24363;
  assign n24841 = n24840 ^ n24365;
  assign n24842 = n24841 ^ n24839;
  assign n24849 = n24848 ^ n24842;
  assign n24865 = n24864 ^ n24849;
  assign n24886 = n24885 ^ n24865;
  assign n24911 = n24910 ^ n24886;
  assign n25106 = n24984 ^ n24911;
  assign n25047 = n25046 ^ n24873;
  assign n25032 = ~n24448 & ~n24456;
  assign n25031 = n24426 & ~n24479;
  assign n25033 = n25032 ^ n25031;
  assign n25034 = n25033 ^ n24856;
  assign n25030 = n24859 ^ n24852;
  assign n25035 = n25034 ^ n25030;
  assign n25028 = n24844 ^ n24837;
  assign n25025 = n24328 & ~n24336;
  assign n25024 = ~n24312 & n24359;
  assign n25026 = n25025 ^ n25024;
  assign n25027 = n25026 ^ n24841;
  assign n25029 = n25028 ^ n25027;
  assign n25036 = n25035 ^ n25029;
  assign n25020 = n24869 ^ n24736;
  assign n25019 = n24742 ^ n24729;
  assign n25021 = n25020 ^ n25019;
  assign n25022 = n25021 ^ n24920;
  assign n24928 = n24517 & n24591;
  assign n24997 = n24928 ^ n24593;
  assign n25016 = n24997 ^ n24876;
  assign n24603 = n24537 & n24602;
  assign n24610 = n24609 ^ n24603;
  assign n25015 = n24877 ^ n24610;
  assign n25017 = n25016 ^ n25015;
  assign n24588 = n24587 ^ n24581;
  assign n24925 = n24924 ^ n24588;
  assign n24922 = n24610 ^ n24594;
  assign n24926 = n24925 ^ n24922;
  assign n25018 = n25017 ^ n24926;
  assign n25023 = n25022 ^ n25018;
  assign n25037 = n25036 ^ n25023;
  assign n25048 = n25047 ^ n25037;
  assign n25080 = n25048 ^ n24984;
  assign n25071 = n25032 ^ n24471;
  assign n24940 = n24428 & ~n24468;
  assign n24942 = n24941 ^ n24940;
  assign n25072 = n25071 ^ n24942;
  assign n25070 = n24860 ^ n24852;
  assign n25073 = n25072 ^ n25070;
  assign n25067 = n25025 ^ n24351;
  assign n24934 = ~n24314 & n24348;
  assign n24936 = n24935 ^ n24934;
  assign n25068 = n25067 ^ n24936;
  assign n25066 = n24845 ^ n24837;
  assign n25069 = n25068 ^ n25066;
  assign n25074 = n25073 ^ n25069;
  assign n25060 = n24526 & n24591;
  assign n25061 = n25060 ^ n24588;
  assign n24998 = n24528 & n24601;
  assign n24999 = n24998 ^ n24997;
  assign n25062 = n25061 ^ n24999;
  assign n25059 = n24881 ^ n24610;
  assign n25063 = n25062 ^ n25059;
  assign n25064 = n25063 ^ n24926;
  assign n25058 = n24920 ^ n24891;
  assign n25065 = n25064 ^ n25058;
  assign n25075 = n25074 ^ n25065;
  assign n24914 = n24867 ^ n24735;
  assign n24915 = n24914 ^ n24706;
  assign n24913 = n24726 ^ n24716;
  assign n24916 = n24915 ^ n24913;
  assign n25056 = n25055 ^ n24916;
  assign n25057 = n25056 ^ n25048;
  assign n25076 = n25075 ^ n25057;
  assign n24740 = n24642 & n24723;
  assign n24744 = n24743 ^ n24740;
  assign n24734 = n24733 ^ n24722;
  assign n24739 = n24738 ^ n24734;
  assign n24745 = n24744 ^ n24739;
  assign n24833 = n24832 ^ n24745;
  assign n24717 = n24716 ^ n24708;
  assign n24730 = n24729 ^ n24717;
  assign n24598 = n24597 ^ n24588;
  assign n24611 = n24610 ^ n24598;
  assign n24731 = n24730 ^ n24611;
  assign n24481 = n24419 & n24480;
  assign n24486 = n24485 ^ n24481;
  assign n24464 = n24463 ^ n24462;
  assign n24475 = n24474 ^ n24464;
  assign n24487 = n24486 ^ n24475;
  assign n24361 = ~n24299 & n24360;
  assign n24366 = n24365 ^ n24361;
  assign n24344 = n24343 ^ n24342;
  assign n24355 = n24354 ^ n24344;
  assign n24367 = n24366 ^ n24355;
  assign n24488 = n24487 ^ n24367;
  assign n24732 = n24731 ^ n24488;
  assign n24834 = n24833 ^ n24732;
  assign n24912 = n24911 ^ n24834;
  assign n25081 = n25076 ^ n24912;
  assign n25103 = ~n25080 & n25081;
  assign n25091 = n25026 ^ n24352;
  assign n25090 = n24839 ^ n24363;
  assign n25092 = n25091 ^ n25090;
  assign n25087 = n25033 ^ n24472;
  assign n25086 = n24854 ^ n24484;
  assign n25088 = n25087 ^ n25086;
  assign n25085 = n25022 ^ n24926;
  assign n25089 = n25088 ^ n25085;
  assign n25093 = n25092 ^ n25089;
  assign n25100 = n25099 ^ n25093;
  assign n25012 = n25011 ^ n24970;
  assign n25001 = n24498 & n24606;
  assign n25002 = n25001 ^ n24879;
  assign n24996 = n24923 ^ n24605;
  assign n25000 = n24999 ^ n24996;
  assign n25003 = n25002 ^ n25000;
  assign n25004 = n25003 ^ n24745;
  assign n24993 = n24858 ^ n24852;
  assign n24943 = n24942 ^ n24470;
  assign n24992 = n24964 ^ n24943;
  assign n24994 = n24993 ^ n24992;
  assign n24990 = n24843 ^ n24837;
  assign n24937 = n24936 ^ n24350;
  assign n24989 = n24960 ^ n24937;
  assign n24991 = n24990 ^ n24989;
  assign n24995 = n24994 ^ n24991;
  assign n25005 = n25004 ^ n24995;
  assign n25013 = n25012 ^ n25005;
  assign n25084 = n25013 ^ n24834;
  assign n25101 = n25100 ^ n25084;
  assign n25102 = n25048 & ~n25101;
  assign n25104 = n25103 ^ n25102;
  assign n25082 = n25081 ^ n25080;
  assign n24957 = n24956 ^ n24730;
  assign n24944 = n24943 ^ n24860;
  assign n24945 = n24944 ^ n24854;
  assign n24938 = n24937 ^ n24845;
  assign n24939 = n24938 ^ n24839;
  assign n24946 = n24945 ^ n24939;
  assign n24929 = n24928 ^ n24874;
  assign n24930 = n24929 ^ n24596;
  assign n24927 = n24609 ^ n24588;
  assign n24931 = n24930 ^ n24927;
  assign n24932 = n24931 ^ n24926;
  assign n24921 = n24920 ^ n24916;
  assign n24933 = n24932 ^ n24921;
  assign n24947 = n24946 ^ n24933;
  assign n24958 = n24957 ^ n24947;
  assign n24985 = n24984 ^ n24958;
  assign n25014 = n25013 ^ n24911;
  assign n25077 = n25076 ^ n25014;
  assign n25078 = n24985 & n25077;
  assign n24986 = n24985 ^ n24912;
  assign n24987 = n24958 ^ n24911;
  assign n24988 = ~n24986 & n24987;
  assign n25079 = n25078 ^ n24988;
  assign n25083 = n25082 ^ n25079;
  assign n25105 = n25104 ^ n25083;
  assign n25107 = n25076 ^ n24985;
  assign n25132 = n25107 ^ n25014;
  assign n25133 = n25132 ^ n25079;
  assign n25127 = n25101 ^ n25048;
  assign n25128 = n25127 ^ n25106;
  assign n25129 = n25107 ^ n25100;
  assign n25130 = n25128 & n25129;
  assign n25121 = n25080 ^ n24987;
  assign n25122 = ~n25107 & ~n25121;
  assign n25131 = n25130 ^ n25122;
  assign n25134 = n25133 ^ n25131;
  assign n25135 = ~n25105 & n25134;
  assign n25113 = n25101 ^ n25081;
  assign n25111 = n25101 ^ n24958;
  assign n25112 = n25111 ^ n24985;
  assign n25117 = n25113 ^ n25112;
  assign n25114 = ~n25112 & ~n25113;
  assign n25115 = n25114 ^ n25103;
  assign n25108 = n25107 ^ n25084;
  assign n25109 = n25106 & ~n25108;
  assign n25110 = n25109 ^ n25078;
  assign n25116 = n25115 ^ n25110;
  assign n25118 = n25117 ^ n25116;
  assign n25119 = n25118 ^ n25105;
  assign n25150 = n25135 ^ n25119;
  assign n25124 = n25108 ^ n25106;
  assign n25120 = ~n25100 & ~n25111;
  assign n25123 = n25122 ^ n25120;
  assign n25125 = n25124 ^ n25123;
  assign n25126 = n25125 ^ n25110;
  assign n25148 = ~n25105 & ~n25126;
  assign n25149 = ~n25118 & n25148;
  assign n25151 = n25150 ^ n25149;
  assign n25145 = n25126 & n25134;
  assign n25146 = n25118 & n25145;
  assign n25139 = n25134 ^ n25126;
  assign n25144 = n25139 ^ n25135;
  assign n25147 = n25146 ^ n25144;
  assign n25152 = n25151 ^ n25147;
  assign n26417 = n25106 & n25152;
  assign n25140 = n25135 ^ n25118;
  assign n25141 = ~n25139 & n25140;
  assign n25142 = n25141 ^ n25126;
  assign n25156 = n25147 ^ n25142;
  assign n25157 = ~n25080 & n25156;
  assign n25155 = ~n25108 & n25152;
  assign n25158 = n25157 ^ n25155;
  assign n26418 = n26417 ^ n25158;
  assign n25136 = n25135 ^ n25126;
  assign n25137 = ~n25119 & ~n25136;
  assign n25138 = n25137 ^ n25118;
  assign n25143 = n25142 ^ n25138;
  assign n26348 = n25077 & ~n25143;
  assign n25162 = n24985 & ~n25143;
  assign n26415 = n26348 ^ n25162;
  assign n25174 = ~n25100 & n25138;
  assign n25172 = n25151 ^ n25138;
  assign n25173 = ~n25107 & ~n25172;
  assign n25175 = n25174 ^ n25173;
  assign n25171 = ~n25112 & ~n25142;
  assign n25176 = n25175 ^ n25171;
  assign n26416 = n26415 ^ n25176;
  assign n26419 = n26418 ^ n26416;
  assign n23598 = n21867 ^ n21817;
  assign n23599 = n23598 ^ n21827;
  assign n23597 = n22791 ^ n21774;
  assign n23600 = n23599 ^ n23597;
  assign n23595 = n22650 ^ n21552;
  assign n23593 = n21743 ^ n21668;
  assign n21740 = n21739 ^ n21676;
  assign n23594 = n23593 ^ n21740;
  assign n23596 = n23595 ^ n23594;
  assign n23601 = n23600 ^ n23596;
  assign n21669 = n21668 ^ n21157;
  assign n23585 = n21836 ^ n21669;
  assign n23584 = n23583 ^ n22604;
  assign n23586 = n23585 ^ n23584;
  assign n21168 = n21167 ^ n21157;
  assign n23579 = n21743 ^ n21168;
  assign n23580 = n23579 ^ n21429;
  assign n23578 = n23577 ^ n22537;
  assign n23581 = n23580 ^ n23578;
  assign n21657 = n21656 ^ n21645;
  assign n23582 = n23581 ^ n21657;
  assign n23587 = n23586 ^ n23582;
  assign n23602 = n23601 ^ n23587;
  assign n21837 = n21836 ^ n21157;
  assign n23573 = n21837 ^ n21751;
  assign n23574 = n23573 ^ n21842;
  assign n23572 = n23571 ^ n22716;
  assign n23575 = n23574 ^ n23572;
  assign n23569 = n22743 ^ n21805;
  assign n23567 = n21867 ^ n21157;
  assign n21864 = n21863 ^ n21302;
  assign n23568 = n23567 ^ n21864;
  assign n23570 = n23569 ^ n23568;
  assign n23576 = n23575 ^ n23570;
  assign n23588 = n23587 ^ n23576;
  assign n23648 = n23601 ^ n23588;
  assign n23626 = n23596 ^ n23575;
  assign n23606 = n21817 ^ n21751;
  assign n23607 = n23606 ^ n21767;
  assign n23605 = n22690 ^ n21845;
  assign n23608 = n23607 ^ n23605;
  assign n23613 = n23608 ^ n23596;
  assign n23627 = n23613 ^ n23576;
  assign n23628 = n23626 & n23627;
  assign n23603 = n23576 & n23602;
  assign n23629 = n23628 ^ n23603;
  assign n23649 = n23648 ^ n23629;
  assign n21789 = n21788 ^ n21292;
  assign n23590 = n21789 ^ n21168;
  assign n23589 = n22766 ^ n21855;
  assign n23591 = n23590 ^ n23589;
  assign n23592 = n23591 ^ n23588;
  assign n23609 = n23608 ^ n23600;
  assign n23617 = n23609 ^ n23591;
  assign n23644 = n23617 ^ n23581;
  assign n23604 = n23596 ^ n23570;
  assign n23645 = n23644 ^ n23604;
  assign n23646 = n23592 & n23645;
  assign n23615 = n23581 ^ n23570;
  assign n23636 = n23626 ^ n23615;
  assign n23637 = n23588 & n23636;
  assign n23647 = n23646 ^ n23637;
  assign n23650 = n23649 ^ n23647;
  assign n23610 = n23609 ^ n23588;
  assign n23639 = n23610 ^ n23604;
  assign n23619 = n23617 ^ n23575;
  assign n23635 = n23591 & n23619;
  assign n23638 = n23637 ^ n23635;
  assign n23640 = n23639 ^ n23638;
  assign n23611 = n23604 & n23610;
  assign n23612 = n23611 ^ n23603;
  assign n23641 = n23640 ^ n23612;
  assign n23667 = n23650 ^ n23641;
  assign n23632 = ~n23581 & n23617;
  assign n23614 = n23613 ^ n23587;
  assign n23616 = n23614 & n23615;
  assign n23633 = n23632 ^ n23616;
  assign n23630 = n23615 ^ n23614;
  assign n23631 = n23630 ^ n23629;
  assign n23634 = n23633 ^ n23631;
  assign n23651 = n23634 & n23650;
  assign n23620 = n23619 ^ n23576;
  assign n23618 = n23617 ^ n23614;
  assign n23624 = n23620 ^ n23618;
  assign n23621 = n23618 & n23620;
  assign n23622 = n23621 ^ n23616;
  assign n23623 = n23622 ^ n23612;
  assign n23625 = n23624 ^ n23623;
  assign n23673 = n23651 ^ n23625;
  assign n23674 = n23667 & n23673;
  assign n23675 = n23674 ^ n23641;
  assign n23652 = n23634 ^ n23625;
  assign n23656 = n23651 ^ n23641;
  assign n23657 = n23652 & n23656;
  assign n23658 = n23657 ^ n23625;
  assign n23676 = n23675 ^ n23658;
  assign n23992 = n23602 & n23676;
  assign n23668 = n23667 ^ n23651;
  assign n23665 = ~n23641 & n23650;
  assign n23666 = n23625 & n23665;
  assign n23669 = n23668 ^ n23666;
  assign n23653 = n23652 ^ n23651;
  assign n23642 = n23634 & n23641;
  assign n23643 = ~n23625 & n23642;
  assign n23654 = n23653 ^ n23643;
  assign n23678 = n23669 ^ n23654;
  assign n23679 = n23678 ^ n23676;
  assign n23954 = n23627 & n23679;
  assign n24035 = n23992 ^ n23954;
  assign n23670 = n23617 & n23669;
  assign n23664 = n23645 & n23654;
  assign n23671 = n23670 ^ n23664;
  assign n24036 = n24035 ^ n23671;
  assign n23682 = n23675 ^ n23669;
  assign n23683 = n23614 & n23682;
  assign n23680 = n23626 & n23679;
  assign n23677 = n23576 & n23676;
  assign n23681 = n23680 ^ n23677;
  assign n23684 = n23683 ^ n23681;
  assign n23659 = n23658 ^ n23654;
  assign n23660 = n23636 & n23659;
  assign n24034 = n23684 ^ n23660;
  assign n24037 = n24036 ^ n24034;
  assign n24044 = n24043 ^ n24037;
  assign n23465 = n23464 ^ n22683;
  assign n22712 = n22711 ^ n22441;
  assign n23461 = n23460 ^ n22712;
  assign n23463 = n23462 ^ n23461;
  assign n23466 = n23465 ^ n23463;
  assign n23456 = n23455 ^ n22591;
  assign n23453 = n22638 ^ n22207;
  assign n23452 = n22633 ^ n22573;
  assign n23454 = n23453 ^ n23452;
  assign n23457 = n23456 ^ n23454;
  assign n23496 = n23466 ^ n23457;
  assign n23436 = n23435 ^ n22787;
  assign n23434 = n23433 ^ n23432;
  assign n23437 = n23436 ^ n23434;
  assign n23483 = n23457 ^ n23437;
  assign n22592 = n22591 ^ n22441;
  assign n23474 = n23473 ^ n22592;
  assign n23472 = n22580 ^ n22564;
  assign n23475 = n23474 ^ n23472;
  assign n23470 = n23469 ^ n22711;
  assign n23424 = n23423 ^ n22638;
  assign n22452 = n22451 ^ n22441;
  assign n23420 = n23419 ^ n22452;
  assign n23422 = n23421 ^ n23420;
  assign n23425 = n23424 ^ n23422;
  assign n23471 = n23470 ^ n23425;
  assign n23476 = n23475 ^ n23471;
  assign n23484 = n23483 ^ n23476;
  assign n23439 = n22729 ^ n22452;
  assign n23440 = n23439 ^ n22760;
  assign n23441 = n23440 ^ n22082;
  assign n23443 = n23442 ^ n23441;
  assign n23430 = n23429 ^ n22738;
  assign n23428 = n23427 ^ n23426;
  assign n23431 = n23430 ^ n23428;
  assign n23438 = n23437 ^ n23431;
  assign n23444 = n23443 ^ n23438;
  assign n23489 = n23484 ^ n23444;
  assign n23487 = n23466 ^ n23444;
  assign n23450 = n23449 ^ n22441;
  assign n23448 = n23447 ^ n23446;
  assign n23451 = n23450 ^ n23448;
  assign n23467 = n23466 ^ n23451;
  assign n23488 = n23487 ^ n23467;
  assign n23493 = n23489 ^ n23488;
  assign n23490 = ~n23488 & ~n23489;
  assign n23485 = n23451 ^ n23425;
  assign n23486 = n23484 & ~n23485;
  assign n23491 = n23490 ^ n23486;
  assign n23458 = n23457 ^ n23451;
  assign n23479 = n23476 ^ n23467;
  assign n23480 = n23479 ^ n23438;
  assign n23481 = n23458 & ~n23480;
  assign n23468 = n23457 ^ n23431;
  assign n23477 = n23476 ^ n23468;
  assign n23478 = n23467 & n23477;
  assign n23482 = n23481 ^ n23478;
  assign n23492 = n23491 ^ n23482;
  assign n23494 = n23493 ^ n23492;
  assign n23500 = n23480 ^ n23458;
  assign n23497 = n23496 ^ n23485;
  assign n23498 = ~n23479 & ~n23497;
  assign n23495 = ~n23443 & ~n23487;
  assign n23499 = n23498 ^ n23495;
  assign n23501 = n23500 ^ n23499;
  assign n23502 = n23501 ^ n23482;
  assign n23517 = n23479 ^ n23468;
  assign n23504 = n23483 ^ n23467;
  assign n23505 = n23496 & ~n23504;
  assign n23506 = n23505 ^ n23478;
  assign n23518 = n23517 ^ n23506;
  assign n23445 = n23444 ^ n23425;
  assign n23459 = n23458 ^ n23445;
  assign n23514 = n23479 ^ n23443;
  assign n23515 = n23459 & n23514;
  assign n23516 = n23515 ^ n23498;
  assign n23519 = n23518 ^ n23516;
  assign n23526 = n23502 & n23519;
  assign n23527 = n23494 & n23526;
  assign n23524 = n23519 ^ n23502;
  assign n23508 = n23425 & ~n23444;
  assign n23509 = n23508 ^ n23486;
  assign n23503 = n23485 ^ n23484;
  assign n23507 = n23506 ^ n23503;
  assign n23510 = n23509 ^ n23507;
  assign n23520 = ~n23510 & n23519;
  assign n23525 = n23524 ^ n23520;
  assign n23528 = n23527 ^ n23525;
  assign n23513 = n23510 ^ n23494;
  assign n23521 = n23520 ^ n23513;
  assign n23511 = ~n23502 & ~n23510;
  assign n23512 = ~n23494 & n23511;
  assign n23522 = n23521 ^ n23512;
  assign n23539 = n23528 ^ n23522;
  assign n23534 = n23520 ^ n23502;
  assign n23535 = ~n23513 & ~n23534;
  assign n23536 = n23535 ^ n23494;
  assign n23531 = n23520 ^ n23494;
  assign n23532 = ~n23524 & n23531;
  assign n23533 = n23532 ^ n23502;
  assign n23537 = n23536 ^ n23533;
  assign n23540 = n23539 ^ n23537;
  assign n23541 = n23496 & ~n23540;
  assign n23538 = n23467 & ~n23537;
  assign n23542 = n23541 ^ n23538;
  assign n23523 = n23459 & ~n23522;
  assign n24030 = n23542 ^ n23523;
  assign n23548 = n23536 ^ n23522;
  assign n23563 = ~n23479 & ~n23548;
  assign n23549 = ~n23497 & ~n23548;
  assign n23547 = n23514 & ~n23522;
  assign n23550 = n23549 ^ n23547;
  assign n23564 = n23563 ^ n23550;
  assign n23558 = ~n23504 & ~n23540;
  assign n23557 = n23477 & ~n23537;
  assign n23559 = n23558 ^ n23557;
  assign n24029 = n23564 ^ n23559;
  assign n24031 = n24030 ^ n24029;
  assign n23529 = ~n23444 & ~n23528;
  assign n23530 = n23529 ^ n23523;
  assign n23560 = n23559 ^ n23530;
  assign n23553 = n23533 ^ n23528;
  assign n23554 = n23484 & n23553;
  assign n23555 = n23554 ^ n23542;
  assign n23556 = n23555 ^ n23549;
  assign n23561 = n23560 ^ n23556;
  assign n24032 = n24031 ^ n23561;
  assign n23313 = n22901 ^ n17804;
  assign n23311 = n23310 ^ n19955;
  assign n23312 = n23311 ^ n16817;
  assign n23314 = n23313 ^ n23312;
  assign n23300 = n23299 ^ n19799;
  assign n23301 = n23300 ^ n19791;
  assign n23302 = n23301 ^ n19848;
  assign n23303 = n23302 ^ n22881;
  assign n23334 = n23314 ^ n23303;
  assign n19947 = n19946 ^ n19943;
  assign n23328 = n23327 ^ n19947;
  assign n23329 = n23328 ^ n20006;
  assign n23330 = n23329 ^ n22893;
  assign n20000 = n19999 ^ n19900;
  assign n23304 = n20000 ^ n19893;
  assign n23306 = n23305 ^ n23304;
  assign n23307 = n23306 ^ n22884;
  assign n23331 = n23330 ^ n23307;
  assign n23324 = n22896 ^ n17794;
  assign n23322 = n19982 ^ n19951;
  assign n16828 = n16827 ^ n16817;
  assign n23323 = n23322 ^ n16828;
  assign n23325 = n23324 ^ n23323;
  assign n23332 = n23331 ^ n23325;
  assign n23291 = n22889 ^ n19650;
  assign n23289 = n23288 ^ n19642;
  assign n23287 = n19852 ^ n16828;
  assign n23290 = n23289 ^ n23287;
  assign n23292 = n23291 ^ n23290;
  assign n23333 = n23332 ^ n23292;
  assign n23335 = n23334 ^ n23333;
  assign n23308 = n23307 ^ n23303;
  assign n23296 = n23295 ^ n19823;
  assign n19792 = n19791 ^ n16817;
  assign n23294 = n19919 ^ n19792;
  assign n23297 = n23296 ^ n23294;
  assign n23286 = n22887 ^ n19763;
  assign n23293 = n23292 ^ n23286;
  assign n23298 = n23297 ^ n23293;
  assign n23309 = n23308 ^ n23298;
  assign n23369 = n23332 ^ n23309;
  assign n19920 = n19919 ^ n16817;
  assign n19881 = n19880 ^ n19877;
  assign n23315 = n19920 ^ n19881;
  assign n23317 = n23316 ^ n23315;
  assign n23318 = n23317 ^ n19928;
  assign n23319 = n23318 ^ n22879;
  assign n23351 = n23332 ^ n23319;
  assign n23320 = n23319 ^ n23314;
  assign n23368 = n23351 ^ n23320;
  assign n23373 = n23369 ^ n23368;
  assign n23370 = ~n23368 & ~n23369;
  assign n23338 = n23314 ^ n23292;
  assign n23364 = n23309 & ~n23338;
  assign n23371 = n23370 ^ n23364;
  assign n23321 = n23320 ^ n23298;
  assign n23354 = n23331 ^ n23321;
  assign n23357 = n23334 & ~n23354;
  assign n23344 = n23330 ^ n23303;
  assign n23345 = n23344 ^ n23298;
  assign n23346 = n23320 & n23345;
  assign n23358 = n23357 ^ n23346;
  assign n23372 = n23371 ^ n23358;
  assign n23374 = n23373 ^ n23372;
  assign n23363 = n23292 & ~n23332;
  assign n23365 = n23364 ^ n23363;
  assign n23361 = n23338 ^ n23309;
  assign n23337 = n23319 ^ n23303;
  assign n23342 = n23320 ^ n23308;
  assign n23343 = n23337 & ~n23342;
  assign n23347 = n23346 ^ n23343;
  assign n23362 = n23361 ^ n23347;
  assign n23366 = n23365 ^ n23362;
  assign n23384 = n23374 ^ n23366;
  assign n23348 = n23344 ^ n23321;
  assign n23349 = n23348 ^ n23347;
  assign n23339 = n23338 ^ n23337;
  assign n23340 = ~n23321 & ~n23339;
  assign n23326 = n23325 ^ n23321;
  assign n23336 = n23326 & n23335;
  assign n23341 = n23340 ^ n23336;
  assign n23350 = n23349 ^ n23341;
  assign n23367 = n23350 & ~n23366;
  assign n23392 = n23384 ^ n23367;
  assign n23355 = n23354 ^ n23334;
  assign n23352 = ~n23325 & ~n23351;
  assign n23353 = n23352 ^ n23340;
  assign n23356 = n23355 ^ n23353;
  assign n23359 = n23358 ^ n23356;
  assign n23390 = ~n23359 & ~n23366;
  assign n23391 = ~n23374 & n23390;
  assign n23393 = n23392 ^ n23391;
  assign n23402 = n23335 & ~n23393;
  assign n23379 = n23350 & n23359;
  assign n23380 = n23374 & n23379;
  assign n23360 = n23359 ^ n23350;
  assign n23378 = n23367 ^ n23360;
  assign n23381 = n23380 ^ n23378;
  assign n23394 = n23393 ^ n23381;
  assign n23385 = n23367 ^ n23359;
  assign n23386 = ~n23384 & ~n23385;
  assign n23387 = n23386 ^ n23374;
  assign n23375 = n23374 ^ n23367;
  assign n23376 = ~n23360 & n23375;
  assign n23377 = n23376 ^ n23359;
  assign n23388 = n23387 ^ n23377;
  assign n23395 = n23394 ^ n23388;
  assign n23396 = n23337 & ~n23395;
  assign n23389 = n23320 & ~n23388;
  assign n23397 = n23396 ^ n23389;
  assign n24026 = n23402 ^ n23397;
  assign n23399 = n23393 ^ n23387;
  assign n24005 = ~n23321 & ~n23399;
  assign n23414 = n23326 & ~n23393;
  assign n23400 = ~n23339 & ~n23399;
  assign n23415 = n23414 ^ n23400;
  assign n24006 = n24005 ^ n23415;
  assign n23406 = ~n23342 & ~n23395;
  assign n23405 = n23345 & ~n23388;
  assign n23407 = n23406 ^ n23405;
  assign n24025 = n24006 ^ n23407;
  assign n24027 = n24026 ^ n24025;
  assign n23733 = n23732 ^ n20945;
  assign n23731 = n23730 ^ n20765;
  assign n23734 = n23733 ^ n23731;
  assign n23728 = n23727 ^ n20810;
  assign n23726 = n23725 ^ n23724;
  assign n23729 = n23728 ^ n23726;
  assign n23735 = n23734 ^ n23729;
  assign n23713 = n23712 ^ n20875;
  assign n20893 = n20892 ^ n20343;
  assign n23711 = n23710 ^ n20893;
  assign n23714 = n23713 ^ n23711;
  assign n23706 = n23705 ^ n20740;
  assign n20715 = n20714 ^ n20343;
  assign n23703 = n23702 ^ n20715;
  assign n23704 = n23703 ^ n20803;
  assign n23707 = n23706 ^ n23704;
  assign n23709 = n23708 ^ n23707;
  assign n23715 = n23714 ^ n23709;
  assign n23736 = n23735 ^ n23715;
  assign n23742 = n23741 ^ n20852;
  assign n23740 = n23739 ^ n20942;
  assign n23743 = n23742 ^ n23740;
  assign n23753 = n23743 ^ n23734;
  assign n23699 = n23698 ^ n20914;
  assign n20921 = n20920 ^ n20343;
  assign n23696 = n23695 ^ n20921;
  assign n23697 = n23696 ^ n20859;
  assign n23700 = n23699 ^ n23697;
  assign n23693 = n23692 ^ n20783;
  assign n23691 = n23690 ^ n23689;
  assign n23694 = n23693 ^ n23691;
  assign n23701 = n23700 ^ n23694;
  assign n23716 = n23715 ^ n23701;
  assign n23774 = n23753 ^ n23716;
  assign n23761 = n23729 ^ n23694;
  assign n23784 = n23774 ^ n23761;
  assign n23721 = n23720 ^ n20615;
  assign n23719 = n23718 ^ n23717;
  assign n23722 = n23721 ^ n23719;
  assign n23754 = n23753 ^ n23722;
  assign n23769 = n23754 ^ n23700;
  assign n23782 = n23722 & n23769;
  assign n23748 = n23707 ^ n23694;
  assign n23738 = n23729 ^ n23700;
  assign n23758 = n23748 ^ n23738;
  assign n23759 = n23716 & ~n23758;
  assign n23783 = n23782 ^ n23759;
  assign n23785 = n23784 ^ n23783;
  assign n23775 = ~n23761 & ~n23774;
  assign n23737 = ~n23701 & n23736;
  assign n23776 = n23775 ^ n23737;
  assign n23786 = n23785 ^ n23776;
  assign n23765 = n23735 ^ n23716;
  assign n23744 = n23743 ^ n23729;
  assign n23745 = n23744 ^ n23701;
  assign n23746 = n23738 & ~n23745;
  assign n23747 = n23746 ^ n23737;
  assign n23766 = n23765 ^ n23747;
  assign n23723 = n23722 ^ n23716;
  assign n23760 = n23754 ^ n23707;
  assign n23762 = n23761 ^ n23760;
  assign n23763 = n23723 & ~n23762;
  assign n23764 = n23763 ^ n23759;
  assign n23767 = n23766 ^ n23764;
  assign n23802 = n23786 ^ n23767;
  assign n23749 = n23744 ^ n23715;
  assign n23771 = n23754 ^ n23749;
  assign n23770 = n23769 ^ n23701;
  assign n23778 = n23771 ^ n23770;
  assign n23772 = ~n23770 & n23771;
  assign n23752 = ~n23748 & ~n23749;
  assign n23773 = n23772 ^ n23752;
  assign n23777 = n23776 ^ n23773;
  assign n23779 = n23778 ^ n23777;
  assign n23755 = n23707 & ~n23754;
  assign n23756 = n23755 ^ n23752;
  assign n23750 = n23749 ^ n23748;
  assign n23751 = n23750 ^ n23747;
  assign n23757 = n23756 ^ n23751;
  assign n23768 = n23757 & ~n23767;
  assign n23808 = n23779 ^ n23768;
  assign n23809 = ~n23802 & ~n23808;
  assign n23810 = n23809 ^ n23786;
  assign n23780 = n23779 ^ n23757;
  assign n23791 = n23786 ^ n23768;
  assign n23792 = ~n23780 & n23791;
  assign n23793 = n23792 ^ n23779;
  assign n23811 = n23810 ^ n23793;
  assign n23988 = n23736 & ~n23811;
  assign n23803 = n23802 ^ n23768;
  assign n23800 = ~n23767 & ~n23786;
  assign n23801 = ~n23779 & n23800;
  assign n23804 = n23803 ^ n23801;
  assign n23787 = n23757 & n23786;
  assign n23788 = n23779 & n23787;
  assign n23781 = n23780 ^ n23768;
  assign n23789 = n23788 ^ n23781;
  assign n23813 = n23804 ^ n23789;
  assign n23814 = n23813 ^ n23811;
  assign n23913 = ~n23745 & ~n23814;
  assign n24022 = n23988 ^ n23913;
  assign n23805 = ~n23754 & ~n23804;
  assign n23799 = ~n23762 & ~n23789;
  assign n23806 = n23805 ^ n23799;
  assign n24023 = n24022 ^ n23806;
  assign n23817 = n23810 ^ n23804;
  assign n23818 = ~n23749 & ~n23817;
  assign n23815 = n23738 & ~n23814;
  assign n23812 = ~n23701 & ~n23811;
  assign n23816 = n23815 ^ n23812;
  assign n23819 = n23818 ^ n23816;
  assign n23794 = n23793 ^ n23789;
  assign n23795 = ~n23758 & n23794;
  assign n24021 = n23819 ^ n23795;
  assign n24024 = n24023 ^ n24021;
  assign n24028 = n24027 ^ n24024;
  assign n24033 = n24032 ^ n24028;
  assign n24045 = n24044 ^ n24033;
  assign n23961 = n23619 & n23658;
  assign n23962 = n23961 ^ n23671;
  assign n23958 = n23591 & n23658;
  assign n23662 = n23588 & n23659;
  assign n23959 = n23958 ^ n23662;
  assign n23957 = n23620 & n23675;
  assign n23960 = n23959 ^ n23957;
  assign n23963 = n23962 ^ n23960;
  assign n23952 = n23610 & n23678;
  assign n23951 = n23615 & n23682;
  assign n23953 = n23952 ^ n23951;
  assign n23955 = n23954 ^ n23953;
  assign n23956 = n23955 ^ n23684;
  assign n23964 = n23963 ^ n23956;
  assign n23382 = n23381 ^ n23377;
  assign n23945 = ~n23338 & n23382;
  assign n23944 = ~n23354 & n23394;
  assign n23946 = n23945 ^ n23944;
  assign n23947 = n23946 ^ n23406;
  assign n23942 = n23333 & ~n23381;
  assign n23412 = ~n23369 & ~n23377;
  assign n23943 = n23942 ^ n23412;
  assign n23948 = n23947 ^ n23943;
  assign n23403 = ~n23332 & ~n23381;
  assign n23941 = n23403 ^ n23397;
  assign n23949 = n23948 ^ n23941;
  assign n23937 = n23445 & ~n23528;
  assign n23545 = ~n23489 & ~n23533;
  assign n23938 = n23937 ^ n23545;
  assign n23925 = ~n23485 & n23553;
  assign n23924 = ~n23480 & n23539;
  assign n23926 = n23925 ^ n23924;
  assign n23927 = n23926 ^ n23558;
  assign n23939 = n23938 ^ n23927;
  assign n23936 = n23542 ^ n23529;
  assign n23940 = n23939 ^ n23936;
  assign n23950 = n23949 ^ n23940;
  assign n23965 = n23964 ^ n23950;
  assign n23932 = ~n23487 & n23536;
  assign n23933 = n23932 ^ n23530;
  assign n23930 = ~n23488 & ~n23533;
  assign n23544 = ~n23443 & n23536;
  assign n23929 = n23563 ^ n23544;
  assign n23931 = n23930 ^ n23929;
  assign n23934 = n23933 ^ n23931;
  assign n23928 = n23927 ^ n23555;
  assign n23935 = n23934 ^ n23928;
  assign n23966 = n23965 ^ n23935;
  assign n23920 = n23769 & ~n23793;
  assign n23921 = n23920 ^ n23806;
  assign n23917 = n23722 & ~n23793;
  assign n23797 = n23716 & n23794;
  assign n23918 = n23917 ^ n23797;
  assign n23916 = ~n23770 & n23810;
  assign n23919 = n23918 ^ n23916;
  assign n23922 = n23921 ^ n23919;
  assign n23911 = ~n23774 & n23813;
  assign n23910 = ~n23748 & ~n23817;
  assign n23912 = n23911 ^ n23910;
  assign n23914 = n23913 ^ n23912;
  assign n23915 = n23914 ^ n23819;
  assign n23923 = n23922 ^ n23915;
  assign n23967 = n23966 ^ n23923;
  assign n23984 = n23983 ^ n23967;
  assign n24162 = n24045 ^ n23984;
  assign n24095 = n23681 ^ n23670;
  assign n24092 = n23618 & n23675;
  assign n24091 = n23644 & n23669;
  assign n24093 = n24092 ^ n24091;
  assign n24094 = n24093 ^ n23955;
  assign n24096 = n24095 ^ n24094;
  assign n24105 = n24104 ^ n24096;
  assign n24086 = n23938 ^ n23929;
  assign n24085 = n23925 ^ n23555;
  assign n24087 = n24086 ^ n24085;
  assign n24088 = n24087 ^ n23561;
  assign n24089 = n24088 ^ n23940;
  assign n23411 = ~n23325 & n23387;
  assign n24050 = n24005 ^ n23411;
  assign n24081 = n24050 ^ n23943;
  assign n23383 = n23309 & n23382;
  assign n23398 = n23397 ^ n23383;
  assign n24080 = n23945 ^ n23398;
  assign n24082 = n24081 ^ n24080;
  assign n23404 = n23403 ^ n23402;
  assign n23408 = n23407 ^ n23404;
  assign n23401 = n23400 ^ n23398;
  assign n23409 = n23408 ^ n23401;
  assign n24083 = n24082 ^ n23409;
  assign n24078 = n23816 ^ n23805;
  assign n24075 = n23771 & n23810;
  assign n24074 = n23760 & ~n23804;
  assign n24076 = n24075 ^ n24074;
  assign n24077 = n24076 ^ n23914;
  assign n24079 = n24078 ^ n24077;
  assign n24084 = n24083 ^ n24079;
  assign n24090 = n24089 ^ n24084;
  assign n24106 = n24105 ^ n24090;
  assign n24137 = n24106 ^ n24045;
  assign n24130 = n23935 ^ n23561;
  assign n23546 = n23545 ^ n23544;
  assign n23551 = n23550 ^ n23546;
  assign n23543 = n23542 ^ n23530;
  assign n23552 = n23551 ^ n23543;
  assign n24131 = n24130 ^ n23552;
  assign n24124 = ~n23351 & n23387;
  assign n24125 = n24124 ^ n23404;
  assign n24051 = ~n23368 & ~n23377;
  assign n24052 = n24051 ^ n24050;
  assign n24126 = n24125 ^ n24052;
  assign n24123 = n23947 ^ n23398;
  assign n24127 = n24126 ^ n24123;
  assign n24128 = n24127 ^ n23409;
  assign n24120 = n24075 ^ n23917;
  assign n23790 = n23723 & ~n23789;
  assign n23796 = n23795 ^ n23790;
  assign n24121 = n24120 ^ n23796;
  assign n24119 = n23816 ^ n23806;
  assign n24122 = n24121 ^ n24119;
  assign n24129 = n24128 ^ n24122;
  assign n24132 = n24131 ^ n24129;
  assign n24108 = n24092 ^ n23958;
  assign n23655 = n23592 & n23654;
  assign n23661 = n23660 ^ n23655;
  assign n24109 = n24108 ^ n23661;
  assign n24107 = n23681 ^ n23671;
  assign n24110 = n24109 ^ n24107;
  assign n24117 = n24116 ^ n24110;
  assign n24118 = n24117 ^ n24106;
  assign n24133 = n24132 ^ n24118;
  assign n24007 = n24006 ^ n23404;
  assign n24008 = n24007 ^ n23398;
  assign n23565 = n23564 ^ n23530;
  assign n23566 = n23565 ^ n23555;
  assign n24009 = n24008 ^ n23566;
  assign n24000 = n23458 & n23539;
  assign n24001 = n24000 ^ n23926;
  assign n23998 = n23557 ^ n23538;
  assign n23999 = n23998 ^ n23931;
  assign n24002 = n24001 ^ n23999;
  assign n23995 = n23604 & n23678;
  assign n23996 = n23995 ^ n23953;
  assign n23993 = n23992 ^ n23677;
  assign n23994 = n23993 ^ n23960;
  assign n23997 = n23996 ^ n23994;
  assign n24003 = n24002 ^ n23997;
  assign n23989 = n23988 ^ n23812;
  assign n23990 = n23989 ^ n23919;
  assign n23986 = ~n23761 & n23813;
  assign n23987 = n23986 ^ n23912;
  assign n23991 = n23990 ^ n23987;
  assign n24004 = n24003 ^ n23991;
  assign n24010 = n24009 ^ n24004;
  assign n24019 = n24018 ^ n24010;
  assign n24020 = n24019 ^ n23984;
  assign n24138 = n24133 ^ n24020;
  assign n24159 = ~n24137 & n24138;
  assign n24148 = n24093 ^ n23959;
  assign n24147 = n23951 ^ n23684;
  assign n24149 = n24148 ^ n24147;
  assign n24155 = n24154 ^ n24149;
  assign n24143 = n24076 ^ n23918;
  assign n24142 = n23910 ^ n23819;
  assign n24144 = n24143 ^ n24142;
  assign n24145 = n24144 ^ n23409;
  assign n24146 = n24145 ^ n24088;
  assign n24156 = n24155 ^ n24146;
  assign n24064 = n23816 ^ n23799;
  assign n23798 = n23797 ^ n23796;
  assign n24063 = n24022 ^ n23798;
  assign n24065 = n24064 ^ n24063;
  assign n24059 = n23681 ^ n23664;
  assign n23663 = n23662 ^ n23661;
  assign n24058 = n24035 ^ n23663;
  assign n24060 = n24059 ^ n24058;
  assign n24061 = n24060 ^ n24031;
  assign n24054 = n23334 & n23394;
  assign n24055 = n24054 ^ n23946;
  assign n24049 = n23405 ^ n23389;
  assign n24053 = n24052 ^ n24049;
  assign n24056 = n24055 ^ n24053;
  assign n24057 = n24056 ^ n24002;
  assign n24062 = n24061 ^ n24057;
  assign n24066 = n24065 ^ n24062;
  assign n24072 = n24071 ^ n24066;
  assign n24141 = n24072 ^ n24019;
  assign n24157 = n24156 ^ n24141;
  assign n24158 = n24106 & ~n24157;
  assign n24160 = n24159 ^ n24158;
  assign n24139 = n24138 ^ n24137;
  assign n23807 = n23806 ^ n23798;
  assign n23820 = n23819 ^ n23807;
  assign n23672 = n23671 ^ n23663;
  assign n23685 = n23684 ^ n23672;
  assign n23686 = n23685 ^ n23566;
  assign n23562 = n23561 ^ n23552;
  assign n23687 = n23686 ^ n23562;
  assign n23413 = n23412 ^ n23411;
  assign n23416 = n23415 ^ n23413;
  assign n23410 = n23404 ^ n23397;
  assign n23417 = n23416 ^ n23410;
  assign n23418 = n23417 ^ n23409;
  assign n23688 = n23687 ^ n23418;
  assign n23821 = n23820 ^ n23688;
  assign n23909 = n23908 ^ n23821;
  assign n24046 = n24045 ^ n23909;
  assign n24073 = n24072 ^ n23984;
  assign n24134 = n24133 ^ n24073;
  assign n24135 = n24046 & n24134;
  assign n23985 = n23984 ^ n23909;
  assign n24047 = n24046 ^ n24020;
  assign n24048 = n23985 & ~n24047;
  assign n24136 = n24135 ^ n24048;
  assign n24140 = n24139 ^ n24136;
  assign n24161 = n24160 ^ n24140;
  assign n24163 = n24133 ^ n24046;
  assign n24188 = n24163 ^ n24073;
  assign n24189 = n24188 ^ n24136;
  assign n24183 = n24157 ^ n24106;
  assign n24184 = n24183 ^ n24162;
  assign n24185 = n24163 ^ n24156;
  assign n24186 = n24184 & n24185;
  assign n24177 = n24137 ^ n23985;
  assign n24178 = ~n24163 & ~n24177;
  assign n24187 = n24186 ^ n24178;
  assign n24190 = n24189 ^ n24187;
  assign n24191 = ~n24161 & n24190;
  assign n24169 = n24157 ^ n24138;
  assign n24167 = n24157 ^ n23909;
  assign n24168 = n24167 ^ n24046;
  assign n24173 = n24169 ^ n24168;
  assign n24170 = ~n24168 & ~n24169;
  assign n24171 = n24170 ^ n24159;
  assign n24164 = n24163 ^ n24141;
  assign n24165 = n24162 & ~n24164;
  assign n24166 = n24165 ^ n24135;
  assign n24172 = n24171 ^ n24166;
  assign n24174 = n24173 ^ n24172;
  assign n24175 = n24174 ^ n24161;
  assign n24206 = n24191 ^ n24175;
  assign n24180 = n24164 ^ n24162;
  assign n24176 = ~n24156 & ~n24167;
  assign n24179 = n24178 ^ n24176;
  assign n24181 = n24180 ^ n24179;
  assign n24182 = n24181 ^ n24166;
  assign n24204 = ~n24161 & ~n24182;
  assign n24205 = ~n24174 & n24204;
  assign n24207 = n24206 ^ n24205;
  assign n24201 = n24182 & n24190;
  assign n24202 = n24174 & n24201;
  assign n24195 = n24190 ^ n24182;
  assign n24200 = n24195 ^ n24191;
  assign n24203 = n24202 ^ n24200;
  assign n24208 = n24207 ^ n24203;
  assign n26394 = n24162 & n24208;
  assign n24196 = n24191 ^ n24174;
  assign n24197 = ~n24195 & n24196;
  assign n24198 = n24197 ^ n24182;
  assign n24217 = n24203 ^ n24198;
  assign n24218 = ~n24137 & n24217;
  assign n24216 = ~n24164 & n24208;
  assign n24219 = n24218 ^ n24216;
  assign n26395 = n26394 ^ n24219;
  assign n24192 = n24191 ^ n24182;
  assign n24193 = ~n24175 & ~n24192;
  assign n24194 = n24193 ^ n24174;
  assign n24199 = n24198 ^ n24194;
  assign n26244 = n24134 & ~n24199;
  assign n24211 = n24046 & ~n24199;
  assign n26392 = n26244 ^ n24211;
  assign n24236 = n24207 ^ n24194;
  assign n24237 = ~n24163 & ~n24236;
  assign n24235 = ~n24156 & n24194;
  assign n24238 = n24237 ^ n24235;
  assign n24234 = ~n24168 & ~n24198;
  assign n24239 = n24238 ^ n24234;
  assign n26393 = n26392 ^ n24239;
  assign n26396 = n26395 ^ n26393;
  assign n26420 = n26419 ^ n26396;
  assign n23130 = n22899 & n22960;
  assign n23205 = n23130 ^ n22978;
  assign n23076 = n22922 & n22953;
  assign n23078 = n23077 ^ n23076;
  assign n23203 = n23078 ^ n22986;
  assign n23202 = n22965 ^ n21701;
  assign n23204 = n23203 ^ n23202;
  assign n23206 = n23205 ^ n23204;
  assign n22795 = n22794 ^ n22787;
  assign n22774 = n22724 ^ n22663;
  assign n22782 = n22781 ^ n22774;
  assign n22796 = n22795 ^ n22782;
  assign n22694 = n22693 ^ n22683;
  assign n22664 = n22663 ^ n22658;
  assign n22678 = n22677 ^ n22664;
  assign n22695 = n22694 ^ n22678;
  assign n22797 = n22796 ^ n22695;
  assign n22770 = n22769 ^ n22441;
  assign n22762 = n22761 ^ n22091;
  assign n22771 = n22770 ^ n22762;
  assign n22798 = n22797 ^ n22771;
  assign n22654 = n22653 ^ n22638;
  assign n22611 = n22573 ^ n22073;
  assign n22635 = n22634 ^ n22611;
  assign n22655 = n22654 ^ n22635;
  assign n22696 = n22695 ^ n22655;
  assign n22608 = n22607 ^ n22592;
  assign n22581 = n22580 ^ n22574;
  assign n22609 = n22608 ^ n22581;
  assign n22541 = n22540 ^ n22452;
  assign n22092 = n22091 ^ n22073;
  assign n22325 = n22324 ^ n22092;
  assign n22542 = n22541 ^ n22325;
  assign n22566 = n22565 ^ n22542;
  assign n22610 = n22609 ^ n22566;
  assign n22697 = n22696 ^ n22610;
  assign n22830 = n22798 ^ n22697;
  assign n22747 = n22746 ^ n22738;
  assign n22725 = n22724 ^ n22090;
  assign n22735 = n22734 ^ n22725;
  assign n22748 = n22747 ^ n22735;
  assign n22720 = n22719 ^ n22712;
  assign n22699 = n22698 ^ n22658;
  assign n22707 = n22706 ^ n22699;
  assign n22721 = n22720 ^ n22707;
  assign n22749 = n22748 ^ n22721;
  assign n22750 = n22749 ^ n22610;
  assign n22819 = n22797 ^ n22750;
  assign n22773 = n22748 ^ n22655;
  assign n22825 = n22819 ^ n22773;
  assign n22822 = n22798 ^ n22721;
  assign n22823 = ~n22771 & ~n22822;
  assign n22752 = n22721 ^ n22655;
  assign n22751 = n22748 ^ n22542;
  assign n22753 = n22752 ^ n22751;
  assign n22754 = ~n22750 & ~n22753;
  assign n22824 = n22823 ^ n22754;
  assign n22826 = n22825 ^ n22824;
  assign n22820 = n22773 & ~n22819;
  assign n22803 = n22796 ^ n22655;
  assign n22804 = n22803 ^ n22610;
  assign n22805 = n22749 & n22804;
  assign n22821 = n22820 ^ n22805;
  assign n22827 = n22826 ^ n22821;
  assign n22809 = n22803 ^ n22750;
  assign n22806 = n22749 ^ n22696;
  assign n22807 = n22752 & ~n22806;
  assign n22808 = n22807 ^ n22805;
  assign n22810 = n22809 ^ n22808;
  assign n22772 = n22771 ^ n22750;
  assign n22799 = n22798 ^ n22542;
  assign n22800 = n22799 ^ n22773;
  assign n22801 = n22772 & n22800;
  assign n22802 = n22801 ^ n22754;
  assign n22811 = n22810 ^ n22802;
  assign n22828 = n22827 ^ n22811;
  assign n22831 = n22822 ^ n22749;
  assign n22835 = n22831 ^ n22830;
  assign n22832 = ~n22830 & ~n22831;
  assign n22814 = n22697 & ~n22751;
  assign n22833 = n22832 ^ n22814;
  assign n22834 = n22833 ^ n22821;
  assign n22836 = n22835 ^ n22834;
  assign n22815 = n22542 & ~n22798;
  assign n22816 = n22815 ^ n22814;
  assign n22812 = n22751 ^ n22697;
  assign n22813 = n22812 ^ n22808;
  assign n22817 = n22816 ^ n22813;
  assign n22818 = n22811 & ~n22817;
  assign n22840 = n22836 ^ n22818;
  assign n22841 = ~n22828 & n22840;
  assign n22842 = n22841 ^ n22827;
  assign n23124 = ~n22830 & ~n22842;
  assign n22845 = n22836 ^ n22817;
  assign n22846 = n22827 ^ n22818;
  assign n22847 = ~n22845 & ~n22846;
  assign n22848 = n22847 ^ n22836;
  assign n22873 = ~n22771 & n22848;
  assign n23199 = n23124 ^ n22873;
  assign n22853 = n22845 ^ n22818;
  assign n22851 = ~n22817 & ~n22827;
  assign n22852 = ~n22836 & n22851;
  assign n22854 = n22853 ^ n22852;
  assign n22871 = n22854 ^ n22848;
  assign n23070 = ~n22753 & ~n22871;
  assign n23069 = n22772 & ~n22854;
  assign n23071 = n23070 ^ n23069;
  assign n23200 = n23199 ^ n23071;
  assign n22868 = n22800 & ~n22854;
  assign n22837 = n22811 & n22827;
  assign n22838 = n22836 & n22837;
  assign n22829 = n22828 ^ n22818;
  assign n22839 = n22838 ^ n22829;
  assign n22867 = ~n22798 & ~n22839;
  assign n22869 = n22868 ^ n22867;
  assign n22855 = n22854 ^ n22839;
  assign n22849 = n22848 ^ n22842;
  assign n22856 = n22855 ^ n22849;
  assign n22857 = n22752 & ~n22856;
  assign n22850 = n22749 & ~n22849;
  assign n22858 = n22857 ^ n22850;
  assign n23198 = n22869 ^ n22858;
  assign n23201 = n23200 ^ n23198;
  assign n23207 = n23206 ^ n23201;
  assign n21849 = n21848 ^ n21845;
  assign n21839 = n21838 ^ n21837;
  assign n21843 = n21842 ^ n21839;
  assign n21850 = n21849 ^ n21843;
  assign n21828 = n21827 ^ n21818;
  assign n21812 = n21811 ^ n21805;
  assign n21829 = n21828 ^ n21812;
  assign n21782 = n21781 ^ n21774;
  assign n21768 = n21767 ^ n21755;
  assign n21783 = n21782 ^ n21768;
  assign n21830 = n21829 ^ n21783;
  assign n21799 = n21798 ^ n21794;
  assign n21791 = n21790 ^ n21789;
  assign n21800 = n21799 ^ n21791;
  assign n21831 = n21830 ^ n21800;
  assign n21851 = n21850 ^ n21831;
  assign n21869 = n21868 ^ n21864;
  assign n21860 = n21859 ^ n21855;
  assign n21870 = n21869 ^ n21860;
  assign n21871 = n21870 ^ n21850;
  assign n21907 = n21871 ^ n21851;
  assign n21745 = n21744 ^ n21740;
  assign n21728 = n21727 ^ n21715;
  assign n21746 = n21745 ^ n21728;
  assign n21784 = n21783 ^ n21746;
  assign n21702 = n21701 ^ n21689;
  assign n21678 = n21677 ^ n21669;
  assign n21703 = n21702 ^ n21678;
  assign n21638 = n21637 ^ n21552;
  assign n21304 = n21303 ^ n21168;
  assign n21430 = n21429 ^ n21304;
  assign n21639 = n21638 ^ n21430;
  assign n21658 = n21657 ^ n21639;
  assign n21704 = n21703 ^ n21658;
  assign n21785 = n21784 ^ n21704;
  assign n21832 = n21831 ^ n21785;
  assign n21911 = n21907 ^ n21832;
  assign n21908 = ~n21832 & ~n21907;
  assign n21874 = n21870 ^ n21639;
  assign n21902 = n21785 & ~n21874;
  assign n21909 = n21908 ^ n21902;
  assign n21883 = n21829 ^ n21746;
  assign n21884 = n21883 ^ n21704;
  assign n21885 = ~n21871 & n21884;
  assign n21872 = n21871 ^ n21704;
  assign n21878 = n21872 ^ n21830;
  assign n21879 = n21870 ^ n21746;
  assign n21882 = ~n21878 & ~n21879;
  assign n21886 = n21885 ^ n21882;
  assign n21910 = n21909 ^ n21886;
  assign n21912 = n21911 ^ n21910;
  assign n21903 = n21639 & ~n21831;
  assign n21904 = n21903 ^ n21902;
  assign n21900 = n21874 ^ n21785;
  assign n21873 = n21850 ^ n21746;
  assign n21894 = n21871 ^ n21784;
  assign n21895 = n21873 & ~n21894;
  assign n21896 = n21895 ^ n21885;
  assign n21901 = n21900 ^ n21896;
  assign n21905 = n21904 ^ n21901;
  assign n21923 = n21912 ^ n21905;
  assign n21893 = n21883 ^ n21872;
  assign n21897 = n21896 ^ n21893;
  assign n21888 = n21831 ^ n21639;
  assign n21889 = n21888 ^ n21879;
  assign n21890 = n21872 ^ n21800;
  assign n21891 = ~n21889 & n21890;
  assign n21875 = n21874 ^ n21873;
  assign n21876 = ~n21872 & ~n21875;
  assign n21892 = n21891 ^ n21876;
  assign n21898 = n21897 ^ n21892;
  assign n21906 = ~n21898 & ~n21905;
  assign n21880 = n21879 ^ n21878;
  assign n21852 = ~n21800 & n21851;
  assign n21877 = n21876 ^ n21852;
  assign n21881 = n21880 ^ n21877;
  assign n21887 = n21886 ^ n21881;
  assign n21924 = n21906 ^ n21887;
  assign n21925 = ~n21923 & n21924;
  assign n21926 = n21925 ^ n21912;
  assign n23192 = n21851 & n21926;
  assign n21930 = n21923 ^ n21906;
  assign n21928 = n21887 & ~n21905;
  assign n21929 = ~n21912 & n21928;
  assign n21931 = n21930 ^ n21929;
  assign n23010 = ~n21889 & ~n21931;
  assign n21899 = n21898 ^ n21887;
  assign n21919 = n21906 ^ n21899;
  assign n21917 = ~n21887 & ~n21898;
  assign n21918 = n21912 & n21917;
  assign n21920 = n21919 ^ n21918;
  assign n21944 = ~n21831 & ~n21920;
  assign n23011 = n23010 ^ n21944;
  assign n23193 = n23192 ^ n23011;
  assign n23050 = ~n21800 & n21926;
  assign n23005 = n21931 ^ n21926;
  assign n23008 = ~n21872 & ~n23005;
  assign n23139 = n23050 ^ n23008;
  assign n21913 = n21912 ^ n21906;
  assign n21914 = ~n21899 & n21913;
  assign n21915 = n21914 ^ n21887;
  assign n23138 = ~n21907 & n21915;
  assign n23140 = n23139 ^ n23138;
  assign n23194 = n23193 ^ n23140;
  assign n21935 = n21920 ^ n21915;
  assign n23013 = n21785 & ~n21935;
  assign n21927 = n21926 ^ n21915;
  assign n21942 = ~n21871 & n21927;
  assign n21932 = n21931 ^ n21920;
  assign n21933 = n21932 ^ n21927;
  assign n21941 = n21873 & n21933;
  assign n21943 = n21942 ^ n21941;
  assign n23014 = n23013 ^ n21943;
  assign n21937 = ~n21878 & n21932;
  assign n21936 = ~n21874 & ~n21935;
  assign n21938 = n21937 ^ n21936;
  assign n21934 = ~n21894 & n21933;
  assign n21939 = n21938 ^ n21934;
  assign n23191 = n23014 ^ n21939;
  assign n23195 = n23194 ^ n23191;
  assign n23055 = n21884 & n21927;
  assign n23056 = n23055 ^ n21934;
  assign n23057 = n23056 ^ n23011;
  assign n23006 = ~n21875 & ~n23005;
  assign n23054 = n23014 ^ n23006;
  assign n23058 = n23057 ^ n23054;
  assign n23196 = n23195 ^ n23058;
  assign n20947 = n20946 ^ n20942;
  assign n20951 = n20950 ^ n20947;
  assign n20957 = n20956 ^ n20951;
  assign n20811 = n20810 ^ n20803;
  assign n20819 = n20818 ^ n20811;
  assign n20827 = n20826 ^ n20819;
  assign n20837 = n20836 ^ n20827;
  assign n20958 = n20957 ^ n20837;
  assign n20906 = n20905 ^ n20904;
  assign n20900 = n20899 ^ n20893;
  assign n20907 = n20906 ^ n20900;
  assign n20884 = n20883 ^ n20875;
  assign n20751 = n20750 ^ n20740;
  assign n20731 = n20730 ^ n20487;
  assign n20724 = n20723 ^ n20715;
  assign n20732 = n20731 ^ n20724;
  assign n20752 = n20751 ^ n20732;
  assign n20885 = n20884 ^ n20752;
  assign n20908 = n20907 ^ n20885;
  assign n20959 = n20958 ^ n20908;
  assign n20794 = n20793 ^ n20783;
  assign n20774 = n20773 ^ n20765;
  assign n20775 = n20774 ^ n20486;
  assign n20795 = n20794 ^ n20775;
  assign n20976 = n20837 ^ n20795;
  assign n20916 = n20915 ^ n20911;
  assign n20922 = n20921 ^ n20916;
  assign n20926 = n20925 ^ n20922;
  assign n20932 = n20931 ^ n20926;
  assign n20934 = n20932 ^ n20795;
  assign n20974 = n20934 ^ n20908;
  assign n20854 = n20853 ^ n20842;
  assign n20860 = n20859 ^ n20854;
  assign n20868 = n20867 ^ n20860;
  assign n20963 = n20957 ^ n20868;
  assign n20975 = n20974 ^ n20963;
  assign n20996 = n20976 ^ n20975;
  assign n20703 = n20702 ^ n20615;
  assign n20344 = n20343 ^ n20220;
  assign n20488 = n20487 ^ n20344;
  assign n20704 = n20703 ^ n20488;
  assign n20964 = n20963 ^ n20704;
  assign n20969 = n20964 ^ n20932;
  assign n20994 = ~n20704 & ~n20969;
  assign n20933 = n20932 ^ n20837;
  assign n20796 = n20795 ^ n20752;
  assign n20987 = n20933 ^ n20796;
  assign n20988 = ~n20974 & ~n20987;
  assign n20995 = n20994 ^ n20988;
  assign n20997 = n20996 ^ n20995;
  assign n20977 = ~n20975 & n20976;
  assign n20960 = n20934 & n20959;
  assign n20978 = n20977 ^ n20960;
  assign n20998 = n20997 ^ n20978;
  assign n20990 = n20974 ^ n20958;
  assign n20869 = n20868 ^ n20837;
  assign n20935 = n20934 ^ n20869;
  assign n20936 = n20933 & ~n20935;
  assign n20961 = n20960 ^ n20936;
  assign n20991 = n20990 ^ n20961;
  assign n20983 = n20964 ^ n20752;
  assign n20984 = n20983 ^ n20976;
  assign n20985 = n20974 ^ n20704;
  assign n20986 = n20984 & n20985;
  assign n20989 = n20988 ^ n20986;
  assign n20992 = n20991 ^ n20989;
  assign n21010 = n20998 ^ n20992;
  assign n20909 = n20908 ^ n20869;
  assign n20966 = ~n20796 & n20909;
  assign n20965 = n20752 & ~n20964;
  assign n20967 = n20966 ^ n20965;
  assign n20910 = n20909 ^ n20796;
  assign n20962 = n20961 ^ n20910;
  assign n20968 = n20967 ^ n20962;
  assign n20993 = ~n20968 & n20992;
  assign n20971 = n20964 ^ n20909;
  assign n20970 = n20969 ^ n20934;
  assign n20980 = n20971 ^ n20970;
  assign n20972 = ~n20970 & ~n20971;
  assign n20973 = n20972 ^ n20966;
  assign n20979 = n20978 ^ n20973;
  assign n20981 = n20980 ^ n20979;
  assign n21011 = n20993 ^ n20981;
  assign n21012 = ~n21010 & n21011;
  assign n21013 = n21012 ^ n20998;
  assign n20982 = n20981 ^ n20968;
  assign n20999 = n20998 ^ n20993;
  assign n21000 = ~n20982 & ~n20999;
  assign n21001 = n21000 ^ n20981;
  assign n21026 = n21013 ^ n21001;
  assign n22991 = n20959 & ~n21026;
  assign n21017 = n20992 & n20998;
  assign n21018 = n20981 & n21017;
  assign n21016 = n21010 ^ n20993;
  assign n21019 = n21018 ^ n21016;
  assign n21005 = n20993 ^ n20982;
  assign n21003 = ~n20968 & ~n20998;
  assign n21004 = ~n20981 & n21003;
  assign n21006 = n21005 ^ n21004;
  assign n21028 = n21019 ^ n21006;
  assign n21029 = n21028 ^ n21026;
  assign n21035 = ~n20935 & ~n21029;
  assign n23045 = n22991 ^ n21035;
  assign n21021 = n20984 & ~n21006;
  assign n21020 = ~n20964 & ~n21019;
  assign n21022 = n21021 ^ n21020;
  assign n23046 = n23045 ^ n21022;
  assign n21007 = n21006 ^ n21001;
  assign n23017 = ~n20987 & ~n21007;
  assign n21032 = n21019 ^ n21013;
  assign n21033 = n20909 & n21032;
  assign n21030 = n20933 & ~n21029;
  assign n21027 = n20934 & ~n21026;
  assign n21031 = n21030 ^ n21027;
  assign n21034 = n21033 ^ n21031;
  assign n23044 = n23017 ^ n21034;
  assign n23047 = n23046 ^ n23044;
  assign n21037 = ~n20975 & n21028;
  assign n21036 = ~n20796 & n21032;
  assign n21038 = n21037 ^ n21036;
  assign n21039 = n21038 ^ n21035;
  assign n21040 = n21039 ^ n21034;
  assign n21023 = ~n20969 & n21001;
  assign n21024 = n21023 ^ n21022;
  assign n21014 = ~n20970 & ~n21013;
  assign n21008 = ~n20974 & ~n21007;
  assign n21002 = ~n20704 & n21001;
  assign n21009 = n21008 ^ n21002;
  assign n21015 = n21014 ^ n21009;
  assign n21025 = n21024 ^ n21015;
  assign n21041 = n21040 ^ n21025;
  assign n23190 = n23047 ^ n21041;
  assign n23197 = n23196 ^ n23190;
  assign n23208 = n23207 ^ n23197;
  assign n23184 = n22984 ^ n22965;
  assign n23129 = n22923 & n22948;
  assign n23131 = n23130 ^ n23129;
  assign n22974 = n22973 ^ n22972;
  assign n23183 = n23131 ^ n22974;
  assign n23185 = n23184 ^ n23183;
  assign n23186 = n23185 ^ n21637;
  assign n23123 = n22799 & ~n22839;
  assign n23125 = n23124 ^ n23123;
  assign n22863 = ~n22806 & ~n22856;
  assign n22843 = n22842 ^ n22839;
  assign n22861 = ~n22751 & n22843;
  assign n22860 = ~n22819 & n22855;
  assign n22862 = n22861 ^ n22860;
  assign n22864 = n22863 ^ n22862;
  assign n23181 = n23125 ^ n22864;
  assign n23180 = n22867 ^ n22858;
  assign n23182 = n23181 ^ n23180;
  assign n23187 = n23186 ^ n23182;
  assign n20017 = n20016 ^ n19943;
  assign n20008 = n20007 ^ n20000;
  assign n20018 = n20017 ^ n20008;
  assign n19912 = n19911 ^ n19900;
  assign n19895 = n19894 ^ n19881;
  assign n19913 = n19912 ^ n19895;
  assign n20019 = n20018 ^ n19913;
  assign n19975 = n17805 ^ n16817;
  assign n19979 = n19978 ^ n19975;
  assign n19983 = n19982 ^ n19979;
  assign n19992 = n19991 ^ n19983;
  assign n20020 = n20019 ^ n19992;
  assign n19871 = n19870 ^ n19799;
  assign n19853 = n19852 ^ n19650;
  assign n19849 = n19848 ^ n19837;
  assign n19854 = n19853 ^ n19849;
  assign n19872 = n19871 ^ n19854;
  assign n19914 = n19913 ^ n19872;
  assign n19824 = n19823 ^ n19812;
  assign n19801 = n19800 ^ n19792;
  assign n19825 = n19824 ^ n19801;
  assign n19780 = n19779 ^ n19763;
  assign n19756 = n19755 ^ n19650;
  assign n17806 = n17805 ^ n16828;
  assign n19644 = n19643 ^ n17806;
  assign n19757 = n19756 ^ n19644;
  assign n19781 = n19780 ^ n19757;
  assign n19826 = n19825 ^ n19781;
  assign n19915 = n19914 ^ n19826;
  assign n20052 = n20020 ^ n19915;
  assign n19967 = n19966 ^ n17804;
  assign n19957 = n19956 ^ n19947;
  assign n19968 = n19967 ^ n19957;
  assign n19939 = n19938 ^ n19880;
  assign n19922 = n19921 ^ n19920;
  assign n19930 = n19929 ^ n19922;
  assign n19940 = n19939 ^ n19930;
  assign n19969 = n19968 ^ n19940;
  assign n19970 = n19969 ^ n19826;
  assign n20041 = n20019 ^ n19970;
  assign n19994 = n19968 ^ n19872;
  assign n20047 = n20041 ^ n19994;
  assign n20044 = n20020 ^ n19940;
  assign n20045 = ~n19992 & ~n20044;
  assign n19972 = n19940 ^ n19872;
  assign n19971 = n19968 ^ n19757;
  assign n19973 = n19972 ^ n19971;
  assign n19974 = ~n19970 & ~n19973;
  assign n20046 = n20045 ^ n19974;
  assign n20048 = n20047 ^ n20046;
  assign n20042 = n19994 & ~n20041;
  assign n20025 = n20018 ^ n19872;
  assign n20026 = n20025 ^ n19826;
  assign n20027 = n19969 & n20026;
  assign n20043 = n20042 ^ n20027;
  assign n20049 = n20048 ^ n20043;
  assign n20031 = n20025 ^ n19970;
  assign n20028 = n19969 ^ n19914;
  assign n20029 = n19972 & ~n20028;
  assign n20030 = n20029 ^ n20027;
  assign n20032 = n20031 ^ n20030;
  assign n19993 = n19992 ^ n19970;
  assign n20021 = n20020 ^ n19757;
  assign n20022 = n20021 ^ n19994;
  assign n20023 = n19993 & n20022;
  assign n20024 = n20023 ^ n19974;
  assign n20033 = n20032 ^ n20024;
  assign n20050 = n20049 ^ n20033;
  assign n20053 = n20044 ^ n19969;
  assign n20057 = n20053 ^ n20052;
  assign n20054 = ~n20052 & ~n20053;
  assign n20036 = n19915 & ~n19971;
  assign n20055 = n20054 ^ n20036;
  assign n20056 = n20055 ^ n20043;
  assign n20058 = n20057 ^ n20056;
  assign n20037 = n19757 & ~n20020;
  assign n20038 = n20037 ^ n20036;
  assign n20034 = n19971 ^ n19915;
  assign n20035 = n20034 ^ n20030;
  assign n20039 = n20038 ^ n20035;
  assign n20040 = n20033 & ~n20039;
  assign n20062 = n20058 ^ n20040;
  assign n20063 = ~n20050 & n20062;
  assign n20064 = n20063 ^ n20049;
  assign n23112 = ~n20052 & ~n20064;
  assign n20059 = n20033 & n20049;
  assign n20060 = n20058 & n20059;
  assign n20051 = n20050 ^ n20040;
  assign n20061 = n20060 ^ n20051;
  assign n23111 = n20021 & ~n20061;
  assign n23113 = n23112 ^ n23111;
  assign n20067 = n20058 ^ n20039;
  assign n20075 = n20067 ^ n20040;
  assign n20073 = ~n20039 & ~n20049;
  assign n20074 = ~n20058 & n20073;
  assign n20076 = n20075 ^ n20074;
  assign n20077 = n20076 ^ n20061;
  assign n20068 = n20049 ^ n20040;
  assign n20069 = ~n20067 & ~n20068;
  assign n20070 = n20069 ^ n20058;
  assign n20071 = n20070 ^ n20064;
  assign n20078 = n20077 ^ n20071;
  assign n20085 = ~n20028 & ~n20078;
  assign n20065 = n20064 ^ n20061;
  assign n20083 = ~n19971 & n20065;
  assign n20082 = ~n20041 & n20077;
  assign n20084 = n20083 ^ n20082;
  assign n20086 = n20085 ^ n20084;
  assign n23176 = n23113 ^ n20086;
  assign n20090 = ~n20020 & ~n20061;
  assign n20079 = n19972 & ~n20078;
  assign n20072 = n19969 & ~n20071;
  assign n20080 = n20079 ^ n20072;
  assign n23175 = n20090 ^ n20080;
  assign n23177 = n23176 ^ n23175;
  assign n21951 = n21031 ^ n21020;
  assign n21948 = n20983 & ~n21019;
  assign n21947 = ~n20971 & ~n21013;
  assign n21949 = n21948 ^ n21947;
  assign n21950 = n21949 ^ n21039;
  assign n21952 = n21951 ^ n21950;
  assign n23178 = n23177 ^ n21952;
  assign n21921 = n21888 & ~n21920;
  assign n21916 = ~n21832 & n21915;
  assign n21922 = n21921 ^ n21916;
  assign n23171 = n23139 ^ n21922;
  assign n23170 = n23014 ^ n21936;
  assign n23172 = n23171 ^ n23170;
  assign n23173 = n23172 ^ n23058;
  assign n23117 = n21949 ^ n21009;
  assign n23116 = n21036 ^ n21034;
  assign n23118 = n23117 ^ n23116;
  assign n23169 = n23118 ^ n23047;
  assign n23174 = n23173 ^ n23169;
  assign n23179 = n23178 ^ n23174;
  assign n23188 = n23187 ^ n23179;
  assign n20095 = ~n19992 & n20070;
  assign n23165 = n23112 ^ n20095;
  assign n20093 = n20076 ^ n20070;
  assign n23062 = ~n19973 & ~n20093;
  assign n23061 = n19993 & ~n20076;
  assign n23063 = n23062 ^ n23061;
  assign n23166 = n23165 ^ n23063;
  assign n20089 = n20022 & ~n20076;
  assign n20091 = n20090 ^ n20089;
  assign n23164 = n20091 ^ n20080;
  assign n23167 = n23166 ^ n23164;
  assign n23042 = n21031 ^ n21022;
  assign n23040 = n21947 ^ n21002;
  assign n23016 = n20985 & ~n21006;
  assign n23018 = n23017 ^ n23016;
  assign n23041 = n23040 ^ n23018;
  assign n23043 = n23042 ^ n23041;
  assign n23168 = n23167 ^ n23043;
  assign n23189 = n23188 ^ n23168;
  assign n23209 = n23208 ^ n23189;
  assign n23024 = n22804 & ~n22849;
  assign n23098 = n23024 ^ n22863;
  assign n23099 = n23098 ^ n22869;
  assign n22844 = n22697 & n22843;
  assign n22859 = n22858 ^ n22844;
  assign n23097 = n23070 ^ n22859;
  assign n23100 = n23099 ^ n23097;
  assign n23106 = n23105 ^ n23100;
  assign n22997 = n20026 & ~n20071;
  assign n23092 = n22997 ^ n20085;
  assign n23093 = n23092 ^ n20091;
  assign n20066 = n19915 & n20065;
  assign n20081 = n20080 ^ n20066;
  assign n23091 = n23062 ^ n20081;
  assign n23094 = n23093 ^ n23091;
  assign n23095 = n23094 ^ n23047;
  assign n23088 = n23010 ^ n21943;
  assign n23004 = n21890 & ~n21931;
  assign n23007 = n23006 ^ n23004;
  assign n23009 = n23008 ^ n23007;
  assign n23087 = n23056 ^ n23009;
  assign n23089 = n23088 ^ n23087;
  assign n23085 = n21031 ^ n21021;
  assign n23019 = n23018 ^ n21008;
  assign n23084 = n23045 ^ n23019;
  assign n23086 = n23085 ^ n23084;
  assign n23090 = n23089 ^ n23086;
  assign n23096 = n23095 ^ n23090;
  assign n23107 = n23106 ^ n23096;
  assign n23079 = n23078 ^ n22977;
  assign n23080 = n23079 ^ n22986;
  assign n23075 = n22968 ^ n21848;
  assign n23081 = n23080 ^ n23075;
  assign n22872 = ~n22750 & ~n22871;
  assign n23072 = n23071 ^ n22872;
  assign n23073 = n23072 ^ n22869;
  assign n23074 = n23073 ^ n22859;
  assign n23082 = n23081 ^ n23074;
  assign n20094 = ~n19970 & ~n20093;
  assign n23064 = n23063 ^ n20094;
  assign n23065 = n23064 ^ n20091;
  assign n23066 = n23065 ^ n20081;
  assign n23020 = n23019 ^ n21022;
  assign n23021 = n23020 ^ n21034;
  assign n23067 = n23066 ^ n23021;
  assign n23051 = n23050 ^ n21916;
  assign n23052 = n23051 ^ n23007;
  assign n23049 = n23011 ^ n21943;
  assign n23053 = n23052 ^ n23049;
  assign n23059 = n23058 ^ n23053;
  assign n23048 = n23047 ^ n23043;
  assign n23060 = n23059 ^ n23048;
  assign n23068 = n23067 ^ n23060;
  assign n23083 = n23082 ^ n23068;
  assign n23108 = n23107 ^ n23083;
  assign n23210 = n23209 ^ n23108;
  assign n23027 = n22773 & n22855;
  assign n23028 = n23027 ^ n22862;
  assign n23025 = n23024 ^ n22850;
  assign n22875 = ~n22831 & ~n22842;
  assign n22874 = n22873 ^ n22872;
  assign n22876 = n22875 ^ n22874;
  assign n23026 = n23025 ^ n22876;
  assign n23029 = n23028 ^ n23026;
  assign n23037 = n23036 ^ n23029;
  assign n23012 = n23011 ^ n23009;
  assign n23015 = n23014 ^ n23012;
  assign n23022 = n23021 ^ n23015;
  assign n23000 = n19994 & n20077;
  assign n23001 = n23000 ^ n20084;
  assign n22998 = n22997 ^ n20072;
  assign n20097 = ~n20053 & ~n20064;
  assign n20096 = n20095 ^ n20094;
  assign n20098 = n20097 ^ n20096;
  assign n22999 = n22998 ^ n20098;
  assign n23002 = n23001 ^ n22999;
  assign n22994 = n20976 & n21028;
  assign n22995 = n22994 ^ n21038;
  assign n22992 = n22991 ^ n21027;
  assign n22993 = n22992 ^ n21015;
  assign n22996 = n22995 ^ n22993;
  assign n23003 = n23002 ^ n22996;
  assign n23023 = n23022 ^ n23003;
  assign n23038 = n23037 ^ n23023;
  assign n22983 = n22900 & n22957;
  assign n22987 = n22986 ^ n22983;
  assign n22981 = n22980 ^ n22974;
  assign n22969 = n22968 ^ n21727;
  assign n22982 = n22981 ^ n22969;
  assign n22988 = n22987 ^ n22982;
  assign n22866 = ~n22822 & n22848;
  assign n22870 = n22869 ^ n22866;
  assign n22877 = n22876 ^ n22870;
  assign n22865 = n22864 ^ n22859;
  assign n22878 = n22877 ^ n22865;
  assign n22989 = n22988 ^ n22878;
  assign n21945 = n21944 ^ n21943;
  assign n21940 = n21939 ^ n21922;
  assign n21946 = n21945 ^ n21940;
  assign n21953 = n21952 ^ n21946;
  assign n20088 = ~n20044 & n20070;
  assign n20092 = n20091 ^ n20088;
  assign n20099 = n20098 ^ n20092;
  assign n20087 = n20086 ^ n20081;
  assign n20100 = n20099 ^ n20087;
  assign n21042 = n21041 ^ n20100;
  assign n21954 = n21953 ^ n21042;
  assign n22990 = n22989 ^ n21954;
  assign n23039 = n23038 ^ n22990;
  assign n23237 = n23209 ^ n23039;
  assign n23155 = n22985 ^ n22965;
  assign n23154 = n23102 ^ n23079;
  assign n23156 = n23155 ^ n23154;
  assign n23157 = n23156 ^ n21811;
  assign n23152 = n22868 ^ n22858;
  assign n23151 = n23098 ^ n23072;
  assign n23153 = n23152 ^ n23151;
  assign n23158 = n23157 ^ n23153;
  assign n23147 = n20089 ^ n20080;
  assign n23146 = n23092 ^ n23064;
  assign n23148 = n23147 ^ n23146;
  assign n23149 = n23148 ^ n23086;
  assign n23142 = ~n21879 & n21932;
  assign n23143 = n23142 ^ n21938;
  assign n23137 = n23055 ^ n21942;
  assign n23141 = n23140 ^ n23137;
  assign n23144 = n23143 ^ n23141;
  assign n23145 = n23144 ^ n22996;
  assign n23150 = n23149 ^ n23145;
  assign n23159 = n23158 ^ n23150;
  assign n23160 = n23159 ^ n23038;
  assign n23132 = n23131 ^ n22979;
  assign n23128 = n22971 ^ n22968;
  assign n23133 = n23132 ^ n23128;
  assign n23134 = n23133 ^ n21798;
  assign n23126 = n23125 ^ n22874;
  assign n23122 = n22861 ^ n22859;
  assign n23127 = n23126 ^ n23122;
  assign n23135 = n23134 ^ n23127;
  assign n23120 = n23058 ^ n23047;
  assign n23114 = n23113 ^ n20096;
  assign n23110 = n20083 ^ n20081;
  assign n23115 = n23114 ^ n23110;
  assign n23119 = n23118 ^ n23115;
  assign n23121 = n23120 ^ n23119;
  assign n23136 = n23135 ^ n23121;
  assign n23161 = n23160 ^ n23136;
  assign n23247 = n23237 ^ n23161;
  assign n23162 = n23161 ^ n23083;
  assign n23246 = n23162 ^ n23108;
  assign n23251 = n23247 ^ n23246;
  assign n23248 = ~n23246 & n23247;
  assign n23212 = n23188 ^ n23107;
  assign n23241 = ~n23212 & n23237;
  assign n23249 = n23248 ^ n23241;
  assign n23216 = n23107 ^ n22990;
  assign n23217 = n23210 ^ n23160;
  assign n23223 = n23216 & ~n23217;
  assign n23220 = n23159 ^ n22990;
  assign n23221 = n23220 ^ n23209;
  assign n23222 = n23108 & n23221;
  assign n23224 = n23223 ^ n23222;
  assign n23250 = n23249 ^ n23224;
  assign n23252 = n23251 ^ n23250;
  assign n23240 = n23161 & ~n23188;
  assign n23242 = n23241 ^ n23240;
  assign n23238 = n23237 ^ n23212;
  assign n23109 = n23108 ^ n23039;
  assign n23211 = n23083 ^ n22990;
  assign n23232 = ~n23109 & n23211;
  assign n23233 = n23232 ^ n23222;
  assign n23239 = n23238 ^ n23233;
  assign n23243 = n23242 ^ n23239;
  assign n23258 = n23252 ^ n23243;
  assign n23231 = n23220 ^ n23210;
  assign n23234 = n23233 ^ n23231;
  assign n23226 = n23188 ^ n23161;
  assign n23227 = n23226 ^ n23216;
  assign n23228 = n23210 ^ n23136;
  assign n23229 = n23227 & ~n23228;
  assign n23213 = n23212 ^ n23211;
  assign n23214 = ~n23210 & ~n23213;
  assign n23230 = n23229 ^ n23214;
  assign n23235 = n23234 ^ n23230;
  assign n23244 = n23235 & ~n23243;
  assign n23218 = n23217 ^ n23216;
  assign n23163 = n23136 & ~n23162;
  assign n23215 = n23214 ^ n23163;
  assign n23219 = n23218 ^ n23215;
  assign n23225 = n23224 ^ n23219;
  assign n23265 = n23244 ^ n23225;
  assign n23266 = n23258 & ~n23265;
  assign n23267 = n23266 ^ n23252;
  assign n23259 = n23258 ^ n23244;
  assign n23256 = ~n23225 & ~n23243;
  assign n23257 = n23252 & n23256;
  assign n23260 = n23259 ^ n23257;
  assign n26223 = n23267 ^ n23260;
  assign n26278 = ~n23210 & ~n26223;
  assign n26224 = ~n23213 & ~n26223;
  assign n26222 = ~n23228 & n23260;
  assign n26225 = n26224 ^ n26222;
  assign n26339 = n26278 ^ n26225;
  assign n26217 = n23227 & n23260;
  assign n23253 = n23225 & n23235;
  assign n23254 = ~n23252 & n23253;
  assign n23236 = n23235 ^ n23225;
  assign n23245 = n23244 ^ n23236;
  assign n23255 = n23254 ^ n23245;
  assign n23283 = n23161 & ~n23255;
  assign n26218 = n26217 ^ n23283;
  assign n26412 = n26339 ^ n26218;
  assign n23262 = n23252 ^ n23244;
  assign n23263 = ~n23236 & ~n23262;
  assign n23264 = n23263 ^ n23225;
  assign n23271 = n23264 ^ n23255;
  assign n26228 = n23237 & n23271;
  assign n23268 = n23267 ^ n23264;
  assign n23281 = n23108 & n23268;
  assign n23261 = n23260 ^ n23255;
  assign n23269 = n23268 ^ n23261;
  assign n23280 = n23211 & ~n23269;
  assign n23282 = n23281 ^ n23280;
  assign n26229 = n26228 ^ n23282;
  assign n26413 = n26412 ^ n26229;
  assign n26239 = ~n24177 & ~n24236;
  assign n26238 = n24185 & ~n24207;
  assign n26240 = n26239 ^ n26238;
  assign n26256 = n26240 ^ n24237;
  assign n24231 = n24184 & ~n24207;
  assign n24213 = ~n24157 & ~n24203;
  assign n24232 = n24231 ^ n24213;
  assign n26257 = n26256 ^ n24232;
  assign n24227 = n24138 & n24217;
  assign n24209 = n24208 ^ n24199;
  assign n24210 = n23985 & ~n24209;
  assign n24212 = n24211 ^ n24210;
  assign n24228 = n24227 ^ n24212;
  assign n26258 = n26257 ^ n24228;
  assign n26414 = n26413 ^ n26258;
  assign n26421 = n26420 ^ n26414;
  assign n26434 = n26433 ^ n26421;
  assign n26407 = n26211 ^ n26191;
  assign n26268 = n26150 & n26179;
  assign n26270 = n26269 ^ n26268;
  assign n26271 = n26270 ^ n26203;
  assign n26406 = n26361 ^ n26271;
  assign n26408 = n26407 ^ n26406;
  assign n26409 = n26408 ^ n23157;
  assign n26094 = n26054 & ~n26077;
  assign n26079 = n26078 ^ n26069;
  assign n26087 = n25909 & ~n26079;
  assign n26089 = n26088 ^ n26087;
  assign n26404 = n26094 ^ n26089;
  assign n26080 = ~n25908 & ~n26079;
  assign n26356 = n26355 ^ n26080;
  assign n26262 = n26055 & ~n26077;
  assign n26261 = ~n26047 & ~n26098;
  assign n26263 = n26262 ^ n26261;
  assign n26264 = n26263 ^ n26099;
  assign n26403 = n26356 ^ n26264;
  assign n26405 = n26404 ^ n26403;
  assign n26410 = n26409 ^ n26405;
  assign n25168 = n25128 & ~n25151;
  assign n25153 = n25152 ^ n25143;
  assign n25161 = n24987 & ~n25153;
  assign n25163 = n25162 ^ n25161;
  assign n26399 = n25168 ^ n25163;
  assign n25154 = ~n24986 & ~n25153;
  assign n26349 = n26348 ^ n25154;
  assign n26251 = n25129 & ~n25151;
  assign n26250 = ~n25121 & ~n25172;
  assign n26252 = n26251 ^ n26250;
  assign n26253 = n26252 ^ n25173;
  assign n26398 = n26349 ^ n26253;
  assign n26400 = n26399 ^ n26398;
  assign n26344 = n24231 ^ n24212;
  assign n24215 = ~n24047 & ~n24209;
  assign n26245 = n26244 ^ n24215;
  assign n26343 = n26256 ^ n26245;
  assign n26345 = n26344 ^ n26343;
  assign n26401 = n26400 ^ n26345;
  assign n26389 = n23216 & ~n23261;
  assign n23273 = ~n23217 & ~n23261;
  assign n23272 = ~n23212 & n23271;
  assign n23274 = n23273 ^ n23272;
  assign n26390 = n26389 ^ n23274;
  assign n26231 = n23221 & n23268;
  assign n26387 = n26231 ^ n23281;
  assign n26320 = ~n23246 & ~n23264;
  assign n26220 = n23136 & ~n23267;
  assign n26279 = n26278 ^ n26220;
  assign n26321 = n26320 ^ n26279;
  assign n26388 = n26387 ^ n26321;
  assign n26391 = n26390 ^ n26388;
  assign n26397 = n26396 ^ n26391;
  assign n26402 = n26401 ^ n26397;
  assign n26411 = n26410 ^ n26402;
  assign n26435 = n26434 ^ n26411;
  assign n26303 = n26125 & n26186;
  assign n26302 = n26148 & n26174;
  assign n26304 = n26303 ^ n26302;
  assign n26382 = n26304 ^ n26205;
  assign n26381 = n26197 ^ n26194;
  assign n26383 = n26382 ^ n26381;
  assign n26384 = n26383 ^ n23134;
  assign n26298 = ~n26039 & ~n26068;
  assign n26297 = n26053 & ~n26073;
  assign n26299 = n26298 ^ n26297;
  assign n26379 = n26299 ^ n26101;
  assign n26086 = n26006 & n26082;
  assign n26090 = n26089 ^ n26086;
  assign n26378 = n26090 ^ n26083;
  assign n26380 = n26379 ^ n26378;
  assign n26385 = n26384 ^ n26380;
  assign n26290 = ~n25113 & ~n25142;
  assign n26289 = n25127 & ~n25147;
  assign n26291 = n26290 ^ n26289;
  assign n26374 = n26291 ^ n25175;
  assign n25160 = n25081 & n25156;
  assign n25164 = n25163 ^ n25160;
  assign n26373 = n25164 ^ n25157;
  assign n26375 = n26374 ^ n26373;
  assign n24222 = n24183 & ~n24203;
  assign n24221 = ~n24169 & ~n24198;
  assign n24223 = n24222 ^ n24221;
  assign n26284 = n24238 ^ n24223;
  assign n26283 = n24228 ^ n24218;
  assign n26285 = n26284 ^ n26283;
  assign n26376 = n26375 ^ n26285;
  assign n26246 = n26245 ^ n24232;
  assign n26243 = n26239 ^ n24228;
  assign n26247 = n26246 ^ n26243;
  assign n23270 = ~n23109 & ~n23269;
  assign n26232 = n26231 ^ n23270;
  assign n26233 = n26232 ^ n26218;
  assign n26230 = n26229 ^ n26224;
  assign n26234 = n26233 ^ n26230;
  assign n26372 = n26247 ^ n26234;
  assign n26377 = n26376 ^ n26372;
  assign n26386 = n26385 ^ n26377;
  assign n26436 = n26435 ^ n26386;
  assign n26209 = n26126 & n26183;
  assign n26213 = n26212 ^ n26209;
  assign n26200 = n26199 ^ n26198;
  assign n26207 = n26206 ^ n26200;
  assign n26195 = n26194 ^ n22988;
  assign n26208 = n26207 ^ n26195;
  assign n26214 = n26213 ^ n26208;
  assign n26093 = ~n26027 & ~n26073;
  assign n26095 = n26094 ^ n26093;
  assign n26092 = ~n26037 & n26064;
  assign n26096 = n26095 ^ n26092;
  assign n26103 = n26102 ^ n26096;
  assign n26085 = n26084 ^ n26080;
  assign n26091 = n26090 ^ n26085;
  assign n26104 = n26103 ^ n26091;
  assign n26215 = n26214 ^ n26104;
  assign n25167 = ~n25101 & ~n25147;
  assign n25169 = n25168 ^ n25167;
  assign n25166 = ~n25111 & n25138;
  assign n25170 = n25169 ^ n25166;
  assign n25177 = n25176 ^ n25170;
  assign n25159 = n25158 ^ n25154;
  assign n25165 = n25164 ^ n25159;
  assign n25178 = n25177 ^ n25165;
  assign n24230 = ~n24167 & n24194;
  assign n24233 = n24232 ^ n24230;
  assign n24240 = n24239 ^ n24233;
  assign n24220 = n24219 ^ n24215;
  assign n24229 = n24228 ^ n24220;
  assign n24241 = n24240 ^ n24229;
  assign n25179 = n25178 ^ n24241;
  assign n24224 = n24223 ^ n24220;
  assign n24214 = n24213 ^ n24212;
  assign n24225 = n24224 ^ n24214;
  assign n23284 = n23283 ^ n23282;
  assign n23277 = n23247 & ~n23264;
  assign n23276 = n23226 & ~n23255;
  assign n23278 = n23277 ^ n23276;
  assign n23275 = n23274 ^ n23270;
  assign n23279 = n23278 ^ n23275;
  assign n23285 = n23284 ^ n23279;
  assign n24226 = n24225 ^ n23285;
  assign n25180 = n25179 ^ n24226;
  assign n26216 = n26215 ^ n25180;
  assign n26450 = n26434 ^ n26216;
  assign n26334 = n26303 ^ n26204;
  assign n26332 = n26270 ^ n26212;
  assign n26331 = n26191 ^ n23206;
  assign n26333 = n26332 ^ n26331;
  assign n26335 = n26334 ^ n26333;
  assign n26328 = n26298 ^ n26100;
  assign n26329 = n26328 ^ n26263;
  assign n26327 = n26095 ^ n26089;
  assign n26330 = n26329 ^ n26327;
  assign n26336 = n26335 ^ n26330;
  assign n26325 = n26247 ^ n24241;
  assign n26318 = ~n23162 & ~n23267;
  assign n26319 = n26318 ^ n26218;
  assign n26322 = n26321 ^ n26319;
  assign n26317 = n26229 ^ n23275;
  assign n26323 = n26322 ^ n26317;
  assign n26324 = n26323 ^ n26234;
  assign n26326 = n26325 ^ n26324;
  assign n26337 = n26336 ^ n26326;
  assign n26312 = n26290 ^ n25174;
  assign n26313 = n26312 ^ n26252;
  assign n26311 = n25169 ^ n25163;
  assign n26314 = n26313 ^ n26311;
  assign n26237 = n24235 ^ n24221;
  assign n26241 = n26240 ^ n26237;
  assign n26236 = n24232 ^ n24212;
  assign n26242 = n26241 ^ n26236;
  assign n26315 = n26314 ^ n26242;
  assign n26306 = n26210 ^ n26191;
  assign n26305 = n26304 ^ n26200;
  assign n26307 = n26306 ^ n26305;
  assign n26308 = n26307 ^ n23186;
  assign n26300 = n26299 ^ n26085;
  assign n26296 = n26093 ^ n26089;
  assign n26301 = n26300 ^ n26296;
  assign n26309 = n26308 ^ n26301;
  assign n26292 = n26291 ^ n25159;
  assign n26288 = n25167 ^ n25163;
  assign n26293 = n26292 ^ n26288;
  assign n26294 = n26293 ^ n24225;
  assign n26286 = n26285 ^ n26247;
  assign n26280 = n26279 ^ n23278;
  assign n26277 = n26229 ^ n23272;
  assign n26281 = n26280 ^ n26277;
  assign n26282 = n26281 ^ n26234;
  assign n26287 = n26286 ^ n26282;
  assign n26295 = n26294 ^ n26287;
  assign n26310 = n26309 ^ n26295;
  assign n26316 = n26315 ^ n26310;
  assign n26338 = n26337 ^ n26316;
  assign n26451 = n26450 ^ n26338;
  assign n26462 = n26451 ^ n26436;
  assign n26272 = n26271 ^ n26212;
  assign n26267 = n26194 ^ n23081;
  assign n26273 = n26272 ^ n26267;
  assign n26265 = n26264 ^ n26095;
  assign n26266 = n26265 ^ n26090;
  assign n26274 = n26273 ^ n26266;
  assign n26254 = n26253 ^ n25169;
  assign n26255 = n26254 ^ n25164;
  assign n26259 = n26258 ^ n26255;
  assign n26248 = n26247 ^ n26242;
  assign n26221 = n26220 ^ n23277;
  assign n26226 = n26225 ^ n26221;
  assign n26219 = n26218 ^ n23282;
  assign n26227 = n26226 ^ n26219;
  assign n26235 = n26234 ^ n26227;
  assign n26249 = n26248 ^ n26235;
  assign n26260 = n26259 ^ n26249;
  assign n26275 = n26274 ^ n26260;
  assign n26437 = n26436 ^ n26275;
  assign n26357 = n26356 ^ n26095;
  assign n26354 = n26261 ^ n26090;
  assign n26358 = n26357 ^ n26354;
  assign n26365 = n26364 ^ n26358;
  assign n26350 = n26349 ^ n25169;
  assign n26347 = n26250 ^ n25164;
  assign n26351 = n26350 ^ n26347;
  assign n26352 = n26351 ^ n26247;
  assign n26341 = n26217 ^ n23282;
  assign n26340 = n26339 ^ n26232;
  assign n26342 = n26341 ^ n26340;
  assign n26346 = n26345 ^ n26342;
  assign n26353 = n26352 ^ n26346;
  assign n26366 = n26365 ^ n26353;
  assign n26367 = n26366 ^ n26275;
  assign n26461 = n26437 ^ n26367;
  assign n26466 = n26462 ^ n26461;
  assign n26463 = ~n26461 & n26462;
  assign n26369 = n26366 ^ n26310;
  assign n26458 = ~n26369 & n26451;
  assign n26464 = n26463 ^ n26458;
  assign n26445 = n26411 ^ n26216;
  assign n26446 = n26445 ^ n26338;
  assign n26447 = ~n26367 & n26446;
  assign n26440 = n26366 ^ n26216;
  assign n26368 = n26367 ^ n26338;
  assign n26441 = n26435 ^ n26368;
  assign n26444 = n26440 & ~n26441;
  assign n26448 = n26447 ^ n26444;
  assign n26465 = n26464 ^ n26448;
  assign n26467 = n26466 ^ n26465;
  assign n26442 = n26441 ^ n26440;
  assign n26438 = n26386 & n26437;
  assign n26276 = n26275 ^ n26216;
  assign n26370 = n26369 ^ n26276;
  assign n26371 = ~n26368 & n26370;
  assign n26439 = n26438 ^ n26371;
  assign n26443 = n26442 ^ n26439;
  assign n26449 = n26448 ^ n26443;
  assign n26476 = n26445 ^ n26368;
  assign n26453 = n26450 ^ n26367;
  assign n26454 = ~n26276 & ~n26453;
  assign n26455 = n26454 ^ n26447;
  assign n26477 = n26476 ^ n26455;
  assign n26471 = n26436 ^ n26310;
  assign n26472 = n26471 ^ n26440;
  assign n26473 = n26386 ^ n26368;
  assign n26474 = n26472 & ~n26473;
  assign n26475 = n26474 ^ n26371;
  assign n26478 = n26477 ^ n26475;
  assign n26484 = n26449 & ~n26478;
  assign n26485 = ~n26467 & n26484;
  assign n26482 = n26478 ^ n26449;
  assign n26457 = ~n26310 & n26436;
  assign n26459 = n26458 ^ n26457;
  assign n26452 = n26451 ^ n26369;
  assign n26456 = n26455 ^ n26452;
  assign n26460 = n26459 ^ n26456;
  assign n26479 = ~n26460 & ~n26478;
  assign n26483 = n26482 ^ n26479;
  assign n26486 = n26485 ^ n26483;
  assign n26509 = n26436 & n26486;
  assign n26468 = n26467 ^ n26460;
  assign n26480 = n26479 ^ n26468;
  assign n26469 = ~n26460 & n26468;
  assign n26470 = ~n26449 & n26469;
  assign n26481 = n26480 ^ n26470;
  assign n26508 = n26472 & n26481;
  assign n26510 = n26509 ^ n26508;
  assign n26491 = n26479 ^ n26449;
  assign n26492 = n26468 & ~n26491;
  assign n26493 = n26492 ^ n26467;
  assign n26488 = n26479 ^ n26467;
  assign n26489 = n26482 & ~n26488;
  assign n26490 = n26489 ^ n26449;
  assign n26494 = n26493 ^ n26490;
  assign n26506 = n26446 & n26494;
  assign n26487 = n26486 ^ n26481;
  assign n26495 = n26494 ^ n26487;
  assign n26505 = ~n26453 & n26495;
  assign n26507 = n26506 ^ n26505;
  assign n26511 = n26510 ^ n26507;
  assign n26502 = n26493 ^ n26481;
  assign n26503 = n26370 & ~n26502;
  assign n26499 = n26490 ^ n26486;
  assign n26500 = n26451 & ~n26499;
  assign n26497 = ~n26367 & n26494;
  assign n26496 = ~n26276 & n26495;
  assign n26498 = n26497 ^ n26496;
  assign n26501 = n26500 ^ n26498;
  assign n26504 = n26503 ^ n26501;
  assign n26512 = n26511 ^ n26504;
  assign n26764 = n26763 ^ n26512;
  assign n26777 = n26759 ^ n26748;
  assign n26774 = ~n26692 & ~n26752;
  assign n26772 = n26721 & ~n26744;
  assign n26773 = n26772 ^ n26753;
  assign n26775 = n26774 ^ n26773;
  assign n26776 = n26775 ^ n26757;
  assign n26778 = n26777 ^ n26776;
  assign n26779 = n26778 ^ n26409;
  assign n26770 = n26508 ^ n26498;
  assign n26767 = ~n26368 & ~n26502;
  assign n26765 = ~n26473 & n26481;
  assign n26766 = n26765 ^ n26503;
  assign n26768 = n26767 ^ n26766;
  assign n26769 = n26768 ^ n26507;
  assign n26771 = n26770 ^ n26769;
  assign n26780 = n26779 ^ n26771;
  assign n26803 = n26755 ^ n26736;
  assign n26800 = n26691 & n26745;
  assign n26801 = n26800 ^ n26432;
  assign n26797 = ~n26688 & n26749;
  assign n26796 = ~n26693 & n26745;
  assign n26798 = n26797 ^ n26796;
  assign n26794 = ~n26657 & ~n26734;
  assign n26792 = ~n26654 & n26730;
  assign n26793 = n26792 ^ n26774;
  assign n26795 = n26794 ^ n26793;
  assign n26799 = n26798 ^ n26795;
  assign n26802 = n26801 ^ n26799;
  assign n26804 = n26803 ^ n26802;
  assign n26805 = n26804 ^ n26497;
  assign n26789 = n26440 & n26487;
  assign n26787 = ~n26369 & ~n26499;
  assign n26786 = ~n26441 & n26487;
  assign n26788 = n26787 ^ n26786;
  assign n26790 = n26789 ^ n26788;
  assign n26783 = ~n26461 & ~n26490;
  assign n26781 = n26386 & ~n26493;
  assign n26782 = n26781 ^ n26767;
  assign n26784 = n26783 ^ n26782;
  assign n26785 = n26784 ^ n26506;
  assign n26791 = n26790 ^ n26785;
  assign n26806 = n26805 ^ n26791;
  assign n26809 = n26775 ^ n26760;
  assign n26808 = n26751 ^ n26273;
  assign n26810 = n26809 ^ n26808;
  assign n26811 = n26810 ^ n26768;
  assign n26807 = n26510 ^ n26501;
  assign n26812 = n26811 ^ n26807;
  assign n26820 = ~n26686 & ~n26734;
  assign n26821 = n26820 ^ n26792;
  assign n26818 = n26773 ^ n26760;
  assign n26817 = n26748 ^ n26335;
  assign n26819 = n26818 ^ n26817;
  assign n26822 = n26821 ^ n26819;
  assign n26816 = n26462 & ~n26490;
  assign n26823 = n26822 ^ n26816;
  assign n26814 = n26781 ^ n26766;
  assign n26813 = n26510 ^ n26498;
  assign n26815 = n26814 ^ n26813;
  assign n26824 = n26823 ^ n26815;
  assign n26835 = n26437 & ~n26493;
  assign n26836 = n26835 ^ n26784;
  assign n26833 = n26788 ^ n26505;
  assign n26829 = ~n26656 & n26730;
  assign n26830 = n26829 ^ n26760;
  assign n26826 = n26798 ^ n26756;
  assign n26827 = n26826 ^ n26795;
  assign n26825 = n26751 ^ n26214;
  assign n26828 = n26827 ^ n26825;
  assign n26831 = n26830 ^ n26828;
  assign n26832 = n26831 ^ n26807;
  assign n26834 = n26833 ^ n26832;
  assign n26837 = n26836 ^ n26834;
  assign n26844 = n26719 & ~n26740;
  assign n26845 = n26844 ^ n26820;
  assign n26846 = n26845 ^ n26826;
  assign n26843 = n26758 ^ n26748;
  assign n26847 = n26846 ^ n26843;
  assign n26848 = n26847 ^ n26308;
  assign n26841 = n26509 ^ n26498;
  assign n26838 = n26471 & n26486;
  assign n26839 = n26838 ^ n26816;
  assign n26840 = n26839 ^ n26833;
  assign n26842 = n26841 ^ n26840;
  assign n26849 = n26848 ^ n26842;
  assign n26854 = n26845 ^ n26793;
  assign n26853 = n26797 ^ n26751;
  assign n26855 = n26854 ^ n26853;
  assign n26856 = n26855 ^ n26384;
  assign n26851 = n26839 ^ n26782;
  assign n26850 = n26787 ^ n26501;
  assign n26852 = n26851 ^ n26850;
  assign n26857 = n26856 ^ n26852;
  assign n27657 = n25934 ^ n25751;
  assign n27664 = n27657 ^ n26024;
  assign n27676 = n27664 ^ n25970;
  assign n27660 = n25934 ^ n25829;
  assign n27655 = n25904 ^ n25877;
  assign n27652 = n25998 ^ n25970;
  assign n27656 = n27655 ^ n27652;
  assign n27683 = n27660 ^ n27656;
  assign n27668 = n25877 ^ n25829;
  assign n27651 = n25829 ^ n25751;
  assign n27680 = n27655 ^ n27651;
  assign n27681 = n27668 & n27680;
  assign n27661 = n27660 ^ n27652;
  assign n27662 = n27655 & n27661;
  assign n27682 = n27681 ^ n27662;
  assign n27684 = n27683 ^ n27682;
  assign n27675 = n27656 ^ n26024;
  assign n27654 = n25904 ^ n25829;
  assign n27677 = n27676 ^ n27654;
  assign n27678 = n27675 & n27677;
  assign n27667 = n25970 ^ n25904;
  assign n27669 = n27668 ^ n27667;
  assign n27670 = n27656 & n27669;
  assign n27679 = n27678 ^ n27670;
  assign n27685 = n27684 ^ n27679;
  assign n27697 = ~n25970 & n27664;
  assign n27653 = n27652 ^ n27651;
  assign n27690 = n27653 & n27667;
  assign n27698 = n27697 ^ n27690;
  assign n27695 = n27667 ^ n27653;
  assign n27696 = n27695 ^ n27682;
  assign n27699 = n27698 ^ n27696;
  assign n27700 = n27685 & n27699;
  assign n27658 = n27657 ^ n27656;
  assign n27672 = n27658 ^ n27654;
  assign n27665 = n27664 ^ n25877;
  assign n27666 = n26024 & n27665;
  assign n27671 = n27670 ^ n27666;
  assign n27673 = n27672 ^ n27671;
  assign n27659 = n27654 & n27658;
  assign n27663 = n27662 ^ n27659;
  assign n27674 = n27673 ^ n27663;
  assign n27686 = n27685 ^ n27674;
  assign n27706 = n27700 ^ n27686;
  assign n27688 = n27664 ^ n27653;
  assign n27687 = n27665 ^ n27655;
  assign n27693 = n27688 ^ n27687;
  assign n27689 = n27687 & n27688;
  assign n27691 = n27690 ^ n27689;
  assign n27692 = n27691 ^ n27663;
  assign n27694 = n27693 ^ n27692;
  assign n27704 = ~n27674 & n27685;
  assign n27705 = n27694 & n27704;
  assign n27707 = n27706 ^ n27705;
  assign n27787 = n27676 & n27707;
  assign n27701 = n27700 ^ n27694;
  assign n27702 = n27686 & n27701;
  assign n27703 = n27702 ^ n27674;
  assign n27781 = n27688 & n27703;
  assign n27788 = n27787 ^ n27781;
  assign n27712 = n27699 ^ n27694;
  assign n27716 = n27700 ^ n27674;
  assign n27717 = n27712 & n27716;
  assign n27718 = n27717 ^ n27694;
  assign n27753 = n26024 & n27718;
  assign n27713 = n27712 ^ n27700;
  assign n27710 = n27674 & n27699;
  assign n27711 = ~n27694 & n27710;
  assign n27714 = n27713 ^ n27711;
  assign n27729 = n27718 ^ n27714;
  assign n27733 = n27656 & n27729;
  assign n27754 = n27753 ^ n27733;
  assign n27807 = n27788 ^ n27754;
  assign n27708 = n27707 ^ n27703;
  assign n27757 = n27667 & n27708;
  assign n27719 = n27718 ^ n27703;
  assign n27722 = n27655 & n27719;
  assign n27715 = n27714 ^ n27707;
  assign n27720 = n27719 ^ n27715;
  assign n27721 = n27668 & n27720;
  assign n27723 = n27722 ^ n27721;
  assign n27709 = n27653 & n27708;
  assign n27724 = n27723 ^ n27709;
  assign n27806 = n27757 ^ n27724;
  assign n27808 = n27807 ^ n27806;
  assign n27809 = n27808 ^ n25097;
  assign n27810 = n27809 ^ n25098;
  assign n27811 = n27810 ^ n25099;
  assign n27812 = n27811 ^ n26533;
  assign n27726 = n27677 & n27714;
  assign n27799 = n27726 ^ n27723;
  assign n27742 = n27680 & n27720;
  assign n27741 = n27661 & n27719;
  assign n27743 = n27742 ^ n27741;
  assign n27731 = n27675 & n27714;
  assign n27730 = n27669 & n27729;
  assign n27732 = n27731 ^ n27730;
  assign n27734 = n27733 ^ n27732;
  assign n27798 = n27743 ^ n27734;
  assign n27800 = n27799 ^ n27798;
  assign n27801 = n27800 ^ n25009;
  assign n27802 = n27801 ^ n25010;
  assign n27803 = n27802 ^ n25011;
  assign n27804 = n27803 ^ n26525;
  assign n27772 = n27741 ^ n27722;
  assign n27769 = n27654 & n27715;
  assign n27770 = n27769 ^ n24830;
  assign n27756 = n27658 & n27715;
  assign n27758 = n27757 ^ n27756;
  assign n27752 = n27687 & n27703;
  assign n27755 = n27754 ^ n27752;
  assign n27768 = n27758 ^ n27755;
  assign n27771 = n27770 ^ n27768;
  assign n27773 = n27772 ^ n27771;
  assign n27774 = n27773 ^ n24831;
  assign n27775 = n27774 ^ n24832;
  assign n27776 = n27775 ^ n26514;
  assign n27805 = n27804 ^ n27776;
  assign n27813 = n27812 ^ n27805;
  assign n27727 = n27664 & n27707;
  assign n27790 = n27727 ^ n27723;
  assign n27759 = n27758 ^ n27742;
  assign n27789 = n27788 ^ n27759;
  assign n27791 = n27790 ^ n27789;
  assign n27792 = n27791 ^ n25044;
  assign n27793 = n27792 ^ n25045;
  assign n27794 = n27793 ^ n25046;
  assign n27795 = n27794 ^ n26517;
  assign n27849 = n27813 ^ n27795;
  assign n27762 = n27665 & n27718;
  assign n27728 = n27727 ^ n27726;
  assign n27763 = n27762 ^ n27728;
  assign n27760 = n27759 ^ n27755;
  assign n27751 = n27724 ^ n24907;
  assign n27761 = n27760 ^ n27751;
  assign n27764 = n27763 ^ n27761;
  assign n27765 = n27764 ^ n24908;
  assign n27766 = n27765 ^ n24909;
  assign n27767 = n27766 ^ n26513;
  assign n27744 = n27743 ^ n27728;
  assign n27740 = n27730 ^ n27724;
  assign n27745 = n27744 ^ n27740;
  assign n27746 = n27745 ^ n24980;
  assign n27747 = n27746 ^ n24981;
  assign n27748 = n27747 ^ n24982;
  assign n27749 = n27748 ^ n26520;
  assign n27821 = n27767 ^ n27749;
  assign n27850 = n27849 ^ n27821;
  assign n27838 = n27795 & ~n27813;
  assign n27782 = n27781 ^ n27753;
  assign n27779 = n27732 ^ n27728;
  assign n27778 = n27723 ^ n25053;
  assign n27780 = n27779 ^ n27778;
  assign n27783 = n27782 ^ n27780;
  assign n27784 = n27783 ^ n25054;
  assign n27785 = n27784 ^ n25055;
  assign n27786 = n27785 ^ n26516;
  assign n27796 = n27795 ^ n27786;
  assign n27777 = n27776 ^ n27767;
  assign n27797 = n27796 ^ n27777;
  assign n27818 = n27795 ^ n27749;
  assign n27819 = n27797 & ~n27818;
  assign n27839 = n27838 ^ n27819;
  assign n27836 = n27818 ^ n27797;
  assign n27735 = n27734 ^ n27728;
  assign n27725 = n27724 ^ n24954;
  assign n27736 = n27735 ^ n27725;
  assign n27737 = n27736 ^ n24955;
  assign n27738 = n27737 ^ n24956;
  assign n27739 = n27738 ^ n26522;
  assign n27832 = n27767 ^ n27739;
  assign n27750 = n27749 ^ n27739;
  assign n27833 = n27777 ^ n27750;
  assign n27834 = n27832 & ~n27833;
  assign n27825 = n27804 ^ n27767;
  assign n27826 = n27825 ^ n27796;
  assign n27827 = n27750 & n27826;
  assign n27835 = n27834 ^ n27827;
  assign n27837 = n27836 ^ n27835;
  assign n27840 = n27839 ^ n27837;
  assign n27822 = n27796 ^ n27750;
  assign n27854 = n27825 ^ n27822;
  assign n27855 = n27854 ^ n27835;
  assign n27851 = n27822 ^ n27812;
  assign n27852 = n27850 & n27851;
  assign n27843 = n27832 ^ n27818;
  assign n27844 = ~n27822 & ~n27843;
  assign n27853 = n27852 ^ n27844;
  assign n27856 = n27855 ^ n27853;
  assign n27857 = ~n27840 & n27856;
  assign n27815 = n27813 ^ n27739;
  assign n27816 = n27815 ^ n27750;
  assign n27814 = n27813 ^ n27797;
  assign n27830 = n27816 ^ n27814;
  assign n27823 = n27822 ^ n27805;
  assign n27824 = n27821 & ~n27823;
  assign n27828 = n27827 ^ n27824;
  assign n27817 = ~n27814 & ~n27816;
  assign n27820 = n27819 ^ n27817;
  assign n27829 = n27828 ^ n27820;
  assign n27831 = n27830 ^ n27829;
  assign n27841 = n27840 ^ n27831;
  assign n27873 = n27857 ^ n27841;
  assign n27846 = n27823 ^ n27821;
  assign n27842 = ~n27812 & ~n27815;
  assign n27845 = n27844 ^ n27842;
  assign n27847 = n27846 ^ n27845;
  assign n27848 = n27847 ^ n27828;
  assign n27871 = ~n27840 & ~n27848;
  assign n27872 = ~n27831 & n27871;
  assign n27874 = n27873 ^ n27872;
  assign n27889 = n27850 & ~n27874;
  assign n27868 = n27848 & n27856;
  assign n27869 = n27831 & n27868;
  assign n27861 = n27856 ^ n27848;
  assign n27867 = n27861 ^ n27857;
  assign n27870 = n27869 ^ n27867;
  assign n27888 = ~n27813 & ~n27870;
  assign n27890 = n27889 ^ n27888;
  assign n27875 = n27874 ^ n27870;
  assign n27862 = n27857 ^ n27831;
  assign n27863 = ~n27861 & n27862;
  assign n27864 = n27863 ^ n27848;
  assign n27858 = n27857 ^ n27848;
  assign n27859 = ~n27841 & ~n27858;
  assign n27860 = n27859 ^ n27831;
  assign n27865 = n27864 ^ n27860;
  assign n27876 = n27875 ^ n27865;
  assign n27886 = ~n27833 & ~n27876;
  assign n27885 = n27826 & ~n27865;
  assign n27887 = n27886 ^ n27885;
  assign n27891 = n27890 ^ n27887;
  assign n27882 = n27874 ^ n27860;
  assign n27883 = ~n27843 & ~n27882;
  assign n27879 = n27870 ^ n27864;
  assign n27880 = n27797 & n27879;
  assign n27877 = n27832 & ~n27876;
  assign n27866 = n27750 & ~n27865;
  assign n27878 = n27877 ^ n27866;
  assign n27881 = n27880 ^ n27878;
  assign n27884 = n27883 ^ n27881;
  assign n27892 = n27891 ^ n27884;
  assign n27893 = n27892 ^ n26616;
  assign n27289 = n23727 ^ n22988;
  assign n27290 = n27289 ^ n23964;
  assign n27287 = n24127 ^ n23935;
  assign n27286 = n24079 ^ n23949;
  assign n27288 = n27287 ^ n27286;
  assign n27291 = n27290 ^ n27288;
  assign n27267 = n23741 ^ n23036;
  assign n27268 = n27267 ^ n23997;
  assign n27265 = n24008 ^ n23820;
  assign n27266 = n27265 ^ n24057;
  assign n27269 = n27268 ^ n27266;
  assign n27292 = n27291 ^ n27269;
  assign n27282 = n23712 ^ n23206;
  assign n27283 = n27282 ^ n24110;
  assign n27280 = n24024 ^ n23923;
  assign n27281 = n27280 ^ n24128;
  assign n27284 = n27283 ^ n27281;
  assign n27278 = n23552 ^ n23417;
  assign n27275 = n23705 ^ n23186;
  assign n27276 = n27275 ^ n24096;
  assign n27272 = n24144 ^ n24024;
  assign n27273 = n27272 ^ n24083;
  assign n27274 = n27273 ^ n23950;
  assign n27277 = n27276 ^ n27274;
  assign n27279 = n27278 ^ n27277;
  assign n27285 = n27284 ^ n27279;
  assign n27293 = n27292 ^ n27285;
  assign n27262 = n23732 ^ n23157;
  assign n27263 = n27262 ^ n24060;
  assign n27260 = n24031 ^ n24027;
  assign n27259 = n24056 ^ n23991;
  assign n27261 = n27260 ^ n27259;
  assign n27264 = n27263 ^ n27261;
  assign n27270 = n27269 ^ n27264;
  assign n27256 = n23720 ^ n23134;
  assign n27257 = n27256 ^ n24149;
  assign n27254 = n24087 ^ n24082;
  assign n27253 = n24024 ^ n23409;
  assign n27255 = n27254 ^ n27253;
  assign n27258 = n27257 ^ n27255;
  assign n27271 = n27270 ^ n27258;
  assign n27294 = n27293 ^ n27271;
  assign n27305 = n23692 ^ n23105;
  assign n27306 = n27305 ^ n24037;
  assign n27303 = n23561 ^ n23409;
  assign n27302 = n24065 ^ n24027;
  assign n27304 = n27303 ^ n27302;
  assign n27307 = n27306 ^ n27304;
  assign n27298 = n23698 ^ n23081;
  assign n27299 = n27298 ^ n23685;
  assign n27295 = n24122 ^ n24024;
  assign n27296 = n27295 ^ n23418;
  assign n27297 = n27296 ^ n24009;
  assign n27300 = n27299 ^ n27297;
  assign n27308 = n27307 ^ n27300;
  assign n27315 = n27308 ^ n27285;
  assign n27316 = n27315 ^ n27270;
  assign n27314 = n27307 ^ n27291;
  assign n27341 = n27316 ^ n27314;
  assign n27301 = n27300 ^ n27271;
  assign n27339 = ~n27258 & n27301;
  assign n27325 = n27300 ^ n27291;
  assign n27311 = n27307 ^ n27277;
  assign n27326 = n27325 ^ n27311;
  assign n27327 = n27315 & ~n27326;
  assign n27340 = n27339 ^ n27327;
  assign n27342 = n27341 ^ n27340;
  assign n27318 = n27291 ^ n27264;
  assign n27319 = n27318 ^ n27285;
  assign n27320 = ~n27308 & n27319;
  assign n27317 = ~n27314 & ~n27316;
  assign n27321 = n27320 ^ n27317;
  assign n27343 = n27342 ^ n27321;
  assign n27336 = n27318 ^ n27315;
  assign n27333 = n27308 ^ n27292;
  assign n27334 = n27325 & ~n27333;
  assign n27335 = n27334 ^ n27320;
  assign n27337 = n27336 ^ n27335;
  assign n27328 = n27277 ^ n27271;
  assign n27329 = n27328 ^ n27314;
  assign n27330 = n27315 ^ n27258;
  assign n27331 = ~n27329 & ~n27330;
  assign n27332 = n27331 ^ n27327;
  assign n27338 = n27337 ^ n27332;
  assign n27352 = n27343 ^ n27338;
  assign n27348 = n27271 & ~n27277;
  assign n27312 = ~n27293 & ~n27311;
  assign n27349 = n27348 ^ n27312;
  assign n27346 = n27311 ^ n27293;
  assign n27347 = n27346 ^ n27335;
  assign n27350 = n27349 ^ n27347;
  assign n27351 = ~n27338 & n27350;
  assign n27309 = n27308 ^ n27301;
  assign n27323 = n27309 ^ n27294;
  assign n27310 = ~n27294 & ~n27309;
  assign n27313 = n27312 ^ n27310;
  assign n27322 = n27321 ^ n27313;
  assign n27324 = n27323 ^ n27322;
  assign n27374 = n27351 ^ n27324;
  assign n27375 = ~n27352 & n27374;
  assign n27376 = n27375 ^ n27343;
  assign n27484 = ~n27294 & n27376;
  assign n27353 = n27352 ^ n27351;
  assign n27344 = ~n27338 & ~n27343;
  assign n27345 = n27324 & n27344;
  assign n27354 = n27353 ^ n27345;
  assign n27483 = n27328 & ~n27354;
  assign n27485 = n27484 ^ n27483;
  assign n27358 = n27350 ^ n27324;
  assign n27363 = n27351 ^ n27343;
  assign n27364 = n27358 & n27363;
  assign n27365 = n27364 ^ n27324;
  assign n27440 = ~n27258 & n27365;
  assign n27359 = n27358 ^ n27351;
  assign n27356 = n27343 & n27350;
  assign n27357 = ~n27324 & n27356;
  assign n27360 = n27359 ^ n27357;
  assign n27366 = n27365 ^ n27360;
  assign n27370 = n27315 & n27366;
  assign n27441 = n27440 ^ n27370;
  assign n27573 = n27485 ^ n27441;
  assign n27382 = n27376 ^ n27354;
  assign n27432 = ~n27311 & ~n27382;
  assign n27383 = ~n27293 & ~n27382;
  assign n27377 = n27376 ^ n27365;
  assign n27380 = ~n27308 & n27377;
  assign n27373 = n27360 ^ n27354;
  assign n27378 = n27377 ^ n27373;
  assign n27379 = n27325 & ~n27378;
  assign n27381 = n27380 ^ n27379;
  assign n27384 = n27383 ^ n27381;
  assign n27572 = n27432 ^ n27384;
  assign n27574 = n27573 ^ n27572;
  assign n27159 = n25035 ^ n24884;
  assign n27160 = n27159 ^ n24891;
  assign n27161 = n27160 ^ n25063;
  assign n27162 = n27161 ^ n24849;
  assign n27163 = n27162 ^ n26107;
  assign n27139 = n24945 ^ n24611;
  assign n27138 = n25004 ^ n24367;
  assign n27140 = n27139 ^ n27138;
  assign n27141 = n27140 ^ n26110;
  assign n27164 = n27163 ^ n27141;
  assign n27127 = n26127 ^ n24920;
  assign n27125 = n24973 ^ n24926;
  assign n27124 = n24994 ^ n24962;
  assign n27126 = n27125 ^ n27124;
  assign n27128 = n27127 ^ n27126;
  assign n27120 = n25073 ^ n24966;
  assign n27119 = n24932 ^ n24731;
  assign n27121 = n27120 ^ n27119;
  assign n27122 = n27121 ^ n24939;
  assign n27123 = n27122 ^ n26105;
  assign n27129 = n27128 ^ n27123;
  assign n27182 = n27164 ^ n27129;
  assign n27134 = n25003 ^ n24487;
  assign n27135 = n27134 ^ n24974;
  assign n27136 = n27135 ^ n24991;
  assign n27137 = n27136 ^ n26119;
  assign n27142 = n27141 ^ n27137;
  assign n27132 = n26122 ^ n25021;
  assign n27130 = n25092 ^ n24966;
  assign n27131 = n27130 ^ n25018;
  assign n27133 = n27132 ^ n27131;
  assign n27143 = n27142 ^ n27133;
  assign n27151 = n26115 ^ n24873;
  assign n27149 = n25018 ^ n24884;
  assign n27147 = n25088 ^ n24966;
  assign n27148 = n27147 ^ n25029;
  assign n27150 = n27149 ^ n27148;
  assign n27152 = n27151 ^ n27150;
  assign n27188 = ~n27143 & n27152;
  assign n27156 = n25064 ^ n24931;
  assign n27154 = n24966 ^ n24864;
  assign n27155 = n27154 ^ n25069;
  assign n27157 = n27156 ^ n27155;
  assign n27146 = n26113 ^ n24916;
  assign n27153 = n27152 ^ n27146;
  assign n27158 = n27157 ^ n27153;
  assign n27165 = n27164 ^ n27158;
  assign n27168 = n27152 ^ n27128;
  assign n27169 = n27165 & ~n27168;
  assign n27189 = n27188 ^ n27169;
  assign n27186 = n27168 ^ n27165;
  assign n27183 = n27163 ^ n27123;
  assign n27184 = ~n27182 & n27183;
  assign n27175 = n27163 ^ n27137;
  assign n27176 = n27175 ^ n27158;
  assign n27177 = n27129 & n27176;
  assign n27185 = n27184 ^ n27177;
  assign n27187 = n27186 ^ n27185;
  assign n27190 = n27189 ^ n27187;
  assign n27172 = n27158 ^ n27129;
  assign n27204 = n27175 ^ n27172;
  assign n27205 = n27204 ^ n27185;
  assign n27199 = n27152 ^ n27143;
  assign n27171 = n27163 ^ n27128;
  assign n27200 = n27199 ^ n27171;
  assign n27201 = n27172 ^ n27133;
  assign n27202 = n27200 & n27201;
  assign n27193 = n27183 ^ n27168;
  assign n27194 = ~n27172 & ~n27193;
  assign n27203 = n27202 ^ n27194;
  assign n27206 = n27205 ^ n27203;
  assign n27207 = ~n27190 & n27206;
  assign n27166 = n27165 ^ n27143;
  assign n27144 = n27143 ^ n27123;
  assign n27145 = n27144 ^ n27129;
  assign n27180 = n27166 ^ n27145;
  assign n27173 = n27172 ^ n27142;
  assign n27174 = n27171 & ~n27173;
  assign n27178 = n27177 ^ n27174;
  assign n27167 = ~n27145 & ~n27166;
  assign n27170 = n27169 ^ n27167;
  assign n27179 = n27178 ^ n27170;
  assign n27181 = n27180 ^ n27179;
  assign n27191 = n27190 ^ n27181;
  assign n27223 = n27207 ^ n27191;
  assign n27196 = n27173 ^ n27171;
  assign n27192 = ~n27133 & ~n27144;
  assign n27195 = n27194 ^ n27192;
  assign n27197 = n27196 ^ n27195;
  assign n27198 = n27197 ^ n27178;
  assign n27221 = ~n27190 & ~n27198;
  assign n27222 = ~n27181 & n27221;
  assign n27224 = n27223 ^ n27222;
  assign n27218 = n27198 & n27206;
  assign n27219 = n27181 & n27218;
  assign n27211 = n27206 ^ n27198;
  assign n27217 = n27211 ^ n27207;
  assign n27220 = n27219 ^ n27217;
  assign n27225 = n27224 ^ n27220;
  assign n27212 = n27207 ^ n27181;
  assign n27213 = ~n27211 & n27212;
  assign n27214 = n27213 ^ n27198;
  assign n27208 = n27207 ^ n27198;
  assign n27209 = ~n27191 & ~n27208;
  assign n27210 = n27209 ^ n27181;
  assign n27215 = n27214 ^ n27210;
  assign n27226 = n27225 ^ n27215;
  assign n27247 = ~n27182 & ~n27226;
  assign n27246 = n27176 & ~n27215;
  assign n27248 = n27247 ^ n27246;
  assign n27230 = n27200 & ~n27224;
  assign n27229 = ~n27143 & ~n27220;
  assign n27231 = n27230 ^ n27229;
  assign n27249 = n27248 ^ n27231;
  assign n27242 = n27220 ^ n27214;
  assign n27243 = n27165 & n27242;
  assign n27227 = n27183 & ~n27226;
  assign n27216 = n27129 & ~n27215;
  assign n27228 = n27227 ^ n27216;
  assign n27244 = n27243 ^ n27228;
  assign n27237 = n27224 ^ n27210;
  assign n27238 = ~n27193 & ~n27237;
  assign n27245 = n27244 ^ n27238;
  assign n27250 = n27249 ^ n27245;
  assign n27575 = n27574 ^ n27250;
  assign n27003 = n25960 ^ n25883;
  assign n27004 = n27003 ^ n26015;
  assign n27005 = n27004 ^ n25940;
  assign n27006 = n27005 ^ n26533;
  assign n26994 = n26517 ^ n25810;
  assign n26992 = n25954 ^ n25761;
  assign n26990 = n26012 ^ n25883;
  assign n26991 = n26990 ^ n25960;
  assign n26993 = n26992 ^ n26991;
  assign n26995 = n26994 ^ n26993;
  assign n27022 = n26514 ^ n25927;
  assign n27020 = n25531 ^ n25411;
  assign n27019 = n25848 ^ n25663;
  assign n27021 = n27020 ^ n27019;
  assign n27023 = n27022 ^ n27021;
  assign n27017 = n26525 ^ n25896;
  assign n27015 = n25916 ^ n25891;
  assign n27014 = n25927 ^ n25295;
  assign n27016 = n27015 ^ n27014;
  assign n27018 = n27017 ^ n27016;
  assign n27024 = n27023 ^ n27018;
  assign n27031 = n27024 ^ n27006;
  assign n27050 = n26995 & ~n27031;
  assign n27011 = n26513 ^ n25989;
  assign n27009 = n25948 ^ n25810;
  assign n27008 = n25797 ^ n25766;
  assign n27010 = n27009 ^ n27008;
  assign n27012 = n27011 ^ n27010;
  assign n27034 = n27023 ^ n27012;
  assign n26999 = n25980 ^ n25836;
  assign n26997 = n25883 ^ n25782;
  assign n26998 = n26997 ^ n25990;
  assign n27000 = n26999 ^ n26998;
  assign n26989 = n26516 ^ n25866;
  assign n26996 = n26995 ^ n26989;
  assign n27001 = n27000 ^ n26996;
  assign n27035 = n27034 ^ n27001;
  assign n26986 = n26520 ^ n25861;
  assign n26984 = n25913 ^ n25896;
  assign n26983 = n25887 ^ n25840;
  assign n26985 = n26984 ^ n26983;
  assign n26987 = n26986 ^ n26985;
  assign n27038 = n26995 ^ n26987;
  assign n27039 = n27035 & ~n27038;
  assign n27051 = n27050 ^ n27039;
  assign n27048 = n27038 ^ n27035;
  assign n26981 = n26522 ^ n25663;
  assign n26979 = n25854 ^ n25545;
  assign n26977 = n25976 ^ n25883;
  assign n26978 = n26977 ^ n25867;
  assign n26980 = n26979 ^ n26978;
  assign n26982 = n26981 ^ n26980;
  assign n27044 = n27012 ^ n26982;
  assign n26988 = n26987 ^ n26982;
  assign n27045 = n27034 ^ n26988;
  assign n27046 = n27044 & ~n27045;
  assign n27027 = n27018 ^ n27012;
  assign n27028 = n27027 ^ n27001;
  assign n27029 = n26988 & n27028;
  assign n27047 = n27046 ^ n27029;
  assign n27049 = n27048 ^ n27047;
  assign n27052 = n27051 ^ n27049;
  assign n27036 = n27035 ^ n27031;
  assign n27032 = n27031 ^ n26982;
  assign n27033 = n27032 ^ n26988;
  assign n27042 = n27036 ^ n27033;
  assign n27037 = ~n27033 & ~n27036;
  assign n27040 = n27039 ^ n27037;
  assign n27013 = n27012 ^ n26987;
  assign n27002 = n27001 ^ n26988;
  assign n27025 = n27024 ^ n27002;
  assign n27026 = n27013 & ~n27025;
  assign n27030 = n27029 ^ n27026;
  assign n27041 = n27040 ^ n27030;
  assign n27043 = n27042 ^ n27041;
  assign n27070 = n27052 ^ n27043;
  assign n27066 = n27027 ^ n27002;
  assign n27067 = n27066 ^ n27047;
  assign n27007 = n27006 ^ n27002;
  assign n27062 = n27031 ^ n26995;
  assign n27063 = n27062 ^ n27013;
  assign n27064 = n27007 & n27063;
  assign n27054 = n27044 ^ n27038;
  assign n27055 = ~n27002 & ~n27054;
  assign n27065 = n27064 ^ n27055;
  assign n27068 = n27067 ^ n27065;
  assign n27069 = ~n27052 & n27068;
  assign n27057 = n27025 ^ n27013;
  assign n27053 = ~n27006 & ~n27032;
  assign n27056 = n27055 ^ n27053;
  assign n27058 = n27057 ^ n27056;
  assign n27059 = n27058 ^ n27030;
  assign n27074 = n27069 ^ n27059;
  assign n27075 = ~n27070 & ~n27074;
  assign n27076 = n27075 ^ n27043;
  assign n27107 = ~n27006 & n27076;
  assign n27071 = n27070 ^ n27069;
  assign n27060 = ~n27052 & ~n27059;
  assign n27061 = ~n27043 & n27060;
  assign n27072 = n27071 ^ n27061;
  assign n27077 = n27076 ^ n27072;
  assign n27080 = ~n27002 & ~n27077;
  assign n27426 = n27107 ^ n27080;
  assign n27084 = n27059 & n27068;
  assign n27085 = n27043 & n27084;
  assign n27082 = n27068 ^ n27059;
  assign n27083 = n27082 ^ n27069;
  assign n27086 = n27085 ^ n27083;
  assign n27407 = n27062 & ~n27086;
  assign n27091 = n27069 ^ n27043;
  assign n27092 = ~n27082 & n27091;
  assign n27093 = n27092 ^ n27059;
  assign n27106 = ~n27036 & ~n27093;
  assign n27408 = n27407 ^ n27106;
  assign n27474 = n27426 ^ n27408;
  assign n27100 = n27093 ^ n27086;
  assign n27404 = ~n27038 & n27100;
  assign n27101 = n27035 & n27100;
  assign n27096 = n27086 ^ n27072;
  assign n27094 = n27093 ^ n27076;
  assign n27097 = n27096 ^ n27094;
  assign n27098 = n27044 & ~n27097;
  assign n27095 = n26988 & ~n27094;
  assign n27099 = n27098 ^ n27095;
  assign n27102 = n27101 ^ n27099;
  assign n27473 = n27404 ^ n27102;
  assign n27475 = n27474 ^ n27473;
  assign n27113 = ~n27045 & ~n27097;
  assign n27112 = n27028 & ~n27094;
  assign n27114 = n27113 ^ n27112;
  assign n27088 = n27063 & ~n27072;
  assign n27087 = ~n27031 & ~n27086;
  assign n27089 = n27088 ^ n27087;
  assign n27115 = n27114 ^ n27089;
  assign n27078 = ~n27054 & ~n27077;
  assign n27111 = n27102 ^ n27078;
  assign n27116 = n27115 ^ n27111;
  assign n27476 = n27475 ^ n27116;
  assign n27576 = n27575 ^ n27476;
  assign n26897 = n25826 ^ n23182;
  assign n26895 = n23195 ^ n21946;
  assign n26896 = n26895 ^ n21042;
  assign n26898 = n26897 ^ n26896;
  assign n26864 = n25748 ^ n23074;
  assign n26862 = n23144 ^ n23015;
  assign n26863 = n26862 ^ n23003;
  assign n26865 = n26864 ^ n26863;
  assign n26907 = n26898 ^ n26865;
  assign n26889 = n23196 ^ n23053;
  assign n26887 = n23100 ^ n22878;
  assign n26888 = n26887 ^ n25995;
  assign n26890 = n26889 ^ n26888;
  assign n26883 = n23127 ^ n23100;
  assign n26884 = n26883 ^ n25967;
  assign n26881 = n23173 ^ n21946;
  assign n26882 = n26881 ^ n23178;
  assign n26885 = n26884 ^ n26882;
  assign n26886 = n26885 ^ n23168;
  assign n26891 = n26890 ^ n26886;
  assign n26917 = n26907 ^ n26891;
  assign n26868 = n26021 ^ n23100;
  assign n26867 = n23173 ^ n23119;
  assign n26869 = n26868 ^ n26867;
  assign n26860 = n25931 ^ n23029;
  assign n26858 = n23144 ^ n23089;
  assign n26859 = n26858 ^ n23149;
  assign n26861 = n26860 ^ n26859;
  assign n26866 = n26865 ^ n26861;
  assign n26870 = n26869 ^ n26866;
  assign n26936 = n26917 ^ n26870;
  assign n26877 = n23201 ^ n23100;
  assign n26878 = n26877 ^ n25874;
  assign n26875 = n23059 ^ n23015;
  assign n26876 = n26875 ^ n23067;
  assign n26879 = n26878 ^ n26876;
  assign n26873 = n25901 ^ n23153;
  assign n26871 = n23089 ^ n23058;
  assign n26872 = n26871 ^ n23095;
  assign n26874 = n26873 ^ n26872;
  assign n26880 = n26879 ^ n26874;
  assign n26892 = n26891 ^ n26880;
  assign n26925 = n26892 ^ n26866;
  assign n26899 = n26898 ^ n26874;
  assign n26931 = n26925 ^ n26899;
  assign n26928 = n26879 ^ n26870;
  assign n26929 = ~n26869 & ~n26928;
  assign n26903 = n26898 ^ n26879;
  assign n26902 = n26885 ^ n26874;
  assign n26904 = n26903 ^ n26902;
  assign n26905 = ~n26892 & ~n26904;
  assign n26930 = n26929 ^ n26905;
  assign n26932 = n26931 ^ n26930;
  assign n26926 = n26899 & ~n26925;
  assign n26910 = n26898 ^ n26861;
  assign n26911 = n26910 ^ n26891;
  assign n26912 = n26880 & n26911;
  assign n26927 = n26926 ^ n26912;
  assign n26933 = n26932 ^ n26927;
  assign n26914 = n26910 ^ n26892;
  assign n26908 = n26907 ^ n26880;
  assign n26909 = n26903 & ~n26908;
  assign n26913 = n26912 ^ n26909;
  assign n26915 = n26914 ^ n26913;
  assign n26893 = n26892 ^ n26869;
  assign n26894 = n26885 ^ n26870;
  assign n26900 = n26899 ^ n26894;
  assign n26901 = n26893 & n26900;
  assign n26906 = n26905 ^ n26901;
  assign n26916 = n26915 ^ n26906;
  assign n26934 = n26933 ^ n26916;
  assign n26937 = n26928 ^ n26880;
  assign n26941 = n26937 ^ n26936;
  assign n26938 = ~n26936 & ~n26937;
  assign n26921 = ~n26902 & n26917;
  assign n26939 = n26938 ^ n26921;
  assign n26940 = n26939 ^ n26927;
  assign n26942 = n26941 ^ n26940;
  assign n26920 = ~n26870 & n26885;
  assign n26922 = n26921 ^ n26920;
  assign n26918 = n26917 ^ n26902;
  assign n26919 = n26918 ^ n26913;
  assign n26923 = n26922 ^ n26919;
  assign n26924 = n26916 & ~n26923;
  assign n26964 = n26942 ^ n26924;
  assign n26965 = ~n26934 & n26964;
  assign n26966 = n26965 ^ n26933;
  assign n27492 = ~n26936 & ~n26966;
  assign n26943 = n26916 & n26933;
  assign n26944 = n26942 & n26943;
  assign n26935 = n26934 ^ n26924;
  assign n26945 = n26944 ^ n26935;
  assign n27491 = n26894 & ~n26945;
  assign n27493 = n27492 ^ n27491;
  assign n26949 = n26942 ^ n26923;
  assign n26954 = n26933 ^ n26924;
  assign n26955 = ~n26949 & ~n26954;
  assign n26956 = n26955 ^ n26942;
  assign n27391 = ~n26869 & n26956;
  assign n26950 = n26949 ^ n26924;
  assign n26947 = ~n26923 & ~n26933;
  assign n26948 = ~n26942 & n26947;
  assign n26951 = n26950 ^ n26948;
  assign n26957 = n26956 ^ n26951;
  assign n26961 = ~n26892 & ~n26957;
  assign n27392 = n27391 ^ n26961;
  assign n27569 = n27493 ^ n27392;
  assign n26973 = n26966 ^ n26945;
  assign n27396 = ~n26902 & n26973;
  assign n26974 = n26917 & n26973;
  assign n26969 = n26951 ^ n26945;
  assign n26967 = n26966 ^ n26956;
  assign n26970 = n26969 ^ n26967;
  assign n26971 = n26903 & ~n26970;
  assign n26968 = n26880 & ~n26967;
  assign n26972 = n26971 ^ n26968;
  assign n26975 = n26974 ^ n26972;
  assign n27568 = n27396 ^ n26975;
  assign n27570 = n27569 ^ n27568;
  assign n27571 = n27570 ^ n26652;
  assign n27577 = n27576 ^ n27571;
  assign n27361 = ~n27329 & n27360;
  assign n27557 = n27381 ^ n27361;
  assign n27458 = n27319 & n27377;
  assign n27434 = ~n27333 & ~n27378;
  assign n27459 = n27458 ^ n27434;
  assign n27368 = ~n27330 & n27360;
  assign n27367 = ~n27326 & n27366;
  assign n27369 = n27368 ^ n27367;
  assign n27371 = n27370 ^ n27369;
  assign n27556 = n27459 ^ n27371;
  assign n27558 = n27557 ^ n27556;
  assign n27551 = n27171 & n27225;
  assign n27413 = ~n27168 & n27242;
  assign n27412 = ~n27173 & n27225;
  assign n27414 = n27413 ^ n27412;
  assign n27552 = n27551 ^ n27414;
  assign n27549 = n27246 ^ n27216;
  assign n27510 = ~n27145 & ~n27214;
  assign n27448 = ~n27172 & ~n27237;
  assign n27234 = ~n27133 & n27210;
  assign n27479 = n27448 ^ n27234;
  assign n27511 = n27510 ^ n27479;
  assign n27550 = n27549 ^ n27511;
  assign n27553 = n27552 ^ n27550;
  assign n27530 = n27013 & n27096;
  assign n27403 = ~n27025 & n27096;
  assign n27405 = n27404 ^ n27403;
  assign n27531 = n27530 ^ n27405;
  assign n27528 = n27112 ^ n27095;
  assign n27425 = ~n27033 & ~n27093;
  assign n27427 = n27426 ^ n27425;
  assign n27529 = n27528 ^ n27427;
  assign n27532 = n27531 ^ n27529;
  assign n27554 = n27553 ^ n27532;
  assign n26952 = n26900 & ~n26951;
  assign n27546 = n26972 ^ n26952;
  assign n27465 = n26911 & ~n26967;
  assign n27398 = ~n26908 & ~n26970;
  assign n27466 = n27465 ^ n27398;
  assign n26959 = n26893 & ~n26951;
  assign n26958 = ~n26904 & ~n26957;
  assign n26960 = n26959 ^ n26958;
  assign n26962 = n26961 ^ n26960;
  assign n27545 = n27466 ^ n26962;
  assign n27547 = n27546 ^ n27545;
  assign n27454 = n27099 ^ n27088;
  assign n27073 = n27007 & ~n27072;
  assign n27079 = n27078 ^ n27073;
  assign n27081 = n27080 ^ n27079;
  assign n27453 = n27114 ^ n27081;
  assign n27455 = n27454 ^ n27453;
  assign n27548 = n27547 ^ n27455;
  assign n27555 = n27554 ^ n27548;
  assign n27559 = n27558 ^ n27555;
  assign n27560 = n27559 ^ n26641;
  assign n27236 = n27201 & ~n27224;
  assign n27239 = n27238 ^ n27236;
  assign n27449 = n27448 ^ n27239;
  assign n27540 = n27449 ^ n27231;
  assign n27541 = n27540 ^ n27244;
  assign n27090 = n27089 ^ n27081;
  assign n27103 = n27102 ^ n27090;
  assign n27542 = n27541 ^ n27103;
  assign n27536 = ~n27314 & ~n27373;
  assign n27431 = ~n27316 & ~n27373;
  assign n27433 = n27432 ^ n27431;
  assign n27537 = n27536 ^ n27433;
  assign n27534 = n27458 ^ n27380;
  assign n27439 = ~n27309 & n27376;
  assign n27442 = n27441 ^ n27439;
  assign n27535 = n27534 ^ n27442;
  assign n27538 = n27537 ^ n27535;
  assign n27525 = n26899 & n26969;
  assign n27395 = ~n26925 & n26969;
  assign n27397 = n27396 ^ n27395;
  assign n27526 = n27525 ^ n27397;
  assign n27523 = n27465 ^ n26968;
  assign n27390 = ~n26937 & ~n26966;
  assign n27393 = n27392 ^ n27390;
  assign n27524 = n27523 ^ n27393;
  assign n27527 = n27526 ^ n27524;
  assign n27533 = n27532 ^ n27527;
  assign n27539 = n27538 ^ n27533;
  assign n27543 = n27542 ^ n27539;
  assign n27544 = n27543 ^ n26634;
  assign n27561 = n27560 ^ n27544;
  assign n27578 = n27577 ^ n27561;
  assign n27437 = n27301 & n27365;
  assign n27355 = n27271 & ~n27354;
  assign n27362 = n27361 ^ n27355;
  assign n27438 = n27437 ^ n27362;
  assign n27443 = n27442 ^ n27438;
  assign n27435 = n27434 ^ n27433;
  assign n27436 = n27435 ^ n27384;
  assign n27444 = n27443 ^ n27436;
  assign n27423 = ~n27032 & n27076;
  assign n27424 = n27423 ^ n27089;
  assign n27428 = n27427 ^ n27424;
  assign n27406 = n27405 ^ n27113;
  assign n27422 = n27406 ^ n27102;
  assign n27429 = n27428 ^ n27422;
  assign n27416 = n27199 & ~n27220;
  assign n27233 = ~n27166 & ~n27214;
  assign n27417 = n27416 ^ n27233;
  assign n27415 = n27414 ^ n27247;
  assign n27418 = n27417 ^ n27415;
  assign n27411 = n27229 ^ n27228;
  assign n27419 = n27418 ^ n27411;
  assign n27409 = n27408 ^ n27406;
  assign n27402 = n27099 ^ n27087;
  assign n27410 = n27409 ^ n27402;
  assign n27420 = n27419 ^ n27410;
  assign n27399 = n27398 ^ n27397;
  assign n27400 = n27399 ^ n26975;
  assign n27388 = ~n26928 & n26956;
  assign n26946 = ~n26870 & ~n26945;
  assign n26953 = n26952 ^ n26946;
  assign n27389 = n27388 ^ n26953;
  assign n27394 = n27393 ^ n27389;
  assign n27401 = n27400 ^ n27394;
  assign n27421 = n27420 ^ n27401;
  assign n27430 = n27429 ^ n27421;
  assign n27445 = n27444 ^ n27430;
  assign n27446 = n27445 ^ n26665;
  assign n27564 = n27560 ^ n27446;
  assign n27516 = n27484 ^ n27440;
  assign n27517 = n27516 ^ n27369;
  assign n27515 = n27381 ^ n27362;
  assign n27518 = n27517 ^ n27515;
  assign n27508 = ~n27144 & n27210;
  assign n27509 = n27508 ^ n27231;
  assign n27512 = n27511 ^ n27509;
  assign n27507 = n27415 ^ n27244;
  assign n27513 = n27512 ^ n27507;
  assign n27514 = n27513 ^ n27250;
  assign n27519 = n27518 ^ n27514;
  assign n27505 = n27429 ^ n27116;
  assign n27108 = n27107 ^ n27106;
  assign n27109 = n27108 ^ n27079;
  assign n27105 = n27099 ^ n27089;
  assign n27110 = n27109 ^ n27105;
  assign n27506 = n27505 ^ n27110;
  assign n27520 = n27519 ^ n27506;
  assign n27501 = n26972 ^ n26953;
  assign n27499 = n27492 ^ n27391;
  assign n27500 = n27499 ^ n26960;
  assign n27502 = n27501 ^ n27500;
  assign n27503 = n27502 ^ n26674;
  assign n27495 = n26972 ^ n26946;
  assign n27494 = n27493 ^ n27399;
  assign n27496 = n27495 ^ n27494;
  assign n27497 = n27496 ^ n26681;
  assign n27487 = n27381 ^ n27355;
  assign n27486 = n27485 ^ n27435;
  assign n27488 = n27487 ^ n27486;
  assign n27480 = n27479 ^ n27417;
  assign n27478 = n27413 ^ n27244;
  assign n27481 = n27480 ^ n27478;
  assign n27482 = n27481 ^ n27250;
  assign n27489 = n27488 ^ n27482;
  assign n27477 = n27476 ^ n27410;
  assign n27490 = n27489 ^ n27477;
  assign n27498 = n27497 ^ n27490;
  assign n27504 = n27503 ^ n27498;
  assign n27521 = n27520 ^ n27504;
  assign n27467 = n27466 ^ n26953;
  assign n27464 = n26975 ^ n26958;
  assign n27468 = n27467 ^ n27464;
  assign n27469 = n27468 ^ n26617;
  assign n27460 = n27459 ^ n27362;
  assign n27457 = n27384 ^ n27367;
  assign n27461 = n27460 ^ n27457;
  assign n27451 = n27230 ^ n27228;
  assign n27450 = n27449 ^ n27248;
  assign n27452 = n27451 ^ n27450;
  assign n27456 = n27455 ^ n27452;
  assign n27462 = n27461 ^ n27456;
  assign n27463 = n27462 ^ n27116;
  assign n27470 = n27469 ^ n27463;
  assign n27372 = n27371 ^ n27362;
  assign n27385 = n27384 ^ n27372;
  assign n27235 = n27234 ^ n27233;
  assign n27240 = n27239 ^ n27235;
  assign n27232 = n27231 ^ n27228;
  assign n27241 = n27240 ^ n27232;
  assign n27251 = n27250 ^ n27241;
  assign n27117 = n27116 ^ n27110;
  assign n26963 = n26962 ^ n26953;
  assign n26976 = n26975 ^ n26963;
  assign n27104 = n27103 ^ n26976;
  assign n27118 = n27117 ^ n27104;
  assign n27252 = n27251 ^ n27118;
  assign n27386 = n27385 ^ n27252;
  assign n27387 = n27386 ^ n26607;
  assign n27472 = n27470 ^ n27387;
  assign n27522 = n27521 ^ n27472;
  assign n27614 = n27564 ^ n27522;
  assign n27447 = n27446 ^ n27387;
  assign n27588 = n27544 ^ n27446;
  assign n27591 = n27588 ^ n27472;
  assign n27592 = n27447 & n27591;
  assign n27565 = n27564 ^ n27521;
  assign n27566 = n27472 & n27565;
  assign n27593 = n27592 ^ n27566;
  assign n27615 = n27614 ^ n27593;
  assign n27609 = n27577 ^ n27522;
  assign n27610 = n27578 ^ n27498;
  assign n27471 = n27470 ^ n27446;
  assign n27611 = n27610 ^ n27471;
  assign n27612 = n27609 & n27611;
  assign n27581 = n27498 ^ n27470;
  assign n27582 = n27581 ^ n27447;
  assign n27583 = n27522 & n27582;
  assign n27613 = n27612 ^ n27583;
  assign n27616 = n27615 ^ n27613;
  assign n27562 = n27561 ^ n27522;
  assign n27585 = n27562 ^ n27471;
  assign n27579 = n27578 ^ n27387;
  assign n27580 = n27577 & n27579;
  assign n27584 = n27583 ^ n27580;
  assign n27586 = n27585 ^ n27584;
  assign n27563 = n27471 & n27562;
  assign n27567 = n27566 ^ n27563;
  assign n27587 = n27586 ^ n27567;
  assign n27622 = n27616 ^ n27587;
  assign n27589 = n27588 ^ n27521;
  assign n27596 = n27581 & n27589;
  assign n27595 = ~n27498 & n27578;
  assign n27597 = n27596 ^ n27595;
  assign n27590 = n27589 ^ n27581;
  assign n27594 = n27593 ^ n27590;
  assign n27598 = n27597 ^ n27594;
  assign n27617 = n27598 & n27616;
  assign n27623 = n27622 ^ n27617;
  assign n27600 = n27579 ^ n27472;
  assign n27599 = n27589 ^ n27578;
  assign n27604 = n27600 ^ n27599;
  assign n27601 = n27599 & n27600;
  assign n27602 = n27601 ^ n27596;
  assign n27603 = n27602 ^ n27567;
  assign n27605 = n27604 ^ n27603;
  assign n27620 = ~n27587 & n27616;
  assign n27621 = n27605 & n27620;
  assign n27624 = n27623 ^ n27621;
  assign n27647 = n27578 & n27624;
  assign n27606 = n27605 ^ n27598;
  assign n27618 = n27617 ^ n27606;
  assign n27607 = n27598 & n27606;
  assign n27608 = n27587 & n27607;
  assign n27619 = n27618 ^ n27608;
  assign n27646 = n27611 & n27619;
  assign n27648 = n27647 ^ n27646;
  assign n27629 = n27617 ^ n27587;
  assign n27630 = n27606 & n27629;
  assign n27631 = n27630 ^ n27605;
  assign n27626 = n27617 ^ n27605;
  assign n27627 = n27622 & n27626;
  assign n27628 = n27627 ^ n27587;
  assign n27632 = n27631 ^ n27628;
  assign n27644 = n27565 & n27632;
  assign n27625 = n27624 ^ n27619;
  assign n27633 = n27632 ^ n27625;
  assign n27643 = n27591 & n27633;
  assign n27645 = n27644 ^ n27643;
  assign n27649 = n27648 ^ n27645;
  assign n27640 = n27631 ^ n27619;
  assign n27641 = n27582 & n27640;
  assign n27637 = n27628 ^ n27624;
  assign n27638 = n27589 & n27637;
  assign n27635 = n27472 & n27632;
  assign n27634 = n27447 & n27633;
  assign n27636 = n27635 ^ n27634;
  assign n27639 = n27638 ^ n27636;
  assign n27642 = n27641 ^ n27639;
  assign n27650 = n27649 ^ n27642;
  assign n27894 = n27893 ^ n27650;
  assign n27907 = n27889 ^ n27878;
  assign n27904 = ~n27822 & ~n27882;
  assign n27902 = n27851 & ~n27874;
  assign n27903 = n27902 ^ n27883;
  assign n27905 = n27904 ^ n27903;
  assign n27906 = n27905 ^ n27887;
  assign n27908 = n27907 ^ n27906;
  assign n27909 = n27908 ^ n26640;
  assign n27900 = n27646 ^ n27636;
  assign n27897 = n27522 & n27640;
  assign n27895 = n27609 & n27619;
  assign n27896 = n27895 ^ n27641;
  assign n27898 = n27897 ^ n27896;
  assign n27899 = n27898 ^ n27645;
  assign n27901 = n27900 ^ n27899;
  assign n27910 = n27909 ^ n27901;
  assign n27933 = n27885 ^ n27866;
  assign n27930 = n27821 & n27875;
  assign n27931 = n27930 ^ n26633;
  assign n27927 = ~n27818 & n27879;
  assign n27926 = ~n27823 & n27875;
  assign n27928 = n27927 ^ n27926;
  assign n27924 = ~n27816 & ~n27864;
  assign n27922 = ~n27812 & n27860;
  assign n27923 = n27922 ^ n27904;
  assign n27925 = n27924 ^ n27923;
  assign n27929 = n27928 ^ n27925;
  assign n27932 = n27931 ^ n27929;
  assign n27934 = n27933 ^ n27932;
  assign n27935 = n27934 ^ n27635;
  assign n27919 = n27471 & n27625;
  assign n27917 = n27581 & n27637;
  assign n27916 = n27562 & n27625;
  assign n27918 = n27917 ^ n27916;
  assign n27920 = n27919 ^ n27918;
  assign n27913 = n27600 & n27628;
  assign n27911 = n27577 & n27631;
  assign n27912 = n27911 ^ n27897;
  assign n27914 = n27913 ^ n27912;
  assign n27915 = n27914 ^ n27644;
  assign n27921 = n27920 ^ n27915;
  assign n27936 = n27935 ^ n27921;
  assign n27939 = n27905 ^ n27890;
  assign n27938 = n27881 ^ n26606;
  assign n27940 = n27939 ^ n27938;
  assign n27941 = n27940 ^ n27898;
  assign n27937 = n27648 ^ n27639;
  assign n27942 = n27941 ^ n27937;
  assign n27950 = ~n27814 & ~n27864;
  assign n27951 = n27950 ^ n27922;
  assign n27948 = n27903 ^ n27890;
  assign n27947 = n27878 ^ n26673;
  assign n27949 = n27948 ^ n27947;
  assign n27952 = n27951 ^ n27949;
  assign n27946 = n27599 & n27628;
  assign n27953 = n27952 ^ n27946;
  assign n27944 = n27911 ^ n27896;
  assign n27943 = n27648 ^ n27636;
  assign n27945 = n27944 ^ n27943;
  assign n27954 = n27953 ^ n27945;
  assign n27964 = ~n27815 & n27860;
  assign n27965 = n27964 ^ n27890;
  assign n27961 = n27928 ^ n27886;
  assign n27962 = n27961 ^ n27925;
  assign n27960 = n27881 ^ n26664;
  assign n27963 = n27962 ^ n27960;
  assign n27966 = n27965 ^ n27963;
  assign n27967 = n27966 ^ n27648;
  assign n27957 = n27579 & n27631;
  assign n27958 = n27957 ^ n27914;
  assign n27955 = n27918 ^ n27643;
  assign n27956 = n27955 ^ n27639;
  assign n27959 = n27958 ^ n27956;
  assign n27968 = n27967 ^ n27959;
  assign n27975 = n27849 & ~n27870;
  assign n27976 = n27975 ^ n27950;
  assign n27977 = n27976 ^ n27961;
  assign n27974 = n27888 ^ n27878;
  assign n27978 = n27977 ^ n27974;
  assign n27979 = n27978 ^ n26680;
  assign n27972 = n27647 ^ n27636;
  assign n27969 = n27610 & n27624;
  assign n27970 = n27969 ^ n27946;
  assign n27971 = n27970 ^ n27955;
  assign n27973 = n27972 ^ n27971;
  assign n27980 = n27979 ^ n27973;
  assign n27985 = n27976 ^ n27923;
  assign n27984 = n27927 ^ n27881;
  assign n27986 = n27985 ^ n27984;
  assign n27987 = n27986 ^ n26651;
  assign n27982 = n27970 ^ n27912;
  assign n27981 = n27917 ^ n27639;
  assign n27983 = n27982 ^ n27981;
  assign n27988 = n27987 ^ n27983;
  assign n28382 = n27262 ^ n24248;
  assign n28778 = n28382 ^ n25418;
  assign n28377 = n27267 ^ n24279;
  assign n28774 = n28377 ^ n25444;
  assign n28779 = n28778 ^ n28774;
  assign n28373 = n27256 ^ n24269;
  assign n28777 = n28373 ^ n25435;
  assign n28780 = n28779 ^ n28777;
  assign n28411 = n27275 ^ n24255;
  assign n28771 = n28411 ^ n25424;
  assign n28781 = n28780 ^ n28771;
  assign n28401 = n27289 ^ n24244;
  assign n28773 = n28401 ^ n25414;
  assign n28775 = n28774 ^ n28773;
  assign n28417 = n27282 ^ n24262;
  assign n28770 = n28417 ^ n25429;
  assign n28772 = n28771 ^ n28770;
  assign n28776 = n28775 ^ n28772;
  assign n28822 = n28780 ^ n28776;
  assign n28390 = n27298 ^ n24275;
  assign n28785 = n28390 ^ n25440;
  assign n28804 = n28785 ^ n28780;
  assign n28396 = n27305 ^ n24288;
  assign n28782 = n28396 ^ n25452;
  assign n28786 = n28785 ^ n28782;
  assign n28821 = n28804 ^ n28786;
  assign n28826 = n28822 ^ n28821;
  assign n28823 = ~n28821 & ~n28822;
  assign n28791 = n28782 ^ n28771;
  assign n28817 = ~n28776 & ~n28791;
  assign n28824 = n28823 ^ n28817;
  assign n28783 = n28782 ^ n28773;
  assign n28787 = n28786 ^ n28772;
  assign n28807 = n28787 ^ n28779;
  assign n28810 = ~n28783 & n28807;
  assign n28797 = n28778 ^ n28773;
  assign n28798 = n28797 ^ n28772;
  assign n28799 = ~n28786 & ~n28798;
  assign n28811 = n28810 ^ n28799;
  assign n28825 = n28824 ^ n28811;
  assign n28827 = n28826 ^ n28825;
  assign n28801 = n28797 ^ n28787;
  assign n28790 = n28785 ^ n28773;
  assign n28795 = n28786 ^ n28775;
  assign n28796 = n28790 & ~n28795;
  assign n28800 = n28799 ^ n28796;
  assign n28802 = n28801 ^ n28800;
  assign n28792 = n28791 ^ n28790;
  assign n28793 = n28787 & ~n28792;
  assign n28784 = n28783 ^ n28781;
  assign n28788 = n28787 ^ n28777;
  assign n28789 = ~n28784 & n28788;
  assign n28794 = n28793 ^ n28789;
  assign n28803 = n28802 ^ n28794;
  assign n28808 = n28807 ^ n28783;
  assign n28805 = n28777 & n28804;
  assign n28806 = n28805 ^ n28793;
  assign n28809 = n28808 ^ n28806;
  assign n28812 = n28811 ^ n28809;
  assign n28832 = n28803 & n28812;
  assign n28833 = n28827 & n28832;
  assign n28816 = ~n28771 & n28780;
  assign n28818 = n28817 ^ n28816;
  assign n28814 = n28791 ^ n28776;
  assign n28815 = n28814 ^ n28800;
  assign n28819 = n28818 ^ n28815;
  assign n28820 = n28803 & n28819;
  assign n28813 = n28812 ^ n28803;
  assign n28831 = n28820 ^ n28813;
  assign n28834 = n28833 ^ n28831;
  assign n28915 = n28781 & ~n28834;
  assign n28828 = n28827 ^ n28820;
  assign n28829 = ~n28813 & n28828;
  assign n28830 = n28829 ^ n28812;
  assign n28908 = ~n28822 & ~n28830;
  assign n28916 = n28915 ^ n28908;
  assign n28837 = n28827 ^ n28819;
  assign n28838 = n28820 ^ n28812;
  assign n28839 = n28837 & ~n28838;
  assign n28840 = n28839 ^ n28827;
  assign n28880 = n28777 & n28840;
  assign n28845 = n28837 ^ n28820;
  assign n28843 = ~n28812 & n28819;
  assign n28844 = ~n28827 & n28843;
  assign n28846 = n28845 ^ n28844;
  assign n28856 = n28846 ^ n28840;
  assign n28860 = n28787 & n28856;
  assign n28881 = n28880 ^ n28860;
  assign n28934 = n28916 ^ n28881;
  assign n28835 = n28834 ^ n28830;
  assign n28884 = ~n28791 & n28835;
  assign n28847 = n28846 ^ n28834;
  assign n28841 = n28840 ^ n28830;
  assign n28848 = n28847 ^ n28841;
  assign n28849 = n28790 & n28848;
  assign n28842 = ~n28786 & ~n28841;
  assign n28850 = n28849 ^ n28842;
  assign n28836 = ~n28776 & n28835;
  assign n28851 = n28850 ^ n28836;
  assign n28933 = n28884 ^ n28851;
  assign n28935 = n28934 ^ n28933;
  assign n28936 = n28935 ^ n26021;
  assign n28937 = n28936 ^ n26022;
  assign n28938 = n28937 ^ n26023;
  assign n28939 = n28938 ^ n26024;
  assign n28853 = ~n28784 & n28846;
  assign n28926 = n28853 ^ n28850;
  assign n28869 = ~n28795 & n28848;
  assign n28868 = ~n28798 & ~n28841;
  assign n28870 = n28869 ^ n28868;
  assign n28858 = n28788 & n28846;
  assign n28857 = ~n28792 & n28856;
  assign n28859 = n28858 ^ n28857;
  assign n28861 = n28860 ^ n28859;
  assign n28925 = n28870 ^ n28861;
  assign n28927 = n28926 ^ n28925;
  assign n28928 = n28927 ^ n25931;
  assign n28929 = n28928 ^ n25932;
  assign n28930 = n28929 ^ n25933;
  assign n28931 = n28930 ^ n25934;
  assign n28899 = n28868 ^ n28842;
  assign n28896 = ~n28783 & ~n28847;
  assign n28897 = n28896 ^ n25748;
  assign n28883 = n28807 & ~n28847;
  assign n28885 = n28884 ^ n28883;
  assign n28879 = ~n28821 & ~n28830;
  assign n28882 = n28881 ^ n28879;
  assign n28895 = n28885 ^ n28882;
  assign n28898 = n28897 ^ n28895;
  assign n28900 = n28899 ^ n28898;
  assign n28901 = n28900 ^ n25749;
  assign n28902 = n28901 ^ n25750;
  assign n28903 = n28902 ^ n25751;
  assign n28932 = n28931 ^ n28903;
  assign n28940 = n28939 ^ n28932;
  assign n28886 = n28885 ^ n28869;
  assign n28917 = n28916 ^ n28886;
  assign n28854 = n28780 & ~n28834;
  assign n28914 = n28854 ^ n28850;
  assign n28918 = n28917 ^ n28914;
  assign n28919 = n28918 ^ n25967;
  assign n28920 = n28919 ^ n25968;
  assign n28921 = n28920 ^ n25969;
  assign n28922 = n28921 ^ n25970;
  assign n28976 = n28940 ^ n28922;
  assign n28889 = n28804 & n28840;
  assign n28855 = n28854 ^ n28853;
  assign n28890 = n28889 ^ n28855;
  assign n28887 = n28886 ^ n28882;
  assign n28878 = n28851 ^ n25826;
  assign n28888 = n28887 ^ n28878;
  assign n28891 = n28890 ^ n28888;
  assign n28892 = n28891 ^ n25827;
  assign n28893 = n28892 ^ n25828;
  assign n28894 = n28893 ^ n25829;
  assign n28871 = n28870 ^ n28855;
  assign n28867 = n28857 ^ n28851;
  assign n28872 = n28871 ^ n28867;
  assign n28873 = n28872 ^ n25901;
  assign n28874 = n28873 ^ n25902;
  assign n28875 = n28874 ^ n25903;
  assign n28876 = n28875 ^ n25904;
  assign n28948 = n28894 ^ n28876;
  assign n28977 = n28976 ^ n28948;
  assign n28965 = n28922 & ~n28940;
  assign n28909 = n28908 ^ n28880;
  assign n28906 = n28859 ^ n28855;
  assign n28905 = n28850 ^ n25995;
  assign n28907 = n28906 ^ n28905;
  assign n28910 = n28909 ^ n28907;
  assign n28911 = n28910 ^ n25996;
  assign n28912 = n28911 ^ n25997;
  assign n28913 = n28912 ^ n25998;
  assign n28923 = n28922 ^ n28913;
  assign n28904 = n28903 ^ n28894;
  assign n28924 = n28923 ^ n28904;
  assign n28945 = n28922 ^ n28876;
  assign n28946 = n28924 & ~n28945;
  assign n28966 = n28965 ^ n28946;
  assign n28963 = n28945 ^ n28924;
  assign n28862 = n28861 ^ n28855;
  assign n28852 = n28851 ^ n25874;
  assign n28863 = n28862 ^ n28852;
  assign n28864 = n28863 ^ n25875;
  assign n28865 = n28864 ^ n25876;
  assign n28866 = n28865 ^ n25877;
  assign n28959 = n28894 ^ n28866;
  assign n28877 = n28876 ^ n28866;
  assign n28960 = n28904 ^ n28877;
  assign n28961 = n28959 & ~n28960;
  assign n28952 = n28931 ^ n28894;
  assign n28953 = n28952 ^ n28923;
  assign n28954 = n28877 & n28953;
  assign n28962 = n28961 ^ n28954;
  assign n28964 = n28963 ^ n28962;
  assign n28967 = n28966 ^ n28964;
  assign n28949 = n28923 ^ n28877;
  assign n28981 = n28952 ^ n28949;
  assign n28982 = n28981 ^ n28962;
  assign n28978 = n28949 ^ n28939;
  assign n28979 = n28977 & n28978;
  assign n28970 = n28959 ^ n28945;
  assign n28971 = ~n28949 & ~n28970;
  assign n28980 = n28979 ^ n28971;
  assign n28983 = n28982 ^ n28980;
  assign n28984 = ~n28967 & n28983;
  assign n28942 = n28940 ^ n28866;
  assign n28943 = n28942 ^ n28877;
  assign n28941 = n28940 ^ n28924;
  assign n28957 = n28943 ^ n28941;
  assign n28950 = n28949 ^ n28932;
  assign n28951 = n28948 & ~n28950;
  assign n28955 = n28954 ^ n28951;
  assign n28944 = ~n28941 & ~n28943;
  assign n28947 = n28946 ^ n28944;
  assign n28956 = n28955 ^ n28947;
  assign n28958 = n28957 ^ n28956;
  assign n28968 = n28967 ^ n28958;
  assign n29000 = n28984 ^ n28968;
  assign n28973 = n28950 ^ n28948;
  assign n28969 = ~n28939 & ~n28942;
  assign n28972 = n28971 ^ n28969;
  assign n28974 = n28973 ^ n28972;
  assign n28975 = n28974 ^ n28955;
  assign n28998 = ~n28967 & ~n28975;
  assign n28999 = ~n28958 & n28998;
  assign n29001 = n29000 ^ n28999;
  assign n29016 = n28977 & ~n29001;
  assign n28995 = n28975 & n28983;
  assign n28996 = n28958 & n28995;
  assign n28988 = n28983 ^ n28975;
  assign n28994 = n28988 ^ n28984;
  assign n28997 = n28996 ^ n28994;
  assign n29015 = ~n28940 & ~n28997;
  assign n29017 = n29016 ^ n29015;
  assign n29002 = n29001 ^ n28997;
  assign n28989 = n28984 ^ n28958;
  assign n28990 = ~n28988 & n28989;
  assign n28991 = n28990 ^ n28975;
  assign n28985 = n28984 ^ n28975;
  assign n28986 = ~n28968 & ~n28985;
  assign n28987 = n28986 ^ n28958;
  assign n28992 = n28991 ^ n28987;
  assign n29003 = n29002 ^ n28992;
  assign n29013 = ~n28960 & ~n29003;
  assign n29012 = n28953 & ~n28992;
  assign n29014 = n29013 ^ n29012;
  assign n29018 = n29017 ^ n29014;
  assign n29009 = n29001 ^ n28987;
  assign n29010 = ~n28970 & ~n29009;
  assign n29006 = n28997 ^ n28991;
  assign n29007 = n28924 & n29006;
  assign n29004 = n28959 & ~n29003;
  assign n28993 = n28877 & ~n28992;
  assign n29005 = n29004 ^ n28993;
  assign n29008 = n29007 ^ n29005;
  assign n29011 = n29010 ^ n29008;
  assign n29019 = n29018 ^ n29011;
  assign n29020 = n29019 ^ n27746;
  assign n28412 = n28411 ^ n24873;
  assign n28408 = n25092 ^ n24962;
  assign n28409 = n28408 ^ n27147;
  assign n28410 = n28409 ^ n27159;
  assign n28413 = n28412 ^ n28410;
  assign n28383 = n28382 ^ n24970;
  assign n28380 = n24994 ^ n24973;
  assign n28381 = n28380 ^ n24488;
  assign n28384 = n28383 ^ n28381;
  assign n28378 = n28377 ^ n24745;
  assign n28376 = n27134 ^ n24946;
  assign n28379 = n28378 ^ n28376;
  assign n28385 = n28384 ^ n28379;
  assign n28374 = n28373 ^ n25021;
  assign n28371 = n25088 ^ n25017;
  assign n28372 = n28371 ^ n24967;
  assign n28375 = n28374 ^ n28372;
  assign n28386 = n28385 ^ n28375;
  assign n28447 = n28413 ^ n28386;
  assign n28418 = n28417 ^ n24916;
  assign n28415 = n24962 ^ n24849;
  assign n28416 = n28415 ^ n27154;
  assign n28419 = n28418 ^ n28416;
  assign n28407 = n25073 ^ n24931;
  assign n28414 = n28413 ^ n28407;
  assign n28420 = n28419 ^ n28414;
  assign n28397 = n28396 ^ n24920;
  assign n28394 = n24966 ^ n24926;
  assign n28395 = n28394 ^ n24995;
  assign n28398 = n28397 ^ n28395;
  assign n28391 = n28390 ^ n24730;
  assign n28387 = n25069 ^ n24962;
  assign n28388 = n28387 ^ n27120;
  assign n28389 = n28388 ^ n27139;
  assign n28392 = n28391 ^ n28389;
  assign n28399 = n28398 ^ n28392;
  assign n28430 = n28420 ^ n28399;
  assign n28403 = n25063 ^ n24864;
  assign n28404 = n28403 ^ n25036;
  assign n28402 = n28401 ^ n24891;
  assign n28405 = n28404 ^ n28402;
  assign n28427 = n28405 ^ n28384;
  assign n28454 = n28430 ^ n28427;
  assign n28438 = n28405 ^ n28392;
  assign n28406 = n28405 ^ n28379;
  assign n28451 = n28406 ^ n28399;
  assign n28452 = ~n28438 & ~n28451;
  assign n28428 = n28427 ^ n28420;
  assign n28429 = ~n28399 & ~n28428;
  assign n28453 = n28452 ^ n28429;
  assign n28455 = n28454 ^ n28453;
  assign n28446 = n28430 ^ n28375;
  assign n28432 = n28405 ^ n28398;
  assign n28448 = n28447 ^ n28432;
  assign n28449 = n28446 & ~n28448;
  assign n28424 = n28413 ^ n28398;
  assign n28439 = n28438 ^ n28424;
  assign n28440 = ~n28430 & ~n28439;
  assign n28450 = n28449 ^ n28440;
  assign n28456 = n28455 ^ n28450;
  assign n28431 = n28430 ^ n28385;
  assign n28443 = n28432 ^ n28431;
  assign n28393 = n28392 ^ n28386;
  assign n28441 = ~n28375 & n28393;
  assign n28442 = n28441 ^ n28440;
  assign n28444 = n28443 ^ n28442;
  assign n28433 = n28431 & n28432;
  assign n28434 = n28433 ^ n28429;
  assign n28445 = n28444 ^ n28434;
  assign n28465 = n28456 ^ n28445;
  assign n28461 = n28386 & n28413;
  assign n28421 = n28420 ^ n28406;
  assign n28425 = n28421 & n28424;
  assign n28462 = n28461 ^ n28425;
  assign n28459 = n28424 ^ n28421;
  assign n28460 = n28459 ^ n28453;
  assign n28463 = n28462 ^ n28460;
  assign n28464 = n28456 & n28463;
  assign n28466 = n28465 ^ n28464;
  assign n28422 = n28421 ^ n28386;
  assign n28400 = n28399 ^ n28393;
  assign n28436 = n28422 ^ n28400;
  assign n28423 = ~n28400 & n28422;
  assign n28426 = n28425 ^ n28423;
  assign n28435 = n28434 ^ n28426;
  assign n28437 = n28436 ^ n28435;
  assign n28457 = ~n28445 & n28456;
  assign n28458 = ~n28437 & n28457;
  assign n28467 = n28466 ^ n28458;
  assign n28611 = ~n28447 & n28467;
  assign n28486 = n28464 ^ n28437;
  assign n28487 = n28465 & ~n28486;
  assign n28488 = n28487 ^ n28445;
  assign n28610 = n28422 & n28488;
  assign n28612 = n28611 ^ n28610;
  assign n28469 = n28463 ^ n28437;
  assign n28477 = n28464 ^ n28445;
  assign n28478 = ~n28469 & n28477;
  assign n28479 = n28478 ^ n28437;
  assign n28558 = ~n28375 & ~n28479;
  assign n28471 = n28445 & n28463;
  assign n28472 = n28437 & n28471;
  assign n28470 = n28469 ^ n28464;
  assign n28473 = n28472 ^ n28470;
  assign n28480 = n28479 ^ n28473;
  assign n28483 = ~n28430 & n28480;
  assign n28559 = n28558 ^ n28483;
  assign n28695 = n28612 ^ n28559;
  assign n28495 = n28488 ^ n28467;
  assign n28551 = n28424 & n28495;
  assign n28496 = n28421 & n28495;
  assign n28491 = n28473 ^ n28467;
  assign n28489 = n28488 ^ n28479;
  assign n28492 = n28491 ^ n28489;
  assign n28493 = ~n28438 & n28492;
  assign n28490 = ~n28399 & ~n28489;
  assign n28494 = n28493 ^ n28490;
  assign n28497 = n28496 ^ n28494;
  assign n28694 = n28551 ^ n28497;
  assign n28696 = n28695 ^ n28694;
  assign n28288 = n25989 ^ n25955;
  assign n28289 = n28288 ^ n25782;
  assign n28290 = n28289 ^ n25766;
  assign n28291 = n28290 ^ n26108;
  assign n28257 = n27014 ^ n25531;
  assign n28258 = n28257 ^ n25855;
  assign n28259 = n28258 ^ n26111;
  assign n28304 = n28291 ^ n28259;
  assign n28282 = n25887 ^ n25797;
  assign n28283 = n28282 ^ n25836;
  assign n28281 = n26997 ^ n25976;
  assign n28284 = n28283 ^ n28281;
  assign n28279 = n26114 ^ n25866;
  assign n28277 = n26116 ^ n25810;
  assign n28274 = n26015 ^ n25887;
  assign n28275 = n28274 ^ n25761;
  assign n28273 = n26990 ^ n25948;
  assign n28276 = n28275 ^ n28273;
  assign n28278 = n28277 ^ n28276;
  assign n28280 = n28279 ^ n28278;
  assign n28285 = n28284 ^ n28280;
  assign n28311 = n28304 ^ n28285;
  assign n28254 = n26984 ^ n25412;
  assign n28255 = n28254 ^ n25891;
  assign n28256 = n28255 ^ n26120;
  assign n28260 = n28259 ^ n28256;
  assign n28252 = n26123 ^ n25959;
  assign n28250 = n25940 ^ n25887;
  assign n28251 = n28250 ^ n26990;
  assign n28253 = n28252 ^ n28251;
  assign n28261 = n28260 ^ n28253;
  assign n28330 = n28311 ^ n28261;
  assign n28270 = n26128 ^ n25861;
  assign n28268 = n25916 ^ n25840;
  assign n28267 = n25913 ^ n25883;
  assign n28269 = n28268 ^ n28267;
  assign n28271 = n28270 ^ n28269;
  assign n28263 = n25980 ^ n25887;
  assign n28262 = n27019 ^ n26977;
  assign n28264 = n28263 ^ n28262;
  assign n28265 = n28264 ^ n25545;
  assign n28266 = n28265 ^ n26106;
  assign n28272 = n28271 ^ n28266;
  assign n28286 = n28285 ^ n28272;
  assign n28319 = n28286 ^ n28260;
  assign n28296 = n28291 ^ n28271;
  assign n28325 = n28319 ^ n28296;
  assign n28322 = n28266 ^ n28261;
  assign n28323 = ~n28253 & ~n28322;
  assign n28292 = n28291 ^ n28266;
  assign n28287 = n28278 ^ n28271;
  assign n28293 = n28292 ^ n28287;
  assign n28294 = ~n28286 & ~n28293;
  assign n28324 = n28323 ^ n28294;
  assign n28326 = n28325 ^ n28324;
  assign n28320 = n28296 & ~n28319;
  assign n28301 = n28291 ^ n28256;
  assign n28302 = n28301 ^ n28285;
  assign n28303 = n28272 & n28302;
  assign n28321 = n28320 ^ n28303;
  assign n28327 = n28326 ^ n28321;
  assign n28308 = n28301 ^ n28286;
  assign n28305 = n28304 ^ n28272;
  assign n28306 = n28292 & ~n28305;
  assign n28307 = n28306 ^ n28303;
  assign n28309 = n28308 ^ n28307;
  assign n28295 = n28286 ^ n28253;
  assign n28297 = n28278 ^ n28261;
  assign n28298 = n28297 ^ n28296;
  assign n28299 = n28295 & n28298;
  assign n28300 = n28299 ^ n28294;
  assign n28310 = n28309 ^ n28300;
  assign n28328 = n28327 ^ n28310;
  assign n28331 = n28322 ^ n28272;
  assign n28335 = n28331 ^ n28330;
  assign n28332 = ~n28330 & ~n28331;
  assign n28314 = ~n28287 & n28311;
  assign n28333 = n28332 ^ n28314;
  assign n28334 = n28333 ^ n28321;
  assign n28336 = n28335 ^ n28334;
  assign n28315 = ~n28261 & n28278;
  assign n28316 = n28315 ^ n28314;
  assign n28312 = n28311 ^ n28287;
  assign n28313 = n28312 ^ n28307;
  assign n28317 = n28316 ^ n28313;
  assign n28318 = n28310 & ~n28317;
  assign n28358 = n28336 ^ n28318;
  assign n28359 = ~n28328 & n28358;
  assign n28360 = n28359 ^ n28327;
  assign n28605 = ~n28330 & ~n28360;
  assign n28337 = n28310 & n28327;
  assign n28338 = n28336 & n28337;
  assign n28329 = n28328 ^ n28318;
  assign n28339 = n28338 ^ n28329;
  assign n28604 = n28297 & ~n28339;
  assign n28606 = n28605 ^ n28604;
  assign n28343 = n28336 ^ n28317;
  assign n28349 = n28327 ^ n28318;
  assign n28350 = ~n28343 & ~n28349;
  assign n28351 = n28350 ^ n28336;
  assign n28544 = ~n28253 & n28351;
  assign n28344 = n28343 ^ n28318;
  assign n28341 = ~n28317 & ~n28327;
  assign n28342 = ~n28336 & n28341;
  assign n28345 = n28344 ^ n28342;
  assign n28352 = n28351 ^ n28345;
  assign n28355 = ~n28286 & ~n28352;
  assign n28545 = n28544 ^ n28355;
  assign n28691 = n28606 ^ n28545;
  assign n28367 = n28360 ^ n28339;
  assign n28537 = ~n28287 & n28367;
  assign n28368 = n28311 & n28367;
  assign n28363 = n28345 ^ n28339;
  assign n28361 = n28360 ^ n28351;
  assign n28364 = n28363 ^ n28361;
  assign n28365 = n28292 & ~n28364;
  assign n28362 = n28272 & ~n28361;
  assign n28366 = n28365 ^ n28362;
  assign n28369 = n28368 ^ n28366;
  assign n28690 = n28537 ^ n28369;
  assign n28692 = n28691 ^ n28690;
  assign n28145 = n24149 ^ n24037;
  assign n28146 = n28145 ^ n25968;
  assign n28143 = n27272 ^ n24079;
  assign n28144 = n28143 ^ n23950;
  assign n28147 = n28146 ^ n28144;
  assign n28131 = n26022 ^ n24037;
  assign n28130 = n27272 ^ n27254;
  assign n28132 = n28131 ^ n28130;
  assign n28127 = n25749 ^ n23685;
  assign n28125 = n23991 ^ n23820;
  assign n28126 = n28125 ^ n24057;
  assign n28128 = n28127 ^ n28126;
  assign n28123 = n25932 ^ n23997;
  assign n28121 = n24065 ^ n23991;
  assign n28122 = n28121 ^ n27260;
  assign n28124 = n28123 ^ n28122;
  assign n28129 = n28128 ^ n28124;
  assign n28133 = n28132 ^ n28129;
  assign n28148 = n28147 ^ n28133;
  assign n28136 = n25827 ^ n24096;
  assign n28134 = n24079 ^ n23923;
  assign n28135 = n28134 ^ n27287;
  assign n28137 = n28136 ^ n28135;
  assign n28170 = n28137 ^ n28128;
  assign n28152 = n24037 ^ n23964;
  assign n28153 = n28152 ^ n25996;
  assign n28151 = n27280 ^ n24122;
  assign n28154 = n28153 ^ n28151;
  assign n28150 = n28147 ^ n27278;
  assign n28155 = n28154 ^ n28150;
  assign n28180 = n28170 ^ n28155;
  assign n28200 = n28180 ^ n28133;
  assign n28158 = n24110 ^ n24037;
  assign n28159 = n28158 ^ n25875;
  assign n28156 = n27295 ^ n23820;
  assign n28157 = n28156 ^ n24009;
  assign n28160 = n28159 ^ n28157;
  assign n28188 = n28160 ^ n28133;
  assign n28140 = n25902 ^ n24060;
  assign n28138 = n24065 ^ n24024;
  assign n28139 = n28138 ^ n27303;
  assign n28141 = n28140 ^ n28139;
  assign n28161 = n28160 ^ n28141;
  assign n28199 = n28188 ^ n28161;
  assign n28204 = n28200 ^ n28199;
  assign n28201 = ~n28199 & ~n28200;
  assign n28166 = n28147 ^ n28141;
  assign n28184 = ~n28166 & n28180;
  assign n28202 = n28201 ^ n28184;
  assign n28142 = n28141 ^ n28137;
  assign n28162 = n28161 ^ n28155;
  assign n28191 = n28162 ^ n28129;
  assign n28194 = n28142 & ~n28191;
  assign n28173 = n28137 ^ n28124;
  assign n28174 = n28173 ^ n28155;
  assign n28175 = n28161 & n28174;
  assign n28195 = n28194 ^ n28175;
  assign n28203 = n28202 ^ n28195;
  assign n28205 = n28204 ^ n28203;
  assign n28177 = n28173 ^ n28162;
  assign n28165 = n28160 ^ n28137;
  assign n28171 = n28170 ^ n28161;
  assign n28172 = n28165 & ~n28171;
  assign n28176 = n28175 ^ n28172;
  assign n28178 = n28177 ^ n28176;
  assign n28167 = n28166 ^ n28165;
  assign n28168 = ~n28162 & ~n28167;
  assign n28149 = n28148 ^ n28142;
  assign n28163 = n28162 ^ n28132;
  assign n28164 = n28149 & n28163;
  assign n28169 = n28168 ^ n28164;
  assign n28179 = n28178 ^ n28169;
  assign n28192 = n28191 ^ n28142;
  assign n28189 = ~n28132 & ~n28188;
  assign n28190 = n28189 ^ n28168;
  assign n28193 = n28192 ^ n28190;
  assign n28196 = n28195 ^ n28193;
  assign n28206 = n28179 & n28196;
  assign n28207 = n28205 & n28206;
  assign n28197 = n28196 ^ n28179;
  assign n28183 = ~n28133 & n28147;
  assign n28185 = n28184 ^ n28183;
  assign n28181 = n28180 ^ n28166;
  assign n28182 = n28181 ^ n28176;
  assign n28186 = n28185 ^ n28182;
  assign n28187 = n28179 & ~n28186;
  assign n28198 = n28197 ^ n28187;
  assign n28208 = n28207 ^ n28198;
  assign n28530 = n28148 & ~n28208;
  assign n28220 = n28205 ^ n28187;
  assign n28221 = ~n28197 & n28220;
  assign n28222 = n28221 ^ n28196;
  assign n28231 = ~n28200 & ~n28222;
  assign n28531 = n28530 ^ n28231;
  assign n28212 = n28205 ^ n28186;
  assign n28217 = n28196 ^ n28187;
  assign n28218 = ~n28212 & ~n28217;
  assign n28219 = n28218 ^ n28205;
  assign n28213 = n28212 ^ n28187;
  assign n28210 = ~n28186 & ~n28196;
  assign n28211 = ~n28205 & n28210;
  assign n28214 = n28213 ^ n28211;
  assign n28234 = n28219 ^ n28214;
  assign n28501 = ~n28162 & ~n28234;
  assign n28230 = ~n28132 & n28219;
  assign n28515 = n28501 ^ n28230;
  assign n28599 = n28531 ^ n28515;
  assign n28239 = n28222 ^ n28208;
  assign n28508 = ~n28166 & n28239;
  assign n28240 = n28180 & n28239;
  assign n28225 = n28214 ^ n28208;
  assign n28223 = n28222 ^ n28219;
  assign n28226 = n28225 ^ n28223;
  assign n28227 = n28165 & ~n28226;
  assign n28224 = n28161 & ~n28223;
  assign n28228 = n28227 ^ n28224;
  assign n28241 = n28240 ^ n28228;
  assign n28598 = n28508 ^ n28241;
  assign n28600 = n28599 ^ n28598;
  assign n28244 = ~n28171 & ~n28226;
  assign n28243 = n28174 & ~n28223;
  assign n28245 = n28244 ^ n28243;
  assign n28215 = n28149 & ~n28214;
  assign n28209 = ~n28133 & ~n28208;
  assign n28216 = n28215 ^ n28209;
  assign n28246 = n28245 ^ n28216;
  assign n28235 = ~n28167 & ~n28234;
  assign n28242 = n28241 ^ n28235;
  assign n28247 = n28246 ^ n28242;
  assign n28601 = n28600 ^ n28247;
  assign n28034 = n24954 ^ n23074;
  assign n28031 = n23167 ^ n23094;
  assign n28032 = n28031 ^ n26877;
  assign n28033 = n28032 ^ n23022;
  assign n28035 = n28034 ^ n28033;
  assign n28027 = n24980 ^ n23100;
  assign n28025 = n23153 ^ n23148;
  assign n28026 = n28025 ^ n23120;
  assign n28028 = n28027 ^ n28026;
  assign n28036 = n28035 ^ n28028;
  assign n28019 = n24907 ^ n22878;
  assign n28017 = n23182 ^ n23177;
  assign n28016 = n23195 ^ n21041;
  assign n28018 = n28017 ^ n28016;
  assign n28020 = n28019 ^ n28018;
  assign n28000 = n24830 ^ n23029;
  assign n27998 = n23074 ^ n23066;
  assign n27999 = n27998 ^ n23145;
  assign n28001 = n28000 ^ n27999;
  assign n28021 = n28020 ^ n28001;
  assign n28045 = n28036 ^ n28021;
  assign n27996 = n25009 ^ n23153;
  assign n27994 = n23029 ^ n23002;
  assign n27995 = n27994 ^ n23090;
  assign n27997 = n27996 ^ n27995;
  assign n28002 = n28001 ^ n27997;
  assign n27992 = n25097 ^ n23127;
  assign n27990 = n23100 ^ n23094;
  assign n27989 = n23172 ^ n23118;
  assign n27991 = n27990 ^ n27989;
  assign n27993 = n27992 ^ n27991;
  assign n28003 = n28002 ^ n27993;
  assign n28054 = n28035 ^ n28003;
  assign n28071 = n28054 ^ n28036;
  assign n28012 = n23094 ^ n20100;
  assign n28013 = n28012 ^ n26887;
  assign n28011 = n23053 ^ n23043;
  assign n28014 = n28013 ^ n28011;
  assign n28008 = n25044 ^ n23182;
  assign n28005 = n23115 ^ n23094;
  assign n28006 = n28005 ^ n26883;
  assign n28007 = n28006 ^ n21953;
  assign n28009 = n28008 ^ n28007;
  assign n28004 = n25053 ^ n23201;
  assign n28010 = n28009 ^ n28004;
  assign n28015 = n28014 ^ n28010;
  assign n28022 = n28021 ^ n28015;
  assign n28023 = n28022 ^ n28003;
  assign n28075 = n28071 ^ n28023;
  assign n28072 = ~n28023 & ~n28071;
  assign n28041 = n28028 ^ n28009;
  assign n28067 = n28022 & ~n28041;
  assign n28073 = n28072 ^ n28067;
  assign n28029 = n28028 ^ n28020;
  assign n28037 = n28036 ^ n28015;
  assign n28057 = n28037 ^ n28002;
  assign n28060 = n28029 & ~n28057;
  assign n28047 = n28020 ^ n27997;
  assign n28048 = n28047 ^ n28015;
  assign n28049 = n28036 & n28048;
  assign n28061 = n28060 ^ n28049;
  assign n28074 = n28073 ^ n28061;
  assign n28076 = n28075 ^ n28074;
  assign n28051 = n28047 ^ n28037;
  assign n28040 = n28035 ^ n28020;
  assign n28046 = n28040 & ~n28045;
  assign n28050 = n28049 ^ n28046;
  assign n28052 = n28051 ^ n28050;
  assign n28042 = n28041 ^ n28040;
  assign n28043 = ~n28037 & ~n28042;
  assign n28024 = n28009 ^ n28003;
  assign n28030 = n28029 ^ n28024;
  assign n28038 = n28037 ^ n27993;
  assign n28039 = n28030 & n28038;
  assign n28044 = n28043 ^ n28039;
  assign n28053 = n28052 ^ n28044;
  assign n28058 = n28057 ^ n28029;
  assign n28055 = ~n27993 & ~n28054;
  assign n28056 = n28055 ^ n28043;
  assign n28059 = n28058 ^ n28056;
  assign n28062 = n28061 ^ n28059;
  assign n28099 = n28053 & n28062;
  assign n28100 = n28076 & n28099;
  assign n28066 = ~n28003 & n28009;
  assign n28068 = n28067 ^ n28066;
  assign n28064 = n28041 ^ n28022;
  assign n28065 = n28064 ^ n28050;
  assign n28069 = n28068 ^ n28065;
  assign n28070 = n28053 & ~n28069;
  assign n28063 = n28062 ^ n28053;
  assign n28098 = n28070 ^ n28063;
  assign n28101 = n28100 ^ n28098;
  assign n28081 = n28076 ^ n28069;
  assign n28089 = n28081 ^ n28070;
  assign n28087 = ~n28062 & ~n28069;
  assign n28088 = ~n28076 & n28087;
  assign n28090 = n28089 ^ n28088;
  assign n28102 = n28101 ^ n28090;
  assign n28082 = n28070 ^ n28062;
  assign n28083 = ~n28081 & ~n28082;
  assign n28084 = n28083 ^ n28076;
  assign n28077 = n28076 ^ n28070;
  assign n28078 = ~n28063 & n28077;
  assign n28079 = n28078 ^ n28062;
  assign n28096 = n28084 ^ n28079;
  assign n28103 = n28102 ^ n28096;
  assign n28116 = ~n28045 & ~n28103;
  assign n28115 = n28048 & ~n28096;
  assign n28117 = n28116 ^ n28115;
  assign n28107 = n28030 & ~n28090;
  assign n28106 = ~n28003 & ~n28101;
  assign n28108 = n28107 ^ n28106;
  assign n28118 = n28117 ^ n28108;
  assign n28111 = n28101 ^ n28079;
  assign n28112 = n28022 & n28111;
  assign n28104 = n28040 & ~n28103;
  assign n28097 = n28036 & ~n28096;
  assign n28105 = n28104 ^ n28097;
  assign n28113 = n28112 ^ n28105;
  assign n28092 = n28090 ^ n28084;
  assign n28093 = ~n28042 & ~n28092;
  assign n28114 = n28113 ^ n28093;
  assign n28119 = n28118 ^ n28114;
  assign n28689 = n28601 ^ n28119;
  assign n28693 = n28692 ^ n28689;
  assign n28697 = n28696 ^ n28693;
  assign n28698 = n28697 ^ n27811;
  assign n28649 = n28142 & n28225;
  assign n28507 = ~n28191 & n28225;
  assign n28509 = n28508 ^ n28507;
  assign n28650 = n28649 ^ n28509;
  assign n28647 = n28243 ^ n28224;
  assign n28514 = ~n28199 & ~n28222;
  assign n28516 = n28515 ^ n28514;
  assign n28648 = n28647 ^ n28516;
  assign n28651 = n28650 ^ n28648;
  assign n28678 = n28651 ^ n27775;
  assign n28673 = n28432 & ~n28491;
  assign n28550 = n28431 & ~n28491;
  assign n28552 = n28551 ^ n28550;
  assign n28674 = n28673 ^ n28552;
  assign n28582 = ~n28428 & ~n28489;
  assign n28671 = n28582 ^ n28490;
  assign n28557 = ~n28400 & n28488;
  assign n28560 = n28559 ^ n28557;
  assign n28672 = n28671 ^ n28560;
  assign n28675 = n28674 ^ n28672;
  assign n28668 = n28296 & n28363;
  assign n28536 = ~n28319 & n28363;
  assign n28538 = n28537 ^ n28536;
  assign n28669 = n28668 ^ n28538;
  assign n28577 = n28302 & ~n28361;
  assign n28666 = n28577 ^ n28362;
  assign n28543 = ~n28331 & ~n28360;
  assign n28546 = n28545 ^ n28543;
  assign n28667 = n28666 ^ n28546;
  assign n28670 = n28669 ^ n28667;
  assign n28676 = n28675 ^ n28670;
  assign n28567 = ~n28037 & ~n28092;
  assign n28091 = n28038 & ~n28090;
  assign n28094 = n28093 ^ n28091;
  assign n28568 = n28567 ^ n28094;
  assign n28663 = n28568 ^ n28108;
  assign n28664 = n28663 ^ n28113;
  assign n28233 = n28163 & ~n28214;
  assign n28236 = n28235 ^ n28233;
  assign n28502 = n28501 ^ n28236;
  assign n28503 = n28502 ^ n28216;
  assign n28504 = n28503 ^ n28241;
  assign n28665 = n28664 ^ n28504;
  assign n28677 = n28676 ^ n28665;
  assign n28679 = n28678 ^ n28677;
  assign n28573 = n28228 ^ n28215;
  assign n28572 = n28502 ^ n28245;
  assign n28574 = n28573 ^ n28572;
  assign n28661 = n28574 ^ n27803;
  assign n28474 = ~n28448 & ~n28473;
  assign n28657 = n28494 ^ n28474;
  assign n28549 = ~n28451 & n28492;
  assign n28583 = n28582 ^ n28549;
  assign n28481 = ~n28439 & n28480;
  assign n28476 = n28446 & ~n28473;
  assign n28482 = n28481 ^ n28476;
  assign n28484 = n28483 ^ n28482;
  assign n28656 = n28583 ^ n28484;
  assign n28658 = n28657 ^ n28656;
  assign n28346 = n28298 & ~n28345;
  assign n28654 = n28366 ^ n28346;
  assign n28535 = ~n28305 & ~n28364;
  assign n28578 = n28577 ^ n28535;
  assign n28353 = ~n28293 & ~n28352;
  assign n28348 = n28295 & ~n28345;
  assign n28354 = n28353 ^ n28348;
  assign n28356 = n28355 ^ n28354;
  assign n28653 = n28578 ^ n28356;
  assign n28655 = n28654 ^ n28653;
  assign n28659 = n28658 ^ n28655;
  assign n28644 = n28029 & n28102;
  assign n28521 = ~n28057 & n28102;
  assign n28520 = ~n28041 & n28111;
  assign n28522 = n28521 ^ n28520;
  assign n28645 = n28644 ^ n28522;
  assign n28642 = n28115 ^ n28097;
  assign n28622 = ~n28071 & ~n28079;
  assign n28085 = ~n27993 & n28084;
  assign n28594 = n28567 ^ n28085;
  assign n28623 = n28622 ^ n28594;
  assign n28643 = n28642 ^ n28623;
  assign n28646 = n28645 ^ n28643;
  assign n28652 = n28651 ^ n28646;
  assign n28660 = n28659 ^ n28652;
  assign n28662 = n28661 ^ n28660;
  assign n28680 = n28679 ^ n28662;
  assign n28699 = n28698 ^ n28680;
  assign n28510 = n28509 ^ n28244;
  assign n28532 = n28531 ^ n28510;
  assign n28529 = n28228 ^ n28209;
  assign n28533 = n28532 ^ n28529;
  assign n28617 = n28533 ^ n27794;
  assign n28553 = n28552 ^ n28549;
  assign n28613 = n28612 ^ n28553;
  assign n28468 = n28386 & n28467;
  assign n28609 = n28494 ^ n28468;
  assign n28614 = n28613 ^ n28609;
  assign n28539 = n28538 ^ n28535;
  assign n28607 = n28606 ^ n28539;
  assign n28340 = ~n28261 & ~n28339;
  assign n28603 = n28366 ^ n28340;
  assign n28608 = n28607 ^ n28603;
  assign n28615 = n28614 ^ n28608;
  assign n28524 = n28024 & ~n28101;
  assign n28080 = ~n28023 & ~n28079;
  assign n28525 = n28524 ^ n28080;
  assign n28595 = n28594 ^ n28525;
  assign n28593 = n28520 ^ n28113;
  assign n28596 = n28595 ^ n28593;
  assign n28597 = n28596 ^ n28119;
  assign n28602 = n28601 ^ n28597;
  assign n28616 = n28615 ^ n28602;
  assign n28618 = n28617 ^ n28616;
  assign n28710 = n28699 ^ n28618;
  assign n28588 = n28247 ^ n27748;
  assign n28475 = n28474 ^ n28468;
  assign n28584 = n28583 ^ n28475;
  assign n28581 = n28497 ^ n28481;
  assign n28585 = n28584 ^ n28581;
  assign n28347 = n28346 ^ n28340;
  assign n28579 = n28578 ^ n28347;
  assign n28576 = n28369 ^ n28353;
  assign n28580 = n28579 ^ n28576;
  assign n28586 = n28585 ^ n28580;
  assign n28570 = n28107 ^ n28105;
  assign n28569 = n28568 ^ n28117;
  assign n28571 = n28570 ^ n28569;
  assign n28575 = n28574 ^ n28571;
  assign n28587 = n28586 ^ n28575;
  assign n28589 = n28588 ^ n28587;
  assign n28555 = n28393 & ~n28479;
  assign n28556 = n28555 ^ n28475;
  assign n28561 = n28560 ^ n28556;
  assign n28554 = n28553 ^ n28497;
  assign n28562 = n28561 ^ n28554;
  assign n28541 = ~n28322 & n28351;
  assign n28542 = n28541 ^ n28347;
  assign n28547 = n28546 ^ n28542;
  assign n28540 = n28539 ^ n28369;
  assign n28548 = n28547 ^ n28540;
  assign n28563 = n28562 ^ n28548;
  assign n28527 = n28106 ^ n28105;
  assign n28523 = n28522 ^ n28116;
  assign n28526 = n28525 ^ n28523;
  assign n28528 = n28527 ^ n28526;
  assign n28534 = n28533 ^ n28528;
  assign n28564 = n28563 ^ n28534;
  assign n28512 = ~n28188 & n28219;
  assign n28513 = n28512 ^ n28216;
  assign n28517 = n28516 ^ n28513;
  assign n28511 = n28510 ^ n28241;
  assign n28518 = n28517 ^ n28511;
  assign n28519 = n28518 ^ n27766;
  assign n28565 = n28564 ^ n28519;
  assign n28590 = n28589 ^ n28565;
  assign n28711 = n28710 ^ n28590;
  assign n28733 = ~n28618 & n28699;
  assign n28687 = n28679 ^ n28565;
  assign n28635 = n28610 ^ n28558;
  assign n28636 = n28635 ^ n28482;
  assign n28634 = n28494 ^ n28475;
  assign n28637 = n28636 ^ n28634;
  assign n28631 = n28605 ^ n28544;
  assign n28632 = n28631 ^ n28354;
  assign n28630 = n28366 ^ n28347;
  assign n28633 = n28632 ^ n28630;
  assign n28638 = n28637 ^ n28633;
  assign n28628 = n28518 ^ n28247;
  assign n28625 = n28523 ^ n28113;
  assign n28620 = ~n28054 & n28084;
  assign n28621 = n28620 ^ n28108;
  assign n28624 = n28623 ^ n28621;
  assign n28626 = n28625 ^ n28624;
  assign n28627 = n28626 ^ n28119;
  assign n28629 = n28628 ^ n28627;
  assign n28639 = n28638 ^ n28629;
  assign n28232 = n28231 ^ n28230;
  assign n28237 = n28236 ^ n28232;
  assign n28229 = n28228 ^ n28216;
  assign n28238 = n28237 ^ n28229;
  assign n28592 = n28238 ^ n27785;
  assign n28619 = n28618 ^ n28592;
  assign n28640 = n28639 ^ n28619;
  assign n28688 = n28687 ^ n28640;
  assign n28704 = n28618 ^ n28589;
  assign n28705 = n28688 & n28704;
  assign n28734 = n28733 ^ n28705;
  assign n28731 = n28704 ^ n28688;
  assign n28505 = n28504 ^ n27738;
  assign n28485 = n28484 ^ n28475;
  assign n28498 = n28497 ^ n28485;
  assign n28357 = n28356 ^ n28347;
  assign n28370 = n28369 ^ n28357;
  assign n28499 = n28498 ^ n28370;
  assign n28248 = n28247 ^ n28238;
  assign n28109 = n28108 ^ n28105;
  assign n28086 = n28085 ^ n28080;
  assign n28095 = n28094 ^ n28086;
  assign n28110 = n28109 ^ n28095;
  assign n28120 = n28119 ^ n28110;
  assign n28249 = n28248 ^ n28120;
  assign n28500 = n28499 ^ n28249;
  assign n28506 = n28505 ^ n28500;
  assign n28566 = n28565 ^ n28506;
  assign n28591 = n28589 ^ n28506;
  assign n28718 = n28687 ^ n28591;
  assign n28719 = n28566 & n28718;
  assign n28683 = n28662 ^ n28565;
  assign n28684 = n28683 ^ n28640;
  assign n28685 = n28591 & n28684;
  assign n28720 = n28719 ^ n28685;
  assign n28732 = n28731 ^ n28720;
  assign n28735 = n28734 ^ n28732;
  assign n28701 = n28699 ^ n28506;
  assign n28702 = n28701 ^ n28591;
  assign n28700 = n28699 ^ n28688;
  assign n28708 = n28702 ^ n28700;
  assign n28703 = n28700 & n28702;
  assign n28706 = n28705 ^ n28703;
  assign n28641 = n28640 ^ n28591;
  assign n28681 = n28680 ^ n28641;
  assign n28682 = n28590 & n28681;
  assign n28686 = n28685 ^ n28682;
  assign n28707 = n28706 ^ n28686;
  assign n28709 = n28708 ^ n28707;
  assign n28741 = n28735 ^ n28709;
  assign n28717 = n28683 ^ n28641;
  assign n28721 = n28720 ^ n28717;
  assign n28714 = n28704 ^ n28566;
  assign n28715 = n28641 & n28714;
  assign n28712 = n28698 ^ n28641;
  assign n28713 = n28711 & n28712;
  assign n28716 = n28715 ^ n28713;
  assign n28722 = n28721 ^ n28716;
  assign n28736 = n28722 & n28735;
  assign n28742 = n28741 ^ n28736;
  assign n28725 = n28681 ^ n28590;
  assign n28723 = n28698 & n28701;
  assign n28724 = n28723 ^ n28715;
  assign n28726 = n28725 ^ n28724;
  assign n28727 = n28726 ^ n28686;
  assign n28739 = n28727 & n28735;
  assign n28740 = ~n28709 & n28739;
  assign n28743 = n28742 ^ n28740;
  assign n28766 = n28711 & n28743;
  assign n28730 = n28727 ^ n28722;
  assign n28737 = n28736 ^ n28730;
  assign n28728 = n28722 & ~n28727;
  assign n28729 = n28709 & n28728;
  assign n28738 = n28737 ^ n28729;
  assign n28765 = n28699 & n28738;
  assign n28767 = n28766 ^ n28765;
  assign n28748 = n28736 ^ n28727;
  assign n28749 = n28741 & n28748;
  assign n28750 = n28749 ^ n28709;
  assign n28745 = n28736 ^ n28709;
  assign n28746 = n28730 & n28745;
  assign n28747 = n28746 ^ n28727;
  assign n28751 = n28750 ^ n28747;
  assign n28763 = n28684 & n28751;
  assign n28744 = n28743 ^ n28738;
  assign n28752 = n28751 ^ n28744;
  assign n28762 = n28718 & n28752;
  assign n28764 = n28763 ^ n28762;
  assign n28768 = n28767 ^ n28764;
  assign n28759 = n28750 ^ n28743;
  assign n28760 = n28714 & n28759;
  assign n28756 = n28747 ^ n28738;
  assign n28757 = n28688 & n28756;
  assign n28754 = n28591 & n28751;
  assign n28753 = n28566 & n28752;
  assign n28755 = n28754 ^ n28753;
  assign n28758 = n28757 ^ n28755;
  assign n28761 = n28760 ^ n28758;
  assign n28769 = n28768 ^ n28761;
  assign n29021 = n29020 ^ n28769;
  assign n29034 = n29016 ^ n29005;
  assign n29031 = ~n28949 & ~n29009;
  assign n29029 = n28978 & ~n29001;
  assign n29030 = n29029 ^ n29010;
  assign n29032 = n29031 ^ n29030;
  assign n29033 = n29032 ^ n29014;
  assign n29035 = n29034 ^ n29033;
  assign n29036 = n29035 ^ n27801;
  assign n29027 = n28766 ^ n28755;
  assign n29024 = n28641 & n28759;
  assign n29022 = n28712 & n28743;
  assign n29023 = n29022 ^ n28760;
  assign n29025 = n29024 ^ n29023;
  assign n29026 = n29025 ^ n28764;
  assign n29028 = n29027 ^ n29026;
  assign n29037 = n29036 ^ n29028;
  assign n29060 = n29012 ^ n28993;
  assign n29057 = n28948 & n29002;
  assign n29058 = n29057 ^ n27773;
  assign n29054 = ~n28945 & n29006;
  assign n29053 = ~n28950 & n29002;
  assign n29055 = n29054 ^ n29053;
  assign n29051 = ~n28943 & ~n28991;
  assign n29049 = ~n28939 & n28987;
  assign n29050 = n29049 ^ n29031;
  assign n29052 = n29051 ^ n29050;
  assign n29056 = n29055 ^ n29052;
  assign n29059 = n29058 ^ n29056;
  assign n29061 = n29060 ^ n29059;
  assign n29062 = n29061 ^ n28754;
  assign n29046 = n28590 & n28744;
  assign n29044 = n28681 & n28744;
  assign n29043 = n28704 & n28756;
  assign n29045 = n29044 ^ n29043;
  assign n29047 = n29046 ^ n29045;
  assign n29040 = n28702 & n28747;
  assign n29038 = n28698 & n28750;
  assign n29039 = n29038 ^ n29024;
  assign n29041 = n29040 ^ n29039;
  assign n29042 = n29041 ^ n28763;
  assign n29048 = n29047 ^ n29042;
  assign n29063 = n29062 ^ n29048;
  assign n29066 = n29032 ^ n29017;
  assign n29065 = n29008 ^ n27736;
  assign n29067 = n29066 ^ n29065;
  assign n29068 = n29067 ^ n29025;
  assign n29064 = n28767 ^ n28758;
  assign n29069 = n29068 ^ n29064;
  assign n29077 = ~n28941 & ~n28991;
  assign n29078 = n29077 ^ n29049;
  assign n29075 = n29030 ^ n29017;
  assign n29074 = n29005 ^ n27783;
  assign n29076 = n29075 ^ n29074;
  assign n29079 = n29078 ^ n29076;
  assign n29073 = n28700 & n28747;
  assign n29080 = n29079 ^ n29073;
  assign n29071 = n29038 ^ n29023;
  assign n29070 = n28767 ^ n28755;
  assign n29072 = n29071 ^ n29070;
  assign n29081 = n29080 ^ n29072;
  assign n29091 = ~n28942 & n28987;
  assign n29092 = n29091 ^ n29017;
  assign n29088 = n29055 ^ n29013;
  assign n29089 = n29088 ^ n29052;
  assign n29087 = n29008 ^ n27764;
  assign n29090 = n29089 ^ n29087;
  assign n29093 = n29092 ^ n29090;
  assign n29094 = n29093 ^ n28767;
  assign n29084 = n28701 & n28750;
  assign n29085 = n29084 ^ n29041;
  assign n29082 = n29045 ^ n28762;
  assign n29083 = n29082 ^ n28758;
  assign n29086 = n29085 ^ n29083;
  assign n29095 = n29094 ^ n29086;
  assign n29102 = n28976 & ~n28997;
  assign n29103 = n29102 ^ n29077;
  assign n29104 = n29103 ^ n29088;
  assign n29101 = n29015 ^ n29005;
  assign n29105 = n29104 ^ n29101;
  assign n29106 = n29105 ^ n27792;
  assign n29099 = n28765 ^ n28755;
  assign n29096 = n28710 & n28738;
  assign n29097 = n29096 ^ n29073;
  assign n29098 = n29097 ^ n29082;
  assign n29100 = n29099 ^ n29098;
  assign n29107 = n29106 ^ n29100;
  assign n29112 = n29103 ^ n29050;
  assign n29111 = n29054 ^ n29008;
  assign n29113 = n29112 ^ n29111;
  assign n29114 = n29113 ^ n27809;
  assign n29109 = n29097 ^ n29039;
  assign n29108 = n29043 ^ n28758;
  assign n29110 = n29109 ^ n29108;
  assign n29115 = n29114 ^ n29110;
  assign n29893 = n27256 ^ n26384;
  assign n29894 = n29893 ^ n28373;
  assign n29895 = n29894 ^ n28777;
  assign n29889 = n27262 ^ n26409;
  assign n29890 = n29889 ^ n28382;
  assign n29891 = n29890 ^ n28778;
  assign n29884 = n27267 ^ n26432;
  assign n29885 = n29884 ^ n28377;
  assign n29886 = n29885 ^ n28774;
  assign n29892 = n29891 ^ n29886;
  assign n29896 = n29895 ^ n29892;
  assign n29877 = n27275 ^ n26308;
  assign n29878 = n29877 ^ n28411;
  assign n29879 = n29878 ^ n28771;
  assign n29932 = n29896 ^ n29879;
  assign n29881 = n27289 ^ n26214;
  assign n29882 = n29881 ^ n28401;
  assign n29883 = n29882 ^ n28773;
  assign n29870 = n27305 ^ n26364;
  assign n29871 = n29870 ^ n28396;
  assign n29872 = n29871 ^ n28782;
  assign n29904 = n29883 ^ n29872;
  assign n29933 = n29932 ^ n29904;
  assign n29921 = ~n29879 & ~n29896;
  assign n29887 = n29886 ^ n29883;
  assign n29874 = n27282 ^ n26335;
  assign n29875 = n29874 ^ n28417;
  assign n29876 = n29875 ^ n28770;
  assign n29880 = n29879 ^ n29876;
  assign n29888 = n29887 ^ n29880;
  assign n29901 = n29879 ^ n29872;
  assign n29902 = n29888 & n29901;
  assign n29922 = n29921 ^ n29902;
  assign n29919 = n29901 ^ n29888;
  assign n29867 = n27298 ^ n26273;
  assign n29868 = n29867 ^ n28390;
  assign n29869 = n29868 ^ n28785;
  assign n29873 = n29872 ^ n29869;
  assign n29915 = n29887 ^ n29873;
  assign n29916 = n29883 ^ n29869;
  assign n29917 = ~n29915 & n29916;
  assign n29908 = n29891 ^ n29883;
  assign n29909 = n29908 ^ n29880;
  assign n29910 = n29873 & n29909;
  assign n29918 = n29917 ^ n29910;
  assign n29920 = n29919 ^ n29918;
  assign n29923 = n29922 ^ n29920;
  assign n29905 = n29880 ^ n29873;
  assign n29937 = n29908 ^ n29905;
  assign n29938 = n29937 ^ n29918;
  assign n29934 = n29905 ^ n29895;
  assign n29935 = ~n29933 & n29934;
  assign n29926 = n29916 ^ n29901;
  assign n29927 = ~n29905 & n29926;
  assign n29936 = n29935 ^ n29927;
  assign n29939 = n29938 ^ n29936;
  assign n29940 = n29923 & n29939;
  assign n29898 = n29896 ^ n29869;
  assign n29899 = n29898 ^ n29873;
  assign n29897 = n29896 ^ n29888;
  assign n29913 = n29899 ^ n29897;
  assign n29906 = n29905 ^ n29892;
  assign n29907 = n29904 & ~n29906;
  assign n29911 = n29910 ^ n29907;
  assign n29900 = ~n29897 & ~n29899;
  assign n29903 = n29902 ^ n29900;
  assign n29912 = n29911 ^ n29903;
  assign n29914 = n29913 ^ n29912;
  assign n29924 = n29923 ^ n29914;
  assign n29956 = n29940 ^ n29924;
  assign n29929 = n29906 ^ n29904;
  assign n29925 = ~n29895 & ~n29898;
  assign n29928 = n29927 ^ n29925;
  assign n29930 = n29929 ^ n29928;
  assign n29931 = n29930 ^ n29911;
  assign n29954 = n29923 & ~n29931;
  assign n29955 = ~n29914 & n29954;
  assign n29957 = n29956 ^ n29955;
  assign n29972 = ~n29933 & n29957;
  assign n29951 = n29931 & n29939;
  assign n29952 = n29914 & n29951;
  assign n29944 = n29939 ^ n29931;
  assign n29950 = n29944 ^ n29940;
  assign n29953 = n29952 ^ n29950;
  assign n29971 = ~n29896 & ~n29953;
  assign n29973 = n29972 ^ n29971;
  assign n29958 = n29957 ^ n29953;
  assign n29945 = n29940 ^ n29914;
  assign n29946 = ~n29944 & n29945;
  assign n29947 = n29946 ^ n29931;
  assign n29941 = n29940 ^ n29931;
  assign n29942 = n29924 & ~n29941;
  assign n29943 = n29942 ^ n29914;
  assign n29948 = n29947 ^ n29943;
  assign n29959 = n29958 ^ n29948;
  assign n29969 = ~n29915 & n29959;
  assign n29968 = n29909 & ~n29948;
  assign n29970 = n29969 ^ n29968;
  assign n29974 = n29973 ^ n29970;
  assign n29965 = n29957 ^ n29943;
  assign n29966 = n29926 & n29965;
  assign n29962 = n29953 ^ n29947;
  assign n29963 = n29888 & n29962;
  assign n29960 = n29916 & n29959;
  assign n29949 = n29873 & ~n29948;
  assign n29961 = n29960 ^ n29949;
  assign n29964 = n29963 ^ n29961;
  assign n29967 = n29966 ^ n29964;
  assign n29975 = n29974 ^ n29967;
  assign n29976 = n29975 ^ n28873;
  assign n29503 = n25828 ^ n24873;
  assign n29501 = n25029 ^ n24849;
  assign n29502 = n29501 ^ n28403;
  assign n29504 = n29503 ^ n29502;
  assign n29495 = n25933 ^ n24745;
  assign n29493 = n24991 ^ n24367;
  assign n29494 = n29493 ^ n28380;
  assign n29496 = n29495 ^ n29494;
  assign n29525 = n29504 ^ n29496;
  assign n29512 = n25997 ^ n25058;
  assign n29511 = n28415 ^ n25069;
  assign n29513 = n29512 ^ n29511;
  assign n29508 = n25969 ^ n25022;
  assign n29506 = n28408 ^ n25029;
  assign n29507 = n29506 ^ n27159;
  assign n29509 = n29508 ^ n29507;
  assign n29510 = n29509 ^ n28407;
  assign n29514 = n29513 ^ n29510;
  assign n29526 = n29525 ^ n29514;
  assign n29483 = n25903 ^ n24970;
  assign n29481 = n24991 ^ n24962;
  assign n29482 = n29481 ^ n28394;
  assign n29484 = n29483 ^ n29482;
  assign n29479 = n25876 ^ n24921;
  assign n29477 = n28387 ^ n24939;
  assign n29478 = n29477 ^ n27139;
  assign n29480 = n29479 ^ n29478;
  assign n29485 = n29484 ^ n29480;
  assign n29522 = n29514 ^ n29485;
  assign n29491 = n25750 ^ n24730;
  assign n29489 = n24939 ^ n24367;
  assign n29490 = n29489 ^ n27134;
  assign n29492 = n29491 ^ n29490;
  assign n29497 = n29496 ^ n29492;
  assign n29523 = n29522 ^ n29497;
  assign n29521 = n29504 ^ n29484;
  assign n29555 = n29523 ^ n29521;
  assign n29487 = n26023 ^ n24920;
  assign n29486 = n28408 ^ n28371;
  assign n29488 = n29487 ^ n29486;
  assign n29498 = n29497 ^ n29488;
  assign n29499 = n29498 ^ n29480;
  assign n29553 = ~n29488 & ~n29499;
  assign n29533 = n29504 ^ n29480;
  assign n29518 = n29509 ^ n29484;
  assign n29542 = n29533 ^ n29518;
  assign n29543 = ~n29522 & ~n29542;
  assign n29554 = n29553 ^ n29543;
  assign n29556 = n29555 ^ n29554;
  assign n29527 = n29485 & n29526;
  assign n29524 = n29521 & ~n29523;
  assign n29528 = n29527 ^ n29524;
  assign n29557 = n29556 ^ n29528;
  assign n29549 = n29525 ^ n29522;
  assign n29505 = n29504 ^ n29492;
  assign n29534 = n29505 ^ n29485;
  assign n29535 = n29533 & ~n29534;
  assign n29536 = n29535 ^ n29527;
  assign n29550 = n29549 ^ n29536;
  assign n29544 = n29509 ^ n29498;
  assign n29545 = n29544 ^ n29521;
  assign n29546 = n29522 ^ n29488;
  assign n29547 = n29545 & n29546;
  assign n29548 = n29547 ^ n29543;
  assign n29551 = n29550 ^ n29548;
  assign n29561 = n29557 ^ n29551;
  assign n29538 = ~n29498 & n29509;
  assign n29515 = n29514 ^ n29505;
  assign n29519 = n29515 & ~n29518;
  assign n29539 = n29538 ^ n29519;
  assign n29532 = n29518 ^ n29515;
  assign n29537 = n29536 ^ n29532;
  assign n29540 = n29539 ^ n29537;
  assign n29552 = ~n29540 & n29551;
  assign n29516 = n29515 ^ n29498;
  assign n29500 = n29499 ^ n29485;
  assign n29530 = n29516 ^ n29500;
  assign n29517 = ~n29500 & ~n29516;
  assign n29520 = n29519 ^ n29517;
  assign n29529 = n29528 ^ n29520;
  assign n29531 = n29530 ^ n29529;
  assign n29562 = n29552 ^ n29531;
  assign n29563 = ~n29561 & n29562;
  assign n29564 = n29563 ^ n29557;
  assign n29541 = n29540 ^ n29531;
  assign n29558 = n29557 ^ n29552;
  assign n29559 = ~n29541 & ~n29558;
  assign n29560 = n29559 ^ n29531;
  assign n29565 = n29564 ^ n29560;
  assign n29597 = n29526 & ~n29565;
  assign n29573 = n29552 ^ n29541;
  assign n29571 = ~n29540 & ~n29557;
  assign n29572 = ~n29531 & n29571;
  assign n29574 = n29573 ^ n29572;
  assign n29568 = n29551 & n29557;
  assign n29569 = n29531 & n29568;
  assign n29567 = n29561 ^ n29552;
  assign n29570 = n29569 ^ n29567;
  assign n29575 = n29574 ^ n29570;
  assign n29576 = n29575 ^ n29565;
  assign n29596 = ~n29534 & ~n29576;
  assign n29598 = n29597 ^ n29596;
  assign n29580 = n29545 & ~n29574;
  assign n29579 = ~n29498 & ~n29570;
  assign n29581 = n29580 ^ n29579;
  assign n29599 = n29598 ^ n29581;
  assign n29592 = n29570 ^ n29564;
  assign n29593 = n29515 & n29592;
  assign n29577 = n29533 & ~n29576;
  assign n29566 = n29485 & ~n29565;
  assign n29578 = n29577 ^ n29566;
  assign n29594 = n29593 ^ n29578;
  assign n29587 = n29574 ^ n29560;
  assign n29588 = ~n29542 & ~n29587;
  assign n29595 = n29594 ^ n29588;
  assign n29600 = n29599 ^ n29595;
  assign n29792 = n29600 ^ n28939;
  assign n29268 = n24908 ^ n23964;
  assign n29266 = n24096 ^ n23940;
  assign n29265 = n24127 ^ n23923;
  assign n29267 = n29266 ^ n29265;
  assign n29269 = n29268 ^ n29267;
  assign n29237 = n24831 ^ n23997;
  assign n29236 = n27259 ^ n23686;
  assign n29238 = n29237 ^ n29236;
  assign n29283 = n29269 ^ n29238;
  assign n29260 = n28152 ^ n24130;
  assign n29259 = n24122 ^ n23417;
  assign n29261 = n29260 ^ n29259;
  assign n29257 = n25054 ^ n24110;
  assign n29255 = n25045 ^ n24096;
  assign n29253 = n28145 ^ n24088;
  assign n29254 = n29253 ^ n27286;
  assign n29256 = n29255 ^ n29254;
  assign n29258 = n29257 ^ n29256;
  assign n29262 = n29261 ^ n29258;
  assign n29289 = n29283 ^ n29262;
  assign n29240 = n28145 ^ n23561;
  assign n29241 = n29240 ^ n24082;
  assign n29242 = n29241 ^ n24144;
  assign n29243 = n29242 ^ n25098;
  assign n29234 = n25010 ^ n24060;
  assign n29233 = n27302 ^ n24003;
  assign n29235 = n29234 ^ n29233;
  assign n29239 = n29238 ^ n29235;
  assign n29244 = n29243 ^ n29239;
  assign n29308 = n29289 ^ n29244;
  assign n29246 = n24981 ^ n24037;
  assign n29245 = n27253 ^ n24061;
  assign n29247 = n29246 ^ n29245;
  assign n29273 = n29269 ^ n29247;
  assign n29250 = n24955 ^ n23685;
  assign n29248 = n28158 ^ n23562;
  assign n29249 = n29248 ^ n27265;
  assign n29251 = n29250 ^ n29249;
  assign n29252 = n29251 ^ n29247;
  assign n29263 = n29262 ^ n29252;
  assign n29300 = n29263 ^ n29239;
  assign n29303 = n29273 & ~n29300;
  assign n29279 = n29269 ^ n29235;
  assign n29281 = n29279 ^ n29262;
  assign n29282 = n29252 & n29281;
  assign n29304 = n29303 ^ n29282;
  assign n29301 = n29300 ^ n29273;
  assign n29297 = n29251 ^ n29244;
  assign n29298 = ~n29243 & ~n29297;
  assign n29270 = n29269 ^ n29251;
  assign n29264 = n29256 ^ n29247;
  assign n29271 = n29270 ^ n29264;
  assign n29272 = ~n29263 & ~n29271;
  assign n29299 = n29298 ^ n29272;
  assign n29302 = n29301 ^ n29299;
  assign n29305 = n29304 ^ n29302;
  assign n29284 = n29283 ^ n29252;
  assign n29285 = n29270 & ~n29284;
  assign n29286 = n29285 ^ n29282;
  assign n29280 = n29279 ^ n29263;
  assign n29287 = n29286 ^ n29280;
  assign n29274 = n29256 ^ n29244;
  assign n29275 = n29274 ^ n29273;
  assign n29276 = n29263 ^ n29243;
  assign n29277 = n29275 & n29276;
  assign n29278 = n29277 ^ n29272;
  assign n29288 = n29287 ^ n29278;
  assign n29306 = n29305 ^ n29288;
  assign n29309 = n29297 ^ n29252;
  assign n29313 = n29309 ^ n29308;
  assign n29310 = ~n29308 & ~n29309;
  assign n29293 = ~n29264 & n29289;
  assign n29311 = n29310 ^ n29293;
  assign n29312 = n29311 ^ n29304;
  assign n29314 = n29313 ^ n29312;
  assign n29292 = ~n29244 & n29256;
  assign n29294 = n29293 ^ n29292;
  assign n29290 = n29289 ^ n29264;
  assign n29291 = n29290 ^ n29286;
  assign n29295 = n29294 ^ n29291;
  assign n29296 = n29288 & ~n29295;
  assign n29336 = n29314 ^ n29296;
  assign n29337 = ~n29306 & n29336;
  assign n29338 = n29337 ^ n29305;
  assign n29697 = ~n29308 & ~n29338;
  assign n29315 = n29288 & n29305;
  assign n29316 = n29314 & n29315;
  assign n29307 = n29306 ^ n29296;
  assign n29317 = n29316 ^ n29307;
  assign n29696 = n29274 & ~n29317;
  assign n29698 = n29697 ^ n29696;
  assign n29321 = n29314 ^ n29295;
  assign n29326 = n29305 ^ n29296;
  assign n29327 = ~n29321 & ~n29326;
  assign n29328 = n29327 ^ n29314;
  assign n29627 = ~n29243 & n29328;
  assign n29322 = n29321 ^ n29296;
  assign n29319 = ~n29295 & ~n29305;
  assign n29320 = ~n29314 & n29319;
  assign n29323 = n29322 ^ n29320;
  assign n29329 = n29328 ^ n29323;
  assign n29333 = ~n29263 & ~n29329;
  assign n29628 = n29627 ^ n29333;
  assign n29788 = n29698 ^ n29628;
  assign n29345 = n29338 ^ n29317;
  assign n29620 = ~n29264 & n29345;
  assign n29346 = n29289 & n29345;
  assign n29341 = n29323 ^ n29317;
  assign n29339 = n29338 ^ n29328;
  assign n29342 = n29341 ^ n29339;
  assign n29343 = n29270 & ~n29342;
  assign n29340 = n29252 & ~n29339;
  assign n29344 = n29343 ^ n29340;
  assign n29347 = n29346 ^ n29344;
  assign n29787 = n29620 ^ n29347;
  assign n29789 = n29788 ^ n29787;
  assign n29150 = n23178 ^ n22878;
  assign n29151 = n29150 ^ n20100;
  assign n29152 = n29151 ^ n23195;
  assign n29153 = n29152 ^ n23982;
  assign n29120 = n27994 ^ n23144;
  assign n29121 = n29120 ^ n24017;
  assign n29122 = n29121 ^ n23067;
  assign n29167 = n29153 ^ n29122;
  assign n29145 = n28012 ^ n23167;
  assign n29144 = n23190 ^ n23053;
  assign n29146 = n29145 ^ n29144;
  assign n29142 = n24115 ^ n23201;
  assign n29140 = n24103 ^ n23182;
  assign n29138 = n28005 ^ n23177;
  assign n29137 = n23169 ^ n21946;
  assign n29139 = n29138 ^ n29137;
  assign n29141 = n29140 ^ n29139;
  assign n29143 = n29142 ^ n29141;
  assign n29147 = n29146 ^ n29143;
  assign n29173 = n29167 ^ n29147;
  assign n29126 = n24153 ^ n23127;
  assign n29124 = n23172 ^ n23047;
  assign n29125 = n29124 ^ n28005;
  assign n29127 = n29126 ^ n29125;
  assign n29118 = n24070 ^ n23153;
  assign n29116 = n23089 ^ n23003;
  assign n29117 = n29116 ^ n23148;
  assign n29119 = n29118 ^ n29117;
  assign n29123 = n29122 ^ n29119;
  assign n29128 = n29127 ^ n29123;
  assign n29192 = n29173 ^ n29128;
  assign n29129 = n23149 ^ n23058;
  assign n29130 = n29129 ^ n27990;
  assign n29131 = n29130 ^ n24042;
  assign n29157 = n29153 ^ n29131;
  assign n29132 = n28031 ^ n27998;
  assign n29133 = n29132 ^ n23048;
  assign n29134 = n29133 ^ n23015;
  assign n29135 = n29134 ^ n23907;
  assign n29136 = n29135 ^ n29131;
  assign n29148 = n29147 ^ n29136;
  assign n29184 = n29148 ^ n29123;
  assign n29187 = n29157 & ~n29184;
  assign n29163 = n29153 ^ n29119;
  assign n29165 = n29163 ^ n29147;
  assign n29166 = n29136 & n29165;
  assign n29188 = n29187 ^ n29166;
  assign n29185 = n29184 ^ n29157;
  assign n29181 = n29135 ^ n29128;
  assign n29182 = ~n29127 & ~n29181;
  assign n29154 = n29153 ^ n29135;
  assign n29149 = n29141 ^ n29131;
  assign n29155 = n29154 ^ n29149;
  assign n29156 = ~n29148 & ~n29155;
  assign n29183 = n29182 ^ n29156;
  assign n29186 = n29185 ^ n29183;
  assign n29189 = n29188 ^ n29186;
  assign n29168 = n29167 ^ n29136;
  assign n29169 = n29154 & ~n29168;
  assign n29170 = n29169 ^ n29166;
  assign n29164 = n29163 ^ n29148;
  assign n29171 = n29170 ^ n29164;
  assign n29158 = n29141 ^ n29128;
  assign n29159 = n29158 ^ n29157;
  assign n29160 = n29148 ^ n29127;
  assign n29161 = n29159 & n29160;
  assign n29162 = n29161 ^ n29156;
  assign n29172 = n29171 ^ n29162;
  assign n29190 = n29189 ^ n29172;
  assign n29193 = n29181 ^ n29136;
  assign n29197 = n29193 ^ n29192;
  assign n29194 = ~n29192 & ~n29193;
  assign n29177 = ~n29149 & n29173;
  assign n29195 = n29194 ^ n29177;
  assign n29196 = n29195 ^ n29188;
  assign n29198 = n29197 ^ n29196;
  assign n29176 = ~n29128 & n29141;
  assign n29178 = n29177 ^ n29176;
  assign n29174 = n29173 ^ n29149;
  assign n29175 = n29174 ^ n29170;
  assign n29179 = n29178 ^ n29175;
  assign n29180 = n29172 & ~n29179;
  assign n29220 = n29198 ^ n29180;
  assign n29221 = ~n29190 & n29220;
  assign n29222 = n29221 ^ n29189;
  assign n29691 = ~n29192 & ~n29222;
  assign n29199 = n29172 & n29189;
  assign n29200 = n29198 & n29199;
  assign n29191 = n29190 ^ n29180;
  assign n29201 = n29200 ^ n29191;
  assign n29690 = n29158 & ~n29201;
  assign n29692 = n29691 ^ n29690;
  assign n29205 = n29198 ^ n29179;
  assign n29210 = n29189 ^ n29180;
  assign n29211 = ~n29205 & ~n29210;
  assign n29212 = n29211 ^ n29198;
  assign n29613 = ~n29127 & n29212;
  assign n29206 = n29205 ^ n29180;
  assign n29203 = ~n29179 & ~n29189;
  assign n29204 = ~n29198 & n29203;
  assign n29207 = n29206 ^ n29204;
  assign n29213 = n29212 ^ n29207;
  assign n29217 = ~n29148 & ~n29213;
  assign n29614 = n29613 ^ n29217;
  assign n29785 = n29692 ^ n29614;
  assign n29229 = n29222 ^ n29201;
  assign n29606 = ~n29149 & n29229;
  assign n29230 = n29173 & n29229;
  assign n29225 = n29207 ^ n29201;
  assign n29223 = n29222 ^ n29212;
  assign n29226 = n29225 ^ n29223;
  assign n29227 = n29154 & ~n29226;
  assign n29224 = n29136 & ~n29223;
  assign n29228 = n29227 ^ n29224;
  assign n29231 = n29230 ^ n29228;
  assign n29784 = n29606 ^ n29231;
  assign n29786 = n29785 ^ n29784;
  assign n29790 = n29789 ^ n29786;
  assign n29377 = n28771 ^ n25810;
  assign n29375 = n28274 ^ n25941;
  assign n29376 = n29375 ^ n25955;
  assign n29378 = n29377 ^ n29376;
  assign n29358 = n28777 ^ n25959;
  assign n29357 = n26983 ^ n26016;
  assign n29359 = n29358 ^ n29357;
  assign n29354 = n28774 ^ n25927;
  assign n29353 = n26979 ^ n25412;
  assign n29355 = n29354 ^ n29353;
  assign n29351 = n28778 ^ n25896;
  assign n29350 = n27020 ^ n25917;
  assign n29352 = n29351 ^ n29350;
  assign n29356 = n29355 ^ n29352;
  assign n29360 = n29359 ^ n29356;
  assign n29404 = n29378 ^ n29360;
  assign n29381 = n28770 ^ n25866;
  assign n29380 = n28282 ^ n25983;
  assign n29382 = n29381 ^ n29380;
  assign n29379 = n29378 ^ n25981;
  assign n29383 = n29382 ^ n29379;
  assign n29367 = n28782 ^ n25861;
  assign n29366 = n27015 ^ n25888;
  assign n29368 = n29367 ^ n29366;
  assign n29363 = n28785 ^ n25663;
  assign n29361 = n28263 ^ n25841;
  assign n29362 = n29361 ^ n25855;
  assign n29364 = n29363 ^ n29362;
  assign n29369 = n29368 ^ n29364;
  assign n29391 = n29383 ^ n29369;
  assign n29392 = n29391 ^ n29356;
  assign n29372 = n28773 ^ n25989;
  assign n29371 = n26992 ^ n25798;
  assign n29373 = n29372 ^ n29371;
  assign n29390 = n29373 ^ n29368;
  assign n29417 = n29392 ^ n29390;
  assign n29365 = n29364 ^ n29360;
  assign n29415 = ~n29359 & ~n29365;
  assign n29401 = n29373 ^ n29364;
  assign n29387 = n29378 ^ n29368;
  assign n29402 = n29401 ^ n29387;
  assign n29403 = ~n29391 & n29402;
  assign n29416 = n29415 ^ n29403;
  assign n29418 = n29417 ^ n29416;
  assign n29394 = n29373 ^ n29352;
  assign n29395 = n29394 ^ n29383;
  assign n29396 = ~n29369 & ~n29395;
  assign n29393 = ~n29390 & ~n29392;
  assign n29397 = n29396 ^ n29393;
  assign n29419 = n29418 ^ n29397;
  assign n29412 = n29394 ^ n29391;
  assign n29374 = n29373 ^ n29355;
  assign n29409 = n29374 ^ n29369;
  assign n29410 = n29401 & n29409;
  assign n29411 = n29410 ^ n29396;
  assign n29413 = n29412 ^ n29411;
  assign n29405 = n29404 ^ n29390;
  assign n29406 = n29391 ^ n29359;
  assign n29407 = ~n29405 & n29406;
  assign n29408 = n29407 ^ n29403;
  assign n29414 = n29413 ^ n29408;
  assign n29428 = n29419 ^ n29414;
  assign n29424 = ~n29360 & n29378;
  assign n29384 = n29383 ^ n29374;
  assign n29388 = ~n29384 & n29387;
  assign n29425 = n29424 ^ n29388;
  assign n29422 = n29387 ^ n29384;
  assign n29423 = n29422 ^ n29411;
  assign n29426 = n29425 ^ n29423;
  assign n29427 = n29414 & ~n29426;
  assign n29429 = n29428 ^ n29427;
  assign n29385 = n29384 ^ n29360;
  assign n29370 = n29369 ^ n29365;
  assign n29399 = n29385 ^ n29370;
  assign n29386 = n29370 & n29385;
  assign n29389 = n29388 ^ n29386;
  assign n29398 = n29397 ^ n29389;
  assign n29400 = n29399 ^ n29398;
  assign n29420 = n29414 & ~n29419;
  assign n29421 = n29400 & n29420;
  assign n29430 = n29429 ^ n29421;
  assign n29645 = n29404 & n29430;
  assign n29443 = n29427 ^ n29400;
  assign n29444 = n29428 & n29443;
  assign n29445 = n29444 ^ n29419;
  assign n29453 = n29385 & n29445;
  assign n29646 = n29645 ^ n29453;
  assign n29434 = n29426 ^ n29400;
  assign n29440 = n29427 ^ n29419;
  assign n29441 = ~n29434 & n29440;
  assign n29442 = n29441 ^ n29400;
  assign n29435 = n29434 ^ n29427;
  assign n29432 = n29419 & ~n29426;
  assign n29433 = ~n29400 & n29432;
  assign n29436 = n29435 ^ n29433;
  assign n29456 = n29442 ^ n29436;
  assign n29471 = ~n29391 & ~n29456;
  assign n29452 = ~n29359 & n29442;
  assign n29641 = n29471 ^ n29452;
  assign n29703 = n29646 ^ n29641;
  assign n29461 = n29445 ^ n29430;
  assign n29634 = n29387 & n29461;
  assign n29462 = ~n29384 & n29461;
  assign n29446 = n29445 ^ n29442;
  assign n29449 = ~n29369 & n29446;
  assign n29439 = n29436 ^ n29430;
  assign n29447 = n29446 ^ n29439;
  assign n29448 = n29401 & ~n29447;
  assign n29450 = n29449 ^ n29448;
  assign n29463 = n29462 ^ n29450;
  assign n29702 = n29634 ^ n29463;
  assign n29704 = n29703 ^ n29702;
  assign n29466 = ~n29395 & n29446;
  assign n29465 = n29409 & ~n29447;
  assign n29467 = n29466 ^ n29465;
  assign n29437 = ~n29405 & ~n29436;
  assign n29431 = ~n29360 & n29430;
  assign n29438 = n29437 ^ n29431;
  assign n29468 = n29467 ^ n29438;
  assign n29457 = n29402 & ~n29456;
  assign n29464 = n29463 ^ n29457;
  assign n29469 = n29468 ^ n29464;
  assign n29705 = n29704 ^ n29469;
  assign n29791 = n29790 ^ n29705;
  assign n29793 = n29792 ^ n29791;
  assign n29680 = ~n29522 & ~n29587;
  assign n29586 = n29546 & ~n29574;
  assign n29589 = n29588 ^ n29586;
  assign n29681 = n29680 ^ n29589;
  assign n29773 = n29681 ^ n29581;
  assign n29774 = n29773 ^ n29594;
  assign n29775 = n29774 ^ n28903;
  assign n29748 = ~n29390 & ~n29439;
  assign n29633 = ~n29392 & ~n29439;
  assign n29635 = n29634 ^ n29633;
  assign n29749 = n29748 ^ n29635;
  assign n29746 = n29466 ^ n29449;
  assign n29640 = n29370 & n29445;
  assign n29642 = n29641 ^ n29640;
  assign n29747 = n29746 ^ n29642;
  assign n29750 = n29749 ^ n29747;
  assign n29455 = n29406 & ~n29436;
  assign n29458 = n29457 ^ n29455;
  assign n29472 = n29471 ^ n29458;
  assign n29473 = n29472 ^ n29438;
  assign n29474 = n29473 ^ n29463;
  assign n29771 = n29750 ^ n29474;
  assign n29767 = n29273 & n29341;
  assign n29619 = ~n29300 & n29341;
  assign n29621 = n29620 ^ n29619;
  assign n29768 = n29767 ^ n29621;
  assign n29670 = n29281 & ~n29339;
  assign n29765 = n29670 ^ n29340;
  assign n29626 = ~n29309 & ~n29338;
  assign n29629 = n29628 ^ n29626;
  assign n29766 = n29765 ^ n29629;
  assign n29769 = n29768 ^ n29766;
  assign n29762 = n29157 & n29225;
  assign n29605 = ~n29184 & n29225;
  assign n29607 = n29606 ^ n29605;
  assign n29763 = n29762 ^ n29607;
  assign n29665 = n29165 & ~n29223;
  assign n29760 = n29665 ^ n29224;
  assign n29612 = ~n29193 & ~n29222;
  assign n29615 = n29614 ^ n29612;
  assign n29761 = n29760 ^ n29615;
  assign n29764 = n29763 ^ n29761;
  assign n29770 = n29769 ^ n29764;
  assign n29772 = n29771 ^ n29770;
  assign n29776 = n29775 ^ n29772;
  assign n29755 = n29521 & n29575;
  assign n29654 = ~n29518 & n29592;
  assign n29653 = ~n29523 & n29575;
  assign n29655 = n29654 ^ n29653;
  assign n29756 = n29755 ^ n29655;
  assign n29753 = n29597 ^ n29566;
  assign n29728 = ~n29500 & ~n29564;
  assign n29584 = ~n29488 & n29560;
  assign n29709 = n29680 ^ n29584;
  assign n29729 = n29728 ^ n29709;
  assign n29754 = n29753 ^ n29729;
  assign n29757 = n29756 ^ n29754;
  assign n29758 = n29757 ^ n28931;
  assign n29676 = n29450 ^ n29437;
  assign n29675 = n29472 ^ n29467;
  assign n29677 = n29676 ^ n29675;
  assign n29751 = n29750 ^ n29677;
  assign n29324 = n29275 & ~n29323;
  assign n29743 = n29344 ^ n29324;
  assign n29618 = ~n29284 & ~n29342;
  assign n29671 = n29670 ^ n29618;
  assign n29331 = n29276 & ~n29323;
  assign n29330 = ~n29271 & ~n29329;
  assign n29332 = n29331 ^ n29330;
  assign n29334 = n29333 ^ n29332;
  assign n29742 = n29671 ^ n29334;
  assign n29744 = n29743 ^ n29742;
  assign n29208 = n29159 & ~n29207;
  assign n29740 = n29228 ^ n29208;
  assign n29604 = ~n29168 & ~n29226;
  assign n29666 = n29665 ^ n29604;
  assign n29215 = n29160 & ~n29207;
  assign n29214 = ~n29155 & ~n29213;
  assign n29216 = n29215 ^ n29214;
  assign n29218 = n29217 ^ n29216;
  assign n29739 = n29666 ^ n29218;
  assign n29741 = n29740 ^ n29739;
  assign n29745 = n29744 ^ n29741;
  assign n29752 = n29751 ^ n29745;
  assign n29759 = n29758 ^ n29752;
  assign n29777 = n29776 ^ n29759;
  assign n29794 = n29793 ^ n29777;
  assign n29657 = n29544 & ~n29570;
  assign n29583 = ~n29516 & ~n29564;
  assign n29658 = n29657 ^ n29583;
  assign n29656 = n29655 ^ n29596;
  assign n29659 = n29658 ^ n29656;
  assign n29652 = n29579 ^ n29578;
  assign n29660 = n29659 ^ n29652;
  assign n29661 = n29660 ^ n28894;
  assign n29648 = n29450 ^ n29431;
  assign n29636 = n29635 ^ n29465;
  assign n29647 = n29646 ^ n29636;
  assign n29649 = n29648 ^ n29647;
  assign n29638 = ~n29365 & n29442;
  assign n29639 = n29638 ^ n29438;
  assign n29643 = n29642 ^ n29639;
  assign n29637 = n29636 ^ n29463;
  assign n29644 = n29643 ^ n29637;
  assign n29650 = n29649 ^ n29644;
  assign n29624 = ~n29297 & n29328;
  assign n29318 = ~n29244 & ~n29317;
  assign n29325 = n29324 ^ n29318;
  assign n29625 = n29624 ^ n29325;
  assign n29630 = n29629 ^ n29625;
  assign n29622 = n29621 ^ n29618;
  assign n29623 = n29622 ^ n29347;
  assign n29631 = n29630 ^ n29623;
  assign n29610 = ~n29181 & n29212;
  assign n29202 = ~n29128 & ~n29201;
  assign n29209 = n29208 ^ n29202;
  assign n29611 = n29610 ^ n29209;
  assign n29616 = n29615 ^ n29611;
  assign n29608 = n29607 ^ n29604;
  assign n29609 = n29608 ^ n29231;
  assign n29617 = n29616 ^ n29609;
  assign n29632 = n29631 ^ n29617;
  assign n29651 = n29650 ^ n29632;
  assign n29662 = n29661 ^ n29651;
  assign n29780 = n29759 ^ n29662;
  assign n29734 = n29644 ^ n29469;
  assign n29454 = n29453 ^ n29452;
  assign n29459 = n29458 ^ n29454;
  assign n29451 = n29450 ^ n29438;
  assign n29460 = n29459 ^ n29451;
  assign n29735 = n29734 ^ n29460;
  assign n29726 = ~n29499 & n29560;
  assign n29727 = n29726 ^ n29581;
  assign n29730 = n29729 ^ n29727;
  assign n29725 = n29656 ^ n29594;
  assign n29731 = n29730 ^ n29725;
  assign n29732 = n29731 ^ n29600;
  assign n29733 = n29732 ^ n28913;
  assign n29736 = n29735 ^ n29733;
  assign n29720 = n29697 ^ n29627;
  assign n29721 = n29720 ^ n29332;
  assign n29719 = n29344 ^ n29325;
  assign n29722 = n29721 ^ n29719;
  assign n29716 = n29691 ^ n29613;
  assign n29717 = n29716 ^ n29216;
  assign n29715 = n29228 ^ n29209;
  assign n29718 = n29717 ^ n29715;
  assign n29723 = n29722 ^ n29718;
  assign n29710 = n29709 ^ n29658;
  assign n29708 = n29654 ^ n29594;
  assign n29711 = n29710 ^ n29708;
  assign n29712 = n29711 ^ n29600;
  assign n29713 = n29712 ^ n28922;
  assign n29706 = n29705 ^ n29649;
  assign n29699 = n29698 ^ n29622;
  assign n29695 = n29344 ^ n29318;
  assign n29700 = n29699 ^ n29695;
  assign n29693 = n29692 ^ n29608;
  assign n29689 = n29228 ^ n29202;
  assign n29694 = n29693 ^ n29689;
  assign n29701 = n29700 ^ n29694;
  assign n29707 = n29706 ^ n29701;
  assign n29714 = n29713 ^ n29707;
  assign n29724 = n29723 ^ n29714;
  assign n29737 = n29736 ^ n29724;
  assign n29683 = n29580 ^ n29578;
  assign n29682 = n29681 ^ n29598;
  assign n29684 = n29683 ^ n29682;
  assign n29685 = n29684 ^ n28876;
  assign n29678 = n29677 ^ n29469;
  assign n29672 = n29671 ^ n29325;
  assign n29669 = n29347 ^ n29330;
  assign n29673 = n29672 ^ n29669;
  assign n29667 = n29666 ^ n29209;
  assign n29664 = n29231 ^ n29214;
  assign n29668 = n29667 ^ n29664;
  assign n29674 = n29673 ^ n29668;
  assign n29679 = n29678 ^ n29674;
  assign n29686 = n29685 ^ n29679;
  assign n29585 = n29584 ^ n29583;
  assign n29590 = n29589 ^ n29585;
  assign n29582 = n29581 ^ n29578;
  assign n29591 = n29590 ^ n29582;
  assign n29601 = n29600 ^ n29591;
  assign n29602 = n29601 ^ n28866;
  assign n29470 = n29469 ^ n29460;
  assign n29475 = n29474 ^ n29470;
  assign n29335 = n29334 ^ n29325;
  assign n29348 = n29347 ^ n29335;
  assign n29219 = n29218 ^ n29209;
  assign n29232 = n29231 ^ n29219;
  assign n29349 = n29348 ^ n29232;
  assign n29476 = n29475 ^ n29349;
  assign n29603 = n29602 ^ n29476;
  assign n29688 = n29686 ^ n29603;
  assign n29738 = n29737 ^ n29688;
  assign n29830 = n29780 ^ n29738;
  assign n29663 = n29662 ^ n29603;
  assign n29804 = n29776 ^ n29662;
  assign n29807 = n29804 ^ n29688;
  assign n29808 = n29663 & n29807;
  assign n29781 = n29780 ^ n29737;
  assign n29782 = n29688 & n29781;
  assign n29809 = n29808 ^ n29782;
  assign n29831 = n29830 ^ n29809;
  assign n29825 = n29794 ^ n29714;
  assign n29687 = n29686 ^ n29662;
  assign n29826 = n29825 ^ n29687;
  assign n29827 = n29793 ^ n29738;
  assign n29828 = n29826 & n29827;
  assign n29797 = n29714 ^ n29686;
  assign n29798 = n29797 ^ n29663;
  assign n29799 = n29738 & n29798;
  assign n29829 = n29828 ^ n29799;
  assign n29832 = n29831 ^ n29829;
  assign n29778 = n29777 ^ n29738;
  assign n29801 = n29778 ^ n29687;
  assign n29795 = n29794 ^ n29603;
  assign n29796 = n29793 & n29795;
  assign n29800 = n29799 ^ n29796;
  assign n29802 = n29801 ^ n29800;
  assign n29779 = n29687 & n29778;
  assign n29783 = n29782 ^ n29779;
  assign n29803 = n29802 ^ n29783;
  assign n29838 = n29832 ^ n29803;
  assign n29812 = ~n29714 & n29794;
  assign n29805 = n29804 ^ n29737;
  assign n29811 = n29797 & n29805;
  assign n29813 = n29812 ^ n29811;
  assign n29806 = n29805 ^ n29797;
  assign n29810 = n29809 ^ n29806;
  assign n29814 = n29813 ^ n29810;
  assign n29833 = n29814 & n29832;
  assign n29839 = n29838 ^ n29833;
  assign n29816 = n29795 ^ n29688;
  assign n29815 = n29805 ^ n29794;
  assign n29820 = n29816 ^ n29815;
  assign n29817 = n29815 & n29816;
  assign n29818 = n29817 ^ n29811;
  assign n29819 = n29818 ^ n29783;
  assign n29821 = n29820 ^ n29819;
  assign n29836 = n29821 & n29832;
  assign n29837 = ~n29803 & n29836;
  assign n29840 = n29839 ^ n29837;
  assign n29863 = n29794 & n29840;
  assign n29822 = n29821 ^ n29814;
  assign n29834 = n29833 ^ n29822;
  assign n29823 = n29814 & n29822;
  assign n29824 = n29803 & n29823;
  assign n29835 = n29834 ^ n29824;
  assign n29862 = n29826 & n29835;
  assign n29864 = n29863 ^ n29862;
  assign n29845 = n29833 ^ n29803;
  assign n29846 = n29822 & n29845;
  assign n29847 = n29846 ^ n29821;
  assign n29842 = n29833 ^ n29821;
  assign n29843 = n29838 & n29842;
  assign n29844 = n29843 ^ n29803;
  assign n29848 = n29847 ^ n29844;
  assign n29860 = n29781 & n29848;
  assign n29841 = n29840 ^ n29835;
  assign n29849 = n29848 ^ n29841;
  assign n29859 = n29807 & n29849;
  assign n29861 = n29860 ^ n29859;
  assign n29865 = n29864 ^ n29861;
  assign n29856 = n29847 ^ n29835;
  assign n29857 = n29798 & n29856;
  assign n29853 = n29844 ^ n29840;
  assign n29854 = n29805 & n29853;
  assign n29851 = n29688 & n29848;
  assign n29850 = n29663 & n29849;
  assign n29852 = n29851 ^ n29850;
  assign n29855 = n29854 ^ n29852;
  assign n29858 = n29857 ^ n29855;
  assign n29866 = n29865 ^ n29858;
  assign n29977 = n29976 ^ n29866;
  assign n29990 = n29972 ^ n29961;
  assign n29987 = ~n29905 & n29965;
  assign n29985 = n29934 & n29957;
  assign n29986 = n29985 ^ n29966;
  assign n29988 = n29987 ^ n29986;
  assign n29989 = n29988 ^ n29970;
  assign n29991 = n29990 ^ n29989;
  assign n29992 = n29991 ^ n28928;
  assign n29983 = n29862 ^ n29852;
  assign n29980 = n29738 & n29856;
  assign n29978 = n29827 & n29835;
  assign n29979 = n29978 ^ n29857;
  assign n29981 = n29980 ^ n29979;
  assign n29982 = n29981 ^ n29861;
  assign n29984 = n29983 ^ n29982;
  assign n29993 = n29992 ^ n29984;
  assign n30016 = n29968 ^ n29949;
  assign n30013 = n29904 & ~n29958;
  assign n30014 = n30013 ^ n28900;
  assign n30010 = n29901 & n29962;
  assign n30009 = ~n29906 & ~n29958;
  assign n30011 = n30010 ^ n30009;
  assign n30007 = ~n29899 & ~n29947;
  assign n30005 = ~n29895 & n29943;
  assign n30006 = n30005 ^ n29987;
  assign n30008 = n30007 ^ n30006;
  assign n30012 = n30011 ^ n30008;
  assign n30015 = n30014 ^ n30012;
  assign n30017 = n30016 ^ n30015;
  assign n30018 = n30017 ^ n29851;
  assign n30002 = n29687 & n29841;
  assign n30000 = n29797 & n29853;
  assign n29999 = n29778 & n29841;
  assign n30001 = n30000 ^ n29999;
  assign n30003 = n30002 ^ n30001;
  assign n29996 = n29816 & n29844;
  assign n29994 = n29793 & n29847;
  assign n29995 = n29994 ^ n29980;
  assign n29997 = n29996 ^ n29995;
  assign n29998 = n29997 ^ n29860;
  assign n30004 = n30003 ^ n29998;
  assign n30019 = n30018 ^ n30004;
  assign n30022 = n29988 ^ n29973;
  assign n30021 = n29964 ^ n28863;
  assign n30023 = n30022 ^ n30021;
  assign n30024 = n30023 ^ n29981;
  assign n30020 = n29864 ^ n29855;
  assign n30025 = n30024 ^ n30020;
  assign n30033 = ~n29897 & ~n29947;
  assign n30034 = n30033 ^ n30005;
  assign n30031 = n29986 ^ n29973;
  assign n30030 = n29961 ^ n28910;
  assign n30032 = n30031 ^ n30030;
  assign n30035 = n30034 ^ n30032;
  assign n30029 = n29815 & n29844;
  assign n30036 = n30035 ^ n30029;
  assign n30027 = n29994 ^ n29979;
  assign n30026 = n29864 ^ n29852;
  assign n30028 = n30027 ^ n30026;
  assign n30037 = n30036 ^ n30028;
  assign n30047 = ~n29898 & n29943;
  assign n30048 = n30047 ^ n29973;
  assign n30044 = n30011 ^ n29969;
  assign n30045 = n30044 ^ n30008;
  assign n30043 = n29964 ^ n28891;
  assign n30046 = n30045 ^ n30043;
  assign n30049 = n30048 ^ n30046;
  assign n30050 = n30049 ^ n29864;
  assign n30040 = n29795 & n29847;
  assign n30041 = n30040 ^ n29997;
  assign n30038 = n30001 ^ n29859;
  assign n30039 = n30038 ^ n29855;
  assign n30042 = n30041 ^ n30039;
  assign n30051 = n30050 ^ n30042;
  assign n30058 = ~n29932 & ~n29953;
  assign n30059 = n30058 ^ n30033;
  assign n30060 = n30059 ^ n30044;
  assign n30057 = n29971 ^ n29961;
  assign n30061 = n30060 ^ n30057;
  assign n30062 = n30061 ^ n28919;
  assign n30055 = n29863 ^ n29852;
  assign n30052 = n29825 & n29840;
  assign n30053 = n30052 ^ n30029;
  assign n30054 = n30053 ^ n30038;
  assign n30056 = n30055 ^ n30054;
  assign n30063 = n30062 ^ n30056;
  assign n30068 = n30059 ^ n30006;
  assign n30067 = n30010 ^ n29964;
  assign n30069 = n30068 ^ n30067;
  assign n30070 = n30069 ^ n28936;
  assign n30065 = n30053 ^ n29995;
  assign n30064 = n30000 ^ n29855;
  assign n30066 = n30065 ^ n30064;
  assign n30071 = n30070 ^ n30066;
  assign n30196 = n29870 ^ n26763;
  assign n30119 = n27461 ^ n27250;
  assign n30118 = n27481 ^ n27475;
  assign n30120 = n30119 ^ n30118;
  assign n30117 = n29893 ^ n27570;
  assign n30121 = n30120 ^ n30117;
  assign n30107 = n27541 ^ n27385;
  assign n30108 = n30107 ^ n27554;
  assign n30106 = n29884 ^ n27527;
  assign n30109 = n30108 ^ n30106;
  assign n30103 = n27553 ^ n27538;
  assign n30104 = n30103 ^ n27456;
  assign n30102 = n29889 ^ n27547;
  assign n30105 = n30104 ^ n30102;
  assign n30110 = n30109 ^ n30105;
  assign n30122 = n30121 ^ n30110;
  assign n30085 = n27488 ^ n27419;
  assign n30084 = n27513 ^ n27429;
  assign n30086 = n30085 ^ n30084;
  assign n30083 = n29881 ^ n27401;
  assign n30087 = n30086 ^ n30083;
  assign n30113 = n30105 ^ n30087;
  assign n30097 = n27461 ^ n27444;
  assign n30098 = n30097 ^ n27514;
  assign n30096 = n29874 ^ n27502;
  assign n30099 = n30098 ^ n30096;
  assign n30094 = n27241 ^ n27110;
  assign n30092 = n29877 ^ n27496;
  assign n30089 = n27574 ^ n27461;
  assign n30090 = n30089 ^ n27482;
  assign n30091 = n30090 ^ n27420;
  assign n30093 = n30092 ^ n30091;
  assign n30095 = n30094 ^ n30093;
  assign n30100 = n30099 ^ n30095;
  assign n30078 = n27518 ^ n27461;
  assign n30079 = n30078 ^ n27251;
  assign n30080 = n30079 ^ n27542;
  assign n30077 = n29867 ^ n26976;
  assign n30081 = n30080 ^ n30077;
  assign n30074 = n27558 ^ n27452;
  assign n30073 = n27250 ^ n27116;
  assign n30075 = n30074 ^ n30073;
  assign n30072 = n29870 ^ n27468;
  assign n30076 = n30075 ^ n30072;
  assign n30082 = n30081 ^ n30076;
  assign n30101 = n30100 ^ n30082;
  assign n30142 = n30113 ^ n30101;
  assign n30126 = n30087 ^ n30081;
  assign n30138 = n30109 ^ n30087;
  assign n30139 = n30138 ^ n30082;
  assign n30140 = ~n30126 & ~n30139;
  assign n30114 = n30113 ^ n30100;
  assign n30115 = n30082 & n30114;
  assign n30141 = n30140 ^ n30115;
  assign n30143 = n30142 ^ n30141;
  assign n30133 = n30121 ^ n30101;
  assign n30134 = n30122 ^ n30093;
  assign n30088 = n30087 ^ n30076;
  assign n30135 = n30134 ^ n30088;
  assign n30136 = n30133 & ~n30135;
  assign n30125 = n30093 ^ n30076;
  assign n30127 = n30126 ^ n30125;
  assign n30128 = n30101 & n30127;
  assign n30137 = n30136 ^ n30128;
  assign n30144 = n30143 ^ n30137;
  assign n30157 = n30093 & ~n30122;
  assign n30146 = n30138 ^ n30100;
  assign n30150 = ~n30125 & ~n30146;
  assign n30158 = n30157 ^ n30150;
  assign n30155 = n30146 ^ n30125;
  assign n30156 = n30155 ^ n30141;
  assign n30159 = n30158 ^ n30156;
  assign n30160 = n30144 & n30159;
  assign n30111 = n30110 ^ n30101;
  assign n30130 = n30111 ^ n30088;
  assign n30123 = n30122 ^ n30081;
  assign n30124 = n30121 & ~n30123;
  assign n30129 = n30128 ^ n30124;
  assign n30131 = n30130 ^ n30129;
  assign n30112 = ~n30088 & ~n30111;
  assign n30116 = n30115 ^ n30112;
  assign n30132 = n30131 ^ n30116;
  assign n30145 = n30144 ^ n30132;
  assign n30176 = n30160 ^ n30145;
  assign n30148 = n30123 ^ n30082;
  assign n30147 = n30146 ^ n30122;
  assign n30153 = n30148 ^ n30147;
  assign n30149 = n30147 & ~n30148;
  assign n30151 = n30150 ^ n30149;
  assign n30152 = n30151 ^ n30116;
  assign n30154 = n30153 ^ n30152;
  assign n30174 = ~n30132 & n30144;
  assign n30175 = ~n30154 & n30174;
  assign n30177 = n30176 ^ n30175;
  assign n30192 = ~n30122 & n30177;
  assign n30171 = n30132 & n30159;
  assign n30172 = n30154 & n30171;
  assign n30164 = n30159 ^ n30154;
  assign n30170 = n30164 ^ n30160;
  assign n30173 = n30172 ^ n30170;
  assign n30191 = ~n30135 & ~n30173;
  assign n30193 = n30192 ^ n30191;
  assign n30178 = n30177 ^ n30173;
  assign n30165 = n30160 ^ n30132;
  assign n30166 = ~n30164 & n30165;
  assign n30167 = n30166 ^ n30154;
  assign n30161 = n30160 ^ n30154;
  assign n30162 = n30145 & ~n30161;
  assign n30163 = n30162 ^ n30132;
  assign n30168 = n30167 ^ n30163;
  assign n30179 = n30178 ^ n30168;
  assign n30189 = ~n30139 & n30179;
  assign n30188 = n30114 & ~n30168;
  assign n30190 = n30189 ^ n30188;
  assign n30194 = n30193 ^ n30190;
  assign n30185 = n30173 ^ n30167;
  assign n30186 = n30127 & n30185;
  assign n30182 = n30177 ^ n30163;
  assign n30183 = ~n30146 & n30182;
  assign n30180 = ~n30126 & n30179;
  assign n30169 = n30082 & ~n30168;
  assign n30181 = n30180 ^ n30169;
  assign n30184 = n30183 ^ n30181;
  assign n30187 = n30186 ^ n30184;
  assign n30195 = n30194 ^ n30187;
  assign n30197 = n30196 ^ n30195;
  assign n30205 = n29889 ^ n26779;
  assign n30203 = n30191 ^ n30181;
  assign n30200 = n30101 & n30185;
  assign n30198 = n30133 & ~n30173;
  assign n30199 = n30198 ^ n30186;
  assign n30201 = n30200 ^ n30199;
  assign n30202 = n30201 ^ n30190;
  assign n30204 = n30203 ^ n30202;
  assign n30206 = n30205 ^ n30204;
  assign n30218 = n29884 ^ n26804;
  assign n30219 = n30218 ^ n30169;
  assign n30215 = ~n30088 & ~n30178;
  assign n30213 = ~n30111 & ~n30178;
  assign n30212 = ~n30125 & n30182;
  assign n30214 = n30213 ^ n30212;
  assign n30216 = n30215 ^ n30214;
  assign n30209 = ~n30148 & n30163;
  assign n30207 = n30121 & ~n30167;
  assign n30208 = n30207 ^ n30200;
  assign n30210 = n30209 ^ n30208;
  assign n30211 = n30210 ^ n30188;
  assign n30217 = n30216 ^ n30211;
  assign n30220 = n30219 ^ n30217;
  assign n30222 = n29867 ^ n26810;
  assign n30223 = n30222 ^ n30201;
  assign n30221 = n30193 ^ n30184;
  assign n30224 = n30223 ^ n30221;
  assign n30229 = n29874 ^ n26822;
  assign n30228 = n30147 & n30163;
  assign n30230 = n30229 ^ n30228;
  assign n30226 = n30207 ^ n30199;
  assign n30225 = n30193 ^ n30181;
  assign n30227 = n30226 ^ n30225;
  assign n30231 = n30230 ^ n30227;
  assign n30237 = n29881 ^ n26831;
  assign n30238 = n30237 ^ n30193;
  assign n30234 = ~n30123 & ~n30167;
  assign n30235 = n30234 ^ n30210;
  assign n30232 = n30214 ^ n30189;
  assign n30233 = n30232 ^ n30184;
  assign n30236 = n30235 ^ n30233;
  assign n30239 = n30238 ^ n30236;
  assign n30245 = n29877 ^ n26848;
  assign n30241 = n30134 & n30177;
  assign n30242 = n30241 ^ n30228;
  assign n30243 = n30242 ^ n30232;
  assign n30240 = n30192 ^ n30181;
  assign n30244 = n30243 ^ n30240;
  assign n30246 = n30245 ^ n30244;
  assign n30250 = n29893 ^ n26856;
  assign n30248 = n30242 ^ n30208;
  assign n30247 = n30212 ^ n30184;
  assign n30249 = n30248 ^ n30247;
  assign n30251 = n30250 ^ n30249;
  assign n30376 = n27893 ^ n26617;
  assign n30272 = n28664 ^ n28370;
  assign n30271 = n28675 ^ n28652;
  assign n30273 = n30272 ^ n30271;
  assign n30274 = n30273 ^ n26635;
  assign n30267 = n28670 ^ n28646;
  assign n30268 = n30267 ^ n28575;
  assign n30269 = n30268 ^ n28658;
  assign n30270 = n30269 ^ n26642;
  assign n30275 = n30274 ^ n30270;
  assign n30265 = n28600 ^ n26653;
  assign n30263 = n28696 ^ n28580;
  assign n30264 = n30263 ^ n28597;
  assign n30266 = n30265 ^ n30264;
  assign n30276 = n30275 ^ n30266;
  assign n30257 = n28608 ^ n28528;
  assign n30258 = n30257 ^ n28518;
  assign n30259 = n30258 ^ n28626;
  assign n30260 = n30259 ^ n28562;
  assign n30261 = n30260 ^ n26666;
  assign n30308 = n30270 ^ n30261;
  assign n30295 = n28247 ^ n26618;
  assign n30293 = n28655 ^ n28585;
  assign n30292 = n28571 ^ n28119;
  assign n30294 = n30293 ^ n30292;
  assign n30296 = n30295 ^ n30294;
  assign n30253 = n28633 ^ n28580;
  assign n30252 = n28665 ^ n28120;
  assign n30254 = n30253 ^ n30252;
  assign n30255 = n30254 ^ n28498;
  assign n30256 = n30255 ^ n26608;
  assign n30297 = n30296 ^ n30256;
  assign n30288 = n28580 ^ n28548;
  assign n30289 = n30288 ^ n28637;
  assign n30287 = n28627 ^ n28110;
  assign n30290 = n30289 ^ n30287;
  assign n30285 = n28238 ^ n26675;
  assign n30283 = n28533 ^ n26682;
  assign n30280 = n28692 ^ n28580;
  assign n30281 = n30280 ^ n28614;
  assign n30279 = n28597 ^ n28528;
  assign n30282 = n30281 ^ n30279;
  assign n30284 = n30283 ^ n30282;
  assign n30286 = n30285 ^ n30284;
  assign n30291 = n30290 ^ n30286;
  assign n30298 = n30297 ^ n30291;
  assign n30339 = n30308 ^ n30298;
  assign n30262 = n30261 ^ n30256;
  assign n30313 = n30274 ^ n30261;
  assign n30316 = n30313 ^ n30297;
  assign n30317 = n30262 & n30316;
  assign n30309 = n30308 ^ n30291;
  assign n30310 = n30297 & n30309;
  assign n30318 = n30317 ^ n30310;
  assign n30340 = n30339 ^ n30318;
  assign n30334 = n30298 ^ n30266;
  assign n30335 = n30284 ^ n30276;
  assign n30304 = n30296 ^ n30261;
  assign n30336 = n30335 ^ n30304;
  assign n30337 = n30334 & n30336;
  assign n30299 = n30296 ^ n30284;
  assign n30300 = n30299 ^ n30262;
  assign n30301 = n30298 & n30300;
  assign n30338 = n30337 ^ n30301;
  assign n30341 = n30340 ^ n30338;
  assign n30303 = n30298 ^ n30275;
  assign n30307 = n30303 & n30304;
  assign n30311 = n30310 ^ n30307;
  assign n30305 = n30304 ^ n30303;
  assign n30277 = n30276 ^ n30256;
  assign n30278 = n30266 & n30277;
  assign n30302 = n30301 ^ n30278;
  assign n30306 = n30305 ^ n30302;
  assign n30312 = n30311 ^ n30306;
  assign n30347 = n30341 ^ n30312;
  assign n30314 = n30313 ^ n30291;
  assign n30321 = n30299 & n30314;
  assign n30320 = n30276 & ~n30284;
  assign n30322 = n30321 ^ n30320;
  assign n30315 = n30314 ^ n30299;
  assign n30319 = n30318 ^ n30315;
  assign n30323 = n30322 ^ n30319;
  assign n30342 = n30323 & n30341;
  assign n30348 = n30347 ^ n30342;
  assign n30325 = n30297 ^ n30277;
  assign n30324 = n30314 ^ n30276;
  assign n30329 = n30325 ^ n30324;
  assign n30326 = n30324 & n30325;
  assign n30327 = n30326 ^ n30321;
  assign n30328 = n30327 ^ n30311;
  assign n30330 = n30329 ^ n30328;
  assign n30345 = ~n30312 & n30341;
  assign n30346 = n30330 & n30345;
  assign n30349 = n30348 ^ n30346;
  assign n30372 = n30276 & n30349;
  assign n30331 = n30330 ^ n30323;
  assign n30343 = n30342 ^ n30331;
  assign n30332 = n30323 & n30331;
  assign n30333 = n30312 & n30332;
  assign n30344 = n30343 ^ n30333;
  assign n30371 = n30336 & n30344;
  assign n30373 = n30372 ^ n30371;
  assign n30354 = n30342 ^ n30312;
  assign n30355 = n30331 & n30354;
  assign n30356 = n30355 ^ n30330;
  assign n30351 = n30342 ^ n30330;
  assign n30352 = n30347 & n30351;
  assign n30353 = n30352 ^ n30312;
  assign n30357 = n30356 ^ n30353;
  assign n30369 = n30309 & n30357;
  assign n30350 = n30349 ^ n30344;
  assign n30358 = n30357 ^ n30350;
  assign n30368 = n30316 & n30358;
  assign n30370 = n30369 ^ n30368;
  assign n30374 = n30373 ^ n30370;
  assign n30365 = n30356 ^ n30344;
  assign n30366 = n30300 & n30365;
  assign n30362 = n30353 ^ n30349;
  assign n30363 = n30314 & n30362;
  assign n30360 = n30297 & n30357;
  assign n30359 = n30262 & n30358;
  assign n30361 = n30360 ^ n30359;
  assign n30364 = n30363 ^ n30361;
  assign n30367 = n30366 ^ n30364;
  assign n30375 = n30374 ^ n30367;
  assign n30377 = n30376 ^ n30375;
  assign n30385 = n27909 ^ n26641;
  assign n30383 = n30371 ^ n30361;
  assign n30380 = n30298 & n30365;
  assign n30378 = n30334 & n30344;
  assign n30379 = n30378 ^ n30366;
  assign n30381 = n30380 ^ n30379;
  assign n30382 = n30381 ^ n30370;
  assign n30384 = n30383 ^ n30382;
  assign n30386 = n30385 ^ n30384;
  assign n30398 = n27934 ^ n26634;
  assign n30399 = n30398 ^ n30360;
  assign n30395 = n30304 & n30350;
  assign n30393 = n30299 & n30362;
  assign n30392 = n30303 & n30350;
  assign n30394 = n30393 ^ n30392;
  assign n30396 = n30395 ^ n30394;
  assign n30389 = n30325 & n30353;
  assign n30387 = n30266 & n30356;
  assign n30388 = n30387 ^ n30380;
  assign n30390 = n30389 ^ n30388;
  assign n30391 = n30390 ^ n30369;
  assign n30397 = n30396 ^ n30391;
  assign n30400 = n30399 ^ n30397;
  assign n30402 = n27940 ^ n26607;
  assign n30403 = n30402 ^ n30381;
  assign n30401 = n30373 ^ n30364;
  assign n30404 = n30403 ^ n30401;
  assign n30409 = n27952 ^ n26674;
  assign n30408 = n30324 & n30353;
  assign n30410 = n30409 ^ n30408;
  assign n30406 = n30387 ^ n30379;
  assign n30405 = n30373 ^ n30361;
  assign n30407 = n30406 ^ n30405;
  assign n30411 = n30410 ^ n30407;
  assign n30417 = n27966 ^ n26665;
  assign n30418 = n30417 ^ n30373;
  assign n30414 = n30277 & n30356;
  assign n30415 = n30414 ^ n30390;
  assign n30412 = n30394 ^ n30368;
  assign n30413 = n30412 ^ n30364;
  assign n30416 = n30415 ^ n30413;
  assign n30419 = n30418 ^ n30416;
  assign n30425 = n27979 ^ n26681;
  assign n30423 = n30372 ^ n30361;
  assign n30420 = n30335 & n30349;
  assign n30421 = n30420 ^ n30408;
  assign n30422 = n30421 ^ n30412;
  assign n30424 = n30423 ^ n30422;
  assign n30426 = n30425 ^ n30424;
  assign n30430 = n27987 ^ n26652;
  assign n30428 = n30421 ^ n30388;
  assign n30427 = n30393 ^ n30364;
  assign n30429 = n30428 ^ n30427;
  assign n30431 = n30430 ^ n30429;
  assign n30559 = n29020 ^ n27747;
  assign n30482 = n29712 ^ n29673;
  assign n30483 = n30482 ^ n29786;
  assign n30484 = n30483 ^ n29704;
  assign n30485 = n30484 ^ n27812;
  assign n30473 = n29757 ^ n27776;
  assign n30471 = n29774 ^ n29348;
  assign n30470 = n29764 ^ n29750;
  assign n30472 = n30471 ^ n30470;
  assign n30474 = n30473 ^ n30472;
  assign n30468 = n29684 ^ n27804;
  assign n30466 = n29769 ^ n29757;
  assign n30465 = n29741 ^ n29677;
  assign n30467 = n30466 ^ n30465;
  assign n30469 = n30468 ^ n30467;
  assign n30475 = n30474 ^ n30469;
  assign n30486 = n30485 ^ n30475;
  assign n30441 = n29731 ^ n27767;
  assign n30439 = n29700 ^ n29660;
  assign n30438 = n29644 ^ n29617;
  assign n30440 = n30439 ^ n30438;
  assign n30442 = n30441 ^ n30440;
  assign n30478 = n30469 ^ n30442;
  assign n30460 = n29673 ^ n29631;
  assign n30461 = n30460 ^ n29732;
  assign n30459 = n29718 ^ n29460;
  assign n30462 = n30461 ^ n30459;
  assign n30457 = n29591 ^ n27786;
  assign n30455 = n29660 ^ n27795;
  assign n30452 = n29789 ^ n29673;
  assign n30453 = n30452 ^ n29712;
  assign n30451 = n29694 ^ n29649;
  assign n30454 = n30453 ^ n30451;
  assign n30456 = n30455 ^ n30454;
  assign n30458 = n30457 ^ n30456;
  assign n30463 = n30462 ^ n30458;
  assign n30447 = n29600 ^ n27749;
  assign n30445 = n29744 ^ n29684;
  assign n30444 = n29668 ^ n29469;
  assign n30446 = n30445 ^ n30444;
  assign n30448 = n30447 ^ n30446;
  assign n30436 = n29774 ^ n27739;
  assign n30433 = n29722 ^ n29673;
  assign n30434 = n30433 ^ n29601;
  assign n30432 = n29474 ^ n29232;
  assign n30435 = n30434 ^ n30432;
  assign n30437 = n30436 ^ n30435;
  assign n30450 = n30448 ^ n30437;
  assign n30464 = n30463 ^ n30450;
  assign n30522 = n30478 ^ n30464;
  assign n30443 = n30442 ^ n30437;
  assign n30496 = n30474 ^ n30442;
  assign n30499 = n30496 ^ n30450;
  assign n30500 = n30443 & n30499;
  assign n30479 = n30478 ^ n30463;
  assign n30480 = n30450 & n30479;
  assign n30501 = n30500 ^ n30480;
  assign n30523 = n30522 ^ n30501;
  assign n30517 = n30486 ^ n30456;
  assign n30449 = n30448 ^ n30442;
  assign n30518 = n30517 ^ n30449;
  assign n30519 = n30485 ^ n30464;
  assign n30520 = n30518 & n30519;
  assign n30489 = n30456 ^ n30448;
  assign n30490 = n30489 ^ n30443;
  assign n30491 = n30464 & n30490;
  assign n30521 = n30520 ^ n30491;
  assign n30524 = n30523 ^ n30521;
  assign n30476 = n30475 ^ n30464;
  assign n30493 = n30476 ^ n30449;
  assign n30487 = n30486 ^ n30437;
  assign n30488 = n30485 & n30487;
  assign n30492 = n30491 ^ n30488;
  assign n30494 = n30493 ^ n30492;
  assign n30477 = n30449 & n30476;
  assign n30481 = n30480 ^ n30477;
  assign n30495 = n30494 ^ n30481;
  assign n30530 = n30524 ^ n30495;
  assign n30504 = ~n30456 & n30486;
  assign n30497 = n30496 ^ n30463;
  assign n30503 = n30489 & n30497;
  assign n30505 = n30504 ^ n30503;
  assign n30498 = n30497 ^ n30489;
  assign n30502 = n30501 ^ n30498;
  assign n30506 = n30505 ^ n30502;
  assign n30525 = n30506 & n30524;
  assign n30531 = n30530 ^ n30525;
  assign n30508 = n30487 ^ n30450;
  assign n30507 = n30497 ^ n30486;
  assign n30512 = n30508 ^ n30507;
  assign n30509 = n30507 & n30508;
  assign n30510 = n30509 ^ n30503;
  assign n30511 = n30510 ^ n30481;
  assign n30513 = n30512 ^ n30511;
  assign n30528 = n30513 & n30524;
  assign n30529 = ~n30495 & n30528;
  assign n30532 = n30531 ^ n30529;
  assign n30555 = n30486 & n30532;
  assign n30514 = n30513 ^ n30506;
  assign n30526 = n30525 ^ n30514;
  assign n30515 = n30506 & n30514;
  assign n30516 = n30495 & n30515;
  assign n30527 = n30526 ^ n30516;
  assign n30554 = n30518 & n30527;
  assign n30556 = n30555 ^ n30554;
  assign n30537 = n30525 ^ n30495;
  assign n30538 = n30514 & n30537;
  assign n30539 = n30538 ^ n30513;
  assign n30534 = n30525 ^ n30513;
  assign n30535 = n30530 & n30534;
  assign n30536 = n30535 ^ n30495;
  assign n30540 = n30539 ^ n30536;
  assign n30552 = n30479 & n30540;
  assign n30533 = n30532 ^ n30527;
  assign n30541 = n30540 ^ n30533;
  assign n30551 = n30499 & n30541;
  assign n30553 = n30552 ^ n30551;
  assign n30557 = n30556 ^ n30553;
  assign n30548 = n30539 ^ n30527;
  assign n30549 = n30490 & n30548;
  assign n30545 = n30536 ^ n30532;
  assign n30546 = n30497 & n30545;
  assign n30543 = n30450 & n30540;
  assign n30542 = n30443 & n30541;
  assign n30544 = n30543 ^ n30542;
  assign n30547 = n30546 ^ n30544;
  assign n30550 = n30549 ^ n30547;
  assign n30558 = n30557 ^ n30550;
  assign n30560 = n30559 ^ n30558;
  assign n30568 = n29036 ^ n27802;
  assign n30566 = n30554 ^ n30544;
  assign n30563 = n30464 & n30548;
  assign n30561 = n30519 & n30527;
  assign n30562 = n30561 ^ n30549;
  assign n30564 = n30563 ^ n30562;
  assign n30565 = n30564 ^ n30553;
  assign n30567 = n30566 ^ n30565;
  assign n30569 = n30568 ^ n30567;
  assign n30581 = n29061 ^ n27774;
  assign n30582 = n30581 ^ n30543;
  assign n30578 = n30449 & n30533;
  assign n30576 = n30489 & n30545;
  assign n30575 = n30476 & n30533;
  assign n30577 = n30576 ^ n30575;
  assign n30579 = n30578 ^ n30577;
  assign n30572 = n30508 & n30536;
  assign n30570 = n30485 & n30539;
  assign n30571 = n30570 ^ n30563;
  assign n30573 = n30572 ^ n30571;
  assign n30574 = n30573 ^ n30552;
  assign n30580 = n30579 ^ n30574;
  assign n30583 = n30582 ^ n30580;
  assign n30585 = n29067 ^ n27737;
  assign n30586 = n30585 ^ n30564;
  assign n30584 = n30556 ^ n30547;
  assign n30587 = n30586 ^ n30584;
  assign n30592 = n29079 ^ n27784;
  assign n30591 = n30507 & n30536;
  assign n30593 = n30592 ^ n30591;
  assign n30589 = n30570 ^ n30562;
  assign n30588 = n30556 ^ n30544;
  assign n30590 = n30589 ^ n30588;
  assign n30594 = n30593 ^ n30590;
  assign n30600 = n29093 ^ n27765;
  assign n30601 = n30600 ^ n30556;
  assign n30597 = n30487 & n30539;
  assign n30598 = n30597 ^ n30573;
  assign n30595 = n30577 ^ n30551;
  assign n30596 = n30595 ^ n30547;
  assign n30599 = n30598 ^ n30596;
  assign n30602 = n30601 ^ n30599;
  assign n30608 = n29106 ^ n27793;
  assign n30606 = n30555 ^ n30544;
  assign n30603 = n30517 & n30532;
  assign n30604 = n30603 ^ n30591;
  assign n30605 = n30604 ^ n30595;
  assign n30607 = n30606 ^ n30605;
  assign n30609 = n30608 ^ n30607;
  assign n30613 = n29114 ^ n27810;
  assign n30611 = n30604 ^ n30571;
  assign n30610 = n30576 ^ n30547;
  assign n30612 = n30611 ^ n30610;
  assign n30614 = n30613 ^ n30612;
  assign n30734 = n29976 ^ n28874;
  assign n30659 = n28936 ^ n26358;
  assign n30658 = n26376 ^ n26282;
  assign n30660 = n30659 ^ n30658;
  assign n30649 = n28900 ^ n26266;
  assign n30647 = n26413 ^ n26391;
  assign n30648 = n30647 ^ n26420;
  assign n30650 = n30649 ^ n30648;
  assign n30645 = n28928 ^ n26426;
  assign n30643 = n26391 ^ n26342;
  assign n30644 = n30643 ^ n26401;
  assign n30646 = n30645 ^ n30644;
  assign n30651 = n30650 ^ n30646;
  assign n30661 = n30660 ^ n30651;
  assign n30622 = n28891 ^ n26301;
  assign n30620 = n26323 ^ n23285;
  assign n30621 = n30620 ^ n25179;
  assign n30623 = n30622 ^ n30621;
  assign n30654 = n30646 ^ n30623;
  assign n30627 = n28873 ^ n26405;
  assign n30625 = n26342 ^ n26234;
  assign n30626 = n30625 ^ n26352;
  assign n30628 = n30627 ^ n30626;
  assign n30617 = n26358 ^ n26330;
  assign n30618 = n30617 ^ n28863;
  assign n30615 = n26413 ^ n26235;
  assign n30616 = n30615 ^ n26259;
  assign n30619 = n30618 ^ n30616;
  assign n30641 = n30628 ^ n30619;
  assign n30637 = n26358 ^ n26104;
  assign n30638 = n30637 ^ n28910;
  assign n30636 = n26324 ^ n26227;
  assign n30639 = n30638 ^ n30636;
  assign n30632 = n26380 ^ n26358;
  assign n30633 = n30632 ^ n28919;
  assign n30630 = n26282 ^ n23285;
  assign n30631 = n30630 ^ n26294;
  assign n30634 = n30633 ^ n30631;
  assign n30635 = n30634 ^ n26315;
  assign n30640 = n30639 ^ n30635;
  assign n30642 = n30641 ^ n30640;
  assign n30697 = n30654 ^ n30642;
  assign n30624 = n30623 ^ n30619;
  assign n30671 = n30650 ^ n30623;
  assign n30674 = n30671 ^ n30641;
  assign n30675 = n30624 & n30674;
  assign n30655 = n30654 ^ n30640;
  assign n30656 = n30641 & n30655;
  assign n30676 = n30675 ^ n30656;
  assign n30698 = n30697 ^ n30676;
  assign n30692 = n30661 ^ n30634;
  assign n30629 = n30628 ^ n30623;
  assign n30693 = n30692 ^ n30629;
  assign n30694 = n30660 ^ n30642;
  assign n30695 = n30693 & n30694;
  assign n30664 = n30634 ^ n30628;
  assign n30665 = n30664 ^ n30624;
  assign n30666 = n30642 & n30665;
  assign n30696 = n30695 ^ n30666;
  assign n30699 = n30698 ^ n30696;
  assign n30652 = n30651 ^ n30642;
  assign n30668 = n30652 ^ n30629;
  assign n30662 = n30661 ^ n30619;
  assign n30663 = n30660 & n30662;
  assign n30667 = n30666 ^ n30663;
  assign n30669 = n30668 ^ n30667;
  assign n30653 = n30629 & n30652;
  assign n30657 = n30656 ^ n30653;
  assign n30670 = n30669 ^ n30657;
  assign n30705 = n30699 ^ n30670;
  assign n30679 = ~n30634 & n30661;
  assign n30672 = n30671 ^ n30640;
  assign n30678 = n30664 & n30672;
  assign n30680 = n30679 ^ n30678;
  assign n30673 = n30672 ^ n30664;
  assign n30677 = n30676 ^ n30673;
  assign n30681 = n30680 ^ n30677;
  assign n30700 = n30681 & n30699;
  assign n30706 = n30705 ^ n30700;
  assign n30683 = n30672 ^ n30661;
  assign n30682 = n30662 ^ n30641;
  assign n30687 = n30683 ^ n30682;
  assign n30684 = n30682 & n30683;
  assign n30685 = n30684 ^ n30678;
  assign n30686 = n30685 ^ n30657;
  assign n30688 = n30687 ^ n30686;
  assign n30703 = ~n30670 & n30699;
  assign n30704 = n30688 & n30703;
  assign n30707 = n30706 ^ n30704;
  assign n30730 = n30661 & n30707;
  assign n30689 = n30688 ^ n30681;
  assign n30701 = n30700 ^ n30689;
  assign n30690 = n30681 & n30689;
  assign n30691 = n30670 & n30690;
  assign n30702 = n30701 ^ n30691;
  assign n30729 = n30693 & n30702;
  assign n30731 = n30730 ^ n30729;
  assign n30712 = n30700 ^ n30670;
  assign n30713 = n30689 & n30712;
  assign n30714 = n30713 ^ n30688;
  assign n30709 = n30700 ^ n30688;
  assign n30710 = n30705 & n30709;
  assign n30711 = n30710 ^ n30670;
  assign n30715 = n30714 ^ n30711;
  assign n30727 = n30655 & n30715;
  assign n30708 = n30707 ^ n30702;
  assign n30716 = n30715 ^ n30708;
  assign n30726 = n30674 & n30716;
  assign n30728 = n30727 ^ n30726;
  assign n30732 = n30731 ^ n30728;
  assign n30723 = n30714 ^ n30702;
  assign n30724 = n30665 & n30723;
  assign n30720 = n30711 ^ n30707;
  assign n30721 = n30672 & n30720;
  assign n30718 = n30641 & n30715;
  assign n30717 = n30624 & n30716;
  assign n30719 = n30718 ^ n30717;
  assign n30722 = n30721 ^ n30719;
  assign n30725 = n30724 ^ n30722;
  assign n30733 = n30732 ^ n30725;
  assign n30735 = n30734 ^ n30733;
  assign n30743 = n29992 ^ n28929;
  assign n30741 = n30729 ^ n30719;
  assign n30738 = n30642 & n30723;
  assign n30736 = n30694 & n30702;
  assign n30737 = n30736 ^ n30724;
  assign n30739 = n30738 ^ n30737;
  assign n30740 = n30739 ^ n30728;
  assign n30742 = n30741 ^ n30740;
  assign n30744 = n30743 ^ n30742;
  assign n30756 = n30017 ^ n28901;
  assign n30757 = n30756 ^ n30718;
  assign n30753 = n30629 & n30708;
  assign n30751 = n30664 & n30720;
  assign n30750 = n30652 & n30708;
  assign n30752 = n30751 ^ n30750;
  assign n30754 = n30753 ^ n30752;
  assign n30747 = n30682 & n30711;
  assign n30745 = n30660 & n30714;
  assign n30746 = n30745 ^ n30738;
  assign n30748 = n30747 ^ n30746;
  assign n30749 = n30748 ^ n30727;
  assign n30755 = n30754 ^ n30749;
  assign n30758 = n30757 ^ n30755;
  assign n30760 = n30023 ^ n28864;
  assign n30761 = n30760 ^ n30739;
  assign n30759 = n30731 ^ n30722;
  assign n30762 = n30761 ^ n30759;
  assign n30767 = n30035 ^ n28911;
  assign n30766 = n30683 & n30711;
  assign n30768 = n30767 ^ n30766;
  assign n30764 = n30745 ^ n30737;
  assign n30763 = n30731 ^ n30719;
  assign n30765 = n30764 ^ n30763;
  assign n30769 = n30768 ^ n30765;
  assign n30775 = n30049 ^ n28892;
  assign n30776 = n30775 ^ n30731;
  assign n30772 = n30662 & n30714;
  assign n30773 = n30772 ^ n30748;
  assign n30770 = n30752 ^ n30726;
  assign n30771 = n30770 ^ n30722;
  assign n30774 = n30773 ^ n30771;
  assign n30777 = n30776 ^ n30774;
  assign n30783 = n30062 ^ n28920;
  assign n30781 = n30730 ^ n30719;
  assign n30778 = n30692 & n30707;
  assign n30779 = n30778 ^ n30766;
  assign n30780 = n30779 ^ n30770;
  assign n30782 = n30781 ^ n30780;
  assign n30784 = n30783 ^ n30782;
  assign n30788 = n30070 ^ n28937;
  assign n30786 = n30779 ^ n30746;
  assign n30785 = n30751 ^ n30722;
  assign n30787 = n30786 ^ n30785;
  assign n30789 = n30788 ^ n30787;
  assign n30910 = n30196 ^ n29871;
  assign n30819 = n29878 ^ n28533;
  assign n30816 = n28696 ^ n28585;
  assign n30817 = n30816 ^ n30280;
  assign n30818 = n30817 ^ n30257;
  assign n30820 = n30819 ^ n30818;
  assign n30810 = n29894 ^ n28600;
  assign n30808 = n28692 ^ n28596;
  assign n30809 = n30808 ^ n28586;
  assign n30811 = n30810 ^ n30809;
  assign n30805 = n29890 ^ n28574;
  assign n30803 = n28655 ^ n28571;
  assign n30804 = n30803 ^ n28676;
  assign n30806 = n30805 ^ n30804;
  assign n30801 = n29885 ^ n28651;
  assign n30800 = n30267 ^ n28499;
  assign n30802 = n30801 ^ n30800;
  assign n30807 = n30806 ^ n30802;
  assign n30812 = n30811 ^ n30807;
  assign n30866 = n30820 ^ n30812;
  assign n30828 = n28626 ^ n28548;
  assign n30829 = n30828 ^ n28615;
  assign n30827 = n29882 ^ n28518;
  assign n30830 = n30829 ^ n30827;
  assign n30797 = n29871 ^ n28247;
  assign n30795 = n28580 ^ n28119;
  assign n30796 = n30795 ^ n28659;
  assign n30798 = n30797 ^ n30796;
  assign n30838 = n30830 ^ n30798;
  assign n30867 = n30866 ^ n30838;
  assign n30855 = n30812 & n30820;
  assign n30831 = n30830 ^ n30802;
  assign n30824 = n29875 ^ n28238;
  assign n30822 = n28585 ^ n28562;
  assign n30823 = n30822 ^ n30288;
  assign n30825 = n30824 ^ n30823;
  assign n30815 = n28633 ^ n28110;
  assign n30821 = n30820 ^ n30815;
  assign n30826 = n30825 ^ n30821;
  assign n30832 = n30831 ^ n30826;
  assign n30835 = n30820 ^ n30798;
  assign n30836 = ~n30832 & n30835;
  assign n30856 = n30855 ^ n30836;
  assign n30853 = n30835 ^ n30832;
  assign n30793 = n29868 ^ n28504;
  assign n30790 = n28637 ^ n28585;
  assign n30791 = n30790 ^ n30253;
  assign n30792 = n30791 ^ n30272;
  assign n30794 = n30793 ^ n30792;
  assign n30849 = n30830 ^ n30794;
  assign n30799 = n30798 ^ n30794;
  assign n30850 = n30831 ^ n30799;
  assign n30851 = n30849 & ~n30850;
  assign n30842 = n30830 ^ n30806;
  assign n30843 = n30842 ^ n30826;
  assign n30844 = ~n30799 & ~n30843;
  assign n30852 = n30851 ^ n30844;
  assign n30854 = n30853 ^ n30852;
  assign n30857 = n30856 ^ n30854;
  assign n30839 = n30826 ^ n30799;
  assign n30871 = n30842 ^ n30839;
  assign n30872 = n30871 ^ n30852;
  assign n30868 = n30839 ^ n30811;
  assign n30869 = n30867 & n30868;
  assign n30860 = n30849 ^ n30835;
  assign n30861 = n30839 & n30860;
  assign n30870 = n30869 ^ n30861;
  assign n30873 = n30872 ^ n30870;
  assign n30874 = ~n30857 & n30873;
  assign n30833 = n30832 ^ n30812;
  assign n30813 = n30812 ^ n30794;
  assign n30814 = n30813 ^ n30799;
  assign n30847 = n30833 ^ n30814;
  assign n30840 = n30839 ^ n30807;
  assign n30841 = ~n30838 & n30840;
  assign n30845 = n30844 ^ n30841;
  assign n30834 = ~n30814 & ~n30833;
  assign n30837 = n30836 ^ n30834;
  assign n30846 = n30845 ^ n30837;
  assign n30848 = n30847 ^ n30846;
  assign n30858 = n30857 ^ n30848;
  assign n30890 = n30874 ^ n30858;
  assign n30863 = n30840 ^ n30838;
  assign n30859 = n30811 & n30813;
  assign n30862 = n30861 ^ n30859;
  assign n30864 = n30863 ^ n30862;
  assign n30865 = n30864 ^ n30845;
  assign n30888 = ~n30857 & ~n30865;
  assign n30889 = ~n30848 & n30888;
  assign n30891 = n30890 ^ n30889;
  assign n30906 = n30867 & ~n30891;
  assign n30885 = n30865 & n30873;
  assign n30886 = n30848 & n30885;
  assign n30878 = n30873 ^ n30865;
  assign n30884 = n30878 ^ n30874;
  assign n30887 = n30886 ^ n30884;
  assign n30905 = n30812 & ~n30887;
  assign n30907 = n30906 ^ n30905;
  assign n30892 = n30891 ^ n30887;
  assign n30879 = n30874 ^ n30848;
  assign n30880 = ~n30878 & n30879;
  assign n30881 = n30880 ^ n30865;
  assign n30875 = n30874 ^ n30865;
  assign n30876 = ~n30858 & ~n30875;
  assign n30877 = n30876 ^ n30848;
  assign n30882 = n30881 ^ n30877;
  assign n30893 = n30892 ^ n30882;
  assign n30903 = ~n30850 & ~n30893;
  assign n30902 = ~n30843 & ~n30882;
  assign n30904 = n30903 ^ n30902;
  assign n30908 = n30907 ^ n30904;
  assign n30899 = n30891 ^ n30877;
  assign n30900 = n30860 & ~n30899;
  assign n30896 = n30887 ^ n30881;
  assign n30897 = ~n30832 & n30896;
  assign n30894 = n30849 & ~n30893;
  assign n30883 = ~n30799 & ~n30882;
  assign n30895 = n30894 ^ n30883;
  assign n30898 = n30897 ^ n30895;
  assign n30901 = n30900 ^ n30898;
  assign n30909 = n30908 ^ n30901;
  assign n30911 = n30910 ^ n30909;
  assign n30919 = n30205 ^ n29890;
  assign n30917 = n30906 ^ n30895;
  assign n30914 = n30839 & ~n30899;
  assign n30912 = n30868 & ~n30891;
  assign n30913 = n30912 ^ n30900;
  assign n30915 = n30914 ^ n30913;
  assign n30916 = n30915 ^ n30904;
  assign n30918 = n30917 ^ n30916;
  assign n30920 = n30919 ^ n30918;
  assign n30932 = n30218 ^ n29885;
  assign n30933 = n30932 ^ n30883;
  assign n30929 = ~n30838 & n30892;
  assign n30927 = n30835 & n30896;
  assign n30926 = n30840 & n30892;
  assign n30928 = n30927 ^ n30926;
  assign n30930 = n30929 ^ n30928;
  assign n30923 = ~n30814 & ~n30881;
  assign n30921 = n30811 & n30877;
  assign n30922 = n30921 ^ n30914;
  assign n30924 = n30923 ^ n30922;
  assign n30925 = n30924 ^ n30902;
  assign n30931 = n30930 ^ n30925;
  assign n30934 = n30933 ^ n30931;
  assign n30936 = n30222 ^ n29868;
  assign n30937 = n30936 ^ n30915;
  assign n30935 = n30907 ^ n30898;
  assign n30938 = n30937 ^ n30935;
  assign n30943 = n30229 ^ n29875;
  assign n30942 = ~n30833 & ~n30881;
  assign n30944 = n30943 ^ n30942;
  assign n30940 = n30921 ^ n30913;
  assign n30939 = n30907 ^ n30895;
  assign n30941 = n30940 ^ n30939;
  assign n30945 = n30944 ^ n30941;
  assign n30951 = n30237 ^ n29882;
  assign n30952 = n30951 ^ n30907;
  assign n30948 = n30813 & n30877;
  assign n30949 = n30948 ^ n30924;
  assign n30946 = n30928 ^ n30903;
  assign n30947 = n30946 ^ n30898;
  assign n30950 = n30949 ^ n30947;
  assign n30953 = n30952 ^ n30950;
  assign n30959 = n30245 ^ n29878;
  assign n30955 = ~n30866 & ~n30887;
  assign n30956 = n30955 ^ n30942;
  assign n30957 = n30956 ^ n30946;
  assign n30954 = n30905 ^ n30895;
  assign n30958 = n30957 ^ n30954;
  assign n30960 = n30959 ^ n30958;
  assign n30964 = n30250 ^ n29894;
  assign n30962 = n30956 ^ n30922;
  assign n30961 = n30927 ^ n30898;
  assign n30963 = n30962 ^ n30961;
  assign n30965 = n30964 ^ n30963;
  assign n31086 = n30376 ^ n26618;
  assign n31011 = n29711 ^ n26654;
  assign n31009 = n29704 ^ n29668;
  assign n31010 = n31009 ^ n30452;
  assign n31012 = n31011 ^ n31010;
  assign n30999 = n30466 ^ n29750;
  assign n31000 = n30999 ^ n29349;
  assign n31001 = n31000 ^ n26636;
  assign n30996 = n30445 ^ n29770;
  assign n30997 = n30996 ^ n29677;
  assign n30998 = n30997 ^ n26643;
  assign n31002 = n31001 ^ n30998;
  assign n31013 = n31012 ^ n31002;
  assign n30971 = n29731 ^ n29701;
  assign n30972 = n30971 ^ n29631;
  assign n30973 = n30972 ^ n29644;
  assign n30974 = n30973 ^ n26667;
  assign n31005 = n30998 ^ n30974;
  assign n30978 = n29600 ^ n26619;
  assign n30976 = n29745 ^ n29469;
  assign n30977 = n30976 ^ n29673;
  assign n30979 = n30978 ^ n30977;
  assign n30967 = n30471 ^ n30433;
  assign n30966 = n29718 ^ n29668;
  assign n30968 = n30967 ^ n30966;
  assign n30969 = n30968 ^ n29474;
  assign n30970 = n30969 ^ n26609;
  assign n30994 = n30979 ^ n30970;
  assign n30991 = n30460 ^ n29722;
  assign n30989 = n29668 ^ n29617;
  assign n30990 = n30989 ^ n29460;
  assign n30992 = n30991 ^ n30990;
  assign n30987 = n29591 ^ n26676;
  assign n30985 = n29660 ^ n26683;
  assign n30983 = n30452 ^ n29700;
  assign n30981 = n29786 ^ n29668;
  assign n30982 = n30981 ^ n29649;
  assign n30984 = n30983 ^ n30982;
  assign n30986 = n30985 ^ n30984;
  assign n30988 = n30987 ^ n30986;
  assign n30993 = n30992 ^ n30988;
  assign n30995 = n30994 ^ n30993;
  assign n31049 = n31005 ^ n30995;
  assign n30975 = n30974 ^ n30970;
  assign n31023 = n31001 ^ n30974;
  assign n31026 = n31023 ^ n30994;
  assign n31027 = n30975 & n31026;
  assign n31006 = n31005 ^ n30993;
  assign n31007 = n30994 & n31006;
  assign n31028 = n31027 ^ n31007;
  assign n31050 = n31049 ^ n31028;
  assign n31044 = n31012 ^ n30995;
  assign n31045 = n31013 ^ n30986;
  assign n30980 = n30979 ^ n30974;
  assign n31046 = n31045 ^ n30980;
  assign n31047 = n31044 & n31046;
  assign n31016 = n30986 ^ n30979;
  assign n31017 = n31016 ^ n30975;
  assign n31018 = n30995 & n31017;
  assign n31048 = n31047 ^ n31018;
  assign n31051 = n31050 ^ n31048;
  assign n31003 = n31002 ^ n30995;
  assign n31020 = n31003 ^ n30980;
  assign n31014 = n31013 ^ n30970;
  assign n31015 = n31012 & n31014;
  assign n31019 = n31018 ^ n31015;
  assign n31021 = n31020 ^ n31019;
  assign n31004 = n30980 & n31003;
  assign n31008 = n31007 ^ n31004;
  assign n31022 = n31021 ^ n31008;
  assign n31057 = n31051 ^ n31022;
  assign n31031 = ~n30986 & n31013;
  assign n31024 = n31023 ^ n30993;
  assign n31030 = n31016 & n31024;
  assign n31032 = n31031 ^ n31030;
  assign n31025 = n31024 ^ n31016;
  assign n31029 = n31028 ^ n31025;
  assign n31033 = n31032 ^ n31029;
  assign n31052 = n31033 & n31051;
  assign n31058 = n31057 ^ n31052;
  assign n31035 = n31014 ^ n30994;
  assign n31034 = n31024 ^ n31013;
  assign n31039 = n31035 ^ n31034;
  assign n31036 = n31034 & n31035;
  assign n31037 = n31036 ^ n31030;
  assign n31038 = n31037 ^ n31008;
  assign n31040 = n31039 ^ n31038;
  assign n31055 = n31040 & n31051;
  assign n31056 = ~n31022 & n31055;
  assign n31059 = n31058 ^ n31056;
  assign n31082 = n31013 & n31059;
  assign n31041 = n31040 ^ n31033;
  assign n31053 = n31052 ^ n31041;
  assign n31042 = n31033 & n31041;
  assign n31043 = n31022 & n31042;
  assign n31054 = n31053 ^ n31043;
  assign n31081 = n31046 & n31054;
  assign n31083 = n31082 ^ n31081;
  assign n31064 = n31052 ^ n31022;
  assign n31065 = n31041 & n31064;
  assign n31066 = n31065 ^ n31040;
  assign n31061 = n31052 ^ n31040;
  assign n31062 = n31057 & n31061;
  assign n31063 = n31062 ^ n31022;
  assign n31067 = n31066 ^ n31063;
  assign n31079 = n31006 & n31067;
  assign n31060 = n31059 ^ n31054;
  assign n31068 = n31067 ^ n31060;
  assign n31078 = n31026 & n31068;
  assign n31080 = n31079 ^ n31078;
  assign n31084 = n31083 ^ n31080;
  assign n31075 = n31066 ^ n31054;
  assign n31076 = n31017 & n31075;
  assign n31072 = n31063 ^ n31059;
  assign n31073 = n31024 & n31072;
  assign n31070 = n30994 & n31067;
  assign n31069 = n30975 & n31068;
  assign n31071 = n31070 ^ n31069;
  assign n31074 = n31073 ^ n31071;
  assign n31077 = n31076 ^ n31074;
  assign n31085 = n31084 ^ n31077;
  assign n31087 = n31086 ^ n31085;
  assign n31095 = n30385 ^ n26642;
  assign n31093 = n31081 ^ n31071;
  assign n31090 = n30995 & n31075;
  assign n31088 = n31044 & n31054;
  assign n31089 = n31088 ^ n31076;
  assign n31091 = n31090 ^ n31089;
  assign n31092 = n31091 ^ n31080;
  assign n31094 = n31093 ^ n31092;
  assign n31096 = n31095 ^ n31094;
  assign n31108 = n30398 ^ n26635;
  assign n31109 = n31108 ^ n31070;
  assign n31105 = n30980 & n31060;
  assign n31103 = n31016 & n31072;
  assign n31102 = n31003 & n31060;
  assign n31104 = n31103 ^ n31102;
  assign n31106 = n31105 ^ n31104;
  assign n31099 = n31035 & n31063;
  assign n31097 = n31012 & n31066;
  assign n31098 = n31097 ^ n31090;
  assign n31100 = n31099 ^ n31098;
  assign n31101 = n31100 ^ n31079;
  assign n31107 = n31106 ^ n31101;
  assign n31110 = n31109 ^ n31107;
  assign n31112 = n30402 ^ n26608;
  assign n31113 = n31112 ^ n31091;
  assign n31111 = n31083 ^ n31074;
  assign n31114 = n31113 ^ n31111;
  assign n31119 = n30409 ^ n26675;
  assign n31118 = n31034 & n31063;
  assign n31120 = n31119 ^ n31118;
  assign n31116 = n31097 ^ n31089;
  assign n31115 = n31083 ^ n31071;
  assign n31117 = n31116 ^ n31115;
  assign n31121 = n31120 ^ n31117;
  assign n31127 = n30417 ^ n26666;
  assign n31128 = n31127 ^ n31083;
  assign n31124 = n31014 & n31066;
  assign n31125 = n31124 ^ n31100;
  assign n31122 = n31104 ^ n31078;
  assign n31123 = n31122 ^ n31074;
  assign n31126 = n31125 ^ n31123;
  assign n31129 = n31128 ^ n31126;
  assign n31135 = n30425 ^ n26682;
  assign n31133 = n31082 ^ n31071;
  assign n31130 = n31045 & n31059;
  assign n31131 = n31130 ^ n31118;
  assign n31132 = n31131 ^ n31122;
  assign n31134 = n31133 ^ n31132;
  assign n31136 = n31135 ^ n31134;
  assign n31140 = n30430 ^ n26653;
  assign n31138 = n31131 ^ n31098;
  assign n31137 = n31103 ^ n31074;
  assign n31139 = n31138 ^ n31137;
  assign n31141 = n31140 ^ n31139;
  assign n31265 = n30559 ^ n27748;
  assign n31190 = n27809 ^ n26380;
  assign n31188 = n26358 ^ n26351;
  assign n31187 = n26285 ^ n26281;
  assign n31189 = n31188 ^ n31187;
  assign n31191 = n31190 ^ n31189;
  assign n31178 = n27773 ^ n26426;
  assign n31176 = n26266 ^ n26255;
  assign n31177 = n31176 ^ n26397;
  assign n31179 = n31178 ^ n31177;
  assign n31174 = n27801 ^ n26405;
  assign n31172 = n26426 ^ n26419;
  assign n31173 = n31172 ^ n26346;
  assign n31175 = n31174 ^ n31173;
  assign n31180 = n31179 ^ n31175;
  assign n31192 = n31191 ^ n31180;
  assign n31150 = n27764 ^ n26104;
  assign n31148 = n26301 ^ n26293;
  assign n31147 = n26323 ^ n24241;
  assign n31149 = n31148 ^ n31147;
  assign n31151 = n31150 ^ n31149;
  assign n31183 = n31175 ^ n31151;
  assign n31167 = n26351 ^ n25178;
  assign n31168 = n31167 ^ n30637;
  assign n31166 = n26242 ^ n26227;
  assign n31169 = n31168 ^ n31166;
  assign n31164 = n27783 ^ n26330;
  assign n31162 = n27792 ^ n26301;
  assign n31159 = n26375 ^ n26351;
  assign n31160 = n31159 ^ n30632;
  assign n31161 = n31160 ^ n24226;
  assign n31163 = n31162 ^ n31161;
  assign n31165 = n31164 ^ n31163;
  assign n31170 = n31169 ^ n31165;
  assign n31155 = n27746 ^ n26358;
  assign n31153 = n26405 ^ n26400;
  assign n31154 = n31153 ^ n26372;
  assign n31156 = n31155 ^ n31154;
  assign n31145 = n27736 ^ n26266;
  assign n31142 = n26351 ^ n26314;
  assign n31143 = n31142 ^ n30617;
  assign n31144 = n31143 ^ n26414;
  assign n31146 = n31145 ^ n31144;
  assign n31158 = n31156 ^ n31146;
  assign n31171 = n31170 ^ n31158;
  assign n31228 = n31183 ^ n31171;
  assign n31152 = n31151 ^ n31146;
  assign n31202 = n31179 ^ n31151;
  assign n31205 = n31202 ^ n31158;
  assign n31206 = n31152 & n31205;
  assign n31184 = n31183 ^ n31170;
  assign n31185 = n31158 & n31184;
  assign n31207 = n31206 ^ n31185;
  assign n31229 = n31228 ^ n31207;
  assign n31223 = n31191 ^ n31171;
  assign n31224 = n31192 ^ n31163;
  assign n31157 = n31156 ^ n31151;
  assign n31225 = n31224 ^ n31157;
  assign n31226 = n31223 & n31225;
  assign n31195 = n31163 ^ n31156;
  assign n31196 = n31195 ^ n31152;
  assign n31197 = n31171 & n31196;
  assign n31227 = n31226 ^ n31197;
  assign n31230 = n31229 ^ n31227;
  assign n31181 = n31180 ^ n31171;
  assign n31199 = n31181 ^ n31157;
  assign n31193 = n31192 ^ n31146;
  assign n31194 = n31191 & n31193;
  assign n31198 = n31197 ^ n31194;
  assign n31200 = n31199 ^ n31198;
  assign n31182 = n31157 & n31181;
  assign n31186 = n31185 ^ n31182;
  assign n31201 = n31200 ^ n31186;
  assign n31236 = n31230 ^ n31201;
  assign n31210 = ~n31163 & n31192;
  assign n31203 = n31202 ^ n31170;
  assign n31209 = n31195 & n31203;
  assign n31211 = n31210 ^ n31209;
  assign n31204 = n31203 ^ n31195;
  assign n31208 = n31207 ^ n31204;
  assign n31212 = n31211 ^ n31208;
  assign n31231 = n31212 & n31230;
  assign n31237 = n31236 ^ n31231;
  assign n31214 = n31193 ^ n31158;
  assign n31213 = n31203 ^ n31192;
  assign n31218 = n31214 ^ n31213;
  assign n31215 = n31213 & n31214;
  assign n31216 = n31215 ^ n31209;
  assign n31217 = n31216 ^ n31186;
  assign n31219 = n31218 ^ n31217;
  assign n31234 = ~n31201 & n31230;
  assign n31235 = n31219 & n31234;
  assign n31238 = n31237 ^ n31235;
  assign n31261 = n31192 & n31238;
  assign n31220 = n31219 ^ n31212;
  assign n31232 = n31231 ^ n31220;
  assign n31221 = n31212 & n31220;
  assign n31222 = n31201 & n31221;
  assign n31233 = n31232 ^ n31222;
  assign n31260 = n31225 & n31233;
  assign n31262 = n31261 ^ n31260;
  assign n31243 = n31231 ^ n31201;
  assign n31244 = n31220 & n31243;
  assign n31245 = n31244 ^ n31219;
  assign n31240 = n31231 ^ n31219;
  assign n31241 = n31236 & n31240;
  assign n31242 = n31241 ^ n31201;
  assign n31246 = n31245 ^ n31242;
  assign n31258 = n31184 & n31246;
  assign n31239 = n31238 ^ n31233;
  assign n31247 = n31246 ^ n31239;
  assign n31257 = n31205 & n31247;
  assign n31259 = n31258 ^ n31257;
  assign n31263 = n31262 ^ n31259;
  assign n31254 = n31245 ^ n31233;
  assign n31255 = n31196 & n31254;
  assign n31251 = n31242 ^ n31238;
  assign n31252 = n31203 & n31251;
  assign n31249 = n31158 & n31246;
  assign n31248 = n31152 & n31247;
  assign n31250 = n31249 ^ n31248;
  assign n31253 = n31252 ^ n31250;
  assign n31256 = n31255 ^ n31253;
  assign n31264 = n31263 ^ n31256;
  assign n31266 = n31265 ^ n31264;
  assign n31274 = n30568 ^ n27803;
  assign n31272 = n31260 ^ n31250;
  assign n31269 = n31171 & n31254;
  assign n31267 = n31223 & n31233;
  assign n31268 = n31267 ^ n31255;
  assign n31270 = n31269 ^ n31268;
  assign n31271 = n31270 ^ n31259;
  assign n31273 = n31272 ^ n31271;
  assign n31275 = n31274 ^ n31273;
  assign n31287 = n30581 ^ n27775;
  assign n31288 = n31287 ^ n31249;
  assign n31284 = n31157 & n31239;
  assign n31282 = n31195 & n31251;
  assign n31281 = n31181 & n31239;
  assign n31283 = n31282 ^ n31281;
  assign n31285 = n31284 ^ n31283;
  assign n31278 = n31214 & n31242;
  assign n31276 = n31191 & n31245;
  assign n31277 = n31276 ^ n31269;
  assign n31279 = n31278 ^ n31277;
  assign n31280 = n31279 ^ n31258;
  assign n31286 = n31285 ^ n31280;
  assign n31289 = n31288 ^ n31286;
  assign n31291 = n30585 ^ n27738;
  assign n31292 = n31291 ^ n31270;
  assign n31290 = n31262 ^ n31253;
  assign n31293 = n31292 ^ n31290;
  assign n31298 = n30592 ^ n27785;
  assign n31297 = n31213 & n31242;
  assign n31299 = n31298 ^ n31297;
  assign n31295 = n31276 ^ n31268;
  assign n31294 = n31262 ^ n31250;
  assign n31296 = n31295 ^ n31294;
  assign n31300 = n31299 ^ n31296;
  assign n31306 = n30600 ^ n27766;
  assign n31307 = n31306 ^ n31262;
  assign n31303 = n31193 & n31245;
  assign n31304 = n31303 ^ n31279;
  assign n31301 = n31283 ^ n31257;
  assign n31302 = n31301 ^ n31253;
  assign n31305 = n31304 ^ n31302;
  assign n31308 = n31307 ^ n31305;
  assign n31314 = n30608 ^ n27794;
  assign n31312 = n31261 ^ n31250;
  assign n31309 = n31224 & n31238;
  assign n31310 = n31309 ^ n31297;
  assign n31311 = n31310 ^ n31301;
  assign n31313 = n31312 ^ n31311;
  assign n31315 = n31314 ^ n31313;
  assign n31319 = n30613 ^ n27811;
  assign n31317 = n31310 ^ n31277;
  assign n31316 = n31282 ^ n31253;
  assign n31318 = n31317 ^ n31316;
  assign n31320 = n31319 ^ n31318;
  assign n31440 = n30734 ^ n28875;
  assign n31365 = n30118 ^ n30089;
  assign n31364 = n28937 ^ n27468;
  assign n31366 = n31365 ^ n31364;
  assign n31354 = n27538 ^ n27385;
  assign n31355 = n31354 ^ n27554;
  assign n31353 = n28901 ^ n26976;
  assign n31356 = n31355 ^ n31353;
  assign n31350 = n27558 ^ n27538;
  assign n31351 = n31350 ^ n27456;
  assign n31349 = n28929 ^ n27527;
  assign n31352 = n31351 ^ n31349;
  assign n31357 = n31356 ^ n31352;
  assign n31367 = n31366 ^ n31357;
  assign n31328 = n28892 ^ n27496;
  assign n31326 = n27488 ^ n27444;
  assign n31327 = n31326 ^ n30084;
  assign n31329 = n31328 ^ n31327;
  assign n31360 = n31352 ^ n31329;
  assign n31332 = n27558 ^ n27461;
  assign n31333 = n31332 ^ n30073;
  assign n31331 = n28874 ^ n27547;
  assign n31334 = n31333 ^ n31331;
  assign n31323 = n30078 ^ n27385;
  assign n31324 = n31323 ^ n27542;
  assign n31321 = n27502 ^ n27468;
  assign n31322 = n31321 ^ n28864;
  assign n31325 = n31324 ^ n31322;
  assign n31347 = n31334 ^ n31325;
  assign n31344 = n30097 ^ n27518;
  assign n31342 = n27468 ^ n27401;
  assign n31343 = n31342 ^ n28911;
  assign n31345 = n31344 ^ n31343;
  assign n31338 = n30089 ^ n27488;
  assign n31339 = n31338 ^ n27420;
  assign n31336 = n27570 ^ n27468;
  assign n31337 = n31336 ^ n28920;
  assign n31340 = n31339 ^ n31337;
  assign n31341 = n31340 ^ n30094;
  assign n31346 = n31345 ^ n31341;
  assign n31348 = n31347 ^ n31346;
  assign n31403 = n31360 ^ n31348;
  assign n31330 = n31329 ^ n31325;
  assign n31377 = n31356 ^ n31329;
  assign n31380 = n31377 ^ n31347;
  assign n31381 = n31330 & n31380;
  assign n31361 = n31360 ^ n31346;
  assign n31362 = n31347 & n31361;
  assign n31382 = n31381 ^ n31362;
  assign n31404 = n31403 ^ n31382;
  assign n31398 = n31366 ^ n31348;
  assign n31399 = n31367 ^ n31340;
  assign n31335 = n31334 ^ n31329;
  assign n31400 = n31399 ^ n31335;
  assign n31401 = n31398 & n31400;
  assign n31370 = n31340 ^ n31334;
  assign n31371 = n31370 ^ n31330;
  assign n31372 = n31348 & n31371;
  assign n31402 = n31401 ^ n31372;
  assign n31405 = n31404 ^ n31402;
  assign n31358 = n31357 ^ n31348;
  assign n31374 = n31358 ^ n31335;
  assign n31368 = n31367 ^ n31325;
  assign n31369 = n31366 & n31368;
  assign n31373 = n31372 ^ n31369;
  assign n31375 = n31374 ^ n31373;
  assign n31359 = n31335 & n31358;
  assign n31363 = n31362 ^ n31359;
  assign n31376 = n31375 ^ n31363;
  assign n31411 = n31405 ^ n31376;
  assign n31385 = ~n31340 & n31367;
  assign n31378 = n31377 ^ n31346;
  assign n31384 = n31370 & n31378;
  assign n31386 = n31385 ^ n31384;
  assign n31379 = n31378 ^ n31370;
  assign n31383 = n31382 ^ n31379;
  assign n31387 = n31386 ^ n31383;
  assign n31406 = n31387 & n31405;
  assign n31412 = n31411 ^ n31406;
  assign n31389 = n31368 ^ n31347;
  assign n31388 = n31378 ^ n31367;
  assign n31393 = n31389 ^ n31388;
  assign n31390 = n31388 & n31389;
  assign n31391 = n31390 ^ n31384;
  assign n31392 = n31391 ^ n31363;
  assign n31394 = n31393 ^ n31392;
  assign n31409 = n31394 & n31405;
  assign n31410 = ~n31376 & n31409;
  assign n31413 = n31412 ^ n31410;
  assign n31436 = n31367 & n31413;
  assign n31395 = n31394 ^ n31387;
  assign n31407 = n31406 ^ n31395;
  assign n31396 = n31387 & n31395;
  assign n31397 = n31376 & n31396;
  assign n31408 = n31407 ^ n31397;
  assign n31435 = n31400 & n31408;
  assign n31437 = n31436 ^ n31435;
  assign n31418 = n31406 ^ n31376;
  assign n31419 = n31395 & n31418;
  assign n31420 = n31419 ^ n31394;
  assign n31415 = n31406 ^ n31394;
  assign n31416 = n31411 & n31415;
  assign n31417 = n31416 ^ n31376;
  assign n31421 = n31420 ^ n31417;
  assign n31433 = n31361 & n31421;
  assign n31414 = n31413 ^ n31408;
  assign n31422 = n31421 ^ n31414;
  assign n31432 = n31380 & n31422;
  assign n31434 = n31433 ^ n31432;
  assign n31438 = n31437 ^ n31434;
  assign n31429 = n31420 ^ n31408;
  assign n31430 = n31371 & n31429;
  assign n31426 = n31417 ^ n31413;
  assign n31427 = n31378 & n31426;
  assign n31424 = n31347 & n31421;
  assign n31423 = n31330 & n31422;
  assign n31425 = n31424 ^ n31423;
  assign n31428 = n31427 ^ n31425;
  assign n31431 = n31430 ^ n31428;
  assign n31439 = n31438 ^ n31431;
  assign n31441 = n31440 ^ n31439;
  assign n31449 = n30743 ^ n28930;
  assign n31447 = n31435 ^ n31425;
  assign n31444 = n31348 & n31429;
  assign n31442 = n31398 & n31408;
  assign n31443 = n31442 ^ n31430;
  assign n31445 = n31444 ^ n31443;
  assign n31446 = n31445 ^ n31434;
  assign n31448 = n31447 ^ n31446;
  assign n31450 = n31449 ^ n31448;
  assign n31462 = n30756 ^ n28902;
  assign n31463 = n31462 ^ n31424;
  assign n31459 = n31335 & n31414;
  assign n31457 = n31370 & n31426;
  assign n31456 = n31358 & n31414;
  assign n31458 = n31457 ^ n31456;
  assign n31460 = n31459 ^ n31458;
  assign n31453 = n31389 & n31417;
  assign n31451 = n31366 & n31420;
  assign n31452 = n31451 ^ n31444;
  assign n31454 = n31453 ^ n31452;
  assign n31455 = n31454 ^ n31433;
  assign n31461 = n31460 ^ n31455;
  assign n31464 = n31463 ^ n31461;
  assign n31466 = n30760 ^ n28865;
  assign n31467 = n31466 ^ n31445;
  assign n31465 = n31437 ^ n31428;
  assign n31468 = n31467 ^ n31465;
  assign n31473 = n30767 ^ n28912;
  assign n31472 = n31388 & n31417;
  assign n31474 = n31473 ^ n31472;
  assign n31470 = n31451 ^ n31443;
  assign n31469 = n31437 ^ n31425;
  assign n31471 = n31470 ^ n31469;
  assign n31475 = n31474 ^ n31471;
  assign n31481 = n30775 ^ n28893;
  assign n31482 = n31481 ^ n31437;
  assign n31478 = n31368 & n31420;
  assign n31479 = n31478 ^ n31454;
  assign n31476 = n31458 ^ n31432;
  assign n31477 = n31476 ^ n31428;
  assign n31480 = n31479 ^ n31477;
  assign n31483 = n31482 ^ n31480;
  assign n31489 = n30783 ^ n28921;
  assign n31487 = n31436 ^ n31425;
  assign n31484 = n31399 & n31413;
  assign n31485 = n31484 ^ n31472;
  assign n31486 = n31485 ^ n31476;
  assign n31488 = n31487 ^ n31486;
  assign n31490 = n31489 ^ n31488;
  assign n31494 = n30788 ^ n28938;
  assign n31492 = n31485 ^ n31452;
  assign n31491 = n31457 ^ n31428;
  assign n31493 = n31492 ^ n31491;
  assign n31495 = n31494 ^ n31493;
  assign n31608 = n30910 ^ n29872;
  assign n31533 = n29895 ^ n29711;
  assign n31532 = n30444 ^ n29790;
  assign n31534 = n31533 ^ n31532;
  assign n31523 = n29886 ^ n29757;
  assign n31522 = n30432 ^ n29770;
  assign n31524 = n31523 ^ n31522;
  assign n31520 = n29891 ^ n29684;
  assign n31519 = n30470 ^ n29745;
  assign n31521 = n31520 ^ n31519;
  assign n31525 = n31524 ^ n31521;
  assign n31535 = n31534 ^ n31525;
  assign n31501 = n29883 ^ n29731;
  assign n31500 = n30451 ^ n29632;
  assign n31502 = n31501 ^ n31500;
  assign n31528 = n31521 ^ n31502;
  assign n31505 = n29872 ^ n29600;
  assign n31504 = n30465 ^ n29674;
  assign n31506 = n31505 ^ n31504;
  assign n31498 = n29869 ^ n29774;
  assign n31496 = n30966 ^ n29470;
  assign n31497 = n31496 ^ n29349;
  assign n31499 = n31498 ^ n31497;
  assign n31517 = n31506 ^ n31499;
  assign n31514 = n29876 ^ n29591;
  assign n31513 = n30989 ^ n29734;
  assign n31515 = n31514 ^ n31513;
  assign n31510 = n29879 ^ n29660;
  assign n31508 = n30981 ^ n29705;
  assign n31509 = n31508 ^ n29701;
  assign n31511 = n31510 ^ n31509;
  assign n31512 = n31511 ^ n29723;
  assign n31516 = n31515 ^ n31512;
  assign n31518 = n31517 ^ n31516;
  assign n31571 = n31528 ^ n31518;
  assign n31503 = n31502 ^ n31499;
  assign n31545 = n31524 ^ n31502;
  assign n31548 = n31545 ^ n31517;
  assign n31549 = n31503 & n31548;
  assign n31529 = n31528 ^ n31516;
  assign n31530 = n31517 & n31529;
  assign n31550 = n31549 ^ n31530;
  assign n31572 = n31571 ^ n31550;
  assign n31566 = n31535 ^ n31511;
  assign n31507 = n31506 ^ n31502;
  assign n31567 = n31566 ^ n31507;
  assign n31568 = n31534 ^ n31518;
  assign n31569 = ~n31567 & n31568;
  assign n31538 = n31511 ^ n31506;
  assign n31539 = n31538 ^ n31503;
  assign n31540 = n31518 & ~n31539;
  assign n31570 = n31569 ^ n31540;
  assign n31573 = n31572 ^ n31570;
  assign n31526 = n31525 ^ n31518;
  assign n31542 = n31526 ^ n31507;
  assign n31536 = n31535 ^ n31499;
  assign n31537 = n31534 & n31536;
  assign n31541 = n31540 ^ n31537;
  assign n31543 = n31542 ^ n31541;
  assign n31527 = n31507 & n31526;
  assign n31531 = n31530 ^ n31527;
  assign n31544 = n31543 ^ n31531;
  assign n31579 = n31573 ^ n31544;
  assign n31553 = n31511 & n31535;
  assign n31546 = n31545 ^ n31516;
  assign n31552 = ~n31538 & n31546;
  assign n31554 = n31553 ^ n31552;
  assign n31547 = n31546 ^ n31538;
  assign n31551 = n31550 ^ n31547;
  assign n31555 = n31554 ^ n31551;
  assign n31574 = ~n31555 & n31573;
  assign n31580 = n31579 ^ n31574;
  assign n31557 = n31546 ^ n31535;
  assign n31556 = n31536 ^ n31517;
  assign n31561 = n31557 ^ n31556;
  assign n31558 = n31556 & n31557;
  assign n31559 = n31558 ^ n31552;
  assign n31560 = n31559 ^ n31531;
  assign n31562 = n31561 ^ n31560;
  assign n31577 = ~n31544 & n31573;
  assign n31578 = n31562 & n31577;
  assign n31581 = n31580 ^ n31578;
  assign n31604 = n31535 & n31581;
  assign n31563 = n31562 ^ n31555;
  assign n31575 = n31574 ^ n31563;
  assign n31564 = ~n31555 & ~n31563;
  assign n31565 = n31544 & n31564;
  assign n31576 = n31575 ^ n31565;
  assign n31603 = ~n31567 & ~n31576;
  assign n31605 = n31604 ^ n31603;
  assign n31586 = n31574 ^ n31562;
  assign n31587 = n31579 & n31586;
  assign n31588 = n31587 ^ n31544;
  assign n31583 = n31574 ^ n31544;
  assign n31584 = ~n31563 & n31583;
  assign n31585 = n31584 ^ n31562;
  assign n31589 = n31588 ^ n31585;
  assign n31601 = n31529 & n31589;
  assign n31582 = n31581 ^ n31576;
  assign n31590 = n31589 ^ n31582;
  assign n31600 = n31548 & ~n31590;
  assign n31602 = n31601 ^ n31600;
  assign n31606 = n31605 ^ n31602;
  assign n31597 = n31585 ^ n31576;
  assign n31598 = ~n31539 & ~n31597;
  assign n31594 = n31588 ^ n31581;
  assign n31595 = n31546 & n31594;
  assign n31592 = n31517 & n31589;
  assign n31591 = n31503 & ~n31590;
  assign n31593 = n31592 ^ n31591;
  assign n31596 = n31595 ^ n31593;
  assign n31599 = n31598 ^ n31596;
  assign n31607 = n31606 ^ n31599;
  assign n31609 = n31608 ^ n31607;
  assign n31617 = n30919 ^ n29891;
  assign n31615 = n31603 ^ n31593;
  assign n31612 = n31518 & ~n31597;
  assign n31610 = n31568 & ~n31576;
  assign n31611 = n31610 ^ n31598;
  assign n31613 = n31612 ^ n31611;
  assign n31614 = n31613 ^ n31602;
  assign n31616 = n31615 ^ n31614;
  assign n31618 = n31617 ^ n31616;
  assign n31629 = n31507 & ~n31582;
  assign n31627 = ~n31538 & n31594;
  assign n31626 = n31526 & ~n31582;
  assign n31628 = n31627 ^ n31626;
  assign n31630 = n31629 ^ n31628;
  assign n31631 = n31630 ^ n30932;
  assign n31624 = n31592 ^ n29886;
  assign n31621 = n31556 & n31588;
  assign n31619 = n31534 & n31585;
  assign n31620 = n31619 ^ n31612;
  assign n31622 = n31621 ^ n31620;
  assign n31623 = n31622 ^ n31601;
  assign n31625 = n31624 ^ n31623;
  assign n31632 = n31631 ^ n31625;
  assign n31635 = n30936 ^ n29869;
  assign n31633 = n31613 ^ n31605;
  assign n31634 = n31633 ^ n31596;
  assign n31636 = n31635 ^ n31634;
  assign n31640 = n31557 & n31588;
  assign n31641 = n31640 ^ n29876;
  assign n31639 = n31619 ^ n31611;
  assign n31642 = n31641 ^ n31639;
  assign n31637 = n31605 ^ n31593;
  assign n31638 = n31637 ^ n30943;
  assign n31643 = n31642 ^ n31638;
  assign n31649 = n31605 ^ n29883;
  assign n31647 = n31536 & n31585;
  assign n31648 = n31647 ^ n31622;
  assign n31650 = n31649 ^ n31648;
  assign n31644 = n31628 ^ n31600;
  assign n31645 = n31644 ^ n31596;
  assign n31646 = n31645 ^ n30951;
  assign n31651 = n31650 ^ n31646;
  assign n31657 = n30959 ^ n29879;
  assign n31655 = n31604 ^ n31593;
  assign n31652 = ~n31566 & n31581;
  assign n31653 = n31652 ^ n31640;
  assign n31654 = n31653 ^ n31644;
  assign n31656 = n31655 ^ n31654;
  assign n31658 = n31657 ^ n31656;
  assign n31662 = n30964 ^ n29895;
  assign n31660 = n31653 ^ n31620;
  assign n31659 = n31627 ^ n31596;
  assign n31661 = n31660 ^ n31659;
  assign n31663 = n31662 ^ n31661;
  assign n31781 = n31086 ^ n26619;
  assign n31708 = n26651 ^ n26380;
  assign n31706 = n26281 ^ n26247;
  assign n31707 = n31706 ^ n31159;
  assign n31709 = n31708 ^ n31707;
  assign n31694 = n31172 ^ n26391;
  assign n31695 = n31694 ^ n26633;
  assign n31696 = n31695 ^ n26259;
  assign n31692 = n26640 ^ n26405;
  assign n31690 = n26420 ^ n26342;
  assign n31691 = n31690 ^ n26400;
  assign n31693 = n31692 ^ n31691;
  assign n31697 = n31696 ^ n31693;
  assign n31710 = n31709 ^ n31697;
  assign n31682 = n26680 ^ n26301;
  assign n31680 = n31159 ^ n26293;
  assign n31679 = n26286 ^ n23285;
  assign n31681 = n31680 ^ n31679;
  assign n31683 = n31682 ^ n31681;
  assign n31721 = n31710 ^ n31683;
  assign n31673 = n26401 ^ n26234;
  assign n31674 = n31673 ^ n31188;
  assign n31675 = n31674 ^ n26616;
  assign n31668 = n26294 ^ n26104;
  assign n31669 = n31668 ^ n25178;
  assign n31670 = n31669 ^ n26323;
  assign n31671 = n31670 ^ n26664;
  assign n31676 = n31675 ^ n31671;
  assign n31722 = n31721 ^ n31676;
  assign n31744 = ~n31683 & n31710;
  assign n31704 = n31696 ^ n31671;
  assign n31686 = n31167 ^ n26314;
  assign n31685 = n26325 ^ n26227;
  assign n31687 = n31686 ^ n31685;
  assign n31678 = n26673 ^ n26330;
  assign n31684 = n31683 ^ n31678;
  assign n31688 = n31687 ^ n31684;
  assign n31705 = n31704 ^ n31688;
  assign n31715 = n31683 ^ n31675;
  assign n31716 = n31705 & n31715;
  assign n31745 = n31744 ^ n31716;
  assign n31742 = n31715 ^ n31705;
  assign n31664 = n31176 ^ n31142;
  assign n31665 = n31664 ^ n26248;
  assign n31666 = n31665 ^ n26413;
  assign n31667 = n31666 ^ n26606;
  assign n31672 = n31671 ^ n31667;
  assign n31677 = n31675 ^ n31667;
  assign n31729 = n31704 ^ n31677;
  assign n31730 = n31672 & n31729;
  assign n31700 = n31693 ^ n31671;
  assign n31701 = n31700 ^ n31688;
  assign n31702 = n31677 & n31701;
  assign n31731 = n31730 ^ n31702;
  assign n31743 = n31742 ^ n31731;
  assign n31746 = n31745 ^ n31743;
  assign n31712 = n31710 ^ n31667;
  assign n31713 = n31712 ^ n31677;
  assign n31711 = n31710 ^ n31705;
  assign n31719 = n31713 ^ n31711;
  assign n31714 = n31711 & n31713;
  assign n31717 = n31716 ^ n31714;
  assign n31689 = n31688 ^ n31677;
  assign n31698 = n31697 ^ n31689;
  assign n31699 = n31676 & n31698;
  assign n31703 = n31702 ^ n31699;
  assign n31718 = n31717 ^ n31703;
  assign n31720 = n31719 ^ n31718;
  assign n31752 = n31746 ^ n31720;
  assign n31728 = n31700 ^ n31689;
  assign n31732 = n31731 ^ n31728;
  assign n31725 = n31715 ^ n31672;
  assign n31726 = n31689 & n31725;
  assign n31723 = n31709 ^ n31689;
  assign n31724 = n31722 & n31723;
  assign n31727 = n31726 ^ n31724;
  assign n31733 = n31732 ^ n31727;
  assign n31747 = n31733 & n31746;
  assign n31753 = n31752 ^ n31747;
  assign n31736 = n31698 ^ n31676;
  assign n31734 = n31709 & n31712;
  assign n31735 = n31734 ^ n31726;
  assign n31737 = n31736 ^ n31735;
  assign n31738 = n31737 ^ n31703;
  assign n31750 = n31738 & n31746;
  assign n31751 = ~n31720 & n31750;
  assign n31754 = n31753 ^ n31751;
  assign n31777 = n31722 & n31754;
  assign n31741 = n31738 ^ n31733;
  assign n31748 = n31747 ^ n31741;
  assign n31739 = n31733 & ~n31738;
  assign n31740 = n31720 & n31739;
  assign n31749 = n31748 ^ n31740;
  assign n31776 = n31710 & n31749;
  assign n31778 = n31777 ^ n31776;
  assign n31759 = n31747 ^ n31738;
  assign n31760 = n31752 & n31759;
  assign n31761 = n31760 ^ n31720;
  assign n31756 = n31747 ^ n31720;
  assign n31757 = n31741 & n31756;
  assign n31758 = n31757 ^ n31738;
  assign n31762 = n31761 ^ n31758;
  assign n31774 = n31701 & n31762;
  assign n31755 = n31754 ^ n31749;
  assign n31763 = n31762 ^ n31755;
  assign n31773 = n31729 & n31763;
  assign n31775 = n31774 ^ n31773;
  assign n31779 = n31778 ^ n31775;
  assign n31770 = n31761 ^ n31754;
  assign n31771 = n31725 & n31770;
  assign n31767 = n31758 ^ n31749;
  assign n31768 = n31705 & n31767;
  assign n31765 = n31677 & n31762;
  assign n31764 = n31672 & n31763;
  assign n31766 = n31765 ^ n31764;
  assign n31769 = n31768 ^ n31766;
  assign n31772 = n31771 ^ n31769;
  assign n31780 = n31779 ^ n31772;
  assign n31782 = n31781 ^ n31780;
  assign n31790 = n31095 ^ n26643;
  assign n31788 = n31777 ^ n31766;
  assign n31785 = n31689 & n31770;
  assign n31783 = n31723 & n31754;
  assign n31784 = n31783 ^ n31771;
  assign n31786 = n31785 ^ n31784;
  assign n31787 = n31786 ^ n31775;
  assign n31789 = n31788 ^ n31787;
  assign n31791 = n31790 ^ n31789;
  assign n31802 = n31676 & n31755;
  assign n31800 = n31698 & n31755;
  assign n31799 = n31715 & n31767;
  assign n31801 = n31800 ^ n31799;
  assign n31803 = n31802 ^ n31801;
  assign n31804 = n31803 ^ n31108;
  assign n31797 = n31765 ^ n26636;
  assign n31794 = n31713 & n31758;
  assign n31792 = n31709 & n31761;
  assign n31793 = n31792 ^ n31785;
  assign n31795 = n31794 ^ n31793;
  assign n31796 = n31795 ^ n31774;
  assign n31798 = n31797 ^ n31796;
  assign n31805 = n31804 ^ n31798;
  assign n31808 = n31112 ^ n26609;
  assign n31806 = n31786 ^ n31778;
  assign n31807 = n31806 ^ n31769;
  assign n31809 = n31808 ^ n31807;
  assign n31813 = n31711 & n31758;
  assign n31814 = n31813 ^ n26676;
  assign n31812 = n31792 ^ n31784;
  assign n31815 = n31814 ^ n31812;
  assign n31810 = n31778 ^ n31766;
  assign n31811 = n31810 ^ n31119;
  assign n31816 = n31815 ^ n31811;
  assign n31822 = n31778 ^ n26667;
  assign n31820 = n31712 & n31761;
  assign n31821 = n31820 ^ n31795;
  assign n31823 = n31822 ^ n31821;
  assign n31817 = n31801 ^ n31773;
  assign n31818 = n31817 ^ n31769;
  assign n31819 = n31818 ^ n31127;
  assign n31824 = n31823 ^ n31819;
  assign n31830 = n31135 ^ n26683;
  assign n31828 = n31776 ^ n31766;
  assign n31825 = n31721 & n31749;
  assign n31826 = n31825 ^ n31813;
  assign n31827 = n31826 ^ n31817;
  assign n31829 = n31828 ^ n31827;
  assign n31831 = n31830 ^ n31829;
  assign n31835 = n31140 ^ n26654;
  assign n31833 = n31826 ^ n31793;
  assign n31832 = n31799 ^ n31769;
  assign n31834 = n31833 ^ n31832;
  assign n31836 = n31835 ^ n31834;
  assign n31953 = n31265 ^ n27749;
  assign n31876 = n31336 ^ n27116;
  assign n31877 = n31876 ^ n27481;
  assign n31878 = n31877 ^ n27574;
  assign n31879 = n31878 ^ n27810;
  assign n31867 = n30103 ^ n27104;
  assign n31866 = n27774 ^ n27527;
  assign n31868 = n31867 ^ n31866;
  assign n31864 = n30074 ^ n27533;
  assign n31863 = n27802 ^ n27547;
  assign n31865 = n31864 ^ n31863;
  assign n31869 = n31868 ^ n31865;
  assign n31880 = n31879 ^ n31869;
  assign n31843 = n27513 ^ n27444;
  assign n31842 = n27496 ^ n27410;
  assign n31844 = n31843 ^ n31842;
  assign n31841 = n27765 ^ n27401;
  assign n31845 = n31844 ^ n31841;
  assign n31872 = n31865 ^ n31845;
  assign n31848 = n27747 ^ n27468;
  assign n31847 = n30119 ^ n27548;
  assign n31849 = n31848 ^ n31847;
  assign n31839 = n27737 ^ n26976;
  assign n31837 = n31321 ^ n27117;
  assign n31838 = n31837 ^ n30107;
  assign n31840 = n31839 ^ n31838;
  assign n31861 = n31849 ^ n31840;
  assign n31858 = n27518 ^ n27241;
  assign n31857 = n31342 ^ n27505;
  assign n31859 = n31858 ^ n31857;
  assign n31855 = n27784 ^ n27502;
  assign n31853 = n27793 ^ n27496;
  assign n31851 = n31336 ^ n27476;
  assign n31852 = n31851 ^ n30085;
  assign n31854 = n31853 ^ n31852;
  assign n31856 = n31855 ^ n31854;
  assign n31860 = n31859 ^ n31856;
  assign n31862 = n31861 ^ n31860;
  assign n31916 = n31872 ^ n31862;
  assign n31846 = n31845 ^ n31840;
  assign n31890 = n31868 ^ n31845;
  assign n31893 = n31890 ^ n31861;
  assign n31894 = n31846 & n31893;
  assign n31873 = n31872 ^ n31860;
  assign n31874 = n31861 & n31873;
  assign n31895 = n31894 ^ n31874;
  assign n31917 = n31916 ^ n31895;
  assign n31911 = n31880 ^ n31854;
  assign n31850 = n31849 ^ n31845;
  assign n31912 = n31911 ^ n31850;
  assign n31913 = n31879 ^ n31862;
  assign n31914 = n31912 & n31913;
  assign n31883 = n31854 ^ n31849;
  assign n31884 = n31883 ^ n31846;
  assign n31885 = n31862 & n31884;
  assign n31915 = n31914 ^ n31885;
  assign n31918 = n31917 ^ n31915;
  assign n31870 = n31869 ^ n31862;
  assign n31887 = n31870 ^ n31850;
  assign n31881 = n31880 ^ n31840;
  assign n31882 = n31879 & n31881;
  assign n31886 = n31885 ^ n31882;
  assign n31888 = n31887 ^ n31886;
  assign n31871 = n31850 & n31870;
  assign n31875 = n31874 ^ n31871;
  assign n31889 = n31888 ^ n31875;
  assign n31924 = n31918 ^ n31889;
  assign n31898 = ~n31854 & n31880;
  assign n31891 = n31890 ^ n31860;
  assign n31897 = n31883 & n31891;
  assign n31899 = n31898 ^ n31897;
  assign n31892 = n31891 ^ n31883;
  assign n31896 = n31895 ^ n31892;
  assign n31900 = n31899 ^ n31896;
  assign n31919 = n31900 & n31918;
  assign n31925 = n31924 ^ n31919;
  assign n31902 = n31891 ^ n31880;
  assign n31901 = n31881 ^ n31861;
  assign n31906 = n31902 ^ n31901;
  assign n31903 = n31901 & n31902;
  assign n31904 = n31903 ^ n31897;
  assign n31905 = n31904 ^ n31875;
  assign n31907 = n31906 ^ n31905;
  assign n31922 = n31907 & n31918;
  assign n31923 = ~n31889 & n31922;
  assign n31926 = n31925 ^ n31923;
  assign n31949 = n31880 & n31926;
  assign n31908 = n31907 ^ n31900;
  assign n31920 = n31919 ^ n31908;
  assign n31909 = n31900 & n31908;
  assign n31910 = n31889 & n31909;
  assign n31921 = n31920 ^ n31910;
  assign n31948 = n31912 & n31921;
  assign n31950 = n31949 ^ n31948;
  assign n31931 = n31919 ^ n31889;
  assign n31932 = n31908 & n31931;
  assign n31933 = n31932 ^ n31907;
  assign n31928 = n31919 ^ n31907;
  assign n31929 = n31924 & n31928;
  assign n31930 = n31929 ^ n31889;
  assign n31934 = n31933 ^ n31930;
  assign n31946 = n31873 & n31934;
  assign n31927 = n31926 ^ n31921;
  assign n31935 = n31934 ^ n31927;
  assign n31945 = n31893 & n31935;
  assign n31947 = n31946 ^ n31945;
  assign n31951 = n31950 ^ n31947;
  assign n31942 = n31933 ^ n31921;
  assign n31943 = n31884 & n31942;
  assign n31939 = n31930 ^ n31926;
  assign n31940 = n31891 & n31939;
  assign n31937 = n31861 & n31934;
  assign n31936 = n31846 & n31935;
  assign n31938 = n31937 ^ n31936;
  assign n31941 = n31940 ^ n31938;
  assign n31944 = n31943 ^ n31941;
  assign n31952 = n31951 ^ n31944;
  assign n31954 = n31953 ^ n31952;
  assign n31962 = n31274 ^ n27804;
  assign n31960 = n31948 ^ n31938;
  assign n31957 = n31862 & n31942;
  assign n31955 = n31913 & n31921;
  assign n31956 = n31955 ^ n31943;
  assign n31958 = n31957 ^ n31956;
  assign n31959 = n31958 ^ n31947;
  assign n31961 = n31960 ^ n31959;
  assign n31963 = n31962 ^ n31961;
  assign n31974 = n31850 & n31927;
  assign n31972 = n31883 & n31939;
  assign n31971 = n31870 & n31927;
  assign n31973 = n31972 ^ n31971;
  assign n31975 = n31974 ^ n31973;
  assign n31976 = n31975 ^ n31287;
  assign n31969 = n31937 ^ n27776;
  assign n31966 = n31901 & n31930;
  assign n31964 = n31879 & n31933;
  assign n31965 = n31964 ^ n31957;
  assign n31967 = n31966 ^ n31965;
  assign n31968 = n31967 ^ n31946;
  assign n31970 = n31969 ^ n31968;
  assign n31977 = n31976 ^ n31970;
  assign n31980 = n31291 ^ n27739;
  assign n31978 = n31958 ^ n31950;
  assign n31979 = n31978 ^ n31941;
  assign n31981 = n31980 ^ n31979;
  assign n31985 = n31902 & n31930;
  assign n31986 = n31985 ^ n27786;
  assign n31984 = n31964 ^ n31956;
  assign n31987 = n31986 ^ n31984;
  assign n31982 = n31950 ^ n31938;
  assign n31983 = n31982 ^ n31298;
  assign n31988 = n31987 ^ n31983;
  assign n31994 = n31950 ^ n27767;
  assign n31992 = n31881 & n31933;
  assign n31993 = n31992 ^ n31967;
  assign n31995 = n31994 ^ n31993;
  assign n31989 = n31973 ^ n31945;
  assign n31990 = n31989 ^ n31941;
  assign n31991 = n31990 ^ n31306;
  assign n31996 = n31995 ^ n31991;
  assign n32002 = n31314 ^ n27795;
  assign n32000 = n31949 ^ n31938;
  assign n31997 = n31911 & n31926;
  assign n31998 = n31997 ^ n31985;
  assign n31999 = n31998 ^ n31989;
  assign n32001 = n32000 ^ n31999;
  assign n32003 = n32002 ^ n32001;
  assign n32007 = n31319 ^ n27812;
  assign n32005 = n31998 ^ n31965;
  assign n32004 = n31972 ^ n31941;
  assign n32006 = n32005 ^ n32004;
  assign n32008 = n32007 ^ n32006;
  assign n32125 = n31440 ^ n28876;
  assign n32052 = n30816 ^ n30808;
  assign n32051 = n28938 ^ n28247;
  assign n32053 = n32052 ^ n32051;
  assign n32040 = n28902 ^ n28504;
  assign n32038 = n28675 ^ n28498;
  assign n32039 = n32038 ^ n30267;
  assign n32041 = n32040 ^ n32039;
  assign n32036 = n28930 ^ n28651;
  assign n32034 = n28675 ^ n28658;
  assign n32035 = n32034 ^ n30803;
  assign n32037 = n32036 ^ n32035;
  assign n32042 = n32041 ^ n32037;
  assign n32054 = n32053 ^ n32042;
  assign n32025 = n30816 ^ n28614;
  assign n32026 = n32025 ^ n30257;
  assign n32024 = n28921 ^ n28601;
  assign n32027 = n32026 ^ n32024;
  assign n32065 = n32054 ^ n32027;
  assign n32020 = n28875 ^ n28574;
  assign n32018 = n28658 ^ n28585;
  assign n32019 = n32018 ^ n30795;
  assign n32021 = n32020 ^ n32019;
  assign n32015 = n28893 ^ n28533;
  assign n32013 = n28614 ^ n28562;
  assign n32014 = n32013 ^ n30828;
  assign n32016 = n32015 ^ n32014;
  assign n32022 = n32021 ^ n32016;
  assign n32066 = n32065 ^ n32022;
  assign n32088 = ~n32027 & n32054;
  assign n32049 = n32041 ^ n32016;
  assign n32030 = n30822 ^ n28637;
  assign n32029 = n28912 ^ n28628;
  assign n32031 = n32030 ^ n32029;
  assign n32028 = n32027 ^ n30815;
  assign n32032 = n32031 ^ n32028;
  assign n32050 = n32049 ^ n32032;
  assign n32059 = n32027 ^ n32021;
  assign n32060 = n32050 & n32059;
  assign n32089 = n32088 ^ n32060;
  assign n32086 = n32059 ^ n32050;
  assign n32010 = n30790 ^ n28498;
  assign n32011 = n32010 ^ n30272;
  assign n32009 = n28865 ^ n28248;
  assign n32012 = n32011 ^ n32009;
  assign n32017 = n32016 ^ n32012;
  assign n32023 = n32021 ^ n32012;
  assign n32073 = n32049 ^ n32023;
  assign n32074 = n32017 & n32073;
  assign n32045 = n32037 ^ n32016;
  assign n32046 = n32045 ^ n32032;
  assign n32047 = n32023 & n32046;
  assign n32075 = n32074 ^ n32047;
  assign n32087 = n32086 ^ n32075;
  assign n32090 = n32089 ^ n32087;
  assign n32056 = n32054 ^ n32012;
  assign n32057 = n32056 ^ n32023;
  assign n32055 = n32054 ^ n32050;
  assign n32063 = n32057 ^ n32055;
  assign n32058 = n32055 & n32057;
  assign n32061 = n32060 ^ n32058;
  assign n32033 = n32032 ^ n32023;
  assign n32043 = n32042 ^ n32033;
  assign n32044 = n32022 & n32043;
  assign n32048 = n32047 ^ n32044;
  assign n32062 = n32061 ^ n32048;
  assign n32064 = n32063 ^ n32062;
  assign n32096 = n32090 ^ n32064;
  assign n32072 = n32045 ^ n32033;
  assign n32076 = n32075 ^ n32072;
  assign n32069 = n32059 ^ n32017;
  assign n32070 = n32033 & n32069;
  assign n32067 = n32053 ^ n32033;
  assign n32068 = n32066 & n32067;
  assign n32071 = n32070 ^ n32068;
  assign n32077 = n32076 ^ n32071;
  assign n32091 = n32077 & n32090;
  assign n32097 = n32096 ^ n32091;
  assign n32080 = n32043 ^ n32022;
  assign n32078 = n32053 & n32056;
  assign n32079 = n32078 ^ n32070;
  assign n32081 = n32080 ^ n32079;
  assign n32082 = n32081 ^ n32048;
  assign n32094 = n32082 & n32090;
  assign n32095 = ~n32064 & n32094;
  assign n32098 = n32097 ^ n32095;
  assign n32121 = n32066 & n32098;
  assign n32085 = n32082 ^ n32077;
  assign n32092 = n32091 ^ n32085;
  assign n32083 = n32077 & ~n32082;
  assign n32084 = n32064 & n32083;
  assign n32093 = n32092 ^ n32084;
  assign n32120 = n32054 & n32093;
  assign n32122 = n32121 ^ n32120;
  assign n32103 = n32091 ^ n32082;
  assign n32104 = n32096 & n32103;
  assign n32105 = n32104 ^ n32064;
  assign n32100 = n32091 ^ n32064;
  assign n32101 = n32085 & n32100;
  assign n32102 = n32101 ^ n32082;
  assign n32106 = n32105 ^ n32102;
  assign n32118 = n32046 & n32106;
  assign n32099 = n32098 ^ n32093;
  assign n32107 = n32106 ^ n32099;
  assign n32117 = n32073 & n32107;
  assign n32119 = n32118 ^ n32117;
  assign n32123 = n32122 ^ n32119;
  assign n32114 = n32105 ^ n32098;
  assign n32115 = n32069 & n32114;
  assign n32111 = n32102 ^ n32093;
  assign n32112 = n32050 & n32111;
  assign n32109 = n32023 & n32106;
  assign n32108 = n32017 & n32107;
  assign n32110 = n32109 ^ n32108;
  assign n32113 = n32112 ^ n32110;
  assign n32116 = n32115 ^ n32113;
  assign n32124 = n32123 ^ n32116;
  assign n32126 = n32125 ^ n32124;
  assign n32134 = n31449 ^ n28931;
  assign n32132 = n32121 ^ n32110;
  assign n32129 = n32033 & n32114;
  assign n32127 = n32067 & n32098;
  assign n32128 = n32127 ^ n32115;
  assign n32130 = n32129 ^ n32128;
  assign n32131 = n32130 ^ n32119;
  assign n32133 = n32132 ^ n32131;
  assign n32135 = n32134 ^ n32133;
  assign n32146 = n32022 & n32099;
  assign n32144 = n32043 & n32099;
  assign n32143 = n32059 & n32111;
  assign n32145 = n32144 ^ n32143;
  assign n32147 = n32146 ^ n32145;
  assign n32148 = n32147 ^ n31462;
  assign n32141 = n32109 ^ n28903;
  assign n32138 = n32057 & n32102;
  assign n32136 = n32053 & n32105;
  assign n32137 = n32136 ^ n32129;
  assign n32139 = n32138 ^ n32137;
  assign n32140 = n32139 ^ n32118;
  assign n32142 = n32141 ^ n32140;
  assign n32149 = n32148 ^ n32142;
  assign n32152 = n31466 ^ n28866;
  assign n32150 = n32130 ^ n32122;
  assign n32151 = n32150 ^ n32113;
  assign n32153 = n32152 ^ n32151;
  assign n32157 = n32055 & n32102;
  assign n32158 = n32157 ^ n28913;
  assign n32156 = n32136 ^ n32128;
  assign n32159 = n32158 ^ n32156;
  assign n32154 = n32122 ^ n32110;
  assign n32155 = n32154 ^ n31473;
  assign n32160 = n32159 ^ n32155;
  assign n32166 = n32122 ^ n28894;
  assign n32164 = n32056 & n32105;
  assign n32165 = n32164 ^ n32139;
  assign n32167 = n32166 ^ n32165;
  assign n32161 = n32145 ^ n32117;
  assign n32162 = n32161 ^ n32113;
  assign n32163 = n32162 ^ n31481;
  assign n32168 = n32167 ^ n32163;
  assign n32174 = n31489 ^ n28922;
  assign n32172 = n32120 ^ n32110;
  assign n32169 = n32065 & n32093;
  assign n32170 = n32169 ^ n32157;
  assign n32171 = n32170 ^ n32161;
  assign n32173 = n32172 ^ n32171;
  assign n32175 = n32174 ^ n32173;
  assign n32179 = n31494 ^ n28939;
  assign n32177 = n32170 ^ n32137;
  assign n32176 = n32143 ^ n32113;
  assign n32178 = n32177 ^ n32176;
  assign n32180 = n32179 ^ n32178;
  assign y0 = ~n26764;
  assign y1 = n26780;
  assign y2 = ~n26806;
  assign y3 = ~n26812;
  assign y4 = n26824;
  assign y5 = n26837;
  assign y6 = n26849;
  assign y7 = ~n26857;
  assign y8 = n27894;
  assign y9 = ~n27910;
  assign y10 = ~n27936;
  assign y11 = n27942;
  assign y12 = n27954;
  assign y13 = n27968;
  assign y14 = ~n27980;
  assign y15 = ~n27988;
  assign y16 = n29021;
  assign y17 = ~n29037;
  assign y18 = ~n29063;
  assign y19 = n29069;
  assign y20 = n29081;
  assign y21 = n29095;
  assign y22 = ~n29107;
  assign y23 = ~n29115;
  assign y24 = n29977;
  assign y25 = ~n29993;
  assign y26 = ~n30019;
  assign y27 = n30025;
  assign y28 = n30037;
  assign y29 = n30051;
  assign y30 = ~n30063;
  assign y31 = ~n30071;
  assign y32 = ~n30197;
  assign y33 = n30206;
  assign y34 = n30220;
  assign y35 = ~n30224;
  assign y36 = ~n30231;
  assign y37 = ~n30239;
  assign y38 = n30246;
  assign y39 = n30251;
  assign y40 = n30377;
  assign y41 = n30386;
  assign y42 = n30400;
  assign y43 = n30404;
  assign y44 = n30411;
  assign y45 = n30419;
  assign y46 = n30426;
  assign y47 = n30431;
  assign y48 = n30560;
  assign y49 = n30569;
  assign y50 = n30583;
  assign y51 = n30587;
  assign y52 = n30594;
  assign y53 = n30602;
  assign y54 = n30609;
  assign y55 = n30614;
  assign y56 = n30735;
  assign y57 = n30744;
  assign y58 = n30758;
  assign y59 = n30762;
  assign y60 = n30769;
  assign y61 = n30777;
  assign y62 = n30784;
  assign y63 = n30789;
  assign y64 = n30911;
  assign y65 = ~n30920;
  assign y66 = ~n30934;
  assign y67 = ~n30938;
  assign y68 = ~n30945;
  assign y69 = ~n30953;
  assign y70 = n30960;
  assign y71 = ~n30965;
  assign y72 = n31087;
  assign y73 = ~n31096;
  assign y74 = ~n31110;
  assign y75 = n31114;
  assign y76 = n31121;
  assign y77 = n31129;
  assign y78 = ~n31136;
  assign y79 = ~n31141;
  assign y80 = n31266;
  assign y81 = ~n31275;
  assign y82 = ~n31289;
  assign y83 = n31293;
  assign y84 = n31300;
  assign y85 = n31308;
  assign y86 = ~n31315;
  assign y87 = ~n31320;
  assign y88 = n31441;
  assign y89 = ~n31450;
  assign y90 = ~n31464;
  assign y91 = n31468;
  assign y92 = n31475;
  assign y93 = n31483;
  assign y94 = ~n31490;
  assign y95 = ~n31495;
  assign y96 = n31609;
  assign y97 = n31618;
  assign y98 = n31632;
  assign y99 = ~n31636;
  assign y100 = n31643;
  assign y101 = ~n31651;
  assign y102 = n31658;
  assign y103 = n31663;
  assign y104 = n31782;
  assign y105 = n31791;
  assign y106 = n31805;
  assign y107 = n31809;
  assign y108 = n31816;
  assign y109 = n31824;
  assign y110 = n31831;
  assign y111 = n31836;
  assign y112 = n31954;
  assign y113 = n31963;
  assign y114 = n31977;
  assign y115 = n31981;
  assign y116 = n31988;
  assign y117 = n31996;
  assign y118 = n32003;
  assign y119 = n32008;
  assign y120 = n32126;
  assign y121 = n32135;
  assign y122 = n32149;
  assign y123 = n32153;
  assign y124 = n32160;
  assign y125 = n32168;
  assign y126 = n32175;
  assign y127 = n32180;
endmodule
