module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141;
  wire n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079;
  assign n148 = ~x17 & x54;
  assign n150 = ~x8 & ~x10;
  assign n151 = ~x14 & ~x21;
  assign n152 = n150 & n151;
  assign n153 = ~x13 & n152;
  assign n154 = ~x4 & ~x9;
  assign n155 = ~x12 & n154;
  assign n156 = ~x7 & n155;
  assign n157 = n153 & n156;
  assign n159 = x12 & x13;
  assign n158 = x13 ^ x12;
  assign n160 = n159 ^ n158;
  assign n161 = n160 ^ x9;
  assign n164 = x7 ^ x6;
  assign n162 = ~x6 & ~x7;
  assign n163 = ~n159 & n162;
  assign n165 = n164 ^ n163;
  assign n166 = n165 ^ n163;
  assign n167 = ~n160 & n166;
  assign n168 = n167 ^ n163;
  assign n169 = ~n161 & n168;
  assign n170 = n169 ^ n163;
  assign n171 = n157 & ~n170;
  assign n172 = ~x5 & ~x22;
  assign n173 = ~x11 & n172;
  assign n174 = ~x18 & ~x19;
  assign n175 = x16 & n174;
  assign n176 = n175 ^ n174;
  assign n177 = n173 & n176;
  assign n178 = n171 & n177;
  assign n179 = n148 & ~n178;
  assign n149 = n148 ^ x54;
  assign n180 = n179 ^ n149;
  assign n181 = ~x0 & ~n180;
  assign n182 = x7 & ~n153;
  assign n184 = x21 ^ x14;
  assign n185 = x14 ^ x13;
  assign n186 = n184 & n185;
  assign n187 = n186 ^ x14;
  assign n188 = n150 & ~n187;
  assign n183 = x10 ^ x8;
  assign n189 = n188 ^ n183;
  assign n190 = n183 ^ x7;
  assign n191 = ~x13 & n151;
  assign n192 = n191 ^ n183;
  assign n193 = ~n183 & ~n192;
  assign n194 = n193 ^ n183;
  assign n195 = ~n190 & ~n194;
  assign n196 = n195 ^ n193;
  assign n197 = n196 ^ n183;
  assign n198 = n197 ^ n191;
  assign n199 = n189 & ~n198;
  assign n200 = n199 ^ n188;
  assign n201 = ~n182 & n200;
  assign n202 = ~x6 & n176;
  assign n203 = n155 & n202;
  assign n204 = n201 & n203;
  assign n205 = n148 & n173;
  assign n206 = n204 & n205;
  assign n207 = ~x9 & ~x11;
  assign n208 = n207 ^ n172;
  assign n209 = x54 & ~x56;
  assign n210 = n208 & n209;
  assign n211 = ~n206 & ~n210;
  assign n212 = ~n181 & n211;
  assign n213 = ~x3 & ~x129;
  assign n214 = ~n212 & n213;
  assign n215 = ~x1 & n213;
  assign n216 = ~n179 & n215;
  assign n217 = ~x5 & ~n170;
  assign n218 = x54 & n213;
  assign n219 = x17 & n218;
  assign n220 = n219 ^ n218;
  assign n221 = n176 & n220;
  assign n222 = ~x11 & ~x22;
  assign n223 = ~x4 & n222;
  assign n224 = n152 & n223;
  assign n225 = n221 & n224;
  assign n226 = ~n217 & n225;
  assign n228 = ~x5 & n226;
  assign n227 = n171 & n226;
  assign n229 = n228 ^ n227;
  assign n230 = ~n216 & ~n229;
  assign n231 = ~x15 & ~x20;
  assign n232 = x82 & ~n231;
  assign n236 = ~x42 & ~x44;
  assign n237 = ~x40 & n236;
  assign n238 = ~x38 & ~x50;
  assign n239 = n237 & n238;
  assign n240 = ~x41 & ~x46;
  assign n241 = ~x47 & ~x48;
  assign n242 = n240 & n241;
  assign n243 = ~x43 & n242;
  assign n244 = n239 & n243;
  assign n245 = ~x24 & ~x49;
  assign n246 = ~x45 & n245;
  assign n247 = n244 & n246;
  assign n248 = x82 & ~n247;
  assign n233 = x122 & x127;
  assign n234 = ~x82 & ~n233;
  assign n235 = n234 ^ x82;
  assign n249 = n248 ^ n235;
  assign n250 = ~n232 & n249;
  assign n251 = x2 & ~n250;
  assign n252 = ~x2 & n231;
  assign n253 = n246 & n252;
  assign n254 = n243 & n253;
  assign n255 = x82 & ~n254;
  assign n256 = x82 & ~n238;
  assign n257 = ~n255 & ~n256;
  assign n258 = x82 & ~n237;
  assign n259 = n257 & ~n258;
  assign n260 = n233 & n259;
  assign n261 = n260 ^ n259;
  assign n262 = ~x65 & n261;
  assign n263 = ~n251 & ~n262;
  assign n264 = ~x129 & ~n263;
  assign n265 = ~x17 & n178;
  assign n266 = ~x61 & ~x118;
  assign n267 = ~x129 & n266;
  assign n268 = ~n265 & n267;
  assign n269 = x0 & ~x113;
  assign n270 = x123 & ~x129;
  assign n271 = n270 ^ x129;
  assign n272 = n269 & ~n271;
  assign n273 = ~n268 & ~n272;
  assign n277 = n218 ^ n213;
  assign n278 = x4 & n277;
  assign n274 = n173 & n220;
  assign n275 = n204 & n274;
  assign n276 = x10 & n275;
  assign n279 = n278 ^ n276;
  assign n280 = ~x29 & ~x59;
  assign n281 = n174 & n280;
  assign n282 = n171 & n274;
  assign n283 = ~x16 & n282;
  assign n284 = n281 & n283;
  assign n285 = ~x25 & ~x28;
  assign n286 = n285 ^ x25;
  assign n287 = n284 & ~n286;
  assign n288 = x5 & n277;
  assign n289 = ~n287 & ~n288;
  assign n290 = n285 ^ x28;
  assign n291 = n284 & ~n290;
  assign n292 = x6 & n277;
  assign n293 = ~n291 & ~n292;
  assign n295 = x7 & n277;
  assign n294 = x8 & n275;
  assign n296 = n295 ^ n294;
  assign n298 = x8 & n277;
  assign n297 = x21 & n275;
  assign n299 = n298 ^ n297;
  assign n301 = ~x5 & n221;
  assign n302 = n171 & n301;
  assign n303 = x11 & n302;
  assign n304 = ~x22 & n303;
  assign n300 = x9 & n277;
  assign n305 = n304 ^ n300;
  assign n307 = x10 & n277;
  assign n306 = x14 & n275;
  assign n308 = n307 ^ n306;
  assign n309 = x22 & n302;
  assign n310 = n309 ^ n277;
  assign n311 = ~x11 & n310;
  assign n312 = n311 ^ n277;
  assign n314 = ~x18 & n283;
  assign n315 = n314 ^ n283;
  assign n316 = ~x19 & n315;
  assign n313 = x12 & n277;
  assign n317 = n316 ^ n313;
  assign n319 = x29 & x54;
  assign n320 = ~x59 & n319;
  assign n321 = n285 & n320;
  assign n322 = n265 & n321;
  assign n323 = n213 & n322;
  assign n318 = x13 & n277;
  assign n324 = n323 ^ n318;
  assign n326 = x14 & n277;
  assign n325 = x13 & n275;
  assign n327 = n326 ^ n325;
  assign n328 = x15 & ~n249;
  assign n330 = ~x70 & ~n233;
  assign n329 = ~x15 & n247;
  assign n331 = n330 ^ n329;
  assign n332 = ~x82 & n331;
  assign n333 = n332 ^ n329;
  assign n334 = ~n328 & ~n333;
  assign n335 = n252 & ~n330;
  assign n336 = ~x129 & ~n335;
  assign n337 = ~n334 & n336;
  assign n339 = x16 & n277;
  assign n338 = x6 & n229;
  assign n340 = n339 ^ n338;
  assign n342 = ~x29 & n285;
  assign n343 = n178 & n342;
  assign n344 = x59 & n220;
  assign n345 = n343 & n344;
  assign n341 = x17 & n277;
  assign n346 = n345 ^ n341;
  assign n348 = n175 & n282;
  assign n347 = x18 & n277;
  assign n349 = n348 ^ n347;
  assign n351 = x19 & n277;
  assign n350 = n178 & n219;
  assign n352 = n351 ^ n350;
  assign n353 = n329 ^ x20;
  assign n354 = x82 & ~n353;
  assign n357 = x71 ^ x20;
  assign n358 = ~n233 & ~n357;
  assign n360 = n358 ^ x82;
  assign n355 = x20 ^ x2;
  assign n356 = ~x20 & n355;
  assign n361 = n356 ^ x20;
  assign n362 = ~n360 & ~n361;
  assign n359 = n358 ^ n356;
  assign n363 = n362 ^ n359;
  assign n364 = ~x82 & n363;
  assign n365 = n364 ^ n356;
  assign n366 = n365 ^ n362;
  assign n367 = n366 ^ x20;
  assign n368 = ~x129 & n367;
  assign n369 = ~n354 & n368;
  assign n371 = x19 & n314;
  assign n370 = x21 & n277;
  assign n372 = n371 ^ n370;
  assign n373 = x22 & n277;
  assign n374 = n373 ^ n227;
  assign n375 = ~x23 & x55;
  assign n376 = x61 & ~x129;
  assign n377 = ~n375 & n376;
  assign n378 = x63 & n261;
  assign n379 = x82 & n244;
  assign n380 = ~x45 & n379;
  assign n381 = n380 ^ x82;
  assign n382 = n381 ^ n260;
  assign n383 = n382 ^ n380;
  assign n384 = ~x24 & n383;
  assign n385 = n384 ^ n380;
  assign n386 = ~x129 & ~n385;
  assign n387 = ~n378 & n386;
  assign n391 = ~x53 & ~x58;
  assign n396 = ~x85 & n391;
  assign n388 = ~x26 & x27;
  assign n389 = n388 ^ x26;
  assign n399 = n389 ^ x27;
  assign n400 = n399 ^ x26;
  assign n401 = n396 & ~n400;
  assign n397 = ~n389 & n396;
  assign n390 = x58 ^ x53;
  assign n392 = n391 ^ n390;
  assign n393 = ~x85 & n392;
  assign n394 = n393 ^ n391;
  assign n395 = ~n389 & n394;
  assign n398 = n397 ^ n395;
  assign n402 = n401 ^ n398;
  assign n403 = ~x116 & n402;
  assign n409 = ~x39 & ~x52;
  assign n410 = ~x51 & n409;
  assign n411 = x26 & x116;
  assign n412 = n410 & n411;
  assign n413 = n401 & ~n412;
  assign n404 = ~x95 & ~x100;
  assign n405 = ~x97 & n404;
  assign n406 = ~x110 & ~n405;
  assign n407 = n397 & ~n406;
  assign n408 = n407 ^ n397;
  assign n414 = n413 ^ n408;
  assign n415 = ~n403 & ~n414;
  assign n416 = x27 & x116;
  assign n417 = ~n410 & n416;
  assign n418 = n213 & ~n417;
  assign n419 = x116 & n389;
  assign n420 = ~x25 & ~n419;
  assign n421 = n418 & ~n420;
  assign n422 = ~n415 & n421;
  assign n423 = ~x96 & ~x110;
  assign n424 = n423 ^ x116;
  assign n425 = ~x85 & n424;
  assign n426 = n425 ^ x116;
  assign n427 = x100 & n426;
  assign n428 = n213 & ~n389;
  assign n429 = n391 & n428;
  assign n430 = n427 & n429;
  assign n431 = ~n422 & ~n430;
  assign n432 = x116 & n410;
  assign n433 = n396 & ~n432;
  assign n434 = n213 & n399;
  assign n435 = n433 & n434;
  assign n436 = n435 ^ n430;
  assign n437 = n388 & n433;
  assign n438 = x85 & x116;
  assign n439 = ~x95 & ~n438;
  assign n440 = ~n389 & n391;
  assign n441 = ~n439 & n440;
  assign n442 = ~x100 & n441;
  assign n443 = n426 & n442;
  assign n444 = ~n437 & ~n443;
  assign n445 = n213 & ~n444;
  assign n446 = ~x27 & n396;
  assign n447 = ~x26 & ~n406;
  assign n448 = x28 & n447;
  assign n449 = n448 ^ n412;
  assign n450 = n446 & n449;
  assign n451 = n445 ^ x28;
  assign n452 = n403 & n451;
  assign n453 = n452 ^ n445;
  assign n454 = ~n450 & ~n453;
  assign n455 = n213 & ~n454;
  assign n456 = n407 ^ n403;
  assign n457 = x53 & x116;
  assign n458 = n393 & ~n457;
  assign n459 = n428 & n458;
  assign n460 = ~x53 & x97;
  assign n461 = n404 & n423;
  assign n462 = n461 ^ x116;
  assign n463 = n460 ^ x58;
  assign n464 = n462 & ~n463;
  assign n465 = n464 ^ n461;
  assign n466 = n460 & n465;
  assign n467 = n466 ^ x53;
  assign n468 = n459 & n467;
  assign n469 = n468 ^ x29;
  assign n470 = ~n456 & n469;
  assign n471 = n470 ^ x29;
  assign n472 = n213 & n471;
  assign n473 = x60 ^ x30;
  assign n474 = x109 & n473;
  assign n475 = n474 ^ x30;
  assign n476 = n475 ^ x88;
  assign n477 = ~x106 & n476;
  assign n478 = n477 ^ x88;
  assign n479 = ~x129 & n478;
  assign n480 = x31 ^ x30;
  assign n481 = ~x109 & n480;
  assign n482 = n481 ^ x30;
  assign n483 = n482 ^ x89;
  assign n484 = ~x106 & n483;
  assign n485 = n484 ^ x89;
  assign n486 = ~x129 & n485;
  assign n487 = x32 ^ x31;
  assign n488 = ~x109 & n487;
  assign n489 = n488 ^ x31;
  assign n490 = n489 ^ x99;
  assign n491 = ~x106 & n490;
  assign n492 = n491 ^ x99;
  assign n493 = ~x129 & n492;
  assign n494 = x33 ^ x32;
  assign n495 = ~x109 & n494;
  assign n496 = n495 ^ x32;
  assign n497 = n496 ^ x90;
  assign n498 = ~x106 & n497;
  assign n499 = n498 ^ x90;
  assign n500 = ~x129 & n499;
  assign n501 = x34 ^ x33;
  assign n502 = ~x109 & n501;
  assign n503 = n502 ^ x33;
  assign n504 = n503 ^ x91;
  assign n505 = ~x106 & n504;
  assign n506 = n505 ^ x91;
  assign n507 = ~x129 & n506;
  assign n508 = x35 ^ x34;
  assign n509 = ~x109 & n508;
  assign n510 = n509 ^ x34;
  assign n511 = n510 ^ x92;
  assign n512 = ~x106 & n511;
  assign n513 = n512 ^ x92;
  assign n514 = ~x129 & n513;
  assign n515 = x36 ^ x35;
  assign n516 = ~x109 & n515;
  assign n517 = n516 ^ x35;
  assign n518 = n517 ^ x98;
  assign n519 = ~x106 & n518;
  assign n520 = n519 ^ x98;
  assign n521 = ~x129 & n520;
  assign n522 = x37 ^ x36;
  assign n523 = ~x109 & n522;
  assign n524 = n523 ^ x36;
  assign n525 = n524 ^ x93;
  assign n526 = ~x106 & n525;
  assign n527 = n526 ^ x93;
  assign n528 = ~x129 & n527;
  assign n529 = x74 ^ x38;
  assign n530 = ~n233 & ~n529;
  assign n531 = n530 ^ x38;
  assign n532 = n257 & ~n531;
  assign n533 = n237 ^ x38;
  assign n534 = x82 & ~n533;
  assign n535 = ~x129 & ~n534;
  assign n536 = ~n532 & n535;
  assign n537 = ~x51 & x109;
  assign n538 = ~x52 & n537;
  assign n539 = n538 ^ x39;
  assign n540 = ~x106 & ~n539;
  assign n541 = ~x129 & ~n540;
  assign n542 = ~x73 & ~n233;
  assign n543 = n257 & ~n542;
  assign n544 = ~n258 & ~n543;
  assign n545 = x82 & ~n236;
  assign n546 = n545 ^ n235;
  assign n547 = x40 & ~n546;
  assign n548 = ~n544 & ~n547;
  assign n549 = ~x129 & ~n548;
  assign n550 = ~x46 & n239;
  assign n551 = n550 ^ x41;
  assign n552 = x82 & ~n551;
  assign n553 = ~x129 & ~n552;
  assign n554 = x76 ^ x41;
  assign n555 = ~n233 & ~n554;
  assign n556 = n555 ^ x41;
  assign n557 = ~n255 & ~n556;
  assign n558 = n553 & ~n557;
  assign n561 = x72 & n259;
  assign n562 = ~n260 & ~n561;
  assign n560 = x44 & x82;
  assign n563 = n562 ^ n560;
  assign n559 = x42 & ~n234;
  assign n564 = n563 ^ n559;
  assign n565 = ~x129 & n564;
  assign n566 = n239 & n240;
  assign n567 = n566 ^ x43;
  assign n568 = x82 & ~n567;
  assign n569 = ~x129 & ~n568;
  assign n570 = x77 ^ x43;
  assign n571 = ~n233 & ~n570;
  assign n572 = n571 ^ x43;
  assign n573 = ~n255 & ~n572;
  assign n574 = n569 & ~n573;
  assign n575 = x67 ^ x44;
  assign n576 = ~n233 & ~n575;
  assign n577 = n576 ^ x44;
  assign n578 = n259 & ~n577;
  assign n579 = ~x129 & ~n560;
  assign n580 = ~n578 & n579;
  assign n581 = x82 & ~n253;
  assign n582 = ~x68 & ~n233;
  assign n583 = ~n581 & ~n582;
  assign n584 = ~n381 & ~n583;
  assign n585 = x45 & ~n234;
  assign n586 = ~n379 & n585;
  assign n587 = ~n584 & ~n586;
  assign n588 = ~x129 & ~n587;
  assign n589 = x75 ^ x46;
  assign n590 = ~n233 & ~n589;
  assign n591 = n590 ^ x46;
  assign n592 = n259 & ~n591;
  assign n593 = n239 ^ x46;
  assign n594 = x82 & ~n593;
  assign n595 = ~x129 & ~n594;
  assign n596 = ~n592 & n595;
  assign n597 = ~x43 & n566;
  assign n598 = n597 ^ x47;
  assign n599 = x82 & ~n598;
  assign n600 = x64 ^ x47;
  assign n601 = ~n233 & ~n600;
  assign n602 = n601 ^ x47;
  assign n603 = ~n255 & ~n602;
  assign n604 = ~x129 & ~n603;
  assign n605 = ~n599 & n604;
  assign n606 = ~x47 & n597;
  assign n607 = n606 ^ x48;
  assign n608 = x82 & ~n607;
  assign n609 = x48 & ~n234;
  assign n610 = ~x62 & ~n233;
  assign n611 = ~n609 & ~n610;
  assign n612 = ~n581 & n611;
  assign n613 = ~x129 & ~n612;
  assign n614 = ~n608 & n613;
  assign n617 = ~x69 & ~n233;
  assign n618 = n617 ^ n380;
  assign n619 = n259 & n618;
  assign n616 = ~x24 & n380;
  assign n620 = n619 ^ n616;
  assign n615 = x49 & ~n234;
  assign n621 = n620 ^ n615;
  assign n622 = ~x129 & n621;
  assign n623 = ~x66 & ~n233;
  assign n624 = n254 & ~n623;
  assign n625 = n256 ^ n235;
  assign n626 = ~n258 & n625;
  assign n627 = ~n624 & n626;
  assign n628 = ~x50 & ~n627;
  assign n629 = ~x38 & n237;
  assign n630 = n256 & n629;
  assign n631 = x66 & n234;
  assign n632 = ~x129 & ~n631;
  assign n633 = ~n630 & n632;
  assign n634 = ~n628 & n633;
  assign n635 = x109 ^ x51;
  assign n636 = ~x106 & ~n635;
  assign n637 = ~x129 & ~n636;
  assign n638 = n537 ^ x52;
  assign n639 = ~x106 & ~n638;
  assign n640 = ~x129 & ~n639;
  assign n641 = ~x129 & ~n261;
  assign n642 = ~x114 & ~x122;
  assign n643 = n642 ^ x122;
  assign n644 = ~n271 & ~n643;
  assign n645 = n401 ^ n395;
  assign n646 = n213 & n645;
  assign n647 = ~x37 & ~x58;
  assign n648 = n647 ^ x94;
  assign n649 = x58 & x116;
  assign n650 = n649 ^ x58;
  assign n651 = n650 ^ n411;
  assign n652 = ~n648 & ~n651;
  assign n653 = n652 ^ x94;
  assign n654 = n646 & n653;
  assign n655 = x60 ^ x57;
  assign n656 = n649 & n655;
  assign n657 = n656 ^ x57;
  assign n658 = n646 & n657;
  assign n659 = n410 & n419;
  assign n660 = n659 ^ n650;
  assign n661 = n646 & n660;
  assign n663 = x96 & n408;
  assign n662 = x59 & n456;
  assign n664 = n663 ^ n662;
  assign n665 = n213 & n664;
  assign n666 = ~x117 & ~x122;
  assign n667 = x123 ^ x60;
  assign n668 = n666 & n667;
  assign n669 = n668 ^ x60;
  assign n670 = n270 & n642;
  assign n671 = x132 & x133;
  assign n672 = x131 & n671;
  assign n673 = ~x138 & n672;
  assign n674 = x136 & x137;
  assign n675 = n674 ^ x136;
  assign n676 = n673 & n675;
  assign n677 = x140 ^ x62;
  assign n678 = n676 & ~n677;
  assign n679 = n678 ^ x62;
  assign n680 = ~x129 & n679;
  assign n681 = x142 ^ x63;
  assign n682 = n676 & ~n681;
  assign n683 = n682 ^ x63;
  assign n684 = ~x129 & n683;
  assign n685 = x139 ^ x64;
  assign n686 = n676 & ~n685;
  assign n687 = n686 ^ x64;
  assign n688 = ~x129 & n687;
  assign n689 = x146 ^ x65;
  assign n690 = n676 & ~n689;
  assign n691 = n690 ^ x65;
  assign n692 = ~x129 & n691;
  assign n693 = n674 ^ x137;
  assign n694 = n693 ^ x136;
  assign n695 = n673 & ~n694;
  assign n696 = x143 ^ x66;
  assign n697 = n695 & ~n696;
  assign n698 = n697 ^ x66;
  assign n699 = ~x129 & n698;
  assign n700 = x139 ^ x67;
  assign n701 = n695 & ~n700;
  assign n702 = n701 ^ x67;
  assign n703 = ~x129 & n702;
  assign n704 = x141 ^ x68;
  assign n705 = n676 & ~n704;
  assign n706 = n705 ^ x68;
  assign n707 = ~x129 & n706;
  assign n708 = x143 ^ x69;
  assign n709 = n676 & ~n708;
  assign n710 = n709 ^ x69;
  assign n711 = ~x129 & n710;
  assign n712 = x144 ^ x70;
  assign n713 = n676 & ~n712;
  assign n714 = n713 ^ x70;
  assign n715 = ~x129 & n714;
  assign n716 = x145 ^ x71;
  assign n717 = n676 & ~n716;
  assign n718 = n717 ^ x71;
  assign n719 = ~x129 & n718;
  assign n720 = x140 ^ x72;
  assign n721 = n695 & ~n720;
  assign n722 = n721 ^ x72;
  assign n723 = ~x129 & n722;
  assign n724 = x141 ^ x73;
  assign n725 = n695 & ~n724;
  assign n726 = n725 ^ x73;
  assign n727 = ~x129 & n726;
  assign n728 = x142 ^ x74;
  assign n729 = n695 & ~n728;
  assign n730 = n729 ^ x74;
  assign n731 = ~x129 & n730;
  assign n732 = x144 ^ x75;
  assign n733 = n695 & ~n732;
  assign n734 = n733 ^ x75;
  assign n735 = ~x129 & n734;
  assign n736 = x145 ^ x76;
  assign n737 = n695 & ~n736;
  assign n738 = n737 ^ x76;
  assign n739 = ~x129 & n738;
  assign n740 = x146 ^ x77;
  assign n741 = n695 & ~n740;
  assign n742 = n741 ^ x77;
  assign n743 = ~x129 & n742;
  assign n744 = n673 & n693;
  assign n745 = x142 ^ x78;
  assign n746 = n744 & n745;
  assign n747 = n746 ^ x78;
  assign n748 = ~x129 & n747;
  assign n749 = x143 ^ x79;
  assign n750 = n744 & n749;
  assign n751 = n750 ^ x79;
  assign n752 = ~x129 & n751;
  assign n753 = x144 ^ x80;
  assign n754 = n744 & n753;
  assign n755 = n754 ^ x80;
  assign n756 = ~x129 & n755;
  assign n757 = x145 ^ x81;
  assign n758 = n744 & n757;
  assign n759 = n758 ^ x81;
  assign n760 = ~x129 & n759;
  assign n761 = x146 ^ x82;
  assign n762 = n744 & n761;
  assign n763 = n762 ^ x82;
  assign n764 = ~x129 & n763;
  assign n779 = x115 ^ x87;
  assign n780 = ~x138 & ~n779;
  assign n781 = n780 ^ x115;
  assign n776 = x119 ^ x72;
  assign n777 = ~x138 & ~n776;
  assign n778 = n777 ^ x119;
  assign n782 = n781 ^ n778;
  assign n783 = ~x137 & ~n782;
  assign n784 = n783 ^ n781;
  assign n765 = x138 ^ x136;
  assign n768 = x62 ^ x31;
  assign n769 = ~x137 & ~n768;
  assign n770 = n769 ^ x31;
  assign n766 = x137 ^ x89;
  assign n767 = ~x137 & ~n766;
  assign n771 = n770 ^ n767;
  assign n772 = n771 ^ x137;
  assign n773 = n765 & ~n772;
  assign n774 = n773 ^ n767;
  assign n775 = n774 ^ x137;
  assign n785 = n784 ^ n775;
  assign n786 = ~x136 & n785;
  assign n787 = n786 ^ n775;
  assign n788 = x141 ^ x84;
  assign n789 = n744 & n788;
  assign n790 = n789 ^ x84;
  assign n791 = ~x129 & n790;
  assign n792 = x96 & n406;
  assign n793 = n792 ^ x116;
  assign n794 = ~x85 & ~n793;
  assign n795 = n794 ^ x116;
  assign n796 = n429 & ~n795;
  assign n797 = x139 ^ x86;
  assign n798 = n744 & n797;
  assign n799 = n798 ^ x86;
  assign n800 = ~x129 & n799;
  assign n801 = x140 ^ x87;
  assign n802 = n744 & n801;
  assign n803 = n802 ^ x87;
  assign n804 = ~x129 & n803;
  assign n805 = n673 & n674;
  assign n806 = x139 ^ x88;
  assign n807 = n805 & n806;
  assign n808 = n807 ^ x88;
  assign n809 = ~x129 & n808;
  assign n810 = x140 ^ x89;
  assign n811 = n805 & n810;
  assign n812 = n811 ^ x89;
  assign n813 = ~x129 & n812;
  assign n814 = x142 ^ x90;
  assign n815 = n805 & n814;
  assign n816 = n815 ^ x90;
  assign n817 = ~x129 & n816;
  assign n818 = x143 ^ x91;
  assign n819 = n805 & n818;
  assign n820 = n819 ^ x91;
  assign n821 = ~x129 & n820;
  assign n822 = x144 ^ x92;
  assign n823 = n805 & n822;
  assign n824 = n823 ^ x92;
  assign n825 = ~x129 & n824;
  assign n826 = x146 ^ x93;
  assign n827 = n805 & n826;
  assign n828 = n827 ^ x93;
  assign n829 = ~x129 & n828;
  assign n830 = x82 & x138;
  assign n831 = ~n694 & n830;
  assign n832 = n672 & n831;
  assign n833 = x142 ^ x94;
  assign n834 = n832 & n833;
  assign n835 = n834 ^ x94;
  assign n836 = ~x129 & n835;
  assign n837 = ~x3 & ~x110;
  assign n838 = ~n672 & ~n837;
  assign n839 = x95 & ~n838;
  assign n840 = n839 ^ x143;
  assign n841 = ~n832 & n840;
  assign n842 = n841 ^ x143;
  assign n843 = ~x129 & n842;
  assign n844 = x96 & ~n838;
  assign n845 = n844 ^ x146;
  assign n846 = ~n832 & n845;
  assign n847 = n846 ^ x146;
  assign n848 = ~x129 & n847;
  assign n849 = x97 & ~n838;
  assign n850 = n849 ^ x145;
  assign n851 = ~n832 & n850;
  assign n852 = n851 ^ x145;
  assign n853 = ~x129 & n852;
  assign n854 = x145 ^ x98;
  assign n855 = n805 & n854;
  assign n856 = n855 ^ x98;
  assign n857 = ~x129 & n856;
  assign n858 = x141 ^ x99;
  assign n859 = n805 & n858;
  assign n860 = n859 ^ x99;
  assign n861 = ~x129 & n860;
  assign n862 = x100 & ~n838;
  assign n863 = n862 ^ x144;
  assign n864 = ~n832 & n863;
  assign n865 = n864 ^ x144;
  assign n866 = ~x129 & n865;
  assign n867 = x137 ^ x136;
  assign n868 = n867 ^ x138;
  assign n869 = x96 ^ x93;
  assign n870 = ~x137 & n869;
  assign n871 = n870 ^ x96;
  assign n872 = n871 ^ n867;
  assign n873 = n868 & n872;
  assign n874 = n873 ^ n870;
  assign n875 = n874 ^ x96;
  assign n876 = n875 ^ x138;
  assign n877 = n867 & n876;
  assign n878 = n877 ^ n867;
  assign n879 = n878 ^ x138;
  assign n883 = x136 ^ x65;
  assign n884 = ~x65 & ~n883;
  assign n880 = x82 ^ x37;
  assign n881 = x136 & n880;
  assign n882 = n881 ^ x82;
  assign n885 = n884 ^ n882;
  assign n886 = n885 ^ x65;
  assign n887 = x138 ^ x137;
  assign n888 = ~n886 & n887;
  assign n889 = n888 ^ n884;
  assign n890 = n889 ^ x65;
  assign n891 = ~x138 & ~n890;
  assign n892 = n891 ^ x138;
  assign n893 = ~n879 & n892;
  assign n894 = x124 ^ x77;
  assign n895 = ~x138 & ~n894;
  assign n896 = n895 ^ x124;
  assign n897 = ~n694 & n896;
  assign n898 = ~n893 & ~n897;
  assign n899 = x69 ^ x66;
  assign n900 = ~x136 & n899;
  assign n901 = n900 ^ x69;
  assign n902 = ~x137 & ~n901;
  assign n903 = x79 ^ x34;
  assign n904 = ~x136 & n903;
  assign n905 = n904 ^ x34;
  assign n906 = n905 ^ x138;
  assign n907 = ~n887 & ~n906;
  assign n908 = n907 ^ n904;
  assign n909 = n908 ^ x34;
  assign n910 = n909 ^ x137;
  assign n911 = ~x138 & n910;
  assign n912 = n911 ^ x138;
  assign n913 = n912 ^ x138;
  assign n914 = ~n902 & n913;
  assign n915 = x95 ^ x91;
  assign n916 = ~x137 & n915;
  assign n917 = n916 ^ x95;
  assign n918 = n917 ^ n867;
  assign n919 = n868 & n918;
  assign n920 = n919 ^ n916;
  assign n921 = n920 ^ x95;
  assign n922 = n921 ^ x138;
  assign n923 = n867 & n922;
  assign n924 = n923 ^ n867;
  assign n925 = n924 ^ x138;
  assign n926 = ~n914 & ~n925;
  assign n927 = x78 & n693;
  assign n928 = ~x138 & ~n927;
  assign n930 = x63 ^ x33;
  assign n931 = x137 & ~n930;
  assign n932 = n931 ^ x63;
  assign n929 = ~x74 & ~x137;
  assign n933 = n932 ^ n929;
  assign n934 = ~x136 & ~n933;
  assign n935 = n934 ^ n932;
  assign n936 = n928 & n935;
  assign n937 = x94 ^ x90;
  assign n938 = ~x137 & n937;
  assign n939 = n938 ^ x94;
  assign n940 = n939 ^ n867;
  assign n941 = n868 & n940;
  assign n942 = n941 ^ n938;
  assign n943 = n942 ^ x94;
  assign n944 = n943 ^ x138;
  assign n945 = n867 & n944;
  assign n946 = n945 ^ n867;
  assign n947 = n946 ^ x138;
  assign n948 = ~n936 & ~n947;
  assign n949 = x73 ^ x68;
  assign n950 = ~x136 & n949;
  assign n951 = n950 ^ x68;
  assign n952 = n951 ^ x138;
  assign n953 = n887 & n952;
  assign n954 = n953 ^ n950;
  assign n955 = n954 ^ x68;
  assign n956 = n955 ^ x137;
  assign n957 = ~x138 & n956;
  assign n958 = n957 ^ x138;
  assign n959 = n958 ^ x138;
  assign n960 = x84 ^ x32;
  assign n961 = x136 & n960;
  assign n962 = n961 ^ x84;
  assign n963 = x137 & n962;
  assign n964 = n959 & ~n963;
  assign n965 = x112 ^ x99;
  assign n966 = ~x137 & ~n965;
  assign n967 = n966 ^ x112;
  assign n968 = n967 ^ n867;
  assign n969 = n868 & ~n968;
  assign n970 = n969 ^ n966;
  assign n971 = n970 ^ x112;
  assign n972 = n971 ^ x138;
  assign n973 = n867 & ~n972;
  assign n974 = n973 ^ n867;
  assign n975 = n974 ^ x138;
  assign n976 = ~n964 & ~n975;
  assign n987 = x125 ^ x100;
  assign n988 = x137 & n987;
  assign n989 = n988 ^ x125;
  assign n986 = x92 & ~x137;
  assign n990 = n989 ^ n986;
  assign n991 = x136 & n990;
  assign n992 = n991 ^ n989;
  assign n980 = x80 ^ x75;
  assign n981 = ~x137 & ~n980;
  assign n982 = n981 ^ x80;
  assign n977 = x70 ^ x35;
  assign n978 = x137 & ~n977;
  assign n979 = n978 ^ x70;
  assign n983 = n982 ^ n979;
  assign n984 = x136 & ~n983;
  assign n985 = n984 ^ n982;
  assign n993 = n992 ^ n985;
  assign n994 = x138 & n993;
  assign n995 = n994 ^ n985;
  assign n996 = n438 ^ n408;
  assign n997 = n213 & n996;
  assign n1008 = x71 ^ x36;
  assign n1009 = ~x137 & ~n1008;
  assign n1010 = n1009 ^ x36;
  assign n1007 = x98 & ~x137;
  assign n1011 = n1010 ^ n1007;
  assign n1012 = x138 & n1011;
  assign n1013 = n1012 ^ n1010;
  assign n1001 = x76 ^ x23;
  assign n1002 = x138 & ~n1001;
  assign n1003 = n1002 ^ x76;
  assign n998 = x97 ^ x81;
  assign n999 = ~x138 & n998;
  assign n1000 = n999 ^ x97;
  assign n1004 = n1003 ^ n1000;
  assign n1005 = x137 & ~n1004;
  assign n1006 = n1005 ^ n1003;
  assign n1014 = n1013 ^ n1006;
  assign n1015 = ~x136 & ~n1014;
  assign n1016 = n1015 ^ n1013;
  assign n1030 = x120 ^ x67;
  assign n1031 = ~x138 & ~n1030;
  assign n1032 = n1031 ^ x120;
  assign n1027 = x111 ^ x86;
  assign n1028 = ~x138 & n1027;
  assign n1029 = n1028 ^ x111;
  assign n1033 = n1032 ^ n1029;
  assign n1034 = x137 & n1033;
  assign n1035 = n1034 ^ n1032;
  assign n1019 = x64 ^ x30;
  assign n1020 = ~x137 & ~n1019;
  assign n1021 = n1020 ^ x30;
  assign n1017 = x137 ^ x88;
  assign n1018 = ~x137 & ~n1017;
  assign n1022 = n1021 ^ n1018;
  assign n1023 = n1022 ^ x137;
  assign n1024 = n765 & ~n1023;
  assign n1025 = n1024 ^ n1018;
  assign n1026 = n1025 ^ x137;
  assign n1036 = n1035 ^ n1026;
  assign n1037 = ~x136 & ~n1036;
  assign n1038 = n1037 ^ n1026;
  assign n1039 = x116 & n213;
  assign n1040 = n388 & ~n410;
  assign n1041 = n1040 ^ n399;
  assign n1042 = n1039 & n1041;
  assign n1043 = n390 & ~n460;
  assign n1044 = n1039 & n1043;
  assign n1045 = ~x129 & n672;
  assign n1046 = x139 ^ x111;
  assign n1047 = ~n831 & n1046;
  assign n1048 = n1047 ^ x139;
  assign n1049 = n1045 & n1048;
  assign n1050 = x141 ^ x112;
  assign n1051 = ~n831 & ~n1050;
  assign n1052 = n1051 ^ x141;
  assign n1053 = n1045 & n1052;
  assign n1054 = n222 ^ x113;
  assign n1055 = x54 & n1054;
  assign n1056 = n1055 ^ x113;
  assign n1057 = n213 & ~n1056;
  assign n1058 = x140 ^ x115;
  assign n1059 = ~n831 & ~n1058;
  assign n1060 = n1059 ^ x140;
  assign n1061 = n1045 & n1060;
  assign n1062 = ~n156 & n218;
  assign n1063 = x122 & ~x129;
  assign n1064 = ~x54 & x118;
  assign n1065 = n1064 ^ n321;
  assign n1066 = ~x129 & n1065;
  assign n1067 = ~x129 & ~n404;
  assign n1068 = ~x120 & n837;
  assign n1069 = ~x111 & ~x129;
  assign n1070 = ~n1068 & n1069;
  assign n1071 = x81 & x120;
  assign n1072 = ~x129 & n1071;
  assign n1073 = ~x129 & ~x134;
  assign n1074 = ~x129 & ~x135;
  assign n1075 = x57 & ~x129;
  assign n1076 = ~x96 & x125;
  assign n1077 = ~x3 & ~n1076;
  assign n1078 = ~x129 & ~n1077;
  assign n1079 = ~x126 & n671;
  assign y0 = x108;
  assign y1 = x83;
  assign y2 = x104;
  assign y3 = x103;
  assign y4 = x102;
  assign y5 = x105;
  assign y6 = x107;
  assign y7 = x101;
  assign y8 = x126;
  assign y9 = x121;
  assign y10 = x1;
  assign y11 = x0;
  assign y12 = ~1'b0;
  assign y13 = x130;
  assign y14 = x128;
  assign y15 = ~n214;
  assign y16 = n230;
  assign y17 = n264;
  assign y18 = ~n273;
  assign y19 = n279;
  assign y20 = ~n289;
  assign y21 = ~n293;
  assign y22 = n296;
  assign y23 = n299;
  assign y24 = n305;
  assign y25 = n308;
  assign y26 = n312;
  assign y27 = n317;
  assign y28 = n324;
  assign y29 = n327;
  assign y30 = n337;
  assign y31 = n340;
  assign y32 = n346;
  assign y33 = n349;
  assign y34 = n352;
  assign y35 = n369;
  assign y36 = n372;
  assign y37 = n374;
  assign y38 = n377;
  assign y39 = n387;
  assign y40 = ~n431;
  assign y41 = n436;
  assign y42 = n445;
  assign y43 = n455;
  assign y44 = n472;
  assign y45 = n479;
  assign y46 = n486;
  assign y47 = n493;
  assign y48 = n500;
  assign y49 = n507;
  assign y50 = n514;
  assign y51 = n521;
  assign y52 = n528;
  assign y53 = n536;
  assign y54 = n541;
  assign y55 = n549;
  assign y56 = n558;
  assign y57 = n565;
  assign y58 = n574;
  assign y59 = n580;
  assign y60 = n588;
  assign y61 = n596;
  assign y62 = n605;
  assign y63 = n614;
  assign y64 = n622;
  assign y65 = n634;
  assign y66 = n637;
  assign y67 = n640;
  assign y68 = n468;
  assign y69 = ~n641;
  assign y70 = n644;
  assign y71 = n654;
  assign y72 = n658;
  assign y73 = n661;
  assign y74 = n665;
  assign y75 = n669;
  assign y76 = n670;
  assign y77 = ~n680;
  assign y78 = ~n684;
  assign y79 = ~n688;
  assign y80 = ~n692;
  assign y81 = ~n699;
  assign y82 = ~n703;
  assign y83 = ~n707;
  assign y84 = ~n711;
  assign y85 = ~n715;
  assign y86 = ~n719;
  assign y87 = ~n723;
  assign y88 = ~n727;
  assign y89 = ~n731;
  assign y90 = ~n735;
  assign y91 = ~n739;
  assign y92 = ~n743;
  assign y93 = n748;
  assign y94 = n752;
  assign y95 = n756;
  assign y96 = n760;
  assign y97 = n764;
  assign y98 = ~n787;
  assign y99 = n791;
  assign y100 = n796;
  assign y101 = n800;
  assign y102 = n804;
  assign y103 = n809;
  assign y104 = n813;
  assign y105 = n817;
  assign y106 = n821;
  assign y107 = n825;
  assign y108 = n829;
  assign y109 = n836;
  assign y110 = n843;
  assign y111 = n848;
  assign y112 = n853;
  assign y113 = n857;
  assign y114 = n861;
  assign y115 = n866;
  assign y116 = ~n898;
  assign y117 = n926;
  assign y118 = n948;
  assign y119 = n976;
  assign y120 = n995;
  assign y121 = n997;
  assign y122 = n1016;
  assign y123 = ~n1038;
  assign y124 = n1042;
  assign y125 = n1044;
  assign y126 = n1049;
  assign y127 = n1053;
  assign y128 = n1057;
  assign y129 = n271;
  assign y130 = n1061;
  assign y131 = n1062;
  assign y132 = ~n1063;
  assign y133 = n1066;
  assign y134 = n1067;
  assign y135 = n1070;
  assign y136 = n1072;
  assign y137 = ~n1073;
  assign y138 = ~n1074;
  assign y139 = n1075;
  assign y140 = n1078;
  assign y141 = n1079;
endmodule
