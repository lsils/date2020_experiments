module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , x233 , x234 , x235 , x236 , x237 , x238 , x239 , x240 , x241 , x242 , x243 , x244 , x245 , x246 , x247 , x248 , x249 , x250 , x251 , x252 , x253 , x254 , x255 , x256 , x257 , x258 , x259 , x260 , x261 , x262 , x263 , x264 , x265 , x266 , x267 , x268 , x269 , x270 , x271 , x272 , x273 , x274 , x275 , x276 , x277 , x278 , x279 , x280 , x281 , x282 , x283 , x284 , x285 , x286 , x287 , x288 , x289 , x290 , x291 , x292 , x293 , x294 , x295 , x296 , x297 , x298 , x299 , x300 , x301 , x302 , x303 , x304 , x305 , x306 , x307 , x308 , x309 , x310 , x311 , x312 , x313 , x314 , x315 , x316 , x317 , x318 , x319 , x320 , x321 , x322 , x323 , x324 , x325 , x326 , x327 , x328 , x329 , x330 , x331 , x332 , x333 , x334 , x335 , x336 , x337 , x338 , x339 , x340 , x341 , x342 , x343 , x344 , x345 , x346 , x347 , x348 , x349 , x350 , x351 , x352 , x353 , x354 , x355 , x356 , x357 , x358 , x359 , x360 , x361 , x362 , x363 , x364 , x365 , x366 , x367 , x368 , x369 , x370 , x371 , x372 , x373 , x374 , x375 , x376 , x377 , x378 , x379 , x380 , x381 , x382 , x383 , x384 , x385 , x386 , x387 , x388 , x389 , x390 , x391 , x392 , x393 , x394 , x395 , x396 , x397 , x398 , x399 , x400 , x401 , x402 , x403 , x404 , x405 , x406 , x407 , x408 , x409 , x410 , x411 , x412 , x413 , x414 , x415 , x416 , x417 , x418 , x419 , x420 , x421 , x422 , x423 , x424 , x425 , x426 , x427 , x428 , x429 , x430 , x431 , x432 , x433 , x434 , x435 , x436 , x437 , x438 , x439 , x440 , x441 , x442 , x443 , x444 , x445 , x446 , x447 , x448 , x449 , x450 , x451 , x452 , x453 , x454 , x455 , x456 , x457 , x458 , x459 , x460 , x461 , x462 , x463 , x464 , x465 , x466 , x467 , x468 , x469 , x470 , x471 , x472 , x473 , x474 , x475 , x476 , x477 , x478 , x479 , x480 , x481 , x482 , x483 , x484 , x485 , x486 , x487 , x488 , x489 , x490 , x491 , x492 , x493 , x494 , x495 , x496 , x497 , x498 , x499 , x500 , x501 , x502 , x503 , x504 , x505 , x506 , x507 , x508 , x509 , x510 , x511 , x512 , x513 , x514 , x515 , x516 , x517 , x518 , x519 , x520 , x521 , x522 , x523 , x524 , x525 , x526 , x527 , x528 , x529 , x530 , x531 , x532 , x533 , x534 , x535 , x536 , x537 , x538 , x539 , x540 , x541 , x542 , x543 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 ;
  wire n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 ;
  assign n634 = x541 ^ x29 ;
  assign n633 = x542 ^ x30 ;
  assign n635 = n634 ^ n633 ;
  assign n632 = x543 ^ x31 ;
  assign n667 = n633 ^ n632 ;
  assign n668 = n635 & ~n667 ;
  assign n669 = n668 ^ n634 ;
  assign n637 = x537 ^ x25 ;
  assign n636 = n635 ^ n632 ;
  assign n638 = n637 ^ n636 ;
  assign n629 = x539 ^ x27 ;
  assign n628 = x538 ^ x26 ;
  assign n630 = n629 ^ n628 ;
  assign n627 = x540 ^ x28 ;
  assign n631 = n630 ^ n627 ;
  assign n664 = n636 ^ n631 ;
  assign n665 = n638 & ~n664 ;
  assign n666 = n665 ^ n637 ;
  assign n670 = n669 ^ n666 ;
  assign n661 = n628 ^ n627 ;
  assign n662 = n630 & ~n661 ;
  assign n663 = n662 ^ n629 ;
  assign n685 = n666 ^ n663 ;
  assign n686 = n670 & ~n685 ;
  assign n687 = n686 ^ n669 ;
  assign n671 = n670 ^ n663 ;
  assign n639 = n638 ^ n631 ;
  assign n626 = x529 ^ x17 ;
  assign n640 = n639 ^ n626 ;
  assign n621 = x535 ^ x23 ;
  assign n620 = x534 ^ x22 ;
  assign n622 = n621 ^ n620 ;
  assign n619 = x536 ^ x24 ;
  assign n623 = n622 ^ n619 ;
  assign n618 = x530 ^ x18 ;
  assign n624 = n623 ^ n618 ;
  assign n615 = x532 ^ x20 ;
  assign n614 = x531 ^ x19 ;
  assign n616 = n615 ^ n614 ;
  assign n613 = x533 ^ x21 ;
  assign n617 = n616 ^ n613 ;
  assign n625 = n624 ^ n617 ;
  assign n658 = n626 ^ n625 ;
  assign n659 = n640 & ~n658 ;
  assign n660 = n659 ^ n639 ;
  assign n672 = n671 ^ n660 ;
  assign n653 = n618 ^ n617 ;
  assign n654 = n624 & ~n653 ;
  assign n655 = n654 ^ n623 ;
  assign n650 = n620 ^ n619 ;
  assign n651 = n622 & ~n650 ;
  assign n652 = n651 ^ n621 ;
  assign n656 = n655 ^ n652 ;
  assign n647 = n614 ^ n613 ;
  assign n648 = n616 & ~n647 ;
  assign n649 = n648 ^ n615 ;
  assign n657 = n656 ^ n649 ;
  assign n682 = n671 ^ n657 ;
  assign n683 = n672 & ~n682 ;
  assign n684 = n683 ^ n660 ;
  assign n688 = n687 ^ n684 ;
  assign n679 = n652 ^ n649 ;
  assign n680 = n656 & ~n679 ;
  assign n681 = n680 ^ n655 ;
  assign n695 = n684 ^ n681 ;
  assign n696 = n688 & ~n695 ;
  assign n697 = n696 ^ n687 ;
  assign n689 = n688 ^ n681 ;
  assign n673 = n672 ^ n657 ;
  assign n641 = n640 ^ n625 ;
  assign n612 = x513 ^ x1 ;
  assign n642 = n641 ^ n612 ;
  assign n582 = x517 ^ x5 ;
  assign n581 = x516 ^ x4 ;
  assign n583 = n582 ^ n581 ;
  assign n580 = x518 ^ x6 ;
  assign n584 = n583 ^ n580 ;
  assign n576 = x520 ^ x8 ;
  assign n575 = x519 ^ x7 ;
  assign n577 = n576 ^ n575 ;
  assign n574 = x521 ^ x9 ;
  assign n578 = n577 ^ n574 ;
  assign n573 = x515 ^ x3 ;
  assign n579 = n578 ^ n573 ;
  assign n585 = n584 ^ n579 ;
  assign n571 = x514 ^ x2 ;
  assign n557 = x524 ^ x12 ;
  assign n556 = x523 ^ x11 ;
  assign n558 = n557 ^ n556 ;
  assign n555 = x525 ^ x13 ;
  assign n559 = n558 ^ n555 ;
  assign n548 = x528 ^ x16 ;
  assign n546 = x527 ^ x15 ;
  assign n545 = x526 ^ x14 ;
  assign n547 = n546 ^ n545 ;
  assign n553 = n548 ^ n547 ;
  assign n552 = x522 ^ x10 ;
  assign n554 = n553 ^ n552 ;
  assign n570 = n559 ^ n554 ;
  assign n572 = n571 ^ n570 ;
  assign n643 = n585 ^ n572 ;
  assign n644 = n643 ^ n612 ;
  assign n645 = n642 & ~n644 ;
  assign n646 = n645 ^ n641 ;
  assign n674 = n673 ^ n646 ;
  assign n597 = n575 ^ n574 ;
  assign n598 = n577 & ~n597 ;
  assign n599 = n598 ^ n576 ;
  assign n594 = n584 ^ n578 ;
  assign n595 = ~n579 & n594 ;
  assign n596 = n595 ^ n584 ;
  assign n600 = n599 ^ n596 ;
  assign n591 = n581 ^ n580 ;
  assign n592 = n583 & ~n591 ;
  assign n593 = n592 ^ n582 ;
  assign n601 = n600 ^ n593 ;
  assign n564 = n556 ^ n555 ;
  assign n565 = n558 & ~n564 ;
  assign n566 = n565 ^ n557 ;
  assign n560 = n559 ^ n552 ;
  assign n561 = n554 & ~n560 ;
  assign n562 = n561 ^ n553 ;
  assign n549 = n548 ^ n545 ;
  assign n550 = n547 & ~n549 ;
  assign n551 = n550 ^ n546 ;
  assign n563 = n562 ^ n551 ;
  assign n589 = n566 ^ n563 ;
  assign n586 = n585 ^ n570 ;
  assign n587 = n572 & ~n586 ;
  assign n588 = n587 ^ n571 ;
  assign n590 = n589 ^ n588 ;
  assign n675 = n601 ^ n590 ;
  assign n676 = n675 ^ n673 ;
  assign n677 = n674 & ~n676 ;
  assign n678 = n677 ^ n646 ;
  assign n690 = n689 ^ n678 ;
  assign n606 = n596 ^ n593 ;
  assign n607 = n600 & ~n606 ;
  assign n608 = n607 ^ n599 ;
  assign n602 = n601 ^ n589 ;
  assign n603 = n590 & ~n602 ;
  assign n604 = n603 ^ n588 ;
  assign n567 = n566 ^ n551 ;
  assign n568 = n563 & ~n567 ;
  assign n569 = n568 ^ n562 ;
  assign n605 = n604 ^ n569 ;
  assign n691 = n608 ^ n605 ;
  assign n692 = n691 ^ n678 ;
  assign n693 = n690 & ~n692 ;
  assign n694 = n693 ^ n689 ;
  assign n698 = n697 ^ n694 ;
  assign n609 = n608 ^ n569 ;
  assign n610 = n605 & ~n609 ;
  assign n611 = n610 ^ n604 ;
  assign n699 = n698 ^ n611 ;
  assign n700 = n675 ^ n674 ;
  assign n701 = n643 ^ n642 ;
  assign n702 = x512 ^ x0 ;
  assign n703 = n701 & n702 ;
  assign n704 = n700 & n703 ;
  assign n705 = n691 ^ n690 ;
  assign n706 = n704 & n705 ;
  assign n707 = n699 & n706 ;
  assign n708 = n697 ^ n611 ;
  assign n709 = ~n698 & n708 ;
  assign n710 = n709 ^ n611 ;
  assign n711 = n707 & n710 ;
  assign n968 = x541 ^ x125 ;
  assign n967 = x542 ^ x126 ;
  assign n969 = n968 ^ n967 ;
  assign n966 = x543 ^ x127 ;
  assign n1001 = n967 ^ n966 ;
  assign n1002 = n969 & ~n1001 ;
  assign n1003 = n1002 ^ n968 ;
  assign n971 = x537 ^ x121 ;
  assign n970 = n969 ^ n966 ;
  assign n972 = n971 ^ n970 ;
  assign n963 = x539 ^ x123 ;
  assign n962 = x538 ^ x122 ;
  assign n964 = n963 ^ n962 ;
  assign n961 = x540 ^ x124 ;
  assign n965 = n964 ^ n961 ;
  assign n998 = n970 ^ n965 ;
  assign n999 = n972 & ~n998 ;
  assign n1000 = n999 ^ n971 ;
  assign n1004 = n1003 ^ n1000 ;
  assign n995 = n962 ^ n961 ;
  assign n996 = n964 & ~n995 ;
  assign n997 = n996 ^ n963 ;
  assign n1019 = n1000 ^ n997 ;
  assign n1020 = n1004 & ~n1019 ;
  assign n1021 = n1020 ^ n1003 ;
  assign n1005 = n1004 ^ n997 ;
  assign n973 = n972 ^ n965 ;
  assign n960 = x529 ^ x113 ;
  assign n974 = n973 ^ n960 ;
  assign n955 = x535 ^ x119 ;
  assign n954 = x534 ^ x118 ;
  assign n956 = n955 ^ n954 ;
  assign n953 = x536 ^ x120 ;
  assign n957 = n956 ^ n953 ;
  assign n952 = x530 ^ x114 ;
  assign n958 = n957 ^ n952 ;
  assign n949 = x532 ^ x116 ;
  assign n948 = x531 ^ x115 ;
  assign n950 = n949 ^ n948 ;
  assign n947 = x533 ^ x117 ;
  assign n951 = n950 ^ n947 ;
  assign n959 = n958 ^ n951 ;
  assign n992 = n960 ^ n959 ;
  assign n993 = n974 & ~n992 ;
  assign n994 = n993 ^ n973 ;
  assign n1006 = n1005 ^ n994 ;
  assign n987 = n952 ^ n951 ;
  assign n988 = n958 & ~n987 ;
  assign n989 = n988 ^ n957 ;
  assign n984 = n954 ^ n953 ;
  assign n985 = n956 & ~n984 ;
  assign n986 = n985 ^ n955 ;
  assign n990 = n989 ^ n986 ;
  assign n981 = n948 ^ n947 ;
  assign n982 = n950 & ~n981 ;
  assign n983 = n982 ^ n949 ;
  assign n991 = n990 ^ n983 ;
  assign n1016 = n1005 ^ n991 ;
  assign n1017 = n1006 & ~n1016 ;
  assign n1018 = n1017 ^ n994 ;
  assign n1022 = n1021 ^ n1018 ;
  assign n1013 = n986 ^ n983 ;
  assign n1014 = n990 & ~n1013 ;
  assign n1015 = n1014 ^ n989 ;
  assign n1029 = n1018 ^ n1015 ;
  assign n1030 = n1022 & ~n1029 ;
  assign n1031 = n1030 ^ n1021 ;
  assign n1023 = n1022 ^ n1015 ;
  assign n1007 = n1006 ^ n991 ;
  assign n975 = n974 ^ n959 ;
  assign n946 = x513 ^ x97 ;
  assign n976 = n975 ^ n946 ;
  assign n916 = x517 ^ x101 ;
  assign n915 = x516 ^ x100 ;
  assign n917 = n916 ^ n915 ;
  assign n914 = x518 ^ x102 ;
  assign n918 = n917 ^ n914 ;
  assign n910 = x520 ^ x104 ;
  assign n909 = x519 ^ x103 ;
  assign n911 = n910 ^ n909 ;
  assign n908 = x521 ^ x105 ;
  assign n912 = n911 ^ n908 ;
  assign n907 = x515 ^ x99 ;
  assign n913 = n912 ^ n907 ;
  assign n919 = n918 ^ n913 ;
  assign n905 = x514 ^ x98 ;
  assign n891 = x524 ^ x108 ;
  assign n890 = x523 ^ x107 ;
  assign n892 = n891 ^ n890 ;
  assign n889 = x525 ^ x109 ;
  assign n893 = n892 ^ n889 ;
  assign n882 = x528 ^ x112 ;
  assign n880 = x527 ^ x111 ;
  assign n879 = x526 ^ x110 ;
  assign n881 = n880 ^ n879 ;
  assign n887 = n882 ^ n881 ;
  assign n886 = x522 ^ x106 ;
  assign n888 = n887 ^ n886 ;
  assign n904 = n893 ^ n888 ;
  assign n906 = n905 ^ n904 ;
  assign n977 = n919 ^ n906 ;
  assign n978 = n977 ^ n946 ;
  assign n979 = n976 & ~n978 ;
  assign n980 = n979 ^ n975 ;
  assign n1008 = n1007 ^ n980 ;
  assign n931 = n909 ^ n908 ;
  assign n932 = n911 & ~n931 ;
  assign n933 = n932 ^ n910 ;
  assign n928 = n918 ^ n912 ;
  assign n929 = ~n913 & n928 ;
  assign n930 = n929 ^ n918 ;
  assign n934 = n933 ^ n930 ;
  assign n925 = n915 ^ n914 ;
  assign n926 = n917 & ~n925 ;
  assign n927 = n926 ^ n916 ;
  assign n935 = n934 ^ n927 ;
  assign n898 = n890 ^ n889 ;
  assign n899 = n892 & ~n898 ;
  assign n900 = n899 ^ n891 ;
  assign n894 = n893 ^ n886 ;
  assign n895 = n888 & ~n894 ;
  assign n896 = n895 ^ n887 ;
  assign n883 = n882 ^ n879 ;
  assign n884 = n881 & ~n883 ;
  assign n885 = n884 ^ n880 ;
  assign n897 = n896 ^ n885 ;
  assign n923 = n900 ^ n897 ;
  assign n920 = n919 ^ n904 ;
  assign n921 = n906 & ~n920 ;
  assign n922 = n921 ^ n905 ;
  assign n924 = n923 ^ n922 ;
  assign n1009 = n935 ^ n924 ;
  assign n1010 = n1009 ^ n1007 ;
  assign n1011 = n1008 & ~n1010 ;
  assign n1012 = n1011 ^ n980 ;
  assign n1024 = n1023 ^ n1012 ;
  assign n940 = n930 ^ n927 ;
  assign n941 = n934 & ~n940 ;
  assign n942 = n941 ^ n933 ;
  assign n936 = n935 ^ n923 ;
  assign n937 = n924 & ~n936 ;
  assign n938 = n937 ^ n922 ;
  assign n901 = n900 ^ n885 ;
  assign n902 = n897 & ~n901 ;
  assign n903 = n902 ^ n896 ;
  assign n939 = n938 ^ n903 ;
  assign n1025 = n942 ^ n939 ;
  assign n1026 = n1025 ^ n1012 ;
  assign n1027 = n1024 & ~n1026 ;
  assign n1028 = n1027 ^ n1023 ;
  assign n1032 = n1031 ^ n1028 ;
  assign n943 = n942 ^ n903 ;
  assign n944 = n939 & ~n943 ;
  assign n945 = n944 ^ n938 ;
  assign n1033 = n1032 ^ n945 ;
  assign n1034 = n1009 ^ n1008 ;
  assign n1035 = n977 ^ n976 ;
  assign n1036 = x512 ^ x96 ;
  assign n1037 = n1035 & n1036 ;
  assign n1038 = n1034 & n1037 ;
  assign n1039 = n1025 ^ n1024 ;
  assign n1040 = n1038 & n1039 ;
  assign n1041 = n1033 & n1040 ;
  assign n1042 = n1031 ^ n945 ;
  assign n1043 = ~n1032 & n1042 ;
  assign n1044 = n1043 ^ n945 ;
  assign n1045 = n1041 & n1044 ;
  assign n3025 = x541 ^ x189 ;
  assign n3024 = x542 ^ x190 ;
  assign n3026 = n3025 ^ n3024 ;
  assign n3023 = x543 ^ x191 ;
  assign n3058 = n3024 ^ n3023 ;
  assign n3059 = n3026 & ~n3058 ;
  assign n3060 = n3059 ^ n3025 ;
  assign n3028 = x537 ^ x185 ;
  assign n3027 = n3026 ^ n3023 ;
  assign n3029 = n3028 ^ n3027 ;
  assign n3020 = x539 ^ x187 ;
  assign n3019 = x538 ^ x186 ;
  assign n3021 = n3020 ^ n3019 ;
  assign n3018 = x540 ^ x188 ;
  assign n3022 = n3021 ^ n3018 ;
  assign n3055 = n3027 ^ n3022 ;
  assign n3056 = n3029 & ~n3055 ;
  assign n3057 = n3056 ^ n3028 ;
  assign n3061 = n3060 ^ n3057 ;
  assign n3052 = n3019 ^ n3018 ;
  assign n3053 = n3021 & ~n3052 ;
  assign n3054 = n3053 ^ n3020 ;
  assign n3076 = n3057 ^ n3054 ;
  assign n3077 = n3061 & ~n3076 ;
  assign n3078 = n3077 ^ n3060 ;
  assign n3062 = n3061 ^ n3054 ;
  assign n3030 = n3029 ^ n3022 ;
  assign n3017 = x529 ^ x177 ;
  assign n3031 = n3030 ^ n3017 ;
  assign n3012 = x535 ^ x183 ;
  assign n3011 = x534 ^ x182 ;
  assign n3013 = n3012 ^ n3011 ;
  assign n3010 = x536 ^ x184 ;
  assign n3014 = n3013 ^ n3010 ;
  assign n3009 = x530 ^ x178 ;
  assign n3015 = n3014 ^ n3009 ;
  assign n3006 = x532 ^ x180 ;
  assign n3005 = x531 ^ x179 ;
  assign n3007 = n3006 ^ n3005 ;
  assign n3004 = x533 ^ x181 ;
  assign n3008 = n3007 ^ n3004 ;
  assign n3016 = n3015 ^ n3008 ;
  assign n3049 = n3017 ^ n3016 ;
  assign n3050 = n3031 & ~n3049 ;
  assign n3051 = n3050 ^ n3030 ;
  assign n3063 = n3062 ^ n3051 ;
  assign n3044 = n3009 ^ n3008 ;
  assign n3045 = n3015 & ~n3044 ;
  assign n3046 = n3045 ^ n3014 ;
  assign n3041 = n3011 ^ n3010 ;
  assign n3042 = n3013 & ~n3041 ;
  assign n3043 = n3042 ^ n3012 ;
  assign n3047 = n3046 ^ n3043 ;
  assign n3038 = n3005 ^ n3004 ;
  assign n3039 = n3007 & ~n3038 ;
  assign n3040 = n3039 ^ n3006 ;
  assign n3048 = n3047 ^ n3040 ;
  assign n3073 = n3062 ^ n3048 ;
  assign n3074 = n3063 & ~n3073 ;
  assign n3075 = n3074 ^ n3051 ;
  assign n3079 = n3078 ^ n3075 ;
  assign n3070 = n3043 ^ n3040 ;
  assign n3071 = n3047 & ~n3070 ;
  assign n3072 = n3071 ^ n3046 ;
  assign n3086 = n3075 ^ n3072 ;
  assign n3087 = n3079 & ~n3086 ;
  assign n3088 = n3087 ^ n3078 ;
  assign n3080 = n3079 ^ n3072 ;
  assign n3064 = n3063 ^ n3048 ;
  assign n3032 = n3031 ^ n3016 ;
  assign n3003 = x513 ^ x161 ;
  assign n3033 = n3032 ^ n3003 ;
  assign n2973 = x517 ^ x165 ;
  assign n2972 = x516 ^ x164 ;
  assign n2974 = n2973 ^ n2972 ;
  assign n2971 = x518 ^ x166 ;
  assign n2975 = n2974 ^ n2971 ;
  assign n2967 = x520 ^ x168 ;
  assign n2966 = x519 ^ x167 ;
  assign n2968 = n2967 ^ n2966 ;
  assign n2965 = x521 ^ x169 ;
  assign n2969 = n2968 ^ n2965 ;
  assign n2964 = x515 ^ x163 ;
  assign n2970 = n2969 ^ n2964 ;
  assign n2976 = n2975 ^ n2970 ;
  assign n2962 = x514 ^ x162 ;
  assign n2948 = x524 ^ x172 ;
  assign n2947 = x523 ^ x171 ;
  assign n2949 = n2948 ^ n2947 ;
  assign n2946 = x525 ^ x173 ;
  assign n2950 = n2949 ^ n2946 ;
  assign n2939 = x528 ^ x176 ;
  assign n2937 = x527 ^ x175 ;
  assign n2936 = x526 ^ x174 ;
  assign n2938 = n2937 ^ n2936 ;
  assign n2944 = n2939 ^ n2938 ;
  assign n2943 = x522 ^ x170 ;
  assign n2945 = n2944 ^ n2943 ;
  assign n2961 = n2950 ^ n2945 ;
  assign n2963 = n2962 ^ n2961 ;
  assign n3034 = n2976 ^ n2963 ;
  assign n3035 = n3034 ^ n3003 ;
  assign n3036 = n3033 & ~n3035 ;
  assign n3037 = n3036 ^ n3032 ;
  assign n3065 = n3064 ^ n3037 ;
  assign n2988 = n2966 ^ n2965 ;
  assign n2989 = n2968 & ~n2988 ;
  assign n2990 = n2989 ^ n2967 ;
  assign n2985 = n2975 ^ n2969 ;
  assign n2986 = ~n2970 & n2985 ;
  assign n2987 = n2986 ^ n2975 ;
  assign n2991 = n2990 ^ n2987 ;
  assign n2982 = n2972 ^ n2971 ;
  assign n2983 = n2974 & ~n2982 ;
  assign n2984 = n2983 ^ n2973 ;
  assign n2992 = n2991 ^ n2984 ;
  assign n2955 = n2947 ^ n2946 ;
  assign n2956 = n2949 & ~n2955 ;
  assign n2957 = n2956 ^ n2948 ;
  assign n2951 = n2950 ^ n2943 ;
  assign n2952 = n2945 & ~n2951 ;
  assign n2953 = n2952 ^ n2944 ;
  assign n2940 = n2939 ^ n2936 ;
  assign n2941 = n2938 & ~n2940 ;
  assign n2942 = n2941 ^ n2937 ;
  assign n2954 = n2953 ^ n2942 ;
  assign n2980 = n2957 ^ n2954 ;
  assign n2977 = n2976 ^ n2961 ;
  assign n2978 = n2963 & ~n2977 ;
  assign n2979 = n2978 ^ n2962 ;
  assign n2981 = n2980 ^ n2979 ;
  assign n3066 = n2992 ^ n2981 ;
  assign n3067 = n3066 ^ n3064 ;
  assign n3068 = n3065 & ~n3067 ;
  assign n3069 = n3068 ^ n3037 ;
  assign n3081 = n3080 ^ n3069 ;
  assign n2997 = n2987 ^ n2984 ;
  assign n2998 = n2991 & ~n2997 ;
  assign n2999 = n2998 ^ n2990 ;
  assign n2993 = n2992 ^ n2980 ;
  assign n2994 = n2981 & ~n2993 ;
  assign n2995 = n2994 ^ n2979 ;
  assign n2958 = n2957 ^ n2942 ;
  assign n2959 = n2954 & ~n2958 ;
  assign n2960 = n2959 ^ n2953 ;
  assign n2996 = n2995 ^ n2960 ;
  assign n3082 = n2999 ^ n2996 ;
  assign n3083 = n3082 ^ n3069 ;
  assign n3084 = n3081 & ~n3083 ;
  assign n3085 = n3084 ^ n3080 ;
  assign n3089 = n3088 ^ n3085 ;
  assign n3000 = n2999 ^ n2960 ;
  assign n3001 = n2996 & ~n3000 ;
  assign n3002 = n3001 ^ n2995 ;
  assign n3090 = n3089 ^ n3002 ;
  assign n3091 = n3066 ^ n3065 ;
  assign n3092 = n3034 ^ n3033 ;
  assign n3093 = x512 ^ x160 ;
  assign n3094 = n3092 & n3093 ;
  assign n3095 = n3091 & n3094 ;
  assign n3096 = n3082 ^ n3081 ;
  assign n3097 = n3095 & n3096 ;
  assign n3098 = n3090 & n3097 ;
  assign n3099 = n3088 ^ n3002 ;
  assign n3100 = ~n3089 & n3099 ;
  assign n3101 = n3100 ^ n3002 ;
  assign n3102 = n3098 & n3101 ;
  assign n1302 = x541 ^ x221 ;
  assign n1301 = x542 ^ x222 ;
  assign n1303 = n1302 ^ n1301 ;
  assign n1300 = x543 ^ x223 ;
  assign n1335 = n1301 ^ n1300 ;
  assign n1336 = n1303 & ~n1335 ;
  assign n1337 = n1336 ^ n1302 ;
  assign n1305 = x537 ^ x217 ;
  assign n1304 = n1303 ^ n1300 ;
  assign n1306 = n1305 ^ n1304 ;
  assign n1297 = x539 ^ x219 ;
  assign n1296 = x538 ^ x218 ;
  assign n1298 = n1297 ^ n1296 ;
  assign n1295 = x540 ^ x220 ;
  assign n1299 = n1298 ^ n1295 ;
  assign n1332 = n1304 ^ n1299 ;
  assign n1333 = n1306 & ~n1332 ;
  assign n1334 = n1333 ^ n1305 ;
  assign n1338 = n1337 ^ n1334 ;
  assign n1329 = n1296 ^ n1295 ;
  assign n1330 = n1298 & ~n1329 ;
  assign n1331 = n1330 ^ n1297 ;
  assign n1353 = n1334 ^ n1331 ;
  assign n1354 = n1338 & ~n1353 ;
  assign n1355 = n1354 ^ n1337 ;
  assign n1339 = n1338 ^ n1331 ;
  assign n1307 = n1306 ^ n1299 ;
  assign n1294 = x529 ^ x209 ;
  assign n1308 = n1307 ^ n1294 ;
  assign n1289 = x535 ^ x215 ;
  assign n1288 = x534 ^ x214 ;
  assign n1290 = n1289 ^ n1288 ;
  assign n1287 = x536 ^ x216 ;
  assign n1291 = n1290 ^ n1287 ;
  assign n1286 = x530 ^ x210 ;
  assign n1292 = n1291 ^ n1286 ;
  assign n1283 = x532 ^ x212 ;
  assign n1282 = x531 ^ x211 ;
  assign n1284 = n1283 ^ n1282 ;
  assign n1281 = x533 ^ x213 ;
  assign n1285 = n1284 ^ n1281 ;
  assign n1293 = n1292 ^ n1285 ;
  assign n1326 = n1294 ^ n1293 ;
  assign n1327 = n1308 & ~n1326 ;
  assign n1328 = n1327 ^ n1307 ;
  assign n1340 = n1339 ^ n1328 ;
  assign n1321 = n1286 ^ n1285 ;
  assign n1322 = n1292 & ~n1321 ;
  assign n1323 = n1322 ^ n1291 ;
  assign n1318 = n1288 ^ n1287 ;
  assign n1319 = n1290 & ~n1318 ;
  assign n1320 = n1319 ^ n1289 ;
  assign n1324 = n1323 ^ n1320 ;
  assign n1315 = n1282 ^ n1281 ;
  assign n1316 = n1284 & ~n1315 ;
  assign n1317 = n1316 ^ n1283 ;
  assign n1325 = n1324 ^ n1317 ;
  assign n1350 = n1339 ^ n1325 ;
  assign n1351 = n1340 & ~n1350 ;
  assign n1352 = n1351 ^ n1328 ;
  assign n1356 = n1355 ^ n1352 ;
  assign n1347 = n1320 ^ n1317 ;
  assign n1348 = n1324 & ~n1347 ;
  assign n1349 = n1348 ^ n1323 ;
  assign n1363 = n1352 ^ n1349 ;
  assign n1364 = n1356 & ~n1363 ;
  assign n1365 = n1364 ^ n1355 ;
  assign n1357 = n1356 ^ n1349 ;
  assign n1341 = n1340 ^ n1325 ;
  assign n1309 = n1308 ^ n1293 ;
  assign n1280 = x513 ^ x193 ;
  assign n1310 = n1309 ^ n1280 ;
  assign n1250 = x517 ^ x197 ;
  assign n1249 = x516 ^ x196 ;
  assign n1251 = n1250 ^ n1249 ;
  assign n1248 = x518 ^ x198 ;
  assign n1252 = n1251 ^ n1248 ;
  assign n1244 = x520 ^ x200 ;
  assign n1243 = x519 ^ x199 ;
  assign n1245 = n1244 ^ n1243 ;
  assign n1242 = x521 ^ x201 ;
  assign n1246 = n1245 ^ n1242 ;
  assign n1241 = x515 ^ x195 ;
  assign n1247 = n1246 ^ n1241 ;
  assign n1253 = n1252 ^ n1247 ;
  assign n1239 = x514 ^ x194 ;
  assign n1225 = x524 ^ x204 ;
  assign n1224 = x523 ^ x203 ;
  assign n1226 = n1225 ^ n1224 ;
  assign n1223 = x525 ^ x205 ;
  assign n1227 = n1226 ^ n1223 ;
  assign n1216 = x528 ^ x208 ;
  assign n1214 = x527 ^ x207 ;
  assign n1213 = x526 ^ x206 ;
  assign n1215 = n1214 ^ n1213 ;
  assign n1221 = n1216 ^ n1215 ;
  assign n1220 = x522 ^ x202 ;
  assign n1222 = n1221 ^ n1220 ;
  assign n1238 = n1227 ^ n1222 ;
  assign n1240 = n1239 ^ n1238 ;
  assign n1311 = n1253 ^ n1240 ;
  assign n1312 = n1311 ^ n1280 ;
  assign n1313 = n1310 & ~n1312 ;
  assign n1314 = n1313 ^ n1309 ;
  assign n1342 = n1341 ^ n1314 ;
  assign n1265 = n1243 ^ n1242 ;
  assign n1266 = n1245 & ~n1265 ;
  assign n1267 = n1266 ^ n1244 ;
  assign n1262 = n1252 ^ n1246 ;
  assign n1263 = ~n1247 & n1262 ;
  assign n1264 = n1263 ^ n1252 ;
  assign n1268 = n1267 ^ n1264 ;
  assign n1259 = n1249 ^ n1248 ;
  assign n1260 = n1251 & ~n1259 ;
  assign n1261 = n1260 ^ n1250 ;
  assign n1269 = n1268 ^ n1261 ;
  assign n1232 = n1224 ^ n1223 ;
  assign n1233 = n1226 & ~n1232 ;
  assign n1234 = n1233 ^ n1225 ;
  assign n1228 = n1227 ^ n1220 ;
  assign n1229 = n1222 & ~n1228 ;
  assign n1230 = n1229 ^ n1221 ;
  assign n1217 = n1216 ^ n1213 ;
  assign n1218 = n1215 & ~n1217 ;
  assign n1219 = n1218 ^ n1214 ;
  assign n1231 = n1230 ^ n1219 ;
  assign n1257 = n1234 ^ n1231 ;
  assign n1254 = n1253 ^ n1238 ;
  assign n1255 = n1240 & ~n1254 ;
  assign n1256 = n1255 ^ n1239 ;
  assign n1258 = n1257 ^ n1256 ;
  assign n1343 = n1269 ^ n1258 ;
  assign n1344 = n1343 ^ n1341 ;
  assign n1345 = n1342 & ~n1344 ;
  assign n1346 = n1345 ^ n1314 ;
  assign n1358 = n1357 ^ n1346 ;
  assign n1274 = n1264 ^ n1261 ;
  assign n1275 = n1268 & ~n1274 ;
  assign n1276 = n1275 ^ n1267 ;
  assign n1270 = n1269 ^ n1257 ;
  assign n1271 = n1258 & ~n1270 ;
  assign n1272 = n1271 ^ n1256 ;
  assign n1235 = n1234 ^ n1219 ;
  assign n1236 = n1231 & ~n1235 ;
  assign n1237 = n1236 ^ n1230 ;
  assign n1273 = n1272 ^ n1237 ;
  assign n1359 = n1276 ^ n1273 ;
  assign n1360 = n1359 ^ n1346 ;
  assign n1361 = n1358 & ~n1360 ;
  assign n1362 = n1361 ^ n1357 ;
  assign n1366 = n1365 ^ n1362 ;
  assign n1277 = n1276 ^ n1237 ;
  assign n1278 = n1273 & ~n1277 ;
  assign n1279 = n1278 ^ n1272 ;
  assign n1367 = n1366 ^ n1279 ;
  assign n1368 = n1343 ^ n1342 ;
  assign n1369 = n1311 ^ n1310 ;
  assign n1370 = x512 ^ x192 ;
  assign n1371 = n1369 & n1370 ;
  assign n1372 = n1368 & n1371 ;
  assign n1373 = n1359 ^ n1358 ;
  assign n1374 = n1372 & n1373 ;
  assign n1375 = n1367 & n1374 ;
  assign n1376 = n1365 ^ n1279 ;
  assign n1377 = ~n1366 & n1376 ;
  assign n1378 = n1377 ^ n1279 ;
  assign n1379 = n1375 & n1378 ;
  assign n2840 = x541 ^ x285 ;
  assign n2839 = x542 ^ x286 ;
  assign n2841 = n2840 ^ n2839 ;
  assign n2838 = x543 ^ x287 ;
  assign n2873 = n2839 ^ n2838 ;
  assign n2874 = n2841 & ~n2873 ;
  assign n2875 = n2874 ^ n2840 ;
  assign n2843 = x537 ^ x281 ;
  assign n2842 = n2841 ^ n2838 ;
  assign n2844 = n2843 ^ n2842 ;
  assign n2835 = x539 ^ x283 ;
  assign n2834 = x538 ^ x282 ;
  assign n2836 = n2835 ^ n2834 ;
  assign n2833 = x540 ^ x284 ;
  assign n2837 = n2836 ^ n2833 ;
  assign n2870 = n2842 ^ n2837 ;
  assign n2871 = n2844 & ~n2870 ;
  assign n2872 = n2871 ^ n2843 ;
  assign n2876 = n2875 ^ n2872 ;
  assign n2867 = n2834 ^ n2833 ;
  assign n2868 = n2836 & ~n2867 ;
  assign n2869 = n2868 ^ n2835 ;
  assign n2891 = n2872 ^ n2869 ;
  assign n2892 = n2876 & ~n2891 ;
  assign n2893 = n2892 ^ n2875 ;
  assign n2877 = n2876 ^ n2869 ;
  assign n2845 = n2844 ^ n2837 ;
  assign n2832 = x529 ^ x273 ;
  assign n2846 = n2845 ^ n2832 ;
  assign n2827 = x535 ^ x279 ;
  assign n2826 = x534 ^ x278 ;
  assign n2828 = n2827 ^ n2826 ;
  assign n2825 = x536 ^ x280 ;
  assign n2829 = n2828 ^ n2825 ;
  assign n2824 = x530 ^ x274 ;
  assign n2830 = n2829 ^ n2824 ;
  assign n2821 = x532 ^ x276 ;
  assign n2820 = x531 ^ x275 ;
  assign n2822 = n2821 ^ n2820 ;
  assign n2819 = x533 ^ x277 ;
  assign n2823 = n2822 ^ n2819 ;
  assign n2831 = n2830 ^ n2823 ;
  assign n2864 = n2832 ^ n2831 ;
  assign n2865 = n2846 & ~n2864 ;
  assign n2866 = n2865 ^ n2845 ;
  assign n2878 = n2877 ^ n2866 ;
  assign n2859 = n2824 ^ n2823 ;
  assign n2860 = n2830 & ~n2859 ;
  assign n2861 = n2860 ^ n2829 ;
  assign n2856 = n2826 ^ n2825 ;
  assign n2857 = n2828 & ~n2856 ;
  assign n2858 = n2857 ^ n2827 ;
  assign n2862 = n2861 ^ n2858 ;
  assign n2853 = n2820 ^ n2819 ;
  assign n2854 = n2822 & ~n2853 ;
  assign n2855 = n2854 ^ n2821 ;
  assign n2863 = n2862 ^ n2855 ;
  assign n2888 = n2877 ^ n2863 ;
  assign n2889 = n2878 & ~n2888 ;
  assign n2890 = n2889 ^ n2866 ;
  assign n2894 = n2893 ^ n2890 ;
  assign n2885 = n2858 ^ n2855 ;
  assign n2886 = n2862 & ~n2885 ;
  assign n2887 = n2886 ^ n2861 ;
  assign n2901 = n2890 ^ n2887 ;
  assign n2902 = n2894 & ~n2901 ;
  assign n2903 = n2902 ^ n2893 ;
  assign n2895 = n2894 ^ n2887 ;
  assign n2879 = n2878 ^ n2863 ;
  assign n2847 = n2846 ^ n2831 ;
  assign n2818 = x513 ^ x257 ;
  assign n2848 = n2847 ^ n2818 ;
  assign n2788 = x517 ^ x261 ;
  assign n2787 = x516 ^ x260 ;
  assign n2789 = n2788 ^ n2787 ;
  assign n2786 = x518 ^ x262 ;
  assign n2790 = n2789 ^ n2786 ;
  assign n2782 = x520 ^ x264 ;
  assign n2781 = x519 ^ x263 ;
  assign n2783 = n2782 ^ n2781 ;
  assign n2780 = x521 ^ x265 ;
  assign n2784 = n2783 ^ n2780 ;
  assign n2779 = x515 ^ x259 ;
  assign n2785 = n2784 ^ n2779 ;
  assign n2791 = n2790 ^ n2785 ;
  assign n2777 = x514 ^ x258 ;
  assign n2763 = x524 ^ x268 ;
  assign n2762 = x523 ^ x267 ;
  assign n2764 = n2763 ^ n2762 ;
  assign n2761 = x525 ^ x269 ;
  assign n2765 = n2764 ^ n2761 ;
  assign n2754 = x528 ^ x272 ;
  assign n2752 = x527 ^ x271 ;
  assign n2751 = x526 ^ x270 ;
  assign n2753 = n2752 ^ n2751 ;
  assign n2759 = n2754 ^ n2753 ;
  assign n2758 = x522 ^ x266 ;
  assign n2760 = n2759 ^ n2758 ;
  assign n2776 = n2765 ^ n2760 ;
  assign n2778 = n2777 ^ n2776 ;
  assign n2849 = n2791 ^ n2778 ;
  assign n2850 = n2849 ^ n2818 ;
  assign n2851 = n2848 & ~n2850 ;
  assign n2852 = n2851 ^ n2847 ;
  assign n2880 = n2879 ^ n2852 ;
  assign n2803 = n2781 ^ n2780 ;
  assign n2804 = n2783 & ~n2803 ;
  assign n2805 = n2804 ^ n2782 ;
  assign n2800 = n2790 ^ n2784 ;
  assign n2801 = ~n2785 & n2800 ;
  assign n2802 = n2801 ^ n2790 ;
  assign n2806 = n2805 ^ n2802 ;
  assign n2797 = n2787 ^ n2786 ;
  assign n2798 = n2789 & ~n2797 ;
  assign n2799 = n2798 ^ n2788 ;
  assign n2807 = n2806 ^ n2799 ;
  assign n2770 = n2762 ^ n2761 ;
  assign n2771 = n2764 & ~n2770 ;
  assign n2772 = n2771 ^ n2763 ;
  assign n2766 = n2765 ^ n2758 ;
  assign n2767 = n2760 & ~n2766 ;
  assign n2768 = n2767 ^ n2759 ;
  assign n2755 = n2754 ^ n2751 ;
  assign n2756 = n2753 & ~n2755 ;
  assign n2757 = n2756 ^ n2752 ;
  assign n2769 = n2768 ^ n2757 ;
  assign n2795 = n2772 ^ n2769 ;
  assign n2792 = n2791 ^ n2776 ;
  assign n2793 = n2778 & ~n2792 ;
  assign n2794 = n2793 ^ n2777 ;
  assign n2796 = n2795 ^ n2794 ;
  assign n2881 = n2807 ^ n2796 ;
  assign n2882 = n2881 ^ n2879 ;
  assign n2883 = n2880 & ~n2882 ;
  assign n2884 = n2883 ^ n2852 ;
  assign n2896 = n2895 ^ n2884 ;
  assign n2812 = n2802 ^ n2799 ;
  assign n2813 = n2806 & ~n2812 ;
  assign n2814 = n2813 ^ n2805 ;
  assign n2808 = n2807 ^ n2795 ;
  assign n2809 = n2796 & ~n2808 ;
  assign n2810 = n2809 ^ n2794 ;
  assign n2773 = n2772 ^ n2757 ;
  assign n2774 = n2769 & ~n2773 ;
  assign n2775 = n2774 ^ n2768 ;
  assign n2811 = n2810 ^ n2775 ;
  assign n2897 = n2814 ^ n2811 ;
  assign n2898 = n2897 ^ n2884 ;
  assign n2899 = n2896 & ~n2898 ;
  assign n2900 = n2899 ^ n2895 ;
  assign n2904 = n2903 ^ n2900 ;
  assign n2815 = n2814 ^ n2775 ;
  assign n2816 = n2811 & ~n2815 ;
  assign n2817 = n2816 ^ n2810 ;
  assign n2905 = n2904 ^ n2817 ;
  assign n2906 = n2881 ^ n2880 ;
  assign n2907 = n2849 ^ n2848 ;
  assign n2908 = x512 ^ x256 ;
  assign n2909 = n2907 & n2908 ;
  assign n2910 = n2906 & n2909 ;
  assign n2911 = n2897 ^ n2896 ;
  assign n2912 = n2910 & n2911 ;
  assign n2913 = n2905 & n2912 ;
  assign n2914 = n2903 ^ n2817 ;
  assign n2915 = ~n2904 & n2914 ;
  assign n2916 = n2915 ^ n2817 ;
  assign n2917 = n2913 & n2916 ;
  assign n1636 = x541 ^ x317 ;
  assign n1635 = x542 ^ x318 ;
  assign n1637 = n1636 ^ n1635 ;
  assign n1634 = x543 ^ x319 ;
  assign n1669 = n1635 ^ n1634 ;
  assign n1670 = n1637 & ~n1669 ;
  assign n1671 = n1670 ^ n1636 ;
  assign n1639 = x537 ^ x313 ;
  assign n1638 = n1637 ^ n1634 ;
  assign n1640 = n1639 ^ n1638 ;
  assign n1631 = x539 ^ x315 ;
  assign n1630 = x538 ^ x314 ;
  assign n1632 = n1631 ^ n1630 ;
  assign n1629 = x540 ^ x316 ;
  assign n1633 = n1632 ^ n1629 ;
  assign n1666 = n1638 ^ n1633 ;
  assign n1667 = n1640 & ~n1666 ;
  assign n1668 = n1667 ^ n1639 ;
  assign n1672 = n1671 ^ n1668 ;
  assign n1663 = n1630 ^ n1629 ;
  assign n1664 = n1632 & ~n1663 ;
  assign n1665 = n1664 ^ n1631 ;
  assign n1687 = n1668 ^ n1665 ;
  assign n1688 = n1672 & ~n1687 ;
  assign n1689 = n1688 ^ n1671 ;
  assign n1673 = n1672 ^ n1665 ;
  assign n1641 = n1640 ^ n1633 ;
  assign n1628 = x529 ^ x305 ;
  assign n1642 = n1641 ^ n1628 ;
  assign n1623 = x535 ^ x311 ;
  assign n1622 = x534 ^ x310 ;
  assign n1624 = n1623 ^ n1622 ;
  assign n1621 = x536 ^ x312 ;
  assign n1625 = n1624 ^ n1621 ;
  assign n1620 = x530 ^ x306 ;
  assign n1626 = n1625 ^ n1620 ;
  assign n1617 = x532 ^ x308 ;
  assign n1616 = x531 ^ x307 ;
  assign n1618 = n1617 ^ n1616 ;
  assign n1615 = x533 ^ x309 ;
  assign n1619 = n1618 ^ n1615 ;
  assign n1627 = n1626 ^ n1619 ;
  assign n1660 = n1628 ^ n1627 ;
  assign n1661 = n1642 & ~n1660 ;
  assign n1662 = n1661 ^ n1641 ;
  assign n1674 = n1673 ^ n1662 ;
  assign n1655 = n1620 ^ n1619 ;
  assign n1656 = n1626 & ~n1655 ;
  assign n1657 = n1656 ^ n1625 ;
  assign n1652 = n1622 ^ n1621 ;
  assign n1653 = n1624 & ~n1652 ;
  assign n1654 = n1653 ^ n1623 ;
  assign n1658 = n1657 ^ n1654 ;
  assign n1649 = n1616 ^ n1615 ;
  assign n1650 = n1618 & ~n1649 ;
  assign n1651 = n1650 ^ n1617 ;
  assign n1659 = n1658 ^ n1651 ;
  assign n1684 = n1673 ^ n1659 ;
  assign n1685 = n1674 & ~n1684 ;
  assign n1686 = n1685 ^ n1662 ;
  assign n1690 = n1689 ^ n1686 ;
  assign n1681 = n1654 ^ n1651 ;
  assign n1682 = n1658 & ~n1681 ;
  assign n1683 = n1682 ^ n1657 ;
  assign n1697 = n1686 ^ n1683 ;
  assign n1698 = n1690 & ~n1697 ;
  assign n1699 = n1698 ^ n1689 ;
  assign n1691 = n1690 ^ n1683 ;
  assign n1675 = n1674 ^ n1659 ;
  assign n1643 = n1642 ^ n1627 ;
  assign n1614 = x513 ^ x289 ;
  assign n1644 = n1643 ^ n1614 ;
  assign n1584 = x517 ^ x293 ;
  assign n1583 = x516 ^ x292 ;
  assign n1585 = n1584 ^ n1583 ;
  assign n1582 = x518 ^ x294 ;
  assign n1586 = n1585 ^ n1582 ;
  assign n1578 = x520 ^ x296 ;
  assign n1577 = x519 ^ x295 ;
  assign n1579 = n1578 ^ n1577 ;
  assign n1576 = x521 ^ x297 ;
  assign n1580 = n1579 ^ n1576 ;
  assign n1575 = x515 ^ x291 ;
  assign n1581 = n1580 ^ n1575 ;
  assign n1587 = n1586 ^ n1581 ;
  assign n1573 = x514 ^ x290 ;
  assign n1559 = x524 ^ x300 ;
  assign n1558 = x523 ^ x299 ;
  assign n1560 = n1559 ^ n1558 ;
  assign n1557 = x525 ^ x301 ;
  assign n1561 = n1560 ^ n1557 ;
  assign n1550 = x528 ^ x304 ;
  assign n1548 = x527 ^ x303 ;
  assign n1547 = x526 ^ x302 ;
  assign n1549 = n1548 ^ n1547 ;
  assign n1555 = n1550 ^ n1549 ;
  assign n1554 = x522 ^ x298 ;
  assign n1556 = n1555 ^ n1554 ;
  assign n1572 = n1561 ^ n1556 ;
  assign n1574 = n1573 ^ n1572 ;
  assign n1645 = n1587 ^ n1574 ;
  assign n1646 = n1645 ^ n1614 ;
  assign n1647 = n1644 & ~n1646 ;
  assign n1648 = n1647 ^ n1643 ;
  assign n1676 = n1675 ^ n1648 ;
  assign n1599 = n1577 ^ n1576 ;
  assign n1600 = n1579 & ~n1599 ;
  assign n1601 = n1600 ^ n1578 ;
  assign n1596 = n1586 ^ n1580 ;
  assign n1597 = ~n1581 & n1596 ;
  assign n1598 = n1597 ^ n1586 ;
  assign n1602 = n1601 ^ n1598 ;
  assign n1593 = n1583 ^ n1582 ;
  assign n1594 = n1585 & ~n1593 ;
  assign n1595 = n1594 ^ n1584 ;
  assign n1603 = n1602 ^ n1595 ;
  assign n1566 = n1558 ^ n1557 ;
  assign n1567 = n1560 & ~n1566 ;
  assign n1568 = n1567 ^ n1559 ;
  assign n1562 = n1561 ^ n1554 ;
  assign n1563 = n1556 & ~n1562 ;
  assign n1564 = n1563 ^ n1555 ;
  assign n1551 = n1550 ^ n1547 ;
  assign n1552 = n1549 & ~n1551 ;
  assign n1553 = n1552 ^ n1548 ;
  assign n1565 = n1564 ^ n1553 ;
  assign n1591 = n1568 ^ n1565 ;
  assign n1588 = n1587 ^ n1572 ;
  assign n1589 = n1574 & ~n1588 ;
  assign n1590 = n1589 ^ n1573 ;
  assign n1592 = n1591 ^ n1590 ;
  assign n1677 = n1603 ^ n1592 ;
  assign n1678 = n1677 ^ n1675 ;
  assign n1679 = n1676 & ~n1678 ;
  assign n1680 = n1679 ^ n1648 ;
  assign n1692 = n1691 ^ n1680 ;
  assign n1608 = n1598 ^ n1595 ;
  assign n1609 = n1602 & ~n1608 ;
  assign n1610 = n1609 ^ n1601 ;
  assign n1604 = n1603 ^ n1591 ;
  assign n1605 = n1592 & ~n1604 ;
  assign n1606 = n1605 ^ n1590 ;
  assign n1569 = n1568 ^ n1553 ;
  assign n1570 = n1565 & ~n1569 ;
  assign n1571 = n1570 ^ n1564 ;
  assign n1607 = n1606 ^ n1571 ;
  assign n1693 = n1610 ^ n1607 ;
  assign n1694 = n1693 ^ n1680 ;
  assign n1695 = n1692 & ~n1694 ;
  assign n1696 = n1695 ^ n1691 ;
  assign n1700 = n1699 ^ n1696 ;
  assign n1611 = n1610 ^ n1571 ;
  assign n1612 = n1607 & ~n1611 ;
  assign n1613 = n1612 ^ n1606 ;
  assign n1701 = n1700 ^ n1613 ;
  assign n1702 = n1677 ^ n1676 ;
  assign n1703 = n1645 ^ n1644 ;
  assign n1704 = x512 ^ x288 ;
  assign n1705 = n1703 & n1704 ;
  assign n1706 = n1702 & n1705 ;
  assign n1707 = n1693 ^ n1692 ;
  assign n1708 = n1706 & n1707 ;
  assign n1709 = n1701 & n1708 ;
  assign n1710 = n1699 ^ n1613 ;
  assign n1711 = ~n1700 & n1710 ;
  assign n1712 = n1711 ^ n1613 ;
  assign n1713 = n1709 & n1712 ;
  assign n2655 = x541 ^ x381 ;
  assign n2654 = x542 ^ x382 ;
  assign n2656 = n2655 ^ n2654 ;
  assign n2653 = x543 ^ x383 ;
  assign n2688 = n2654 ^ n2653 ;
  assign n2689 = n2656 & ~n2688 ;
  assign n2690 = n2689 ^ n2655 ;
  assign n2658 = x537 ^ x377 ;
  assign n2657 = n2656 ^ n2653 ;
  assign n2659 = n2658 ^ n2657 ;
  assign n2650 = x539 ^ x379 ;
  assign n2649 = x538 ^ x378 ;
  assign n2651 = n2650 ^ n2649 ;
  assign n2648 = x540 ^ x380 ;
  assign n2652 = n2651 ^ n2648 ;
  assign n2685 = n2657 ^ n2652 ;
  assign n2686 = n2659 & ~n2685 ;
  assign n2687 = n2686 ^ n2658 ;
  assign n2691 = n2690 ^ n2687 ;
  assign n2682 = n2649 ^ n2648 ;
  assign n2683 = n2651 & ~n2682 ;
  assign n2684 = n2683 ^ n2650 ;
  assign n2706 = n2687 ^ n2684 ;
  assign n2707 = n2691 & ~n2706 ;
  assign n2708 = n2707 ^ n2690 ;
  assign n2692 = n2691 ^ n2684 ;
  assign n2660 = n2659 ^ n2652 ;
  assign n2647 = x529 ^ x369 ;
  assign n2661 = n2660 ^ n2647 ;
  assign n2642 = x535 ^ x375 ;
  assign n2641 = x534 ^ x374 ;
  assign n2643 = n2642 ^ n2641 ;
  assign n2640 = x536 ^ x376 ;
  assign n2644 = n2643 ^ n2640 ;
  assign n2639 = x530 ^ x370 ;
  assign n2645 = n2644 ^ n2639 ;
  assign n2636 = x532 ^ x372 ;
  assign n2635 = x531 ^ x371 ;
  assign n2637 = n2636 ^ n2635 ;
  assign n2634 = x533 ^ x373 ;
  assign n2638 = n2637 ^ n2634 ;
  assign n2646 = n2645 ^ n2638 ;
  assign n2679 = n2647 ^ n2646 ;
  assign n2680 = n2661 & ~n2679 ;
  assign n2681 = n2680 ^ n2660 ;
  assign n2693 = n2692 ^ n2681 ;
  assign n2674 = n2639 ^ n2638 ;
  assign n2675 = n2645 & ~n2674 ;
  assign n2676 = n2675 ^ n2644 ;
  assign n2671 = n2641 ^ n2640 ;
  assign n2672 = n2643 & ~n2671 ;
  assign n2673 = n2672 ^ n2642 ;
  assign n2677 = n2676 ^ n2673 ;
  assign n2668 = n2635 ^ n2634 ;
  assign n2669 = n2637 & ~n2668 ;
  assign n2670 = n2669 ^ n2636 ;
  assign n2678 = n2677 ^ n2670 ;
  assign n2703 = n2692 ^ n2678 ;
  assign n2704 = n2693 & ~n2703 ;
  assign n2705 = n2704 ^ n2681 ;
  assign n2709 = n2708 ^ n2705 ;
  assign n2700 = n2673 ^ n2670 ;
  assign n2701 = n2677 & ~n2700 ;
  assign n2702 = n2701 ^ n2676 ;
  assign n2716 = n2705 ^ n2702 ;
  assign n2717 = n2709 & ~n2716 ;
  assign n2718 = n2717 ^ n2708 ;
  assign n2710 = n2709 ^ n2702 ;
  assign n2694 = n2693 ^ n2678 ;
  assign n2662 = n2661 ^ n2646 ;
  assign n2633 = x513 ^ x353 ;
  assign n2663 = n2662 ^ n2633 ;
  assign n2603 = x517 ^ x357 ;
  assign n2602 = x516 ^ x356 ;
  assign n2604 = n2603 ^ n2602 ;
  assign n2601 = x518 ^ x358 ;
  assign n2605 = n2604 ^ n2601 ;
  assign n2597 = x520 ^ x360 ;
  assign n2596 = x519 ^ x359 ;
  assign n2598 = n2597 ^ n2596 ;
  assign n2595 = x521 ^ x361 ;
  assign n2599 = n2598 ^ n2595 ;
  assign n2594 = x515 ^ x355 ;
  assign n2600 = n2599 ^ n2594 ;
  assign n2606 = n2605 ^ n2600 ;
  assign n2592 = x514 ^ x354 ;
  assign n2578 = x524 ^ x364 ;
  assign n2577 = x523 ^ x363 ;
  assign n2579 = n2578 ^ n2577 ;
  assign n2576 = x525 ^ x365 ;
  assign n2580 = n2579 ^ n2576 ;
  assign n2569 = x528 ^ x368 ;
  assign n2567 = x527 ^ x367 ;
  assign n2566 = x526 ^ x366 ;
  assign n2568 = n2567 ^ n2566 ;
  assign n2574 = n2569 ^ n2568 ;
  assign n2573 = x522 ^ x362 ;
  assign n2575 = n2574 ^ n2573 ;
  assign n2591 = n2580 ^ n2575 ;
  assign n2593 = n2592 ^ n2591 ;
  assign n2664 = n2606 ^ n2593 ;
  assign n2665 = n2664 ^ n2633 ;
  assign n2666 = n2663 & ~n2665 ;
  assign n2667 = n2666 ^ n2662 ;
  assign n2695 = n2694 ^ n2667 ;
  assign n2618 = n2596 ^ n2595 ;
  assign n2619 = n2598 & ~n2618 ;
  assign n2620 = n2619 ^ n2597 ;
  assign n2615 = n2605 ^ n2599 ;
  assign n2616 = ~n2600 & n2615 ;
  assign n2617 = n2616 ^ n2605 ;
  assign n2621 = n2620 ^ n2617 ;
  assign n2612 = n2602 ^ n2601 ;
  assign n2613 = n2604 & ~n2612 ;
  assign n2614 = n2613 ^ n2603 ;
  assign n2622 = n2621 ^ n2614 ;
  assign n2585 = n2577 ^ n2576 ;
  assign n2586 = n2579 & ~n2585 ;
  assign n2587 = n2586 ^ n2578 ;
  assign n2581 = n2580 ^ n2573 ;
  assign n2582 = n2575 & ~n2581 ;
  assign n2583 = n2582 ^ n2574 ;
  assign n2570 = n2569 ^ n2566 ;
  assign n2571 = n2568 & ~n2570 ;
  assign n2572 = n2571 ^ n2567 ;
  assign n2584 = n2583 ^ n2572 ;
  assign n2610 = n2587 ^ n2584 ;
  assign n2607 = n2606 ^ n2591 ;
  assign n2608 = n2593 & ~n2607 ;
  assign n2609 = n2608 ^ n2592 ;
  assign n2611 = n2610 ^ n2609 ;
  assign n2696 = n2622 ^ n2611 ;
  assign n2697 = n2696 ^ n2694 ;
  assign n2698 = n2695 & ~n2697 ;
  assign n2699 = n2698 ^ n2667 ;
  assign n2711 = n2710 ^ n2699 ;
  assign n2627 = n2617 ^ n2614 ;
  assign n2628 = n2621 & ~n2627 ;
  assign n2629 = n2628 ^ n2620 ;
  assign n2623 = n2622 ^ n2610 ;
  assign n2624 = n2611 & ~n2623 ;
  assign n2625 = n2624 ^ n2609 ;
  assign n2588 = n2587 ^ n2572 ;
  assign n2589 = n2584 & ~n2588 ;
  assign n2590 = n2589 ^ n2583 ;
  assign n2626 = n2625 ^ n2590 ;
  assign n2712 = n2629 ^ n2626 ;
  assign n2713 = n2712 ^ n2699 ;
  assign n2714 = n2711 & ~n2713 ;
  assign n2715 = n2714 ^ n2710 ;
  assign n2719 = n2718 ^ n2715 ;
  assign n2630 = n2629 ^ n2590 ;
  assign n2631 = n2626 & ~n2630 ;
  assign n2632 = n2631 ^ n2625 ;
  assign n2720 = n2719 ^ n2632 ;
  assign n2721 = n2696 ^ n2695 ;
  assign n2722 = n2664 ^ n2663 ;
  assign n2723 = x512 ^ x352 ;
  assign n2724 = n2722 & n2723 ;
  assign n2725 = n2721 & n2724 ;
  assign n2726 = n2712 ^ n2711 ;
  assign n2727 = n2725 & n2726 ;
  assign n2728 = n2720 & n2727 ;
  assign n2729 = n2718 ^ n2632 ;
  assign n2730 = ~n2719 & n2729 ;
  assign n2731 = n2730 ^ n2632 ;
  assign n2732 = n2728 & n2731 ;
  assign n1970 = x541 ^ x413 ;
  assign n1969 = x542 ^ x414 ;
  assign n1971 = n1970 ^ n1969 ;
  assign n1968 = x543 ^ x415 ;
  assign n2003 = n1969 ^ n1968 ;
  assign n2004 = n1971 & ~n2003 ;
  assign n2005 = n2004 ^ n1970 ;
  assign n1973 = x537 ^ x409 ;
  assign n1972 = n1971 ^ n1968 ;
  assign n1974 = n1973 ^ n1972 ;
  assign n1965 = x539 ^ x411 ;
  assign n1964 = x538 ^ x410 ;
  assign n1966 = n1965 ^ n1964 ;
  assign n1963 = x540 ^ x412 ;
  assign n1967 = n1966 ^ n1963 ;
  assign n2000 = n1972 ^ n1967 ;
  assign n2001 = n1974 & ~n2000 ;
  assign n2002 = n2001 ^ n1973 ;
  assign n2006 = n2005 ^ n2002 ;
  assign n1997 = n1964 ^ n1963 ;
  assign n1998 = n1966 & ~n1997 ;
  assign n1999 = n1998 ^ n1965 ;
  assign n2021 = n2002 ^ n1999 ;
  assign n2022 = n2006 & ~n2021 ;
  assign n2023 = n2022 ^ n2005 ;
  assign n2007 = n2006 ^ n1999 ;
  assign n1975 = n1974 ^ n1967 ;
  assign n1962 = x529 ^ x401 ;
  assign n1976 = n1975 ^ n1962 ;
  assign n1957 = x535 ^ x407 ;
  assign n1956 = x534 ^ x406 ;
  assign n1958 = n1957 ^ n1956 ;
  assign n1955 = x536 ^ x408 ;
  assign n1959 = n1958 ^ n1955 ;
  assign n1954 = x530 ^ x402 ;
  assign n1960 = n1959 ^ n1954 ;
  assign n1951 = x532 ^ x404 ;
  assign n1950 = x531 ^ x403 ;
  assign n1952 = n1951 ^ n1950 ;
  assign n1949 = x533 ^ x405 ;
  assign n1953 = n1952 ^ n1949 ;
  assign n1961 = n1960 ^ n1953 ;
  assign n1994 = n1962 ^ n1961 ;
  assign n1995 = n1976 & ~n1994 ;
  assign n1996 = n1995 ^ n1975 ;
  assign n2008 = n2007 ^ n1996 ;
  assign n1989 = n1954 ^ n1953 ;
  assign n1990 = n1960 & ~n1989 ;
  assign n1991 = n1990 ^ n1959 ;
  assign n1986 = n1956 ^ n1955 ;
  assign n1987 = n1958 & ~n1986 ;
  assign n1988 = n1987 ^ n1957 ;
  assign n1992 = n1991 ^ n1988 ;
  assign n1983 = n1950 ^ n1949 ;
  assign n1984 = n1952 & ~n1983 ;
  assign n1985 = n1984 ^ n1951 ;
  assign n1993 = n1992 ^ n1985 ;
  assign n2018 = n2007 ^ n1993 ;
  assign n2019 = n2008 & ~n2018 ;
  assign n2020 = n2019 ^ n1996 ;
  assign n2024 = n2023 ^ n2020 ;
  assign n2015 = n1988 ^ n1985 ;
  assign n2016 = n1992 & ~n2015 ;
  assign n2017 = n2016 ^ n1991 ;
  assign n2031 = n2020 ^ n2017 ;
  assign n2032 = n2024 & ~n2031 ;
  assign n2033 = n2032 ^ n2023 ;
  assign n2025 = n2024 ^ n2017 ;
  assign n2009 = n2008 ^ n1993 ;
  assign n1977 = n1976 ^ n1961 ;
  assign n1948 = x513 ^ x385 ;
  assign n1978 = n1977 ^ n1948 ;
  assign n1918 = x517 ^ x389 ;
  assign n1917 = x516 ^ x388 ;
  assign n1919 = n1918 ^ n1917 ;
  assign n1916 = x518 ^ x390 ;
  assign n1920 = n1919 ^ n1916 ;
  assign n1912 = x520 ^ x392 ;
  assign n1911 = x519 ^ x391 ;
  assign n1913 = n1912 ^ n1911 ;
  assign n1910 = x521 ^ x393 ;
  assign n1914 = n1913 ^ n1910 ;
  assign n1909 = x515 ^ x387 ;
  assign n1915 = n1914 ^ n1909 ;
  assign n1921 = n1920 ^ n1915 ;
  assign n1907 = x514 ^ x386 ;
  assign n1893 = x524 ^ x396 ;
  assign n1892 = x523 ^ x395 ;
  assign n1894 = n1893 ^ n1892 ;
  assign n1891 = x525 ^ x397 ;
  assign n1895 = n1894 ^ n1891 ;
  assign n1884 = x528 ^ x400 ;
  assign n1882 = x527 ^ x399 ;
  assign n1881 = x526 ^ x398 ;
  assign n1883 = n1882 ^ n1881 ;
  assign n1889 = n1884 ^ n1883 ;
  assign n1888 = x522 ^ x394 ;
  assign n1890 = n1889 ^ n1888 ;
  assign n1906 = n1895 ^ n1890 ;
  assign n1908 = n1907 ^ n1906 ;
  assign n1979 = n1921 ^ n1908 ;
  assign n1980 = n1979 ^ n1948 ;
  assign n1981 = n1978 & ~n1980 ;
  assign n1982 = n1981 ^ n1977 ;
  assign n2010 = n2009 ^ n1982 ;
  assign n1933 = n1911 ^ n1910 ;
  assign n1934 = n1913 & ~n1933 ;
  assign n1935 = n1934 ^ n1912 ;
  assign n1930 = n1920 ^ n1914 ;
  assign n1931 = ~n1915 & n1930 ;
  assign n1932 = n1931 ^ n1920 ;
  assign n1936 = n1935 ^ n1932 ;
  assign n1927 = n1917 ^ n1916 ;
  assign n1928 = n1919 & ~n1927 ;
  assign n1929 = n1928 ^ n1918 ;
  assign n1937 = n1936 ^ n1929 ;
  assign n1900 = n1892 ^ n1891 ;
  assign n1901 = n1894 & ~n1900 ;
  assign n1902 = n1901 ^ n1893 ;
  assign n1896 = n1895 ^ n1888 ;
  assign n1897 = n1890 & ~n1896 ;
  assign n1898 = n1897 ^ n1889 ;
  assign n1885 = n1884 ^ n1881 ;
  assign n1886 = n1883 & ~n1885 ;
  assign n1887 = n1886 ^ n1882 ;
  assign n1899 = n1898 ^ n1887 ;
  assign n1925 = n1902 ^ n1899 ;
  assign n1922 = n1921 ^ n1906 ;
  assign n1923 = n1908 & ~n1922 ;
  assign n1924 = n1923 ^ n1907 ;
  assign n1926 = n1925 ^ n1924 ;
  assign n2011 = n1937 ^ n1926 ;
  assign n2012 = n2011 ^ n2009 ;
  assign n2013 = n2010 & ~n2012 ;
  assign n2014 = n2013 ^ n1982 ;
  assign n2026 = n2025 ^ n2014 ;
  assign n1942 = n1932 ^ n1929 ;
  assign n1943 = n1936 & ~n1942 ;
  assign n1944 = n1943 ^ n1935 ;
  assign n1938 = n1937 ^ n1925 ;
  assign n1939 = n1926 & ~n1938 ;
  assign n1940 = n1939 ^ n1924 ;
  assign n1903 = n1902 ^ n1887 ;
  assign n1904 = n1899 & ~n1903 ;
  assign n1905 = n1904 ^ n1898 ;
  assign n1941 = n1940 ^ n1905 ;
  assign n2027 = n1944 ^ n1941 ;
  assign n2028 = n2027 ^ n2014 ;
  assign n2029 = n2026 & ~n2028 ;
  assign n2030 = n2029 ^ n2025 ;
  assign n2034 = n2033 ^ n2030 ;
  assign n1945 = n1944 ^ n1905 ;
  assign n1946 = n1941 & ~n1945 ;
  assign n1947 = n1946 ^ n1940 ;
  assign n2035 = n2034 ^ n1947 ;
  assign n2036 = n2011 ^ n2010 ;
  assign n2037 = n1979 ^ n1978 ;
  assign n2038 = x512 ^ x384 ;
  assign n2039 = n2037 & n2038 ;
  assign n2040 = n2036 & n2039 ;
  assign n2041 = n2027 ^ n2026 ;
  assign n2042 = n2040 & n2041 ;
  assign n2043 = n2035 & n2042 ;
  assign n2044 = n2033 ^ n1947 ;
  assign n2045 = ~n2034 & n2044 ;
  assign n2046 = n2045 ^ n1947 ;
  assign n2047 = n2043 & n2046 ;
  assign n2122 = x532 ^ x500 ;
  assign n2121 = x531 ^ x499 ;
  assign n2123 = n2122 ^ n2121 ;
  assign n2120 = x533 ^ x501 ;
  assign n2132 = n2121 ^ n2120 ;
  assign n2133 = n2123 & ~n2132 ;
  assign n2134 = n2133 ^ n2122 ;
  assign n2116 = x535 ^ x503 ;
  assign n2115 = x534 ^ x502 ;
  assign n2117 = n2116 ^ n2115 ;
  assign n2114 = x536 ^ x504 ;
  assign n2128 = n2115 ^ n2114 ;
  assign n2129 = n2117 & ~n2128 ;
  assign n2130 = n2129 ^ n2116 ;
  assign n2118 = n2117 ^ n2114 ;
  assign n2113 = x530 ^ x498 ;
  assign n2119 = n2118 ^ n2113 ;
  assign n2124 = n2123 ^ n2120 ;
  assign n2125 = n2124 ^ n2113 ;
  assign n2126 = n2119 & ~n2125 ;
  assign n2127 = n2126 ^ n2118 ;
  assign n2131 = n2130 ^ n2127 ;
  assign n2172 = n2134 ^ n2131 ;
  assign n2150 = x539 ^ x507 ;
  assign n2149 = x538 ^ x506 ;
  assign n2151 = n2150 ^ n2149 ;
  assign n2148 = x540 ^ x508 ;
  assign n2157 = n2149 ^ n2148 ;
  assign n2158 = n2151 & ~n2157 ;
  assign n2159 = n2158 ^ n2150 ;
  assign n2146 = x537 ^ x505 ;
  assign n2141 = x543 ^ x511 ;
  assign n2139 = x542 ^ x510 ;
  assign n2138 = x541 ^ x509 ;
  assign n2140 = n2139 ^ n2138 ;
  assign n2145 = n2141 ^ n2140 ;
  assign n2147 = n2146 ^ n2145 ;
  assign n2152 = n2151 ^ n2148 ;
  assign n2153 = n2152 ^ n2145 ;
  assign n2154 = n2147 & ~n2153 ;
  assign n2155 = n2154 ^ n2146 ;
  assign n2142 = n2141 ^ n2139 ;
  assign n2143 = ~n2140 & n2142 ;
  assign n2144 = n2143 ^ n2141 ;
  assign n2156 = n2155 ^ n2144 ;
  assign n2170 = n2159 ^ n2156 ;
  assign n2164 = n2152 ^ n2147 ;
  assign n2163 = x529 ^ x497 ;
  assign n2165 = n2164 ^ n2163 ;
  assign n2166 = n2124 ^ n2119 ;
  assign n2167 = n2166 ^ n2163 ;
  assign n2168 = n2165 & ~n2167 ;
  assign n2169 = n2168 ^ n2164 ;
  assign n2171 = n2170 ^ n2169 ;
  assign n2185 = n2172 ^ n2171 ;
  assign n2179 = x513 ^ x481 ;
  assign n2178 = n2166 ^ n2165 ;
  assign n2180 = n2179 ^ n2178 ;
  assign n2057 = x517 ^ x485 ;
  assign n2056 = x516 ^ x484 ;
  assign n2058 = n2057 ^ n2056 ;
  assign n2055 = x518 ^ x486 ;
  assign n2059 = n2058 ^ n2055 ;
  assign n2051 = x520 ^ x488 ;
  assign n2050 = x519 ^ x487 ;
  assign n2052 = n2051 ^ n2050 ;
  assign n2049 = x521 ^ x489 ;
  assign n2053 = n2052 ^ n2049 ;
  assign n2048 = x515 ^ x483 ;
  assign n2054 = n2053 ^ n2048 ;
  assign n2104 = n2059 ^ n2054 ;
  assign n2102 = x514 ^ x482 ;
  assign n2085 = x524 ^ x492 ;
  assign n2084 = x523 ^ x491 ;
  assign n2086 = n2085 ^ n2084 ;
  assign n2083 = x525 ^ x493 ;
  assign n2087 = n2086 ^ n2083 ;
  assign n2081 = x522 ^ x490 ;
  assign n2076 = x528 ^ x496 ;
  assign n2074 = x527 ^ x495 ;
  assign n2073 = x526 ^ x494 ;
  assign n2075 = n2074 ^ n2073 ;
  assign n2080 = n2076 ^ n2075 ;
  assign n2082 = n2081 ^ n2080 ;
  assign n2101 = n2087 ^ n2082 ;
  assign n2103 = n2102 ^ n2101 ;
  assign n2181 = n2104 ^ n2103 ;
  assign n2182 = n2181 ^ n2178 ;
  assign n2183 = n2180 & ~n2182 ;
  assign n2184 = n2183 ^ n2179 ;
  assign n2186 = n2185 ^ n2184 ;
  assign n2105 = n2104 ^ n2102 ;
  assign n2106 = ~n2103 & n2105 ;
  assign n2107 = n2106 ^ n2104 ;
  assign n2092 = n2084 ^ n2083 ;
  assign n2093 = n2086 & ~n2092 ;
  assign n2094 = n2093 ^ n2085 ;
  assign n2088 = n2087 ^ n2080 ;
  assign n2089 = n2082 & ~n2088 ;
  assign n2090 = n2089 ^ n2081 ;
  assign n2077 = n2076 ^ n2074 ;
  assign n2078 = ~n2075 & n2077 ;
  assign n2079 = n2078 ^ n2076 ;
  assign n2091 = n2090 ^ n2079 ;
  assign n2099 = n2094 ^ n2091 ;
  assign n2067 = n2056 ^ n2055 ;
  assign n2068 = n2058 & ~n2067 ;
  assign n2069 = n2068 ^ n2057 ;
  assign n2063 = n2050 ^ n2049 ;
  assign n2064 = n2052 & ~n2063 ;
  assign n2065 = n2064 ^ n2051 ;
  assign n2060 = n2059 ^ n2048 ;
  assign n2061 = n2054 & ~n2060 ;
  assign n2062 = n2061 ^ n2053 ;
  assign n2066 = n2065 ^ n2062 ;
  assign n2098 = n2069 ^ n2066 ;
  assign n2100 = n2099 ^ n2098 ;
  assign n2187 = n2107 ^ n2100 ;
  assign n2188 = n2187 ^ n2185 ;
  assign n2189 = n2186 & ~n2188 ;
  assign n2190 = n2189 ^ n2184 ;
  assign n2173 = n2172 ^ n2170 ;
  assign n2174 = n2171 & ~n2173 ;
  assign n2175 = n2174 ^ n2169 ;
  assign n2160 = n2159 ^ n2155 ;
  assign n2161 = ~n2156 & n2160 ;
  assign n2162 = n2161 ^ n2159 ;
  assign n2176 = n2175 ^ n2162 ;
  assign n2135 = n2134 ^ n2127 ;
  assign n2136 = ~n2131 & n2135 ;
  assign n2137 = n2136 ^ n2134 ;
  assign n2177 = n2176 ^ n2137 ;
  assign n2191 = n2190 ^ n2177 ;
  assign n2108 = n2107 ^ n2098 ;
  assign n2109 = n2100 & ~n2108 ;
  assign n2110 = n2109 ^ n2099 ;
  assign n2095 = n2094 ^ n2090 ;
  assign n2096 = ~n2091 & n2095 ;
  assign n2097 = n2096 ^ n2094 ;
  assign n2111 = n2110 ^ n2097 ;
  assign n2070 = n2069 ^ n2062 ;
  assign n2071 = ~n2066 & n2070 ;
  assign n2072 = n2071 ^ n2069 ;
  assign n2112 = n2111 ^ n2072 ;
  assign n2192 = n2191 ^ n2112 ;
  assign n2193 = n2187 ^ n2186 ;
  assign n2194 = x512 ^ x480 ;
  assign n2195 = n2181 ^ n2180 ;
  assign n2196 = n2194 & n2195 ;
  assign n2197 = n2193 & n2196 ;
  assign n2198 = n2192 & n2197 ;
  assign n2205 = n2177 ^ n2112 ;
  assign n2206 = n2191 & ~n2205 ;
  assign n2207 = n2206 ^ n2190 ;
  assign n2202 = n2162 ^ n2137 ;
  assign n2203 = n2176 & ~n2202 ;
  assign n2204 = n2203 ^ n2175 ;
  assign n2208 = n2207 ^ n2204 ;
  assign n2199 = n2097 ^ n2072 ;
  assign n2200 = n2111 & ~n2199 ;
  assign n2201 = n2200 ^ n2110 ;
  assign n2209 = n2208 ^ n2201 ;
  assign n2210 = n2198 & n2209 ;
  assign n2211 = n2204 ^ n2201 ;
  assign n2212 = n2208 & ~n2211 ;
  assign n2213 = n2212 ^ n2207 ;
  assign n2214 = n2210 & n2213 ;
  assign n2237 = x541 ^ x477 ;
  assign n2236 = x542 ^ x478 ;
  assign n2238 = n2237 ^ n2236 ;
  assign n2235 = x543 ^ x479 ;
  assign n2298 = n2236 ^ n2235 ;
  assign n2299 = n2238 & ~n2298 ;
  assign n2300 = n2299 ^ n2237 ;
  assign n2239 = n2238 ^ n2235 ;
  assign n2234 = x537 ^ x473 ;
  assign n2240 = n2239 ^ n2234 ;
  assign n2231 = x539 ^ x475 ;
  assign n2230 = x538 ^ x474 ;
  assign n2232 = n2231 ^ n2230 ;
  assign n2229 = x540 ^ x476 ;
  assign n2233 = n2232 ^ n2229 ;
  assign n2295 = n2234 ^ n2233 ;
  assign n2296 = n2240 & ~n2295 ;
  assign n2297 = n2296 ^ n2239 ;
  assign n2301 = n2300 ^ n2297 ;
  assign n2292 = n2230 ^ n2229 ;
  assign n2293 = n2232 & ~n2292 ;
  assign n2294 = n2293 ^ n2231 ;
  assign n2342 = n2297 ^ n2294 ;
  assign n2343 = n2301 & ~n2342 ;
  assign n2344 = n2343 ^ n2300 ;
  assign n2302 = n2301 ^ n2294 ;
  assign n2241 = n2240 ^ n2233 ;
  assign n2228 = x529 ^ x465 ;
  assign n2242 = n2241 ^ n2228 ;
  assign n2225 = x533 ^ x469 ;
  assign n2223 = x531 ^ x467 ;
  assign n2222 = x532 ^ x468 ;
  assign n2224 = n2223 ^ n2222 ;
  assign n2226 = n2225 ^ n2224 ;
  assign n2220 = x530 ^ x466 ;
  assign n2218 = x536 ^ x472 ;
  assign n2216 = x534 ^ x470 ;
  assign n2215 = x535 ^ x471 ;
  assign n2217 = n2216 ^ n2215 ;
  assign n2219 = n2218 ^ n2217 ;
  assign n2221 = n2220 ^ n2219 ;
  assign n2227 = n2226 ^ n2221 ;
  assign n2289 = n2228 ^ n2227 ;
  assign n2290 = n2242 & ~n2289 ;
  assign n2291 = n2290 ^ n2241 ;
  assign n2303 = n2302 ^ n2291 ;
  assign n2284 = n2218 ^ n2215 ;
  assign n2285 = n2217 & ~n2284 ;
  assign n2286 = n2285 ^ n2216 ;
  assign n2281 = n2226 ^ n2219 ;
  assign n2282 = n2221 & ~n2281 ;
  assign n2283 = n2282 ^ n2220 ;
  assign n2287 = n2286 ^ n2283 ;
  assign n2278 = n2225 ^ n2222 ;
  assign n2279 = n2224 & ~n2278 ;
  assign n2280 = n2279 ^ n2223 ;
  assign n2288 = n2287 ^ n2280 ;
  assign n2339 = n2302 ^ n2288 ;
  assign n2340 = ~n2303 & n2339 ;
  assign n2341 = n2340 ^ n2288 ;
  assign n2345 = n2344 ^ n2341 ;
  assign n2336 = n2283 ^ n2280 ;
  assign n2337 = ~n2287 & n2336 ;
  assign n2338 = n2337 ^ n2280 ;
  assign n2369 = n2341 ^ n2338 ;
  assign n2370 = n2345 & ~n2369 ;
  assign n2371 = n2370 ^ n2344 ;
  assign n2346 = n2345 ^ n2338 ;
  assign n2304 = n2303 ^ n2288 ;
  assign n2244 = x513 ^ x449 ;
  assign n2243 = n2242 ^ n2227 ;
  assign n2245 = n2244 ^ n2243 ;
  assign n2270 = x522 ^ x458 ;
  assign n2268 = x528 ^ x464 ;
  assign n2266 = x527 ^ x463 ;
  assign n2265 = x526 ^ x462 ;
  assign n2267 = n2266 ^ n2265 ;
  assign n2269 = n2268 ^ n2267 ;
  assign n2271 = n2270 ^ n2269 ;
  assign n2262 = x524 ^ x460 ;
  assign n2261 = x523 ^ x459 ;
  assign n2263 = n2262 ^ n2261 ;
  assign n2260 = x525 ^ x461 ;
  assign n2264 = n2263 ^ n2260 ;
  assign n2272 = n2271 ^ n2264 ;
  assign n2259 = x514 ^ x450 ;
  assign n2273 = n2272 ^ n2259 ;
  assign n2254 = x520 ^ x456 ;
  assign n2253 = x519 ^ x455 ;
  assign n2255 = n2254 ^ n2253 ;
  assign n2252 = x521 ^ x457 ;
  assign n2256 = n2255 ^ n2252 ;
  assign n2251 = x515 ^ x451 ;
  assign n2257 = n2256 ^ n2251 ;
  assign n2248 = x517 ^ x453 ;
  assign n2247 = x516 ^ x452 ;
  assign n2249 = n2248 ^ n2247 ;
  assign n2246 = x518 ^ x454 ;
  assign n2250 = n2249 ^ n2246 ;
  assign n2258 = n2257 ^ n2250 ;
  assign n2274 = n2273 ^ n2258 ;
  assign n2275 = n2274 ^ n2243 ;
  assign n2276 = n2245 & ~n2275 ;
  assign n2277 = n2276 ^ n2244 ;
  assign n2305 = n2304 ^ n2277 ;
  assign n2326 = n2269 ^ n2264 ;
  assign n2327 = n2271 & ~n2326 ;
  assign n2328 = n2327 ^ n2270 ;
  assign n2323 = n2268 ^ n2266 ;
  assign n2324 = ~n2267 & n2323 ;
  assign n2325 = n2324 ^ n2268 ;
  assign n2329 = n2328 ^ n2325 ;
  assign n2320 = n2261 ^ n2260 ;
  assign n2321 = n2263 & ~n2320 ;
  assign n2322 = n2321 ^ n2262 ;
  assign n2330 = n2329 ^ n2322 ;
  assign n2315 = n2253 ^ n2252 ;
  assign n2316 = n2255 & ~n2315 ;
  assign n2317 = n2316 ^ n2254 ;
  assign n2312 = n2251 ^ n2250 ;
  assign n2313 = n2257 & ~n2312 ;
  assign n2314 = n2313 ^ n2256 ;
  assign n2318 = n2317 ^ n2314 ;
  assign n2309 = n2247 ^ n2246 ;
  assign n2310 = n2249 & ~n2309 ;
  assign n2311 = n2310 ^ n2248 ;
  assign n2319 = n2318 ^ n2311 ;
  assign n2331 = n2330 ^ n2319 ;
  assign n2306 = n2259 ^ n2258 ;
  assign n2307 = n2273 & ~n2306 ;
  assign n2308 = n2307 ^ n2272 ;
  assign n2332 = n2331 ^ n2308 ;
  assign n2333 = n2332 ^ n2304 ;
  assign n2334 = n2305 & ~n2333 ;
  assign n2335 = n2334 ^ n2277 ;
  assign n2347 = n2346 ^ n2335 ;
  assign n2354 = n2330 ^ n2308 ;
  assign n2355 = ~n2331 & n2354 ;
  assign n2356 = n2355 ^ n2308 ;
  assign n2351 = n2328 ^ n2322 ;
  assign n2352 = ~n2329 & n2351 ;
  assign n2353 = n2352 ^ n2322 ;
  assign n2357 = n2356 ^ n2353 ;
  assign n2348 = n2314 ^ n2311 ;
  assign n2349 = ~n2318 & n2348 ;
  assign n2350 = n2349 ^ n2311 ;
  assign n2358 = n2357 ^ n2350 ;
  assign n2366 = n2358 ^ n2346 ;
  assign n2367 = ~n2347 & n2366 ;
  assign n2368 = n2367 ^ n2358 ;
  assign n2372 = n2371 ^ n2368 ;
  assign n2373 = n2353 ^ n2350 ;
  assign n2374 = n2357 & ~n2373 ;
  assign n2375 = n2374 ^ n2356 ;
  assign n2378 = n2375 ^ n2368 ;
  assign n2379 = n2372 & ~n2378 ;
  assign n2380 = n2379 ^ n2371 ;
  assign n2359 = n2358 ^ n2347 ;
  assign n2360 = n2332 ^ n2305 ;
  assign n2361 = x512 ^ x448 ;
  assign n2362 = n2274 ^ n2245 ;
  assign n2363 = n2361 & n2362 ;
  assign n2364 = n2360 & n2363 ;
  assign n2365 = n2359 & n2364 ;
  assign n2376 = n2375 ^ n2372 ;
  assign n2377 = n2365 & n2376 ;
  assign n2382 = n2380 ^ n2377 ;
  assign n2381 = ~n2377 & ~n2380 ;
  assign n2383 = n2382 ^ n2381 ;
  assign n2384 = ~n2214 & ~n2383 ;
  assign n2385 = n2384 ^ n2214 ;
  assign n2555 = n2385 ^ n2383 ;
  assign n2556 = n2555 ^ n2214 ;
  assign n2475 = x541 ^ x445 ;
  assign n2474 = x542 ^ x446 ;
  assign n2476 = n2475 ^ n2474 ;
  assign n2473 = x543 ^ x447 ;
  assign n2508 = n2474 ^ n2473 ;
  assign n2509 = n2476 & ~n2508 ;
  assign n2510 = n2509 ^ n2475 ;
  assign n2478 = x537 ^ x441 ;
  assign n2477 = n2476 ^ n2473 ;
  assign n2479 = n2478 ^ n2477 ;
  assign n2470 = x539 ^ x443 ;
  assign n2469 = x538 ^ x442 ;
  assign n2471 = n2470 ^ n2469 ;
  assign n2468 = x540 ^ x444 ;
  assign n2472 = n2471 ^ n2468 ;
  assign n2505 = n2477 ^ n2472 ;
  assign n2506 = n2479 & ~n2505 ;
  assign n2507 = n2506 ^ n2478 ;
  assign n2511 = n2510 ^ n2507 ;
  assign n2502 = n2469 ^ n2468 ;
  assign n2503 = n2471 & ~n2502 ;
  assign n2504 = n2503 ^ n2470 ;
  assign n2526 = n2507 ^ n2504 ;
  assign n2527 = n2511 & ~n2526 ;
  assign n2528 = n2527 ^ n2510 ;
  assign n2512 = n2511 ^ n2504 ;
  assign n2480 = n2479 ^ n2472 ;
  assign n2467 = x529 ^ x433 ;
  assign n2481 = n2480 ^ n2467 ;
  assign n2462 = x535 ^ x439 ;
  assign n2461 = x534 ^ x438 ;
  assign n2463 = n2462 ^ n2461 ;
  assign n2460 = x536 ^ x440 ;
  assign n2464 = n2463 ^ n2460 ;
  assign n2459 = x530 ^ x434 ;
  assign n2465 = n2464 ^ n2459 ;
  assign n2456 = x532 ^ x436 ;
  assign n2455 = x531 ^ x435 ;
  assign n2457 = n2456 ^ n2455 ;
  assign n2454 = x533 ^ x437 ;
  assign n2458 = n2457 ^ n2454 ;
  assign n2466 = n2465 ^ n2458 ;
  assign n2499 = n2467 ^ n2466 ;
  assign n2500 = n2481 & ~n2499 ;
  assign n2501 = n2500 ^ n2480 ;
  assign n2513 = n2512 ^ n2501 ;
  assign n2494 = n2459 ^ n2458 ;
  assign n2495 = n2465 & ~n2494 ;
  assign n2496 = n2495 ^ n2464 ;
  assign n2491 = n2461 ^ n2460 ;
  assign n2492 = n2463 & ~n2491 ;
  assign n2493 = n2492 ^ n2462 ;
  assign n2497 = n2496 ^ n2493 ;
  assign n2488 = n2455 ^ n2454 ;
  assign n2489 = n2457 & ~n2488 ;
  assign n2490 = n2489 ^ n2456 ;
  assign n2498 = n2497 ^ n2490 ;
  assign n2523 = n2512 ^ n2498 ;
  assign n2524 = n2513 & ~n2523 ;
  assign n2525 = n2524 ^ n2501 ;
  assign n2529 = n2528 ^ n2525 ;
  assign n2520 = n2493 ^ n2490 ;
  assign n2521 = n2497 & ~n2520 ;
  assign n2522 = n2521 ^ n2496 ;
  assign n2536 = n2525 ^ n2522 ;
  assign n2537 = n2529 & ~n2536 ;
  assign n2538 = n2537 ^ n2528 ;
  assign n2530 = n2529 ^ n2522 ;
  assign n2514 = n2513 ^ n2498 ;
  assign n2482 = n2481 ^ n2466 ;
  assign n2453 = x513 ^ x417 ;
  assign n2483 = n2482 ^ n2453 ;
  assign n2423 = x517 ^ x421 ;
  assign n2422 = x516 ^ x420 ;
  assign n2424 = n2423 ^ n2422 ;
  assign n2421 = x518 ^ x422 ;
  assign n2425 = n2424 ^ n2421 ;
  assign n2417 = x520 ^ x424 ;
  assign n2416 = x519 ^ x423 ;
  assign n2418 = n2417 ^ n2416 ;
  assign n2415 = x521 ^ x425 ;
  assign n2419 = n2418 ^ n2415 ;
  assign n2414 = x515 ^ x419 ;
  assign n2420 = n2419 ^ n2414 ;
  assign n2426 = n2425 ^ n2420 ;
  assign n2412 = x514 ^ x418 ;
  assign n2398 = x524 ^ x428 ;
  assign n2397 = x523 ^ x427 ;
  assign n2399 = n2398 ^ n2397 ;
  assign n2396 = x525 ^ x429 ;
  assign n2400 = n2399 ^ n2396 ;
  assign n2389 = x528 ^ x432 ;
  assign n2387 = x527 ^ x431 ;
  assign n2386 = x526 ^ x430 ;
  assign n2388 = n2387 ^ n2386 ;
  assign n2394 = n2389 ^ n2388 ;
  assign n2393 = x522 ^ x426 ;
  assign n2395 = n2394 ^ n2393 ;
  assign n2411 = n2400 ^ n2395 ;
  assign n2413 = n2412 ^ n2411 ;
  assign n2484 = n2426 ^ n2413 ;
  assign n2485 = n2484 ^ n2453 ;
  assign n2486 = n2483 & ~n2485 ;
  assign n2487 = n2486 ^ n2482 ;
  assign n2515 = n2514 ^ n2487 ;
  assign n2438 = n2416 ^ n2415 ;
  assign n2439 = n2418 & ~n2438 ;
  assign n2440 = n2439 ^ n2417 ;
  assign n2435 = n2425 ^ n2419 ;
  assign n2436 = ~n2420 & n2435 ;
  assign n2437 = n2436 ^ n2425 ;
  assign n2441 = n2440 ^ n2437 ;
  assign n2432 = n2422 ^ n2421 ;
  assign n2433 = n2424 & ~n2432 ;
  assign n2434 = n2433 ^ n2423 ;
  assign n2442 = n2441 ^ n2434 ;
  assign n2405 = n2397 ^ n2396 ;
  assign n2406 = n2399 & ~n2405 ;
  assign n2407 = n2406 ^ n2398 ;
  assign n2401 = n2400 ^ n2393 ;
  assign n2402 = n2395 & ~n2401 ;
  assign n2403 = n2402 ^ n2394 ;
  assign n2390 = n2389 ^ n2386 ;
  assign n2391 = n2388 & ~n2390 ;
  assign n2392 = n2391 ^ n2387 ;
  assign n2404 = n2403 ^ n2392 ;
  assign n2430 = n2407 ^ n2404 ;
  assign n2427 = n2426 ^ n2411 ;
  assign n2428 = n2413 & ~n2427 ;
  assign n2429 = n2428 ^ n2412 ;
  assign n2431 = n2430 ^ n2429 ;
  assign n2516 = n2442 ^ n2431 ;
  assign n2517 = n2516 ^ n2514 ;
  assign n2518 = n2515 & ~n2517 ;
  assign n2519 = n2518 ^ n2487 ;
  assign n2531 = n2530 ^ n2519 ;
  assign n2447 = n2437 ^ n2434 ;
  assign n2448 = n2441 & ~n2447 ;
  assign n2449 = n2448 ^ n2440 ;
  assign n2443 = n2442 ^ n2430 ;
  assign n2444 = n2431 & ~n2443 ;
  assign n2445 = n2444 ^ n2429 ;
  assign n2408 = n2407 ^ n2392 ;
  assign n2409 = n2404 & ~n2408 ;
  assign n2410 = n2409 ^ n2403 ;
  assign n2446 = n2445 ^ n2410 ;
  assign n2532 = n2449 ^ n2446 ;
  assign n2533 = n2532 ^ n2519 ;
  assign n2534 = n2531 & ~n2533 ;
  assign n2535 = n2534 ^ n2530 ;
  assign n2539 = n2538 ^ n2535 ;
  assign n2450 = n2449 ^ n2410 ;
  assign n2451 = n2446 & ~n2450 ;
  assign n2452 = n2451 ^ n2445 ;
  assign n2540 = n2539 ^ n2452 ;
  assign n2541 = n2516 ^ n2515 ;
  assign n2542 = n2484 ^ n2483 ;
  assign n2543 = x512 ^ x416 ;
  assign n2544 = n2542 & n2543 ;
  assign n2545 = n2541 & n2544 ;
  assign n2546 = n2532 ^ n2531 ;
  assign n2547 = n2545 & n2546 ;
  assign n2548 = n2540 & n2547 ;
  assign n2549 = n2538 ^ n2452 ;
  assign n2550 = ~n2539 & n2549 ;
  assign n2551 = n2550 ^ n2452 ;
  assign n2552 = n2548 & n2551 ;
  assign n2553 = n2385 & ~n2552 ;
  assign n2554 = n2553 ^ n2385 ;
  assign n2558 = n2556 ^ n2554 ;
  assign n2557 = n2554 & n2556 ;
  assign n2559 = n2558 ^ n2557 ;
  assign n2560 = n2559 ^ n2554 ;
  assign n2561 = ~n2047 & ~n2560 ;
  assign n2562 = n2561 ^ n2560 ;
  assign n2563 = n2559 ^ n2556 ;
  assign n2564 = ~n2562 & ~n2563 ;
  assign n2565 = n2564 ^ n2562 ;
  assign n2733 = n2565 ^ n2563 ;
  assign n2734 = n2733 ^ n2562 ;
  assign n2735 = ~n2732 & n2734 ;
  assign n2736 = n2735 ^ n2734 ;
  assign n2740 = n2736 ^ n2565 ;
  assign n1803 = x541 ^ x349 ;
  assign n1802 = x542 ^ x350 ;
  assign n1804 = n1803 ^ n1802 ;
  assign n1801 = x543 ^ x351 ;
  assign n1836 = n1802 ^ n1801 ;
  assign n1837 = n1804 & ~n1836 ;
  assign n1838 = n1837 ^ n1803 ;
  assign n1806 = x537 ^ x345 ;
  assign n1805 = n1804 ^ n1801 ;
  assign n1807 = n1806 ^ n1805 ;
  assign n1798 = x539 ^ x347 ;
  assign n1797 = x538 ^ x346 ;
  assign n1799 = n1798 ^ n1797 ;
  assign n1796 = x540 ^ x348 ;
  assign n1800 = n1799 ^ n1796 ;
  assign n1833 = n1805 ^ n1800 ;
  assign n1834 = n1807 & ~n1833 ;
  assign n1835 = n1834 ^ n1806 ;
  assign n1839 = n1838 ^ n1835 ;
  assign n1830 = n1797 ^ n1796 ;
  assign n1831 = n1799 & ~n1830 ;
  assign n1832 = n1831 ^ n1798 ;
  assign n1854 = n1835 ^ n1832 ;
  assign n1855 = n1839 & ~n1854 ;
  assign n1856 = n1855 ^ n1838 ;
  assign n1840 = n1839 ^ n1832 ;
  assign n1808 = n1807 ^ n1800 ;
  assign n1795 = x529 ^ x337 ;
  assign n1809 = n1808 ^ n1795 ;
  assign n1790 = x535 ^ x343 ;
  assign n1789 = x534 ^ x342 ;
  assign n1791 = n1790 ^ n1789 ;
  assign n1788 = x536 ^ x344 ;
  assign n1792 = n1791 ^ n1788 ;
  assign n1787 = x530 ^ x338 ;
  assign n1793 = n1792 ^ n1787 ;
  assign n1784 = x532 ^ x340 ;
  assign n1783 = x531 ^ x339 ;
  assign n1785 = n1784 ^ n1783 ;
  assign n1782 = x533 ^ x341 ;
  assign n1786 = n1785 ^ n1782 ;
  assign n1794 = n1793 ^ n1786 ;
  assign n1827 = n1795 ^ n1794 ;
  assign n1828 = n1809 & ~n1827 ;
  assign n1829 = n1828 ^ n1808 ;
  assign n1841 = n1840 ^ n1829 ;
  assign n1822 = n1787 ^ n1786 ;
  assign n1823 = n1793 & ~n1822 ;
  assign n1824 = n1823 ^ n1792 ;
  assign n1819 = n1789 ^ n1788 ;
  assign n1820 = n1791 & ~n1819 ;
  assign n1821 = n1820 ^ n1790 ;
  assign n1825 = n1824 ^ n1821 ;
  assign n1816 = n1783 ^ n1782 ;
  assign n1817 = n1785 & ~n1816 ;
  assign n1818 = n1817 ^ n1784 ;
  assign n1826 = n1825 ^ n1818 ;
  assign n1851 = n1840 ^ n1826 ;
  assign n1852 = n1841 & ~n1851 ;
  assign n1853 = n1852 ^ n1829 ;
  assign n1857 = n1856 ^ n1853 ;
  assign n1848 = n1821 ^ n1818 ;
  assign n1849 = n1825 & ~n1848 ;
  assign n1850 = n1849 ^ n1824 ;
  assign n1864 = n1853 ^ n1850 ;
  assign n1865 = n1857 & ~n1864 ;
  assign n1866 = n1865 ^ n1856 ;
  assign n1858 = n1857 ^ n1850 ;
  assign n1842 = n1841 ^ n1826 ;
  assign n1810 = n1809 ^ n1794 ;
  assign n1781 = x513 ^ x321 ;
  assign n1811 = n1810 ^ n1781 ;
  assign n1751 = x517 ^ x325 ;
  assign n1750 = x516 ^ x324 ;
  assign n1752 = n1751 ^ n1750 ;
  assign n1749 = x518 ^ x326 ;
  assign n1753 = n1752 ^ n1749 ;
  assign n1745 = x520 ^ x328 ;
  assign n1744 = x519 ^ x327 ;
  assign n1746 = n1745 ^ n1744 ;
  assign n1743 = x521 ^ x329 ;
  assign n1747 = n1746 ^ n1743 ;
  assign n1742 = x515 ^ x323 ;
  assign n1748 = n1747 ^ n1742 ;
  assign n1754 = n1753 ^ n1748 ;
  assign n1740 = x514 ^ x322 ;
  assign n1726 = x524 ^ x332 ;
  assign n1725 = x523 ^ x331 ;
  assign n1727 = n1726 ^ n1725 ;
  assign n1724 = x525 ^ x333 ;
  assign n1728 = n1727 ^ n1724 ;
  assign n1717 = x528 ^ x336 ;
  assign n1715 = x527 ^ x335 ;
  assign n1714 = x526 ^ x334 ;
  assign n1716 = n1715 ^ n1714 ;
  assign n1722 = n1717 ^ n1716 ;
  assign n1721 = x522 ^ x330 ;
  assign n1723 = n1722 ^ n1721 ;
  assign n1739 = n1728 ^ n1723 ;
  assign n1741 = n1740 ^ n1739 ;
  assign n1812 = n1754 ^ n1741 ;
  assign n1813 = n1812 ^ n1781 ;
  assign n1814 = n1811 & ~n1813 ;
  assign n1815 = n1814 ^ n1810 ;
  assign n1843 = n1842 ^ n1815 ;
  assign n1766 = n1744 ^ n1743 ;
  assign n1767 = n1746 & ~n1766 ;
  assign n1768 = n1767 ^ n1745 ;
  assign n1763 = n1753 ^ n1747 ;
  assign n1764 = ~n1748 & n1763 ;
  assign n1765 = n1764 ^ n1753 ;
  assign n1769 = n1768 ^ n1765 ;
  assign n1760 = n1750 ^ n1749 ;
  assign n1761 = n1752 & ~n1760 ;
  assign n1762 = n1761 ^ n1751 ;
  assign n1770 = n1769 ^ n1762 ;
  assign n1733 = n1725 ^ n1724 ;
  assign n1734 = n1727 & ~n1733 ;
  assign n1735 = n1734 ^ n1726 ;
  assign n1729 = n1728 ^ n1721 ;
  assign n1730 = n1723 & ~n1729 ;
  assign n1731 = n1730 ^ n1722 ;
  assign n1718 = n1717 ^ n1714 ;
  assign n1719 = n1716 & ~n1718 ;
  assign n1720 = n1719 ^ n1715 ;
  assign n1732 = n1731 ^ n1720 ;
  assign n1758 = n1735 ^ n1732 ;
  assign n1755 = n1754 ^ n1739 ;
  assign n1756 = n1741 & ~n1755 ;
  assign n1757 = n1756 ^ n1740 ;
  assign n1759 = n1758 ^ n1757 ;
  assign n1844 = n1770 ^ n1759 ;
  assign n1845 = n1844 ^ n1842 ;
  assign n1846 = n1843 & ~n1845 ;
  assign n1847 = n1846 ^ n1815 ;
  assign n1859 = n1858 ^ n1847 ;
  assign n1775 = n1765 ^ n1762 ;
  assign n1776 = n1769 & ~n1775 ;
  assign n1777 = n1776 ^ n1768 ;
  assign n1771 = n1770 ^ n1758 ;
  assign n1772 = n1759 & ~n1771 ;
  assign n1773 = n1772 ^ n1757 ;
  assign n1736 = n1735 ^ n1720 ;
  assign n1737 = n1732 & ~n1736 ;
  assign n1738 = n1737 ^ n1731 ;
  assign n1774 = n1773 ^ n1738 ;
  assign n1860 = n1777 ^ n1774 ;
  assign n1861 = n1860 ^ n1847 ;
  assign n1862 = n1859 & ~n1861 ;
  assign n1863 = n1862 ^ n1858 ;
  assign n1867 = n1866 ^ n1863 ;
  assign n1778 = n1777 ^ n1738 ;
  assign n1779 = n1774 & ~n1778 ;
  assign n1780 = n1779 ^ n1773 ;
  assign n1868 = n1867 ^ n1780 ;
  assign n1869 = n1844 ^ n1843 ;
  assign n1870 = n1812 ^ n1811 ;
  assign n1871 = x512 ^ x320 ;
  assign n1872 = n1870 & n1871 ;
  assign n1873 = n1869 & n1872 ;
  assign n1874 = n1860 ^ n1859 ;
  assign n1875 = n1873 & n1874 ;
  assign n1876 = n1868 & n1875 ;
  assign n1877 = n1866 ^ n1780 ;
  assign n1878 = ~n1867 & n1877 ;
  assign n1879 = n1878 ^ n1780 ;
  assign n1880 = n1876 & n1879 ;
  assign n2737 = n2565 & ~n2736 ;
  assign n2738 = ~n1880 & ~n2737 ;
  assign n2743 = n2740 ^ n2738 ;
  assign n2739 = n2738 ^ n2737 ;
  assign n2741 = n2740 ^ n2737 ;
  assign n2742 = ~n2739 & ~n2741 ;
  assign n2744 = n2743 ^ n2742 ;
  assign n2745 = n2744 ^ n2739 ;
  assign n2746 = ~n1713 & n2745 ;
  assign n2747 = n2746 ^ n2745 ;
  assign n2748 = n2744 ^ n2741 ;
  assign n2749 = n2747 & n2748 ;
  assign n2750 = n2749 ^ n2747 ;
  assign n2918 = n2750 ^ n2748 ;
  assign n2919 = n2918 ^ n2747 ;
  assign n2920 = ~n2917 & ~n2919 ;
  assign n2921 = n2920 ^ n2919 ;
  assign n2925 = n2921 ^ n2750 ;
  assign n1469 = x541 ^ x253 ;
  assign n1468 = x542 ^ x254 ;
  assign n1470 = n1469 ^ n1468 ;
  assign n1467 = x543 ^ x255 ;
  assign n1502 = n1468 ^ n1467 ;
  assign n1503 = n1470 & ~n1502 ;
  assign n1504 = n1503 ^ n1469 ;
  assign n1472 = x537 ^ x249 ;
  assign n1471 = n1470 ^ n1467 ;
  assign n1473 = n1472 ^ n1471 ;
  assign n1464 = x539 ^ x251 ;
  assign n1463 = x538 ^ x250 ;
  assign n1465 = n1464 ^ n1463 ;
  assign n1462 = x540 ^ x252 ;
  assign n1466 = n1465 ^ n1462 ;
  assign n1499 = n1471 ^ n1466 ;
  assign n1500 = n1473 & ~n1499 ;
  assign n1501 = n1500 ^ n1472 ;
  assign n1505 = n1504 ^ n1501 ;
  assign n1496 = n1463 ^ n1462 ;
  assign n1497 = n1465 & ~n1496 ;
  assign n1498 = n1497 ^ n1464 ;
  assign n1520 = n1501 ^ n1498 ;
  assign n1521 = n1505 & ~n1520 ;
  assign n1522 = n1521 ^ n1504 ;
  assign n1506 = n1505 ^ n1498 ;
  assign n1474 = n1473 ^ n1466 ;
  assign n1461 = x529 ^ x241 ;
  assign n1475 = n1474 ^ n1461 ;
  assign n1456 = x535 ^ x247 ;
  assign n1455 = x534 ^ x246 ;
  assign n1457 = n1456 ^ n1455 ;
  assign n1454 = x536 ^ x248 ;
  assign n1458 = n1457 ^ n1454 ;
  assign n1453 = x530 ^ x242 ;
  assign n1459 = n1458 ^ n1453 ;
  assign n1450 = x532 ^ x244 ;
  assign n1449 = x531 ^ x243 ;
  assign n1451 = n1450 ^ n1449 ;
  assign n1448 = x533 ^ x245 ;
  assign n1452 = n1451 ^ n1448 ;
  assign n1460 = n1459 ^ n1452 ;
  assign n1493 = n1461 ^ n1460 ;
  assign n1494 = n1475 & ~n1493 ;
  assign n1495 = n1494 ^ n1474 ;
  assign n1507 = n1506 ^ n1495 ;
  assign n1488 = n1453 ^ n1452 ;
  assign n1489 = n1459 & ~n1488 ;
  assign n1490 = n1489 ^ n1458 ;
  assign n1485 = n1455 ^ n1454 ;
  assign n1486 = n1457 & ~n1485 ;
  assign n1487 = n1486 ^ n1456 ;
  assign n1491 = n1490 ^ n1487 ;
  assign n1482 = n1449 ^ n1448 ;
  assign n1483 = n1451 & ~n1482 ;
  assign n1484 = n1483 ^ n1450 ;
  assign n1492 = n1491 ^ n1484 ;
  assign n1517 = n1506 ^ n1492 ;
  assign n1518 = n1507 & ~n1517 ;
  assign n1519 = n1518 ^ n1495 ;
  assign n1523 = n1522 ^ n1519 ;
  assign n1514 = n1487 ^ n1484 ;
  assign n1515 = n1491 & ~n1514 ;
  assign n1516 = n1515 ^ n1490 ;
  assign n1530 = n1519 ^ n1516 ;
  assign n1531 = n1523 & ~n1530 ;
  assign n1532 = n1531 ^ n1522 ;
  assign n1524 = n1523 ^ n1516 ;
  assign n1508 = n1507 ^ n1492 ;
  assign n1476 = n1475 ^ n1460 ;
  assign n1447 = x513 ^ x225 ;
  assign n1477 = n1476 ^ n1447 ;
  assign n1417 = x517 ^ x229 ;
  assign n1416 = x516 ^ x228 ;
  assign n1418 = n1417 ^ n1416 ;
  assign n1415 = x518 ^ x230 ;
  assign n1419 = n1418 ^ n1415 ;
  assign n1411 = x520 ^ x232 ;
  assign n1410 = x519 ^ x231 ;
  assign n1412 = n1411 ^ n1410 ;
  assign n1409 = x521 ^ x233 ;
  assign n1413 = n1412 ^ n1409 ;
  assign n1408 = x515 ^ x227 ;
  assign n1414 = n1413 ^ n1408 ;
  assign n1420 = n1419 ^ n1414 ;
  assign n1406 = x514 ^ x226 ;
  assign n1392 = x524 ^ x236 ;
  assign n1391 = x523 ^ x235 ;
  assign n1393 = n1392 ^ n1391 ;
  assign n1390 = x525 ^ x237 ;
  assign n1394 = n1393 ^ n1390 ;
  assign n1383 = x528 ^ x240 ;
  assign n1381 = x527 ^ x239 ;
  assign n1380 = x526 ^ x238 ;
  assign n1382 = n1381 ^ n1380 ;
  assign n1388 = n1383 ^ n1382 ;
  assign n1387 = x522 ^ x234 ;
  assign n1389 = n1388 ^ n1387 ;
  assign n1405 = n1394 ^ n1389 ;
  assign n1407 = n1406 ^ n1405 ;
  assign n1478 = n1420 ^ n1407 ;
  assign n1479 = n1478 ^ n1447 ;
  assign n1480 = n1477 & ~n1479 ;
  assign n1481 = n1480 ^ n1476 ;
  assign n1509 = n1508 ^ n1481 ;
  assign n1432 = n1410 ^ n1409 ;
  assign n1433 = n1412 & ~n1432 ;
  assign n1434 = n1433 ^ n1411 ;
  assign n1429 = n1419 ^ n1413 ;
  assign n1430 = ~n1414 & n1429 ;
  assign n1431 = n1430 ^ n1419 ;
  assign n1435 = n1434 ^ n1431 ;
  assign n1426 = n1416 ^ n1415 ;
  assign n1427 = n1418 & ~n1426 ;
  assign n1428 = n1427 ^ n1417 ;
  assign n1436 = n1435 ^ n1428 ;
  assign n1399 = n1391 ^ n1390 ;
  assign n1400 = n1393 & ~n1399 ;
  assign n1401 = n1400 ^ n1392 ;
  assign n1395 = n1394 ^ n1387 ;
  assign n1396 = n1389 & ~n1395 ;
  assign n1397 = n1396 ^ n1388 ;
  assign n1384 = n1383 ^ n1380 ;
  assign n1385 = n1382 & ~n1384 ;
  assign n1386 = n1385 ^ n1381 ;
  assign n1398 = n1397 ^ n1386 ;
  assign n1424 = n1401 ^ n1398 ;
  assign n1421 = n1420 ^ n1405 ;
  assign n1422 = n1407 & ~n1421 ;
  assign n1423 = n1422 ^ n1406 ;
  assign n1425 = n1424 ^ n1423 ;
  assign n1510 = n1436 ^ n1425 ;
  assign n1511 = n1510 ^ n1508 ;
  assign n1512 = n1509 & ~n1511 ;
  assign n1513 = n1512 ^ n1481 ;
  assign n1525 = n1524 ^ n1513 ;
  assign n1441 = n1431 ^ n1428 ;
  assign n1442 = n1435 & ~n1441 ;
  assign n1443 = n1442 ^ n1434 ;
  assign n1437 = n1436 ^ n1424 ;
  assign n1438 = n1425 & ~n1437 ;
  assign n1439 = n1438 ^ n1423 ;
  assign n1402 = n1401 ^ n1386 ;
  assign n1403 = n1398 & ~n1402 ;
  assign n1404 = n1403 ^ n1397 ;
  assign n1440 = n1439 ^ n1404 ;
  assign n1526 = n1443 ^ n1440 ;
  assign n1527 = n1526 ^ n1513 ;
  assign n1528 = n1525 & ~n1527 ;
  assign n1529 = n1528 ^ n1524 ;
  assign n1533 = n1532 ^ n1529 ;
  assign n1444 = n1443 ^ n1404 ;
  assign n1445 = n1440 & ~n1444 ;
  assign n1446 = n1445 ^ n1439 ;
  assign n1534 = n1533 ^ n1446 ;
  assign n1535 = n1510 ^ n1509 ;
  assign n1536 = n1478 ^ n1477 ;
  assign n1537 = x512 ^ x224 ;
  assign n1538 = n1536 & n1537 ;
  assign n1539 = n1535 & n1538 ;
  assign n1540 = n1526 ^ n1525 ;
  assign n1541 = n1539 & n1540 ;
  assign n1542 = n1534 & n1541 ;
  assign n1543 = n1532 ^ n1446 ;
  assign n1544 = ~n1533 & n1543 ;
  assign n1545 = n1544 ^ n1446 ;
  assign n1546 = n1542 & n1545 ;
  assign n2922 = ~n2750 & n2921 ;
  assign n2923 = ~n1546 & ~n2922 ;
  assign n2928 = n2925 ^ n2923 ;
  assign n2924 = n2923 ^ n2922 ;
  assign n2926 = n2925 ^ n2922 ;
  assign n2927 = ~n2924 & ~n2926 ;
  assign n2929 = n2928 ^ n2927 ;
  assign n2930 = n2929 ^ n2924 ;
  assign n2931 = ~n1379 & n2930 ;
  assign n2932 = n2931 ^ n2930 ;
  assign n2933 = n2929 ^ n2926 ;
  assign n2934 = n2932 & n2933 ;
  assign n2935 = n2934 ^ n2932 ;
  assign n3103 = n2935 ^ n2933 ;
  assign n3104 = n3103 ^ n2932 ;
  assign n3105 = ~n3102 & ~n3104 ;
  assign n3106 = n3105 ^ n3104 ;
  assign n3110 = n3106 ^ n2935 ;
  assign n1135 = x541 ^ x157 ;
  assign n1134 = x542 ^ x158 ;
  assign n1136 = n1135 ^ n1134 ;
  assign n1133 = x543 ^ x159 ;
  assign n1168 = n1134 ^ n1133 ;
  assign n1169 = n1136 & ~n1168 ;
  assign n1170 = n1169 ^ n1135 ;
  assign n1138 = x537 ^ x153 ;
  assign n1137 = n1136 ^ n1133 ;
  assign n1139 = n1138 ^ n1137 ;
  assign n1130 = x539 ^ x155 ;
  assign n1129 = x538 ^ x154 ;
  assign n1131 = n1130 ^ n1129 ;
  assign n1128 = x540 ^ x156 ;
  assign n1132 = n1131 ^ n1128 ;
  assign n1165 = n1137 ^ n1132 ;
  assign n1166 = n1139 & ~n1165 ;
  assign n1167 = n1166 ^ n1138 ;
  assign n1171 = n1170 ^ n1167 ;
  assign n1162 = n1129 ^ n1128 ;
  assign n1163 = n1131 & ~n1162 ;
  assign n1164 = n1163 ^ n1130 ;
  assign n1186 = n1167 ^ n1164 ;
  assign n1187 = n1171 & ~n1186 ;
  assign n1188 = n1187 ^ n1170 ;
  assign n1172 = n1171 ^ n1164 ;
  assign n1140 = n1139 ^ n1132 ;
  assign n1127 = x529 ^ x145 ;
  assign n1141 = n1140 ^ n1127 ;
  assign n1122 = x535 ^ x151 ;
  assign n1121 = x534 ^ x150 ;
  assign n1123 = n1122 ^ n1121 ;
  assign n1120 = x536 ^ x152 ;
  assign n1124 = n1123 ^ n1120 ;
  assign n1119 = x530 ^ x146 ;
  assign n1125 = n1124 ^ n1119 ;
  assign n1116 = x532 ^ x148 ;
  assign n1115 = x531 ^ x147 ;
  assign n1117 = n1116 ^ n1115 ;
  assign n1114 = x533 ^ x149 ;
  assign n1118 = n1117 ^ n1114 ;
  assign n1126 = n1125 ^ n1118 ;
  assign n1159 = n1127 ^ n1126 ;
  assign n1160 = n1141 & ~n1159 ;
  assign n1161 = n1160 ^ n1140 ;
  assign n1173 = n1172 ^ n1161 ;
  assign n1154 = n1119 ^ n1118 ;
  assign n1155 = n1125 & ~n1154 ;
  assign n1156 = n1155 ^ n1124 ;
  assign n1151 = n1121 ^ n1120 ;
  assign n1152 = n1123 & ~n1151 ;
  assign n1153 = n1152 ^ n1122 ;
  assign n1157 = n1156 ^ n1153 ;
  assign n1148 = n1115 ^ n1114 ;
  assign n1149 = n1117 & ~n1148 ;
  assign n1150 = n1149 ^ n1116 ;
  assign n1158 = n1157 ^ n1150 ;
  assign n1183 = n1172 ^ n1158 ;
  assign n1184 = n1173 & ~n1183 ;
  assign n1185 = n1184 ^ n1161 ;
  assign n1189 = n1188 ^ n1185 ;
  assign n1180 = n1153 ^ n1150 ;
  assign n1181 = n1157 & ~n1180 ;
  assign n1182 = n1181 ^ n1156 ;
  assign n1196 = n1185 ^ n1182 ;
  assign n1197 = n1189 & ~n1196 ;
  assign n1198 = n1197 ^ n1188 ;
  assign n1190 = n1189 ^ n1182 ;
  assign n1174 = n1173 ^ n1158 ;
  assign n1142 = n1141 ^ n1126 ;
  assign n1113 = x513 ^ x129 ;
  assign n1143 = n1142 ^ n1113 ;
  assign n1083 = x517 ^ x133 ;
  assign n1082 = x516 ^ x132 ;
  assign n1084 = n1083 ^ n1082 ;
  assign n1081 = x518 ^ x134 ;
  assign n1085 = n1084 ^ n1081 ;
  assign n1077 = x520 ^ x136 ;
  assign n1076 = x519 ^ x135 ;
  assign n1078 = n1077 ^ n1076 ;
  assign n1075 = x521 ^ x137 ;
  assign n1079 = n1078 ^ n1075 ;
  assign n1074 = x515 ^ x131 ;
  assign n1080 = n1079 ^ n1074 ;
  assign n1086 = n1085 ^ n1080 ;
  assign n1072 = x514 ^ x130 ;
  assign n1058 = x524 ^ x140 ;
  assign n1057 = x523 ^ x139 ;
  assign n1059 = n1058 ^ n1057 ;
  assign n1056 = x525 ^ x141 ;
  assign n1060 = n1059 ^ n1056 ;
  assign n1049 = x528 ^ x144 ;
  assign n1047 = x527 ^ x143 ;
  assign n1046 = x526 ^ x142 ;
  assign n1048 = n1047 ^ n1046 ;
  assign n1054 = n1049 ^ n1048 ;
  assign n1053 = x522 ^ x138 ;
  assign n1055 = n1054 ^ n1053 ;
  assign n1071 = n1060 ^ n1055 ;
  assign n1073 = n1072 ^ n1071 ;
  assign n1144 = n1086 ^ n1073 ;
  assign n1145 = n1144 ^ n1113 ;
  assign n1146 = n1143 & ~n1145 ;
  assign n1147 = n1146 ^ n1142 ;
  assign n1175 = n1174 ^ n1147 ;
  assign n1098 = n1076 ^ n1075 ;
  assign n1099 = n1078 & ~n1098 ;
  assign n1100 = n1099 ^ n1077 ;
  assign n1095 = n1085 ^ n1079 ;
  assign n1096 = ~n1080 & n1095 ;
  assign n1097 = n1096 ^ n1085 ;
  assign n1101 = n1100 ^ n1097 ;
  assign n1092 = n1082 ^ n1081 ;
  assign n1093 = n1084 & ~n1092 ;
  assign n1094 = n1093 ^ n1083 ;
  assign n1102 = n1101 ^ n1094 ;
  assign n1065 = n1057 ^ n1056 ;
  assign n1066 = n1059 & ~n1065 ;
  assign n1067 = n1066 ^ n1058 ;
  assign n1061 = n1060 ^ n1053 ;
  assign n1062 = n1055 & ~n1061 ;
  assign n1063 = n1062 ^ n1054 ;
  assign n1050 = n1049 ^ n1046 ;
  assign n1051 = n1048 & ~n1050 ;
  assign n1052 = n1051 ^ n1047 ;
  assign n1064 = n1063 ^ n1052 ;
  assign n1090 = n1067 ^ n1064 ;
  assign n1087 = n1086 ^ n1071 ;
  assign n1088 = n1073 & ~n1087 ;
  assign n1089 = n1088 ^ n1072 ;
  assign n1091 = n1090 ^ n1089 ;
  assign n1176 = n1102 ^ n1091 ;
  assign n1177 = n1176 ^ n1174 ;
  assign n1178 = n1175 & ~n1177 ;
  assign n1179 = n1178 ^ n1147 ;
  assign n1191 = n1190 ^ n1179 ;
  assign n1107 = n1097 ^ n1094 ;
  assign n1108 = n1101 & ~n1107 ;
  assign n1109 = n1108 ^ n1100 ;
  assign n1103 = n1102 ^ n1090 ;
  assign n1104 = n1091 & ~n1103 ;
  assign n1105 = n1104 ^ n1089 ;
  assign n1068 = n1067 ^ n1052 ;
  assign n1069 = n1064 & ~n1068 ;
  assign n1070 = n1069 ^ n1063 ;
  assign n1106 = n1105 ^ n1070 ;
  assign n1192 = n1109 ^ n1106 ;
  assign n1193 = n1192 ^ n1179 ;
  assign n1194 = n1191 & ~n1193 ;
  assign n1195 = n1194 ^ n1190 ;
  assign n1199 = n1198 ^ n1195 ;
  assign n1110 = n1109 ^ n1070 ;
  assign n1111 = n1106 & ~n1110 ;
  assign n1112 = n1111 ^ n1105 ;
  assign n1200 = n1199 ^ n1112 ;
  assign n1201 = n1176 ^ n1175 ;
  assign n1202 = n1144 ^ n1143 ;
  assign n1203 = x512 ^ x128 ;
  assign n1204 = n1202 & n1203 ;
  assign n1205 = n1201 & n1204 ;
  assign n1206 = n1192 ^ n1191 ;
  assign n1207 = n1205 & n1206 ;
  assign n1208 = n1200 & n1207 ;
  assign n1209 = n1198 ^ n1112 ;
  assign n1210 = ~n1199 & n1209 ;
  assign n1211 = n1210 ^ n1112 ;
  assign n1212 = n1208 & n1211 ;
  assign n3107 = ~n2935 & n3106 ;
  assign n3108 = ~n1212 & ~n3107 ;
  assign n3113 = n3110 ^ n3108 ;
  assign n3109 = n3108 ^ n3107 ;
  assign n3111 = n3110 ^ n3107 ;
  assign n3112 = ~n3109 & ~n3111 ;
  assign n3114 = n3113 ^ n3112 ;
  assign n3115 = n3114 ^ n3109 ;
  assign n3116 = ~n1045 & n3115 ;
  assign n3117 = n3116 ^ n3115 ;
  assign n3118 = n3114 ^ n3111 ;
  assign n3119 = n3117 & n3118 ;
  assign n3120 = n3119 ^ n3117 ;
  assign n801 = x541 ^ x93 ;
  assign n800 = x542 ^ x94 ;
  assign n802 = n801 ^ n800 ;
  assign n799 = x543 ^ x95 ;
  assign n834 = n800 ^ n799 ;
  assign n835 = n802 & ~n834 ;
  assign n836 = n835 ^ n801 ;
  assign n804 = x537 ^ x89 ;
  assign n803 = n802 ^ n799 ;
  assign n805 = n804 ^ n803 ;
  assign n796 = x539 ^ x91 ;
  assign n795 = x538 ^ x90 ;
  assign n797 = n796 ^ n795 ;
  assign n794 = x540 ^ x92 ;
  assign n798 = n797 ^ n794 ;
  assign n831 = n803 ^ n798 ;
  assign n832 = n805 & ~n831 ;
  assign n833 = n832 ^ n804 ;
  assign n837 = n836 ^ n833 ;
  assign n828 = n795 ^ n794 ;
  assign n829 = n797 & ~n828 ;
  assign n830 = n829 ^ n796 ;
  assign n852 = n833 ^ n830 ;
  assign n853 = n837 & ~n852 ;
  assign n854 = n853 ^ n836 ;
  assign n838 = n837 ^ n830 ;
  assign n806 = n805 ^ n798 ;
  assign n793 = x529 ^ x81 ;
  assign n807 = n806 ^ n793 ;
  assign n788 = x535 ^ x87 ;
  assign n787 = x534 ^ x86 ;
  assign n789 = n788 ^ n787 ;
  assign n786 = x536 ^ x88 ;
  assign n790 = n789 ^ n786 ;
  assign n785 = x530 ^ x82 ;
  assign n791 = n790 ^ n785 ;
  assign n782 = x532 ^ x84 ;
  assign n781 = x531 ^ x83 ;
  assign n783 = n782 ^ n781 ;
  assign n780 = x533 ^ x85 ;
  assign n784 = n783 ^ n780 ;
  assign n792 = n791 ^ n784 ;
  assign n825 = n793 ^ n792 ;
  assign n826 = n807 & ~n825 ;
  assign n827 = n826 ^ n806 ;
  assign n839 = n838 ^ n827 ;
  assign n820 = n785 ^ n784 ;
  assign n821 = n791 & ~n820 ;
  assign n822 = n821 ^ n790 ;
  assign n817 = n787 ^ n786 ;
  assign n818 = n789 & ~n817 ;
  assign n819 = n818 ^ n788 ;
  assign n823 = n822 ^ n819 ;
  assign n814 = n781 ^ n780 ;
  assign n815 = n783 & ~n814 ;
  assign n816 = n815 ^ n782 ;
  assign n824 = n823 ^ n816 ;
  assign n849 = n838 ^ n824 ;
  assign n850 = n839 & ~n849 ;
  assign n851 = n850 ^ n827 ;
  assign n855 = n854 ^ n851 ;
  assign n846 = n819 ^ n816 ;
  assign n847 = n823 & ~n846 ;
  assign n848 = n847 ^ n822 ;
  assign n862 = n851 ^ n848 ;
  assign n863 = n855 & ~n862 ;
  assign n864 = n863 ^ n854 ;
  assign n856 = n855 ^ n848 ;
  assign n840 = n839 ^ n824 ;
  assign n808 = n807 ^ n792 ;
  assign n779 = x513 ^ x65 ;
  assign n809 = n808 ^ n779 ;
  assign n749 = x517 ^ x69 ;
  assign n748 = x516 ^ x68 ;
  assign n750 = n749 ^ n748 ;
  assign n747 = x518 ^ x70 ;
  assign n751 = n750 ^ n747 ;
  assign n743 = x520 ^ x72 ;
  assign n742 = x519 ^ x71 ;
  assign n744 = n743 ^ n742 ;
  assign n741 = x521 ^ x73 ;
  assign n745 = n744 ^ n741 ;
  assign n740 = x515 ^ x67 ;
  assign n746 = n745 ^ n740 ;
  assign n752 = n751 ^ n746 ;
  assign n738 = x514 ^ x66 ;
  assign n724 = x524 ^ x76 ;
  assign n723 = x523 ^ x75 ;
  assign n725 = n724 ^ n723 ;
  assign n722 = x525 ^ x77 ;
  assign n726 = n725 ^ n722 ;
  assign n715 = x528 ^ x80 ;
  assign n713 = x527 ^ x79 ;
  assign n712 = x526 ^ x78 ;
  assign n714 = n713 ^ n712 ;
  assign n720 = n715 ^ n714 ;
  assign n719 = x522 ^ x74 ;
  assign n721 = n720 ^ n719 ;
  assign n737 = n726 ^ n721 ;
  assign n739 = n738 ^ n737 ;
  assign n810 = n752 ^ n739 ;
  assign n811 = n810 ^ n779 ;
  assign n812 = n809 & ~n811 ;
  assign n813 = n812 ^ n808 ;
  assign n841 = n840 ^ n813 ;
  assign n764 = n742 ^ n741 ;
  assign n765 = n744 & ~n764 ;
  assign n766 = n765 ^ n743 ;
  assign n761 = n751 ^ n745 ;
  assign n762 = ~n746 & n761 ;
  assign n763 = n762 ^ n751 ;
  assign n767 = n766 ^ n763 ;
  assign n758 = n748 ^ n747 ;
  assign n759 = n750 & ~n758 ;
  assign n760 = n759 ^ n749 ;
  assign n768 = n767 ^ n760 ;
  assign n731 = n723 ^ n722 ;
  assign n732 = n725 & ~n731 ;
  assign n733 = n732 ^ n724 ;
  assign n727 = n726 ^ n719 ;
  assign n728 = n721 & ~n727 ;
  assign n729 = n728 ^ n720 ;
  assign n716 = n715 ^ n712 ;
  assign n717 = n714 & ~n716 ;
  assign n718 = n717 ^ n713 ;
  assign n730 = n729 ^ n718 ;
  assign n756 = n733 ^ n730 ;
  assign n753 = n752 ^ n737 ;
  assign n754 = n739 & ~n753 ;
  assign n755 = n754 ^ n738 ;
  assign n757 = n756 ^ n755 ;
  assign n842 = n768 ^ n757 ;
  assign n843 = n842 ^ n840 ;
  assign n844 = n841 & ~n843 ;
  assign n845 = n844 ^ n813 ;
  assign n857 = n856 ^ n845 ;
  assign n773 = n763 ^ n760 ;
  assign n774 = n767 & ~n773 ;
  assign n775 = n774 ^ n766 ;
  assign n769 = n768 ^ n756 ;
  assign n770 = n757 & ~n769 ;
  assign n771 = n770 ^ n755 ;
  assign n734 = n733 ^ n718 ;
  assign n735 = n730 & ~n734 ;
  assign n736 = n735 ^ n729 ;
  assign n772 = n771 ^ n736 ;
  assign n858 = n775 ^ n772 ;
  assign n859 = n858 ^ n845 ;
  assign n860 = n857 & ~n859 ;
  assign n861 = n860 ^ n856 ;
  assign n865 = n864 ^ n861 ;
  assign n776 = n775 ^ n736 ;
  assign n777 = n772 & ~n776 ;
  assign n778 = n777 ^ n771 ;
  assign n866 = n865 ^ n778 ;
  assign n867 = n842 ^ n841 ;
  assign n868 = n810 ^ n809 ;
  assign n869 = x512 ^ x64 ;
  assign n870 = n868 & n869 ;
  assign n871 = n867 & n870 ;
  assign n872 = n858 ^ n857 ;
  assign n873 = n871 & n872 ;
  assign n874 = n866 & n873 ;
  assign n875 = n864 ^ n778 ;
  assign n876 = ~n865 & n875 ;
  assign n877 = n876 ^ n778 ;
  assign n878 = n874 & n877 ;
  assign n3121 = n3120 ^ n3118 ;
  assign n3122 = n3121 ^ n3117 ;
  assign n3123 = ~n878 & ~n3122 ;
  assign n3124 = n3123 ^ n3122 ;
  assign n3126 = ~n3120 & n3124 ;
  assign n3217 = x541 ^ x61 ;
  assign n3216 = x542 ^ x62 ;
  assign n3218 = n3217 ^ n3216 ;
  assign n3215 = x543 ^ x63 ;
  assign n3250 = n3216 ^ n3215 ;
  assign n3251 = n3218 & ~n3250 ;
  assign n3252 = n3251 ^ n3217 ;
  assign n3220 = x537 ^ x57 ;
  assign n3219 = n3218 ^ n3215 ;
  assign n3221 = n3220 ^ n3219 ;
  assign n3212 = x539 ^ x59 ;
  assign n3211 = x538 ^ x58 ;
  assign n3213 = n3212 ^ n3211 ;
  assign n3210 = x540 ^ x60 ;
  assign n3214 = n3213 ^ n3210 ;
  assign n3247 = n3219 ^ n3214 ;
  assign n3248 = n3221 & ~n3247 ;
  assign n3249 = n3248 ^ n3220 ;
  assign n3253 = n3252 ^ n3249 ;
  assign n3244 = n3211 ^ n3210 ;
  assign n3245 = n3213 & ~n3244 ;
  assign n3246 = n3245 ^ n3212 ;
  assign n3268 = n3249 ^ n3246 ;
  assign n3269 = n3253 & ~n3268 ;
  assign n3270 = n3269 ^ n3252 ;
  assign n3254 = n3253 ^ n3246 ;
  assign n3222 = n3221 ^ n3214 ;
  assign n3209 = x529 ^ x49 ;
  assign n3223 = n3222 ^ n3209 ;
  assign n3204 = x535 ^ x55 ;
  assign n3203 = x534 ^ x54 ;
  assign n3205 = n3204 ^ n3203 ;
  assign n3202 = x536 ^ x56 ;
  assign n3206 = n3205 ^ n3202 ;
  assign n3201 = x530 ^ x50 ;
  assign n3207 = n3206 ^ n3201 ;
  assign n3198 = x532 ^ x52 ;
  assign n3197 = x531 ^ x51 ;
  assign n3199 = n3198 ^ n3197 ;
  assign n3196 = x533 ^ x53 ;
  assign n3200 = n3199 ^ n3196 ;
  assign n3208 = n3207 ^ n3200 ;
  assign n3241 = n3209 ^ n3208 ;
  assign n3242 = n3223 & ~n3241 ;
  assign n3243 = n3242 ^ n3222 ;
  assign n3255 = n3254 ^ n3243 ;
  assign n3236 = n3201 ^ n3200 ;
  assign n3237 = n3207 & ~n3236 ;
  assign n3238 = n3237 ^ n3206 ;
  assign n3233 = n3203 ^ n3202 ;
  assign n3234 = n3205 & ~n3233 ;
  assign n3235 = n3234 ^ n3204 ;
  assign n3239 = n3238 ^ n3235 ;
  assign n3230 = n3197 ^ n3196 ;
  assign n3231 = n3199 & ~n3230 ;
  assign n3232 = n3231 ^ n3198 ;
  assign n3240 = n3239 ^ n3232 ;
  assign n3265 = n3254 ^ n3240 ;
  assign n3266 = n3255 & ~n3265 ;
  assign n3267 = n3266 ^ n3243 ;
  assign n3271 = n3270 ^ n3267 ;
  assign n3262 = n3235 ^ n3232 ;
  assign n3263 = n3239 & ~n3262 ;
  assign n3264 = n3263 ^ n3238 ;
  assign n3278 = n3267 ^ n3264 ;
  assign n3279 = n3271 & ~n3278 ;
  assign n3280 = n3279 ^ n3270 ;
  assign n3272 = n3271 ^ n3264 ;
  assign n3256 = n3255 ^ n3240 ;
  assign n3224 = n3223 ^ n3208 ;
  assign n3195 = x513 ^ x33 ;
  assign n3225 = n3224 ^ n3195 ;
  assign n3165 = x517 ^ x37 ;
  assign n3164 = x516 ^ x36 ;
  assign n3166 = n3165 ^ n3164 ;
  assign n3163 = x518 ^ x38 ;
  assign n3167 = n3166 ^ n3163 ;
  assign n3159 = x520 ^ x40 ;
  assign n3158 = x519 ^ x39 ;
  assign n3160 = n3159 ^ n3158 ;
  assign n3157 = x521 ^ x41 ;
  assign n3161 = n3160 ^ n3157 ;
  assign n3156 = x515 ^ x35 ;
  assign n3162 = n3161 ^ n3156 ;
  assign n3168 = n3167 ^ n3162 ;
  assign n3154 = x514 ^ x34 ;
  assign n3140 = x524 ^ x44 ;
  assign n3139 = x523 ^ x43 ;
  assign n3141 = n3140 ^ n3139 ;
  assign n3138 = x525 ^ x45 ;
  assign n3142 = n3141 ^ n3138 ;
  assign n3131 = x528 ^ x48 ;
  assign n3129 = x527 ^ x47 ;
  assign n3128 = x526 ^ x46 ;
  assign n3130 = n3129 ^ n3128 ;
  assign n3136 = n3131 ^ n3130 ;
  assign n3135 = x522 ^ x42 ;
  assign n3137 = n3136 ^ n3135 ;
  assign n3153 = n3142 ^ n3137 ;
  assign n3155 = n3154 ^ n3153 ;
  assign n3226 = n3168 ^ n3155 ;
  assign n3227 = n3226 ^ n3195 ;
  assign n3228 = n3225 & ~n3227 ;
  assign n3229 = n3228 ^ n3224 ;
  assign n3257 = n3256 ^ n3229 ;
  assign n3180 = n3158 ^ n3157 ;
  assign n3181 = n3160 & ~n3180 ;
  assign n3182 = n3181 ^ n3159 ;
  assign n3177 = n3167 ^ n3161 ;
  assign n3178 = ~n3162 & n3177 ;
  assign n3179 = n3178 ^ n3167 ;
  assign n3183 = n3182 ^ n3179 ;
  assign n3174 = n3164 ^ n3163 ;
  assign n3175 = n3166 & ~n3174 ;
  assign n3176 = n3175 ^ n3165 ;
  assign n3184 = n3183 ^ n3176 ;
  assign n3147 = n3139 ^ n3138 ;
  assign n3148 = n3141 & ~n3147 ;
  assign n3149 = n3148 ^ n3140 ;
  assign n3143 = n3142 ^ n3135 ;
  assign n3144 = n3137 & ~n3143 ;
  assign n3145 = n3144 ^ n3136 ;
  assign n3132 = n3131 ^ n3128 ;
  assign n3133 = n3130 & ~n3132 ;
  assign n3134 = n3133 ^ n3129 ;
  assign n3146 = n3145 ^ n3134 ;
  assign n3172 = n3149 ^ n3146 ;
  assign n3169 = n3168 ^ n3153 ;
  assign n3170 = n3155 & ~n3169 ;
  assign n3171 = n3170 ^ n3154 ;
  assign n3173 = n3172 ^ n3171 ;
  assign n3258 = n3184 ^ n3173 ;
  assign n3259 = n3258 ^ n3256 ;
  assign n3260 = n3257 & ~n3259 ;
  assign n3261 = n3260 ^ n3229 ;
  assign n3273 = n3272 ^ n3261 ;
  assign n3189 = n3179 ^ n3176 ;
  assign n3190 = n3183 & ~n3189 ;
  assign n3191 = n3190 ^ n3182 ;
  assign n3185 = n3184 ^ n3172 ;
  assign n3186 = n3173 & ~n3185 ;
  assign n3187 = n3186 ^ n3171 ;
  assign n3150 = n3149 ^ n3134 ;
  assign n3151 = n3146 & ~n3150 ;
  assign n3152 = n3151 ^ n3145 ;
  assign n3188 = n3187 ^ n3152 ;
  assign n3274 = n3191 ^ n3188 ;
  assign n3275 = n3274 ^ n3261 ;
  assign n3276 = n3273 & ~n3275 ;
  assign n3277 = n3276 ^ n3272 ;
  assign n3281 = n3280 ^ n3277 ;
  assign n3192 = n3191 ^ n3152 ;
  assign n3193 = n3188 & ~n3192 ;
  assign n3194 = n3193 ^ n3187 ;
  assign n3282 = n3281 ^ n3194 ;
  assign n3283 = n3258 ^ n3257 ;
  assign n3284 = n3226 ^ n3225 ;
  assign n3285 = x512 ^ x32 ;
  assign n3286 = n3284 & n3285 ;
  assign n3287 = n3283 & n3286 ;
  assign n3288 = n3274 ^ n3273 ;
  assign n3289 = n3287 & n3288 ;
  assign n3290 = n3282 & n3289 ;
  assign n3291 = n3280 ^ n3194 ;
  assign n3292 = ~n3281 & n3291 ;
  assign n3293 = n3292 ^ n3194 ;
  assign n3294 = n3290 & n3293 ;
  assign n3295 = ~n3126 & ~n3294 ;
  assign n3125 = n3124 ^ n3120 ;
  assign n3298 = n3295 ^ n3125 ;
  assign n3127 = n3126 ^ n3125 ;
  assign n3296 = n3295 ^ n3126 ;
  assign n3297 = ~n3127 & ~n3296 ;
  assign n3299 = n3298 ^ n3297 ;
  assign n3300 = n3299 ^ n3127 ;
  assign n3301 = ~n711 & ~n3300 ;
  assign n4304 = n3293 ^ n3290 ;
  assign n4225 = n877 ^ n874 ;
  assign n4142 = n1044 ^ n1041 ;
  assign n4063 = n1211 ^ n1208 ;
  assign n3984 = n3101 ^ n3098 ;
  assign n3901 = n1378 ^ n1375 ;
  assign n3822 = n1545 ^ n1542 ;
  assign n3743 = n2916 ^ n2913 ;
  assign n3660 = n1712 ^ n1709 ;
  assign n3581 = n1879 ^ n1876 ;
  assign n3497 = n2731 ^ n2728 ;
  assign n3417 = n2046 ^ n2043 ;
  assign n3334 = n2382 ^ n2214 ;
  assign n3302 = n2213 ^ n2210 ;
  assign n3303 = n3302 ^ n2382 ;
  assign n3304 = n2382 & ~n3302 ;
  assign n3305 = n3304 ^ n2384 ;
  assign n3306 = n3304 ^ n3303 ;
  assign n3308 = n2209 ^ n2198 ;
  assign n3307 = n2376 ^ n2365 ;
  assign n3309 = n3308 ^ n3307 ;
  assign n3311 = n2364 ^ n2359 ;
  assign n3310 = n2197 ^ n2192 ;
  assign n3312 = n3311 ^ n3310 ;
  assign n3316 = n2196 ^ n2193 ;
  assign n3313 = n2195 ^ n2194 ;
  assign n3314 = n2362 ^ n2361 ;
  assign n3315 = ~n3313 & n3314 ;
  assign n3317 = n3316 ^ n3315 ;
  assign n3318 = n3315 ^ n2363 ;
  assign n3319 = n3318 ^ n2360 ;
  assign n3320 = ~n3317 & ~n3319 ;
  assign n3321 = n3320 ^ n3316 ;
  assign n3322 = n3321 ^ n3311 ;
  assign n3323 = ~n3312 & n3322 ;
  assign n3324 = n3323 ^ n3310 ;
  assign n3325 = n3324 ^ n3308 ;
  assign n3326 = ~n3309 & n3325 ;
  assign n3327 = n3326 ^ n3308 ;
  assign n3328 = ~n3306 & ~n3327 ;
  assign n3329 = ~n3305 & ~n3328 ;
  assign n3330 = n2555 & ~n3329 ;
  assign n3331 = n3303 & ~n3330 ;
  assign n3335 = n3334 ^ n3331 ;
  assign n3336 = n3335 ^ n2214 ;
  assign n3333 = n2551 ^ n2548 ;
  assign n3337 = n3336 ^ n3333 ;
  assign n3338 = n2544 ^ n2541 ;
  assign n3339 = n2363 ^ n2360 ;
  assign n3340 = n3339 ^ n3316 ;
  assign n3341 = ~n3330 & n3340 ;
  assign n3342 = n3341 ^ n3340 ;
  assign n3343 = n3342 ^ n3316 ;
  assign n3344 = n3338 & ~n3343 ;
  assign n3345 = n2543 ^ n2542 ;
  assign n3346 = n3314 ^ n3313 ;
  assign n3347 = ~n3330 & n3346 ;
  assign n3348 = n3347 ^ n3346 ;
  assign n3349 = n3348 ^ n3313 ;
  assign n3350 = n3345 & ~n3349 ;
  assign n3351 = ~n3344 & ~n3350 ;
  assign n3352 = ~n2541 & n3343 ;
  assign n3356 = n2546 ^ n2545 ;
  assign n3353 = n3312 & ~n3330 ;
  assign n3354 = n3353 ^ n3312 ;
  assign n3355 = n3354 ^ n3310 ;
  assign n3358 = n3356 ^ n3355 ;
  assign n3357 = ~n3355 & n3356 ;
  assign n3359 = n3358 ^ n3357 ;
  assign n3360 = ~n3352 & ~n3359 ;
  assign n3361 = ~n3351 & n3360 ;
  assign n3363 = n3309 & ~n3330 ;
  assign n3364 = n3363 ^ n3307 ;
  assign n3362 = n2547 ^ n2540 ;
  assign n3366 = n3364 ^ n3362 ;
  assign n3365 = ~n3362 & n3364 ;
  assign n3367 = n3366 ^ n3365 ;
  assign n3368 = ~n3357 & ~n3367 ;
  assign n3369 = ~n3361 & n3368 ;
  assign n3370 = ~n3333 & n3336 ;
  assign n3371 = n3370 ^ n2553 ;
  assign n3372 = ~n3365 & ~n3371 ;
  assign n3373 = ~n3369 & n3372 ;
  assign n3374 = n3337 ^ n2552 ;
  assign n3375 = n3374 ^ n3370 ;
  assign n3376 = ~n2385 & n3375 ;
  assign n3377 = ~n3373 & ~n3376 ;
  assign n3378 = n3337 & ~n3377 ;
  assign n3379 = n3378 ^ n3333 ;
  assign n3332 = n3331 ^ n3302 ;
  assign n3380 = n3379 ^ n3332 ;
  assign n3381 = n3332 & ~n3379 ;
  assign n3382 = n3381 ^ n2559 ;
  assign n3383 = n3381 ^ n3380 ;
  assign n3385 = n3366 & n3377 ;
  assign n3386 = n3385 ^ n3364 ;
  assign n3384 = n3363 ^ n3308 ;
  assign n3387 = n3386 ^ n3384 ;
  assign n3389 = n3358 & ~n3377 ;
  assign n3390 = n3389 ^ n3356 ;
  assign n3388 = n3353 ^ n3310 ;
  assign n3391 = n3390 ^ n3388 ;
  assign n3395 = n3341 ^ n3316 ;
  assign n3392 = n3343 ^ n3338 ;
  assign n3393 = ~n3377 & n3392 ;
  assign n3394 = n3393 ^ n3338 ;
  assign n3396 = n3395 ^ n3394 ;
  assign n3397 = n3349 ^ n3345 ;
  assign n3398 = ~n3377 & n3397 ;
  assign n3399 = n3398 ^ n3345 ;
  assign n3400 = n3347 ^ n3313 ;
  assign n3401 = n3399 & ~n3400 ;
  assign n3402 = n3401 ^ n3395 ;
  assign n3403 = ~n3396 & ~n3402 ;
  assign n3404 = n3403 ^ n3395 ;
  assign n3405 = n3404 ^ n3390 ;
  assign n3406 = ~n3391 & ~n3405 ;
  assign n3407 = n3406 ^ n3390 ;
  assign n3408 = n3407 ^ n3386 ;
  assign n3409 = ~n3387 & n3408 ;
  assign n3410 = n3409 ^ n3386 ;
  assign n3411 = ~n3383 & ~n3410 ;
  assign n3412 = n3382 & ~n3411 ;
  assign n3413 = ~n2557 & ~n3412 ;
  assign n3414 = n3380 & n3413 ;
  assign n3416 = n3414 ^ n3379 ;
  assign n3418 = n3417 ^ n3416 ;
  assign n3419 = n2038 ^ n2037 ;
  assign n3420 = n3400 ^ n3399 ;
  assign n3421 = ~n3413 & n3420 ;
  assign n3422 = n3421 ^ n3420 ;
  assign n3423 = n3422 ^ n3399 ;
  assign n3424 = n3419 & ~n3423 ;
  assign n3425 = n2036 & n3424 ;
  assign n3426 = n3396 & ~n3413 ;
  assign n3427 = n3426 ^ n3394 ;
  assign n3428 = n3427 ^ n3395 ;
  assign n3429 = n3428 ^ n3394 ;
  assign n3430 = ~n3425 & n3429 ;
  assign n3431 = n2039 ^ n2036 ;
  assign n3432 = ~n3424 & ~n3431 ;
  assign n3436 = n2041 ^ n2040 ;
  assign n3433 = n3391 & n3413 ;
  assign n3434 = n3433 ^ n3391 ;
  assign n3435 = n3434 ^ n3388 ;
  assign n3438 = n3436 ^ n3435 ;
  assign n3437 = ~n3435 & n3436 ;
  assign n3439 = n3438 ^ n3437 ;
  assign n3440 = ~n3432 & ~n3439 ;
  assign n3441 = ~n3430 & n3440 ;
  assign n3443 = n3387 & n3413 ;
  assign n3444 = n3443 ^ n3386 ;
  assign n3442 = n2042 ^ n2035 ;
  assign n3446 = n3444 ^ n3442 ;
  assign n3445 = ~n3442 & n3444 ;
  assign n3447 = n3446 ^ n3445 ;
  assign n3448 = ~n3437 & ~n3447 ;
  assign n3449 = ~n3441 & n3448 ;
  assign n3450 = n3416 & ~n3417 ;
  assign n3451 = ~n2561 & ~n3445 ;
  assign n3452 = ~n3450 & n3451 ;
  assign n3453 = ~n3449 & n3452 ;
  assign n3454 = n3418 ^ n2047 ;
  assign n3455 = n3454 ^ n3450 ;
  assign n3456 = n2560 & n3455 ;
  assign n3457 = ~n3453 & ~n3456 ;
  assign n3458 = n3418 & ~n3457 ;
  assign n3459 = n3458 ^ n3417 ;
  assign n3415 = n3414 ^ n3332 ;
  assign n3460 = n3459 ^ n3415 ;
  assign n3461 = n2563 ^ n2562 ;
  assign n3463 = n3446 & n3457 ;
  assign n3464 = n3463 ^ n3444 ;
  assign n3462 = n3443 ^ n3384 ;
  assign n3465 = n3464 ^ n3462 ;
  assign n3467 = n3438 & ~n3457 ;
  assign n3468 = n3467 ^ n3436 ;
  assign n3466 = n3433 ^ n3388 ;
  assign n3469 = n3468 ^ n3466 ;
  assign n3470 = n3431 ^ n3429 ;
  assign n3471 = n3457 & n3470 ;
  assign n3472 = n3471 ^ n3429 ;
  assign n3473 = n3472 ^ n3427 ;
  assign n3474 = n3423 ^ n3419 ;
  assign n3475 = ~n3457 & n3474 ;
  assign n3476 = n3475 ^ n3419 ;
  assign n3477 = n3421 ^ n3399 ;
  assign n3478 = n3476 & ~n3477 ;
  assign n3479 = n3478 ^ n3427 ;
  assign n3480 = ~n3473 & ~n3479 ;
  assign n3481 = n3480 ^ n3427 ;
  assign n3482 = n3481 ^ n3468 ;
  assign n3483 = ~n3469 & ~n3482 ;
  assign n3484 = n3483 ^ n3468 ;
  assign n3485 = n3484 ^ n3464 ;
  assign n3486 = ~n3465 & n3485 ;
  assign n3487 = n3486 ^ n3464 ;
  assign n3488 = n3487 ^ n3459 ;
  assign n3489 = ~n3460 & n3488 ;
  assign n3490 = n3489 ^ n3459 ;
  assign n3491 = n3490 ^ n2563 ;
  assign n3492 = n3461 & n3491 ;
  assign n3493 = n3492 ^ n2562 ;
  assign n3494 = n3460 & n3493 ;
  assign n3496 = n3494 ^ n3459 ;
  assign n3498 = n3497 ^ n3496 ;
  assign n3499 = n2724 ^ n2721 ;
  assign n3500 = n3473 & ~n3493 ;
  assign n3501 = n3500 ^ n3472 ;
  assign n3502 = n3501 ^ n3427 ;
  assign n3503 = n3502 ^ n3472 ;
  assign n3504 = n3499 & ~n3503 ;
  assign n3505 = n2723 ^ n2722 ;
  assign n3506 = n3477 ^ n3476 ;
  assign n3507 = ~n3493 & n3506 ;
  assign n3508 = n3507 ^ n3506 ;
  assign n3509 = n3508 ^ n3476 ;
  assign n3510 = n3505 & ~n3509 ;
  assign n3511 = ~n3504 & ~n3510 ;
  assign n3512 = ~n2721 & n3503 ;
  assign n3516 = n2726 ^ n2725 ;
  assign n3513 = n3469 & n3493 ;
  assign n3514 = n3513 ^ n3469 ;
  assign n3515 = n3514 ^ n3466 ;
  assign n3518 = n3516 ^ n3515 ;
  assign n3517 = ~n3515 & n3516 ;
  assign n3519 = n3518 ^ n3517 ;
  assign n3520 = ~n3512 & ~n3519 ;
  assign n3521 = ~n3511 & n3520 ;
  assign n3524 = n2727 ^ n2720 ;
  assign n3522 = n3465 & n3493 ;
  assign n3523 = n3522 ^ n3464 ;
  assign n3526 = n3524 ^ n3523 ;
  assign n3525 = n3523 & ~n3524 ;
  assign n3527 = n3526 ^ n3525 ;
  assign n3528 = ~n3517 & ~n3527 ;
  assign n3529 = ~n3521 & n3528 ;
  assign n3530 = n3496 & ~n3497 ;
  assign n3531 = ~n2735 & ~n3530 ;
  assign n3532 = ~n3525 & n3531 ;
  assign n3533 = ~n3529 & n3532 ;
  assign n3534 = n3498 ^ n2732 ;
  assign n3535 = n3534 ^ n3530 ;
  assign n3536 = ~n2734 & n3535 ;
  assign n3537 = ~n3533 & ~n3536 ;
  assign n3538 = n3498 & ~n3537 ;
  assign n3539 = n3538 ^ n3497 ;
  assign n3495 = n3494 ^ n3415 ;
  assign n3540 = n3539 ^ n3495 ;
  assign n3541 = ~n3495 & n3539 ;
  assign n3542 = n3541 ^ n3540 ;
  assign n3543 = n3542 ^ n2565 ;
  assign n3544 = n3543 ^ n2565 ;
  assign n3546 = n3526 & n3537 ;
  assign n3547 = n3546 ^ n3523 ;
  assign n3545 = n3522 ^ n3462 ;
  assign n3548 = n3547 ^ n3545 ;
  assign n3550 = n3518 & ~n3537 ;
  assign n3551 = n3550 ^ n3516 ;
  assign n3549 = n3513 ^ n3466 ;
  assign n3552 = n3551 ^ n3549 ;
  assign n3553 = n3503 ^ n3499 ;
  assign n3554 = ~n3537 & n3553 ;
  assign n3555 = n3554 ^ n3499 ;
  assign n3556 = n3555 ^ n3501 ;
  assign n3557 = n3509 ^ n3505 ;
  assign n3558 = ~n3537 & n3557 ;
  assign n3559 = n3558 ^ n3505 ;
  assign n3560 = n3507 ^ n3476 ;
  assign n3561 = n3559 & ~n3560 ;
  assign n3562 = n3561 ^ n3501 ;
  assign n3563 = ~n3556 & ~n3562 ;
  assign n3564 = n3563 ^ n3501 ;
  assign n3565 = n3564 ^ n3551 ;
  assign n3566 = ~n3552 & ~n3565 ;
  assign n3567 = n3566 ^ n3551 ;
  assign n3568 = n3567 ^ n3545 ;
  assign n3569 = ~n3548 & ~n3568 ;
  assign n3570 = n3569 ^ n3545 ;
  assign n3571 = ~n3541 & n3570 ;
  assign n3572 = n3571 ^ n2565 ;
  assign n3573 = n3572 ^ n2565 ;
  assign n3574 = ~n3544 & ~n3573 ;
  assign n3575 = n3574 ^ n2565 ;
  assign n3576 = n2740 & ~n3575 ;
  assign n3577 = n3576 ^ n2736 ;
  assign n3578 = n3540 & ~n3577 ;
  assign n3580 = n3578 ^ n3539 ;
  assign n3582 = n3581 ^ n3580 ;
  assign n3583 = n1872 ^ n1869 ;
  assign n3584 = n3556 & n3577 ;
  assign n3585 = n3584 ^ n3556 ;
  assign n3586 = n3585 ^ n3555 ;
  assign n3587 = n3583 & ~n3586 ;
  assign n3588 = n1871 ^ n1870 ;
  assign n3589 = n3560 ^ n3559 ;
  assign n3590 = n3577 & n3589 ;
  assign n3591 = n3590 ^ n3589 ;
  assign n3592 = n3591 ^ n3559 ;
  assign n3593 = n3588 & ~n3592 ;
  assign n3594 = ~n3587 & ~n3593 ;
  assign n3595 = ~n1869 & n3586 ;
  assign n3599 = n1874 ^ n1873 ;
  assign n3596 = n3552 & ~n3577 ;
  assign n3597 = n3596 ^ n3552 ;
  assign n3598 = n3597 ^ n3549 ;
  assign n3601 = n3599 ^ n3598 ;
  assign n3600 = ~n3598 & n3599 ;
  assign n3602 = n3601 ^ n3600 ;
  assign n3603 = ~n3595 & ~n3602 ;
  assign n3604 = ~n3594 & n3603 ;
  assign n3606 = n3548 & ~n3577 ;
  assign n3607 = n3606 ^ n3547 ;
  assign n3605 = n1875 ^ n1868 ;
  assign n3609 = n3607 ^ n3605 ;
  assign n3608 = ~n3605 & n3607 ;
  assign n3610 = n3609 ^ n3608 ;
  assign n3611 = ~n3600 & ~n3610 ;
  assign n3612 = ~n3604 & n3611 ;
  assign n3613 = n3580 & ~n3581 ;
  assign n3614 = ~n2738 & ~n3613 ;
  assign n3615 = ~n3608 & n3614 ;
  assign n3616 = ~n3612 & n3615 ;
  assign n3617 = n3582 ^ n1880 ;
  assign n3618 = n3617 ^ n3613 ;
  assign n3619 = n2737 & n3618 ;
  assign n3620 = ~n3616 & ~n3619 ;
  assign n3621 = n3582 & ~n3620 ;
  assign n3622 = n3621 ^ n3581 ;
  assign n3579 = n3578 ^ n3495 ;
  assign n3623 = n3622 ^ n3579 ;
  assign n3625 = n3609 & n3620 ;
  assign n3626 = n3625 ^ n3607 ;
  assign n3624 = n3606 ^ n3545 ;
  assign n3627 = n3626 ^ n3624 ;
  assign n3629 = n3601 & ~n3620 ;
  assign n3630 = n3629 ^ n3599 ;
  assign n3628 = n3596 ^ n3549 ;
  assign n3631 = n3630 ^ n3628 ;
  assign n3633 = n3586 ^ n3583 ;
  assign n3634 = ~n3620 & n3633 ;
  assign n3635 = n3634 ^ n3583 ;
  assign n3632 = n3584 ^ n3555 ;
  assign n3636 = n3635 ^ n3632 ;
  assign n3637 = n3592 ^ n3588 ;
  assign n3638 = ~n3620 & n3637 ;
  assign n3639 = n3638 ^ n3588 ;
  assign n3640 = n3590 ^ n3559 ;
  assign n3641 = n3639 & ~n3640 ;
  assign n3642 = n3641 ^ n3635 ;
  assign n3643 = ~n3636 & n3642 ;
  assign n3644 = n3643 ^ n3635 ;
  assign n3645 = n3644 ^ n3630 ;
  assign n3646 = ~n3631 & n3645 ;
  assign n3647 = n3646 ^ n3630 ;
  assign n3648 = n3647 ^ n3626 ;
  assign n3649 = ~n3627 & n3648 ;
  assign n3650 = n3649 ^ n3626 ;
  assign n3651 = n3650 ^ n3622 ;
  assign n3652 = ~n3623 & n3651 ;
  assign n3653 = n3652 ^ n3622 ;
  assign n3654 = n3653 ^ n2741 ;
  assign n3655 = ~n2743 & ~n3654 ;
  assign n3656 = n3655 ^ n3653 ;
  assign n3657 = n3623 & ~n3656 ;
  assign n3659 = n3657 ^ n3622 ;
  assign n3661 = n3660 ^ n3659 ;
  assign n3662 = n1705 ^ n1702 ;
  assign n3663 = n3636 & ~n3656 ;
  assign n3664 = n3663 ^ n3632 ;
  assign n3665 = n3664 ^ n3635 ;
  assign n3666 = n3665 ^ n3632 ;
  assign n3667 = n3662 & ~n3666 ;
  assign n3668 = n1704 ^ n1703 ;
  assign n3669 = n3640 ^ n3639 ;
  assign n3670 = n3656 & n3669 ;
  assign n3671 = n3670 ^ n3669 ;
  assign n3672 = n3671 ^ n3639 ;
  assign n3673 = n3668 & ~n3672 ;
  assign n3674 = ~n3667 & ~n3673 ;
  assign n3675 = ~n1702 & n3666 ;
  assign n3679 = n1707 ^ n1706 ;
  assign n3676 = n3631 & ~n3656 ;
  assign n3677 = n3676 ^ n3631 ;
  assign n3678 = n3677 ^ n3628 ;
  assign n3681 = n3679 ^ n3678 ;
  assign n3680 = ~n3678 & n3679 ;
  assign n3682 = n3681 ^ n3680 ;
  assign n3683 = ~n3675 & ~n3682 ;
  assign n3684 = ~n3674 & n3683 ;
  assign n3686 = n3627 & ~n3656 ;
  assign n3687 = n3686 ^ n3626 ;
  assign n3685 = n1708 ^ n1701 ;
  assign n3689 = n3687 ^ n3685 ;
  assign n3688 = ~n3685 & n3687 ;
  assign n3690 = n3689 ^ n3688 ;
  assign n3691 = ~n3680 & ~n3690 ;
  assign n3692 = ~n3684 & n3691 ;
  assign n3693 = n3659 & ~n3660 ;
  assign n3694 = ~n2746 & ~n3693 ;
  assign n3695 = ~n3688 & n3694 ;
  assign n3696 = ~n3692 & n3695 ;
  assign n3697 = n3661 ^ n1713 ;
  assign n3698 = n3697 ^ n3693 ;
  assign n3699 = ~n2745 & n3698 ;
  assign n3700 = ~n3696 & ~n3699 ;
  assign n3701 = n3661 & ~n3700 ;
  assign n3702 = n3701 ^ n3660 ;
  assign n3658 = n3657 ^ n3579 ;
  assign n3703 = n3702 ^ n3658 ;
  assign n3704 = n2748 ^ n2747 ;
  assign n3705 = n3658 & ~n3702 ;
  assign n3706 = n3705 ^ n3703 ;
  assign n3708 = n3689 & n3700 ;
  assign n3709 = n3708 ^ n3687 ;
  assign n3707 = n3686 ^ n3624 ;
  assign n3710 = n3709 ^ n3707 ;
  assign n3712 = n3681 & ~n3700 ;
  assign n3713 = n3712 ^ n3679 ;
  assign n3711 = n3676 ^ n3628 ;
  assign n3714 = n3713 ^ n3711 ;
  assign n3715 = n3666 ^ n3662 ;
  assign n3716 = ~n3700 & n3715 ;
  assign n3717 = n3716 ^ n3662 ;
  assign n3718 = n3717 ^ n3664 ;
  assign n3719 = n3672 ^ n3668 ;
  assign n3720 = ~n3700 & n3719 ;
  assign n3721 = n3720 ^ n3668 ;
  assign n3722 = n3670 ^ n3639 ;
  assign n3723 = n3721 & ~n3722 ;
  assign n3724 = n3723 ^ n3664 ;
  assign n3725 = ~n3718 & ~n3724 ;
  assign n3726 = n3725 ^ n3664 ;
  assign n3727 = n3726 ^ n3713 ;
  assign n3728 = ~n3714 & ~n3727 ;
  assign n3729 = n3728 ^ n3713 ;
  assign n3730 = n3729 ^ n3709 ;
  assign n3731 = ~n3710 & n3730 ;
  assign n3732 = n3731 ^ n3709 ;
  assign n3733 = ~n3706 & ~n3732 ;
  assign n3734 = n3733 ^ n2748 ;
  assign n3735 = n3734 ^ n2748 ;
  assign n3736 = ~n3705 & ~n3735 ;
  assign n3737 = n3736 ^ n2748 ;
  assign n3738 = n3704 & ~n3737 ;
  assign n3739 = n3738 ^ n2747 ;
  assign n3740 = n3703 & ~n3739 ;
  assign n3742 = n3740 ^ n3702 ;
  assign n3744 = n3743 ^ n3742 ;
  assign n3745 = n2909 ^ n2906 ;
  assign n3746 = n3718 & n3739 ;
  assign n3747 = n3746 ^ n3717 ;
  assign n3748 = n3747 ^ n3664 ;
  assign n3749 = n3748 ^ n3717 ;
  assign n3750 = n3745 & ~n3749 ;
  assign n3751 = n2908 ^ n2907 ;
  assign n3752 = n3722 ^ n3721 ;
  assign n3753 = n3739 & n3752 ;
  assign n3754 = n3753 ^ n3752 ;
  assign n3755 = n3754 ^ n3721 ;
  assign n3756 = n3751 & ~n3755 ;
  assign n3757 = ~n3750 & ~n3756 ;
  assign n3758 = ~n2906 & n3749 ;
  assign n3762 = n2911 ^ n2910 ;
  assign n3759 = n3714 & ~n3739 ;
  assign n3760 = n3759 ^ n3714 ;
  assign n3761 = n3760 ^ n3711 ;
  assign n3764 = n3762 ^ n3761 ;
  assign n3763 = ~n3761 & n3762 ;
  assign n3765 = n3764 ^ n3763 ;
  assign n3766 = ~n3758 & ~n3765 ;
  assign n3767 = ~n3757 & n3766 ;
  assign n3770 = n2912 ^ n2905 ;
  assign n3768 = n3710 & ~n3739 ;
  assign n3769 = n3768 ^ n3709 ;
  assign n3772 = n3770 ^ n3769 ;
  assign n3771 = n3769 & ~n3770 ;
  assign n3773 = n3772 ^ n3771 ;
  assign n3774 = ~n3763 & ~n3773 ;
  assign n3775 = ~n3767 & n3774 ;
  assign n3776 = n3742 & ~n3743 ;
  assign n3777 = ~n2920 & ~n3776 ;
  assign n3778 = ~n3771 & n3777 ;
  assign n3779 = ~n3775 & n3778 ;
  assign n3780 = n3744 ^ n2917 ;
  assign n3781 = n3780 ^ n3776 ;
  assign n3782 = n2919 & n3781 ;
  assign n3783 = ~n3779 & ~n3782 ;
  assign n3784 = n3744 & ~n3783 ;
  assign n3785 = n3784 ^ n3743 ;
  assign n3741 = n3740 ^ n3658 ;
  assign n3786 = n3785 ^ n3741 ;
  assign n3788 = n3772 & n3783 ;
  assign n3789 = n3788 ^ n3769 ;
  assign n3787 = n3768 ^ n3707 ;
  assign n3790 = n3789 ^ n3787 ;
  assign n3792 = n3764 & ~n3783 ;
  assign n3793 = n3792 ^ n3762 ;
  assign n3791 = n3759 ^ n3711 ;
  assign n3794 = n3793 ^ n3791 ;
  assign n3795 = n3749 ^ n3745 ;
  assign n3796 = ~n3783 & n3795 ;
  assign n3797 = n3796 ^ n3745 ;
  assign n3798 = n3797 ^ n3747 ;
  assign n3799 = n3755 ^ n3751 ;
  assign n3800 = ~n3783 & n3799 ;
  assign n3801 = n3800 ^ n3751 ;
  assign n3802 = n3753 ^ n3721 ;
  assign n3803 = n3801 & ~n3802 ;
  assign n3804 = n3803 ^ n3747 ;
  assign n3805 = ~n3798 & ~n3804 ;
  assign n3806 = n3805 ^ n3747 ;
  assign n3807 = n3806 ^ n3793 ;
  assign n3808 = ~n3794 & ~n3807 ;
  assign n3809 = n3808 ^ n3793 ;
  assign n3810 = n3809 ^ n3787 ;
  assign n3811 = ~n3790 & ~n3810 ;
  assign n3812 = n3811 ^ n3787 ;
  assign n3813 = n3812 ^ n3741 ;
  assign n3814 = ~n3786 & ~n3813 ;
  assign n3815 = n3814 ^ n3785 ;
  assign n3816 = n3815 ^ n2750 ;
  assign n3817 = n2925 & n3816 ;
  assign n3818 = n3817 ^ n2921 ;
  assign n3819 = n3786 & n3818 ;
  assign n3821 = n3819 ^ n3785 ;
  assign n3823 = n3822 ^ n3821 ;
  assign n3824 = n1538 ^ n1535 ;
  assign n3825 = n3798 & ~n3818 ;
  assign n3826 = n3825 ^ n3798 ;
  assign n3827 = n3826 ^ n3797 ;
  assign n3828 = n3824 & ~n3827 ;
  assign n3829 = n1537 ^ n1536 ;
  assign n3830 = n3802 ^ n3801 ;
  assign n3831 = ~n3818 & n3830 ;
  assign n3832 = n3831 ^ n3830 ;
  assign n3833 = n3832 ^ n3801 ;
  assign n3834 = n3829 & ~n3833 ;
  assign n3835 = ~n3828 & ~n3834 ;
  assign n3836 = ~n1535 & n3827 ;
  assign n3840 = n1540 ^ n1539 ;
  assign n3837 = n3794 & n3818 ;
  assign n3838 = n3837 ^ n3794 ;
  assign n3839 = n3838 ^ n3791 ;
  assign n3842 = n3840 ^ n3839 ;
  assign n3841 = ~n3839 & n3840 ;
  assign n3843 = n3842 ^ n3841 ;
  assign n3844 = ~n3836 & ~n3843 ;
  assign n3845 = ~n3835 & n3844 ;
  assign n3847 = n3790 & n3818 ;
  assign n3848 = n3847 ^ n3789 ;
  assign n3846 = n1541 ^ n1534 ;
  assign n3850 = n3848 ^ n3846 ;
  assign n3849 = ~n3846 & n3848 ;
  assign n3851 = n3850 ^ n3849 ;
  assign n3852 = ~n3841 & ~n3851 ;
  assign n3853 = ~n3845 & n3852 ;
  assign n3854 = n3821 & ~n3822 ;
  assign n3855 = ~n2923 & ~n3854 ;
  assign n3856 = ~n3849 & n3855 ;
  assign n3857 = ~n3853 & n3856 ;
  assign n3858 = n3823 ^ n1546 ;
  assign n3859 = n3858 ^ n3854 ;
  assign n3860 = n2922 & n3859 ;
  assign n3861 = ~n3857 & ~n3860 ;
  assign n3862 = n3823 & ~n3861 ;
  assign n3863 = n3862 ^ n3822 ;
  assign n3820 = n3819 ^ n3741 ;
  assign n3864 = n3863 ^ n3820 ;
  assign n3866 = n3850 & n3861 ;
  assign n3867 = n3866 ^ n3848 ;
  assign n3865 = n3847 ^ n3787 ;
  assign n3868 = n3867 ^ n3865 ;
  assign n3870 = n3842 & ~n3861 ;
  assign n3871 = n3870 ^ n3840 ;
  assign n3869 = n3837 ^ n3791 ;
  assign n3872 = n3871 ^ n3869 ;
  assign n3876 = n3825 ^ n3797 ;
  assign n3873 = n3827 ^ n3824 ;
  assign n3874 = ~n3861 & n3873 ;
  assign n3875 = n3874 ^ n3824 ;
  assign n3877 = n3876 ^ n3875 ;
  assign n3878 = n3833 ^ n3829 ;
  assign n3879 = ~n3861 & n3878 ;
  assign n3880 = n3879 ^ n3829 ;
  assign n3881 = n3831 ^ n3801 ;
  assign n3882 = n3880 & ~n3881 ;
  assign n3883 = n3882 ^ n3876 ;
  assign n3884 = ~n3877 & ~n3883 ;
  assign n3885 = n3884 ^ n3876 ;
  assign n3886 = n3885 ^ n3871 ;
  assign n3887 = ~n3872 & ~n3886 ;
  assign n3888 = n3887 ^ n3871 ;
  assign n3889 = n3888 ^ n3867 ;
  assign n3890 = ~n3868 & n3889 ;
  assign n3891 = n3890 ^ n3867 ;
  assign n3892 = n3891 ^ n3863 ;
  assign n3893 = ~n3864 & n3892 ;
  assign n3894 = n3893 ^ n3863 ;
  assign n3895 = n3894 ^ n2926 ;
  assign n3896 = ~n2928 & ~n3895 ;
  assign n3897 = n3896 ^ n3894 ;
  assign n3898 = n3864 & ~n3897 ;
  assign n3900 = n3898 ^ n3863 ;
  assign n3902 = n3901 ^ n3900 ;
  assign n3903 = n1371 ^ n1368 ;
  assign n3904 = n3877 & n3897 ;
  assign n3905 = n3904 ^ n3875 ;
  assign n3906 = n3905 ^ n3876 ;
  assign n3907 = n3906 ^ n3875 ;
  assign n3908 = n3903 & ~n3907 ;
  assign n3909 = n1370 ^ n1369 ;
  assign n3910 = n3881 ^ n3880 ;
  assign n3911 = n3897 & n3910 ;
  assign n3912 = n3911 ^ n3910 ;
  assign n3913 = n3912 ^ n3880 ;
  assign n3914 = n3909 & ~n3913 ;
  assign n3915 = ~n3908 & ~n3914 ;
  assign n3916 = ~n1368 & n3907 ;
  assign n3920 = n1373 ^ n1372 ;
  assign n3917 = n3872 & ~n3897 ;
  assign n3918 = n3917 ^ n3872 ;
  assign n3919 = n3918 ^ n3869 ;
  assign n3922 = n3920 ^ n3919 ;
  assign n3921 = ~n3919 & n3920 ;
  assign n3923 = n3922 ^ n3921 ;
  assign n3924 = ~n3916 & ~n3923 ;
  assign n3925 = ~n3915 & n3924 ;
  assign n3927 = n3868 & ~n3897 ;
  assign n3928 = n3927 ^ n3867 ;
  assign n3926 = n1374 ^ n1367 ;
  assign n3930 = n3928 ^ n3926 ;
  assign n3929 = ~n3926 & n3928 ;
  assign n3931 = n3930 ^ n3929 ;
  assign n3932 = ~n3921 & ~n3931 ;
  assign n3933 = ~n3925 & n3932 ;
  assign n3934 = n3900 & ~n3901 ;
  assign n3935 = ~n2931 & ~n3934 ;
  assign n3936 = ~n3929 & n3935 ;
  assign n3937 = ~n3933 & n3936 ;
  assign n3938 = n3902 ^ n1379 ;
  assign n3939 = n3938 ^ n3934 ;
  assign n3940 = ~n2930 & n3939 ;
  assign n3941 = ~n3937 & ~n3940 ;
  assign n3942 = n3902 & ~n3941 ;
  assign n3943 = n3942 ^ n3901 ;
  assign n3899 = n3898 ^ n3820 ;
  assign n3944 = n3943 ^ n3899 ;
  assign n3945 = n2933 ^ n2932 ;
  assign n3946 = n3899 & ~n3943 ;
  assign n3947 = n3946 ^ n3944 ;
  assign n3949 = n3930 & n3941 ;
  assign n3950 = n3949 ^ n3928 ;
  assign n3948 = n3927 ^ n3865 ;
  assign n3951 = n3950 ^ n3948 ;
  assign n3953 = n3922 & ~n3941 ;
  assign n3954 = n3953 ^ n3920 ;
  assign n3952 = n3917 ^ n3869 ;
  assign n3955 = n3954 ^ n3952 ;
  assign n3956 = n3907 ^ n3903 ;
  assign n3957 = ~n3941 & n3956 ;
  assign n3958 = n3957 ^ n3903 ;
  assign n3959 = n3958 ^ n3905 ;
  assign n3960 = n3913 ^ n3909 ;
  assign n3961 = ~n3941 & n3960 ;
  assign n3962 = n3961 ^ n3909 ;
  assign n3963 = n3911 ^ n3880 ;
  assign n3964 = n3962 & ~n3963 ;
  assign n3965 = n3964 ^ n3905 ;
  assign n3966 = ~n3959 & ~n3965 ;
  assign n3967 = n3966 ^ n3905 ;
  assign n3968 = n3967 ^ n3954 ;
  assign n3969 = ~n3955 & ~n3968 ;
  assign n3970 = n3969 ^ n3954 ;
  assign n3971 = n3970 ^ n3950 ;
  assign n3972 = ~n3951 & n3971 ;
  assign n3973 = n3972 ^ n3950 ;
  assign n3974 = ~n3947 & ~n3973 ;
  assign n3975 = n3974 ^ n2933 ;
  assign n3976 = n3975 ^ n2933 ;
  assign n3977 = ~n3946 & ~n3976 ;
  assign n3978 = n3977 ^ n2933 ;
  assign n3979 = n3945 & ~n3978 ;
  assign n3980 = n3979 ^ n2932 ;
  assign n3981 = n3944 & ~n3980 ;
  assign n3983 = n3981 ^ n3943 ;
  assign n3985 = n3984 ^ n3983 ;
  assign n3986 = n3094 ^ n3091 ;
  assign n3987 = n3959 & n3980 ;
  assign n3988 = n3987 ^ n3958 ;
  assign n3989 = n3988 ^ n3905 ;
  assign n3990 = n3989 ^ n3958 ;
  assign n3991 = n3986 & ~n3990 ;
  assign n3992 = n3093 ^ n3092 ;
  assign n3993 = n3963 ^ n3962 ;
  assign n3994 = n3980 & n3993 ;
  assign n3995 = n3994 ^ n3993 ;
  assign n3996 = n3995 ^ n3962 ;
  assign n3997 = n3992 & ~n3996 ;
  assign n3998 = ~n3991 & ~n3997 ;
  assign n3999 = ~n3091 & n3990 ;
  assign n4003 = n3096 ^ n3095 ;
  assign n4000 = n3955 & ~n3980 ;
  assign n4001 = n4000 ^ n3955 ;
  assign n4002 = n4001 ^ n3952 ;
  assign n4005 = n4003 ^ n4002 ;
  assign n4004 = ~n4002 & n4003 ;
  assign n4006 = n4005 ^ n4004 ;
  assign n4007 = ~n3999 & ~n4006 ;
  assign n4008 = ~n3998 & n4007 ;
  assign n4011 = n3097 ^ n3090 ;
  assign n4009 = n3951 & ~n3980 ;
  assign n4010 = n4009 ^ n3950 ;
  assign n4013 = n4011 ^ n4010 ;
  assign n4012 = n4010 & ~n4011 ;
  assign n4014 = n4013 ^ n4012 ;
  assign n4015 = ~n4004 & ~n4014 ;
  assign n4016 = ~n4008 & n4015 ;
  assign n4017 = n3983 & ~n3984 ;
  assign n4018 = ~n3105 & ~n4017 ;
  assign n4019 = ~n4012 & n4018 ;
  assign n4020 = ~n4016 & n4019 ;
  assign n4021 = n3985 ^ n3102 ;
  assign n4022 = n4021 ^ n4017 ;
  assign n4023 = n3104 & n4022 ;
  assign n4024 = ~n4020 & ~n4023 ;
  assign n4025 = n3985 & ~n4024 ;
  assign n4026 = n4025 ^ n3984 ;
  assign n3982 = n3981 ^ n3899 ;
  assign n4027 = n4026 ^ n3982 ;
  assign n4029 = n4013 & n4024 ;
  assign n4030 = n4029 ^ n4010 ;
  assign n4028 = n4009 ^ n3948 ;
  assign n4031 = n4030 ^ n4028 ;
  assign n4033 = n4005 & ~n4024 ;
  assign n4034 = n4033 ^ n4003 ;
  assign n4032 = n4000 ^ n3952 ;
  assign n4035 = n4034 ^ n4032 ;
  assign n4036 = n3990 ^ n3986 ;
  assign n4037 = ~n4024 & n4036 ;
  assign n4038 = n4037 ^ n3986 ;
  assign n4039 = n4038 ^ n3988 ;
  assign n4040 = n3996 ^ n3992 ;
  assign n4041 = ~n4024 & n4040 ;
  assign n4042 = n4041 ^ n3992 ;
  assign n4043 = n3994 ^ n3962 ;
  assign n4044 = n4042 & ~n4043 ;
  assign n4045 = n4044 ^ n3988 ;
  assign n4046 = ~n4039 & ~n4045 ;
  assign n4047 = n4046 ^ n3988 ;
  assign n4048 = n4047 ^ n4034 ;
  assign n4049 = ~n4035 & ~n4048 ;
  assign n4050 = n4049 ^ n4034 ;
  assign n4051 = n4050 ^ n4028 ;
  assign n4052 = ~n4031 & ~n4051 ;
  assign n4053 = n4052 ^ n4028 ;
  assign n4054 = n4053 ^ n4026 ;
  assign n4055 = ~n4027 & n4054 ;
  assign n4056 = n4055 ^ n3982 ;
  assign n4057 = n4056 ^ n2935 ;
  assign n4058 = n3110 & ~n4057 ;
  assign n4059 = n4058 ^ n3106 ;
  assign n4060 = n4027 & n4059 ;
  assign n4062 = n4060 ^ n4026 ;
  assign n4064 = n4063 ^ n4062 ;
  assign n4065 = n1204 ^ n1201 ;
  assign n4066 = n4039 & ~n4059 ;
  assign n4067 = n4066 ^ n4039 ;
  assign n4068 = n4067 ^ n4038 ;
  assign n4069 = n4065 & ~n4068 ;
  assign n4070 = n1203 ^ n1202 ;
  assign n4071 = n4043 ^ n4042 ;
  assign n4072 = ~n4059 & n4071 ;
  assign n4073 = n4072 ^ n4071 ;
  assign n4074 = n4073 ^ n4042 ;
  assign n4075 = n4070 & ~n4074 ;
  assign n4076 = ~n4069 & ~n4075 ;
  assign n4077 = ~n1201 & n4068 ;
  assign n4081 = n1206 ^ n1205 ;
  assign n4078 = n4035 & n4059 ;
  assign n4079 = n4078 ^ n4035 ;
  assign n4080 = n4079 ^ n4032 ;
  assign n4083 = n4081 ^ n4080 ;
  assign n4082 = ~n4080 & n4081 ;
  assign n4084 = n4083 ^ n4082 ;
  assign n4085 = ~n4077 & ~n4084 ;
  assign n4086 = ~n4076 & n4085 ;
  assign n4088 = n4031 & n4059 ;
  assign n4089 = n4088 ^ n4030 ;
  assign n4087 = n1207 ^ n1200 ;
  assign n4091 = n4089 ^ n4087 ;
  assign n4090 = ~n4087 & n4089 ;
  assign n4092 = n4091 ^ n4090 ;
  assign n4093 = ~n4082 & ~n4092 ;
  assign n4094 = ~n4086 & n4093 ;
  assign n4095 = n4062 & ~n4063 ;
  assign n4096 = ~n3108 & ~n4095 ;
  assign n4097 = ~n4090 & n4096 ;
  assign n4098 = ~n4094 & n4097 ;
  assign n4099 = n4064 ^ n1212 ;
  assign n4100 = n4099 ^ n4095 ;
  assign n4101 = n3107 & n4100 ;
  assign n4102 = ~n4098 & ~n4101 ;
  assign n4103 = n4064 & ~n4102 ;
  assign n4104 = n4103 ^ n4063 ;
  assign n4061 = n4060 ^ n3982 ;
  assign n4105 = n4104 ^ n4061 ;
  assign n4107 = n4091 & n4102 ;
  assign n4108 = n4107 ^ n4089 ;
  assign n4106 = n4088 ^ n4028 ;
  assign n4109 = n4108 ^ n4106 ;
  assign n4111 = n4083 & ~n4102 ;
  assign n4112 = n4111 ^ n4081 ;
  assign n4110 = n4078 ^ n4032 ;
  assign n4113 = n4112 ^ n4110 ;
  assign n4117 = n4066 ^ n4038 ;
  assign n4114 = n4068 ^ n4065 ;
  assign n4115 = ~n4102 & n4114 ;
  assign n4116 = n4115 ^ n4065 ;
  assign n4118 = n4117 ^ n4116 ;
  assign n4119 = n4074 ^ n4070 ;
  assign n4120 = ~n4102 & n4119 ;
  assign n4121 = n4120 ^ n4070 ;
  assign n4122 = n4072 ^ n4042 ;
  assign n4123 = n4121 & ~n4122 ;
  assign n4124 = n4123 ^ n4117 ;
  assign n4125 = ~n4118 & ~n4124 ;
  assign n4126 = n4125 ^ n4117 ;
  assign n4127 = n4126 ^ n4112 ;
  assign n4128 = ~n4113 & ~n4127 ;
  assign n4129 = n4128 ^ n4112 ;
  assign n4130 = n4129 ^ n4108 ;
  assign n4131 = ~n4109 & n4130 ;
  assign n4132 = n4131 ^ n4108 ;
  assign n4133 = n4132 ^ n4104 ;
  assign n4134 = ~n4105 & n4133 ;
  assign n4135 = n4134 ^ n4104 ;
  assign n4136 = n4135 ^ n3111 ;
  assign n4137 = ~n3113 & ~n4136 ;
  assign n4138 = n4137 ^ n4135 ;
  assign n4139 = n4105 & ~n4138 ;
  assign n4141 = n4139 ^ n4104 ;
  assign n4143 = n4142 ^ n4141 ;
  assign n4144 = n1037 ^ n1034 ;
  assign n4145 = n4118 & n4138 ;
  assign n4146 = n4145 ^ n4116 ;
  assign n4147 = n4146 ^ n4117 ;
  assign n4148 = n4147 ^ n4116 ;
  assign n4149 = n4144 & ~n4148 ;
  assign n4150 = n1036 ^ n1035 ;
  assign n4151 = n4122 ^ n4121 ;
  assign n4152 = n4138 & n4151 ;
  assign n4153 = n4152 ^ n4151 ;
  assign n4154 = n4153 ^ n4121 ;
  assign n4155 = n4150 & ~n4154 ;
  assign n4156 = ~n4149 & ~n4155 ;
  assign n4157 = ~n1034 & n4148 ;
  assign n4161 = n1039 ^ n1038 ;
  assign n4158 = n4113 & ~n4138 ;
  assign n4159 = n4158 ^ n4113 ;
  assign n4160 = n4159 ^ n4110 ;
  assign n4163 = n4161 ^ n4160 ;
  assign n4162 = ~n4160 & n4161 ;
  assign n4164 = n4163 ^ n4162 ;
  assign n4165 = ~n4157 & ~n4164 ;
  assign n4166 = ~n4156 & n4165 ;
  assign n4168 = n4109 & ~n4138 ;
  assign n4169 = n4168 ^ n4108 ;
  assign n4167 = n1040 ^ n1033 ;
  assign n4171 = n4169 ^ n4167 ;
  assign n4170 = ~n4167 & n4169 ;
  assign n4172 = n4171 ^ n4170 ;
  assign n4173 = ~n4162 & ~n4172 ;
  assign n4174 = ~n4166 & n4173 ;
  assign n4175 = n4141 & ~n4142 ;
  assign n4176 = ~n3116 & ~n4175 ;
  assign n4177 = ~n4170 & n4176 ;
  assign n4178 = ~n4174 & n4177 ;
  assign n4179 = n4143 ^ n1045 ;
  assign n4180 = n4179 ^ n4175 ;
  assign n4181 = ~n3115 & n4180 ;
  assign n4182 = ~n4178 & ~n4181 ;
  assign n4183 = n4143 & ~n4182 ;
  assign n4184 = n4183 ^ n4142 ;
  assign n4140 = n4139 ^ n4061 ;
  assign n4185 = n4184 ^ n4140 ;
  assign n4186 = n3118 ^ n3117 ;
  assign n4187 = n4140 & ~n4184 ;
  assign n4188 = n4187 ^ n4185 ;
  assign n4190 = n4171 & n4182 ;
  assign n4191 = n4190 ^ n4169 ;
  assign n4189 = n4168 ^ n4106 ;
  assign n4192 = n4191 ^ n4189 ;
  assign n4194 = n4163 & ~n4182 ;
  assign n4195 = n4194 ^ n4161 ;
  assign n4193 = n4158 ^ n4110 ;
  assign n4196 = n4195 ^ n4193 ;
  assign n4197 = n4148 ^ n4144 ;
  assign n4198 = ~n4182 & n4197 ;
  assign n4199 = n4198 ^ n4144 ;
  assign n4200 = n4199 ^ n4146 ;
  assign n4201 = n4154 ^ n4150 ;
  assign n4202 = ~n4182 & n4201 ;
  assign n4203 = n4202 ^ n4150 ;
  assign n4204 = n4152 ^ n4121 ;
  assign n4205 = n4203 & ~n4204 ;
  assign n4206 = n4205 ^ n4146 ;
  assign n4207 = ~n4200 & ~n4206 ;
  assign n4208 = n4207 ^ n4146 ;
  assign n4209 = n4208 ^ n4195 ;
  assign n4210 = ~n4196 & ~n4209 ;
  assign n4211 = n4210 ^ n4195 ;
  assign n4212 = n4211 ^ n4191 ;
  assign n4213 = ~n4192 & n4212 ;
  assign n4214 = n4213 ^ n4191 ;
  assign n4215 = ~n4188 & ~n4214 ;
  assign n4216 = n4215 ^ n3118 ;
  assign n4217 = n4216 ^ n3118 ;
  assign n4218 = ~n4187 & ~n4217 ;
  assign n4219 = n4218 ^ n3118 ;
  assign n4220 = n4186 & ~n4219 ;
  assign n4221 = n4220 ^ n3117 ;
  assign n4222 = n4185 & ~n4221 ;
  assign n4224 = n4222 ^ n4184 ;
  assign n4226 = n4225 ^ n4224 ;
  assign n4227 = n870 ^ n867 ;
  assign n4228 = n4200 & n4221 ;
  assign n4229 = n4228 ^ n4199 ;
  assign n4230 = n4229 ^ n4146 ;
  assign n4231 = n4230 ^ n4199 ;
  assign n4232 = n4227 & ~n4231 ;
  assign n4233 = n869 ^ n868 ;
  assign n4234 = n4204 ^ n4203 ;
  assign n4235 = n4221 & n4234 ;
  assign n4236 = n4235 ^ n4234 ;
  assign n4237 = n4236 ^ n4203 ;
  assign n4238 = n4233 & ~n4237 ;
  assign n4239 = ~n4232 & ~n4238 ;
  assign n4240 = ~n867 & n4231 ;
  assign n4244 = n872 ^ n871 ;
  assign n4241 = n4196 & ~n4221 ;
  assign n4242 = n4241 ^ n4196 ;
  assign n4243 = n4242 ^ n4193 ;
  assign n4246 = n4244 ^ n4243 ;
  assign n4245 = ~n4243 & n4244 ;
  assign n4247 = n4246 ^ n4245 ;
  assign n4248 = ~n4240 & ~n4247 ;
  assign n4249 = ~n4239 & n4248 ;
  assign n4252 = n873 ^ n866 ;
  assign n4250 = n4192 & ~n4221 ;
  assign n4251 = n4250 ^ n4191 ;
  assign n4254 = n4252 ^ n4251 ;
  assign n4253 = n4251 & ~n4252 ;
  assign n4255 = n4254 ^ n4253 ;
  assign n4256 = ~n4245 & ~n4255 ;
  assign n4257 = ~n4249 & n4256 ;
  assign n4258 = n4224 & ~n4225 ;
  assign n4259 = ~n3123 & ~n4258 ;
  assign n4260 = ~n4253 & n4259 ;
  assign n4261 = ~n4257 & n4260 ;
  assign n4262 = n4226 ^ n878 ;
  assign n4263 = n4262 ^ n4258 ;
  assign n4264 = n3122 & n4263 ;
  assign n4265 = ~n4261 & ~n4264 ;
  assign n4266 = n4226 & ~n4265 ;
  assign n4267 = n4266 ^ n4225 ;
  assign n4223 = n4222 ^ n4140 ;
  assign n4268 = n4267 ^ n4223 ;
  assign n4270 = n4254 & n4265 ;
  assign n4271 = n4270 ^ n4251 ;
  assign n4269 = n4250 ^ n4189 ;
  assign n4272 = n4271 ^ n4269 ;
  assign n4274 = n4246 & ~n4265 ;
  assign n4275 = n4274 ^ n4244 ;
  assign n4273 = n4241 ^ n4193 ;
  assign n4276 = n4275 ^ n4273 ;
  assign n4277 = n4231 ^ n4227 ;
  assign n4278 = ~n4265 & n4277 ;
  assign n4279 = n4278 ^ n4227 ;
  assign n4280 = n4279 ^ n4229 ;
  assign n4281 = n4237 ^ n4233 ;
  assign n4282 = ~n4265 & n4281 ;
  assign n4283 = n4282 ^ n4233 ;
  assign n4284 = n4235 ^ n4203 ;
  assign n4285 = n4283 & ~n4284 ;
  assign n4286 = n4285 ^ n4229 ;
  assign n4287 = ~n4280 & ~n4286 ;
  assign n4288 = n4287 ^ n4229 ;
  assign n4289 = n4288 ^ n4275 ;
  assign n4290 = ~n4276 & ~n4289 ;
  assign n4291 = n4290 ^ n4275 ;
  assign n4292 = n4291 ^ n4269 ;
  assign n4293 = ~n4272 & ~n4292 ;
  assign n4294 = n4293 ^ n4269 ;
  assign n4295 = n4294 ^ n4223 ;
  assign n4296 = ~n4268 & ~n4295 ;
  assign n4297 = n4296 ^ n4267 ;
  assign n4298 = n4297 ^ n3120 ;
  assign n4299 = n3125 & n4298 ;
  assign n4300 = n4299 ^ n3124 ;
  assign n4301 = n4268 & n4300 ;
  assign n4303 = n4301 ^ n4267 ;
  assign n4305 = n4304 ^ n4303 ;
  assign n4306 = n3286 ^ n3283 ;
  assign n4307 = n4280 & ~n4300 ;
  assign n4308 = n4307 ^ n4280 ;
  assign n4309 = n4308 ^ n4279 ;
  assign n4310 = n4306 & ~n4309 ;
  assign n4311 = n3285 ^ n3284 ;
  assign n4312 = n4284 ^ n4283 ;
  assign n4313 = ~n4300 & n4312 ;
  assign n4314 = n4313 ^ n4312 ;
  assign n4315 = n4314 ^ n4283 ;
  assign n4316 = n4311 & ~n4315 ;
  assign n4317 = ~n4310 & ~n4316 ;
  assign n4318 = ~n3283 & n4309 ;
  assign n4322 = n3288 ^ n3287 ;
  assign n4319 = n4276 & n4300 ;
  assign n4320 = n4319 ^ n4276 ;
  assign n4321 = n4320 ^ n4273 ;
  assign n4324 = n4322 ^ n4321 ;
  assign n4323 = ~n4321 & n4322 ;
  assign n4325 = n4324 ^ n4323 ;
  assign n4326 = ~n4318 & ~n4325 ;
  assign n4327 = ~n4317 & n4326 ;
  assign n4329 = n4272 & n4300 ;
  assign n4330 = n4329 ^ n4271 ;
  assign n4328 = n3289 ^ n3282 ;
  assign n4332 = n4330 ^ n4328 ;
  assign n4331 = ~n4328 & n4330 ;
  assign n4333 = n4332 ^ n4331 ;
  assign n4334 = ~n4323 & ~n4333 ;
  assign n4335 = ~n4327 & n4334 ;
  assign n4336 = n4303 & ~n4304 ;
  assign n4337 = ~n3295 & ~n4336 ;
  assign n4338 = ~n4331 & n4337 ;
  assign n4339 = ~n4335 & n4338 ;
  assign n4340 = n4305 ^ n3294 ;
  assign n4341 = n4340 ^ n4336 ;
  assign n4342 = n3126 & n4341 ;
  assign n4343 = ~n4339 & ~n4342 ;
  assign n4344 = n4305 & ~n4343 ;
  assign n4345 = n4344 ^ n4304 ;
  assign n4302 = n4301 ^ n4223 ;
  assign n4346 = n4345 ^ n4302 ;
  assign n4348 = n4332 & n4343 ;
  assign n4349 = n4348 ^ n4330 ;
  assign n4347 = n4329 ^ n4269 ;
  assign n4350 = n4349 ^ n4347 ;
  assign n4352 = n4324 & ~n4343 ;
  assign n4353 = n4352 ^ n4322 ;
  assign n4351 = n4319 ^ n4273 ;
  assign n4354 = n4353 ^ n4351 ;
  assign n4358 = n4307 ^ n4279 ;
  assign n4355 = n4309 ^ n4306 ;
  assign n4356 = ~n4343 & n4355 ;
  assign n4357 = n4356 ^ n4306 ;
  assign n4359 = n4358 ^ n4357 ;
  assign n4360 = n4315 ^ n4311 ;
  assign n4361 = ~n4343 & n4360 ;
  assign n4362 = n4361 ^ n4311 ;
  assign n4363 = n4313 ^ n4283 ;
  assign n4364 = n4362 & ~n4363 ;
  assign n4365 = n4364 ^ n4358 ;
  assign n4366 = ~n4359 & ~n4365 ;
  assign n4367 = n4366 ^ n4358 ;
  assign n4368 = n4367 ^ n4353 ;
  assign n4369 = ~n4354 & ~n4368 ;
  assign n4370 = n4369 ^ n4353 ;
  assign n4371 = n4370 ^ n4349 ;
  assign n4372 = ~n4350 & n4371 ;
  assign n4373 = n4372 ^ n4349 ;
  assign n4374 = n4373 ^ n4345 ;
  assign n4375 = ~n4346 & n4374 ;
  assign n4376 = n4375 ^ n4345 ;
  assign n4377 = n4376 ^ n3296 ;
  assign n4378 = ~n3298 & ~n4377 ;
  assign n4379 = n4378 ^ n4376 ;
  assign n4380 = n4346 & ~n4379 ;
  assign n4383 = n4380 ^ n4345 ;
  assign n4382 = n710 ^ n707 ;
  assign n4384 = n4383 ^ n4382 ;
  assign n4385 = n703 ^ n700 ;
  assign n4386 = n4359 & n4379 ;
  assign n4387 = n4386 ^ n4357 ;
  assign n4388 = n4387 ^ n4358 ;
  assign n4389 = n4388 ^ n4357 ;
  assign n4390 = n4385 & ~n4389 ;
  assign n4391 = n702 ^ n701 ;
  assign n4392 = n4363 ^ n4362 ;
  assign n4393 = n4379 & n4392 ;
  assign n4394 = n4393 ^ n4392 ;
  assign n4395 = n4394 ^ n4362 ;
  assign n4396 = n4391 & ~n4395 ;
  assign n4397 = ~n4390 & ~n4396 ;
  assign n4398 = ~n700 & n4389 ;
  assign n4402 = n705 ^ n704 ;
  assign n4399 = n4354 & ~n4379 ;
  assign n4400 = n4399 ^ n4354 ;
  assign n4401 = n4400 ^ n4351 ;
  assign n4404 = n4402 ^ n4401 ;
  assign n4403 = ~n4401 & n4402 ;
  assign n4405 = n4404 ^ n4403 ;
  assign n4406 = ~n4398 & ~n4405 ;
  assign n4407 = ~n4397 & n4406 ;
  assign n4410 = n706 ^ n699 ;
  assign n4408 = n4350 & ~n4379 ;
  assign n4409 = n4408 ^ n4349 ;
  assign n4412 = n4410 ^ n4409 ;
  assign n4411 = n4409 & ~n4410 ;
  assign n4413 = n4412 ^ n4411 ;
  assign n4414 = ~n4403 & ~n4413 ;
  assign n4415 = ~n4407 & n4414 ;
  assign n4416 = ~n4382 & n4383 ;
  assign n4417 = n3299 ^ n3296 ;
  assign n4418 = ~n711 & n4417 ;
  assign n4419 = ~n4416 & ~n4418 ;
  assign n4420 = ~n4411 & n4419 ;
  assign n4421 = ~n4415 & n4420 ;
  assign n4422 = n4384 ^ n711 ;
  assign n4423 = n4422 ^ n4416 ;
  assign n4424 = ~n4417 & n4423 ;
  assign n4425 = ~n4421 & ~n4424 ;
  assign n4426 = n4384 & n4425 ;
  assign n4427 = n4426 ^ n4383 ;
  assign n4381 = n4380 ^ n4302 ;
  assign n4428 = n4427 ^ n4381 ;
  assign n4430 = n4412 & ~n4425 ;
  assign n4431 = n4430 ^ n4410 ;
  assign n4429 = n4408 ^ n4347 ;
  assign n4432 = n4431 ^ n4429 ;
  assign n4442 = n4389 ^ n4385 ;
  assign n4443 = ~n4425 & n4442 ;
  assign n4444 = n4443 ^ n4385 ;
  assign n4437 = n4393 ^ n4362 ;
  assign n4438 = n4395 ^ n4391 ;
  assign n4439 = n4425 & n4438 ;
  assign n4440 = n4439 ^ n4395 ;
  assign n4441 = ~n4437 & n4440 ;
  assign n4445 = n4444 ^ n4441 ;
  assign n4446 = n4441 ^ n4387 ;
  assign n4447 = n4445 & ~n4446 ;
  assign n4448 = n4447 ^ n4441 ;
  assign n4451 = n4448 ^ n4431 ;
  assign n4434 = n4404 & ~n4425 ;
  assign n4435 = n4434 ^ n4402 ;
  assign n4433 = n4399 ^ n4351 ;
  assign n4436 = n4435 ^ n4433 ;
  assign n4449 = n4448 ^ n4435 ;
  assign n4450 = n4436 & n4449 ;
  assign n4452 = n4451 ^ n4450 ;
  assign n4453 = ~n4432 & ~n4452 ;
  assign n4454 = n4453 ^ n4429 ;
  assign n4455 = n4454 ^ n4427 ;
  assign n4456 = ~n4428 & ~n4455 ;
  assign n4457 = n4456 ^ n4427 ;
  assign n4458 = ~n3301 & n4457 ;
  assign n4459 = n4418 ^ n3298 ;
  assign n4460 = n4459 ^ n3301 ;
  assign n4461 = ~n4458 & n4460 ;
  assign n4462 = x480 ^ x448 ;
  assign n4463 = ~n3330 & n4462 ;
  assign n4466 = n4463 ^ x448 ;
  assign n4467 = n4466 ^ x416 ;
  assign n4468 = ~n3377 & n4467 ;
  assign n4469 = n4468 ^ x416 ;
  assign n4464 = n4463 ^ n4462 ;
  assign n4465 = n4464 ^ x448 ;
  assign n4470 = n4469 ^ n4465 ;
  assign n4471 = ~n3413 & n4470 ;
  assign n4474 = n4471 ^ n4465 ;
  assign n4475 = n4474 ^ x384 ;
  assign n4476 = ~n3457 & n4475 ;
  assign n4477 = n4476 ^ x384 ;
  assign n4472 = n4471 ^ n4470 ;
  assign n4473 = n4472 ^ n4465 ;
  assign n4478 = n4477 ^ n4473 ;
  assign n4479 = ~n3493 & n4478 ;
  assign n4482 = n4479 ^ n4473 ;
  assign n4483 = n4482 ^ x352 ;
  assign n4484 = ~n3537 & n4483 ;
  assign n4485 = n4484 ^ x352 ;
  assign n4480 = n4479 ^ n4478 ;
  assign n4481 = n4480 ^ n4473 ;
  assign n4486 = n4485 ^ n4481 ;
  assign n4487 = n3577 & n4486 ;
  assign n4490 = n4487 ^ n4481 ;
  assign n4491 = n4490 ^ x320 ;
  assign n4492 = ~n3620 & n4491 ;
  assign n4493 = n4492 ^ x320 ;
  assign n4488 = n4487 ^ n4486 ;
  assign n4489 = n4488 ^ n4481 ;
  assign n4494 = n4493 ^ n4489 ;
  assign n4495 = n3656 & n4494 ;
  assign n4498 = n4495 ^ n4489 ;
  assign n4499 = n4498 ^ x288 ;
  assign n4500 = ~n3700 & n4499 ;
  assign n4501 = n4500 ^ x288 ;
  assign n4496 = n4495 ^ n4494 ;
  assign n4497 = n4496 ^ n4489 ;
  assign n4502 = n4501 ^ n4497 ;
  assign n4503 = n3739 & n4502 ;
  assign n4506 = n4503 ^ n4497 ;
  assign n4507 = n4506 ^ x256 ;
  assign n4508 = ~n3783 & n4507 ;
  assign n4509 = n4508 ^ x256 ;
  assign n4504 = n4503 ^ n4502 ;
  assign n4505 = n4504 ^ n4497 ;
  assign n4510 = n4509 ^ n4505 ;
  assign n4511 = ~n3818 & n4510 ;
  assign n4514 = n4511 ^ n4505 ;
  assign n4515 = n4514 ^ x224 ;
  assign n4516 = ~n3861 & n4515 ;
  assign n4517 = n4516 ^ x224 ;
  assign n4512 = n4511 ^ n4510 ;
  assign n4513 = n4512 ^ n4505 ;
  assign n4518 = n4517 ^ n4513 ;
  assign n4519 = n3897 & n4518 ;
  assign n4522 = n4519 ^ n4513 ;
  assign n4523 = n4522 ^ x192 ;
  assign n4524 = ~n3941 & n4523 ;
  assign n4525 = n4524 ^ x192 ;
  assign n4520 = n4519 ^ n4518 ;
  assign n4521 = n4520 ^ n4513 ;
  assign n4526 = n4525 ^ n4521 ;
  assign n4527 = n3980 & n4526 ;
  assign n4530 = n4527 ^ n4521 ;
  assign n4531 = n4530 ^ x160 ;
  assign n4532 = ~n4024 & n4531 ;
  assign n4533 = n4532 ^ x160 ;
  assign n4528 = n4527 ^ n4526 ;
  assign n4529 = n4528 ^ n4521 ;
  assign n4534 = n4533 ^ n4529 ;
  assign n4535 = ~n4059 & n4534 ;
  assign n4538 = n4535 ^ n4529 ;
  assign n4539 = n4538 ^ x128 ;
  assign n4540 = ~n4102 & n4539 ;
  assign n4541 = n4540 ^ x128 ;
  assign n4536 = n4535 ^ n4534 ;
  assign n4537 = n4536 ^ n4529 ;
  assign n4542 = n4541 ^ n4537 ;
  assign n4543 = n4138 & n4542 ;
  assign n4546 = n4543 ^ n4537 ;
  assign n4547 = n4546 ^ x96 ;
  assign n4548 = ~n4182 & n4547 ;
  assign n4549 = n4548 ^ x96 ;
  assign n4544 = n4543 ^ n4542 ;
  assign n4545 = n4544 ^ n4537 ;
  assign n4550 = n4549 ^ n4545 ;
  assign n4551 = n4221 & n4550 ;
  assign n4554 = n4551 ^ n4545 ;
  assign n4555 = n4554 ^ x64 ;
  assign n4556 = ~n4265 & n4555 ;
  assign n4557 = n4556 ^ x64 ;
  assign n4552 = n4551 ^ n4550 ;
  assign n4553 = n4552 ^ n4545 ;
  assign n4558 = n4557 ^ n4553 ;
  assign n4559 = ~n4300 & n4558 ;
  assign n4562 = n4559 ^ n4553 ;
  assign n4563 = n4562 ^ x32 ;
  assign n4564 = ~n4343 & n4563 ;
  assign n4565 = n4564 ^ x32 ;
  assign n4560 = n4559 ^ n4558 ;
  assign n4561 = n4560 ^ n4553 ;
  assign n4566 = n4565 ^ n4561 ;
  assign n4567 = n4379 & n4566 ;
  assign n4570 = n4567 ^ n4561 ;
  assign n4571 = n4570 ^ x0 ;
  assign n4572 = ~n4425 & n4571 ;
  assign n4573 = n4572 ^ x0 ;
  assign n4568 = n4567 ^ n4566 ;
  assign n4569 = n4568 ^ n4561 ;
  assign n4574 = n4573 ^ n4569 ;
  assign n4575 = ~n4461 & n4574 ;
  assign n4576 = n4575 ^ n4574 ;
  assign n4577 = n4576 ^ n4569 ;
  assign n4578 = x481 ^ x449 ;
  assign n4579 = ~n3330 & n4578 ;
  assign n4582 = n4579 ^ x449 ;
  assign n4583 = n4582 ^ x417 ;
  assign n4584 = ~n3377 & n4583 ;
  assign n4585 = n4584 ^ x417 ;
  assign n4580 = n4579 ^ n4578 ;
  assign n4581 = n4580 ^ x449 ;
  assign n4586 = n4585 ^ n4581 ;
  assign n4587 = ~n3413 & n4586 ;
  assign n4590 = n4587 ^ n4581 ;
  assign n4591 = n4590 ^ x385 ;
  assign n4592 = ~n3457 & n4591 ;
  assign n4593 = n4592 ^ x385 ;
  assign n4588 = n4587 ^ n4586 ;
  assign n4589 = n4588 ^ n4581 ;
  assign n4594 = n4593 ^ n4589 ;
  assign n4595 = ~n3493 & n4594 ;
  assign n4598 = n4595 ^ n4589 ;
  assign n4599 = n4598 ^ x353 ;
  assign n4600 = ~n3537 & n4599 ;
  assign n4601 = n4600 ^ x353 ;
  assign n4596 = n4595 ^ n4594 ;
  assign n4597 = n4596 ^ n4589 ;
  assign n4602 = n4601 ^ n4597 ;
  assign n4603 = n3577 & n4602 ;
  assign n4606 = n4603 ^ n4597 ;
  assign n4607 = n4606 ^ x321 ;
  assign n4608 = ~n3620 & n4607 ;
  assign n4609 = n4608 ^ x321 ;
  assign n4604 = n4603 ^ n4602 ;
  assign n4605 = n4604 ^ n4597 ;
  assign n4610 = n4609 ^ n4605 ;
  assign n4611 = n3656 & n4610 ;
  assign n4614 = n4611 ^ n4605 ;
  assign n4615 = n4614 ^ x289 ;
  assign n4616 = ~n3700 & n4615 ;
  assign n4617 = n4616 ^ x289 ;
  assign n4612 = n4611 ^ n4610 ;
  assign n4613 = n4612 ^ n4605 ;
  assign n4618 = n4617 ^ n4613 ;
  assign n4619 = n3739 & n4618 ;
  assign n4622 = n4619 ^ n4613 ;
  assign n4623 = n4622 ^ x257 ;
  assign n4624 = ~n3783 & n4623 ;
  assign n4625 = n4624 ^ x257 ;
  assign n4620 = n4619 ^ n4618 ;
  assign n4621 = n4620 ^ n4613 ;
  assign n4626 = n4625 ^ n4621 ;
  assign n4627 = ~n3818 & n4626 ;
  assign n4630 = n4627 ^ n4621 ;
  assign n4631 = n4630 ^ x225 ;
  assign n4632 = ~n3861 & n4631 ;
  assign n4633 = n4632 ^ x225 ;
  assign n4628 = n4627 ^ n4626 ;
  assign n4629 = n4628 ^ n4621 ;
  assign n4634 = n4633 ^ n4629 ;
  assign n4635 = n3897 & n4634 ;
  assign n4638 = n4635 ^ n4629 ;
  assign n4639 = n4638 ^ x193 ;
  assign n4640 = ~n3941 & n4639 ;
  assign n4641 = n4640 ^ x193 ;
  assign n4636 = n4635 ^ n4634 ;
  assign n4637 = n4636 ^ n4629 ;
  assign n4642 = n4641 ^ n4637 ;
  assign n4643 = n3980 & n4642 ;
  assign n4646 = n4643 ^ n4637 ;
  assign n4647 = n4646 ^ x161 ;
  assign n4648 = ~n4024 & n4647 ;
  assign n4649 = n4648 ^ x161 ;
  assign n4644 = n4643 ^ n4642 ;
  assign n4645 = n4644 ^ n4637 ;
  assign n4650 = n4649 ^ n4645 ;
  assign n4651 = ~n4059 & n4650 ;
  assign n4654 = n4651 ^ n4645 ;
  assign n4655 = n4654 ^ x129 ;
  assign n4656 = ~n4102 & n4655 ;
  assign n4657 = n4656 ^ x129 ;
  assign n4652 = n4651 ^ n4650 ;
  assign n4653 = n4652 ^ n4645 ;
  assign n4658 = n4657 ^ n4653 ;
  assign n4659 = n4138 & n4658 ;
  assign n4662 = n4659 ^ n4653 ;
  assign n4663 = n4662 ^ x97 ;
  assign n4664 = ~n4182 & n4663 ;
  assign n4665 = n4664 ^ x97 ;
  assign n4660 = n4659 ^ n4658 ;
  assign n4661 = n4660 ^ n4653 ;
  assign n4666 = n4665 ^ n4661 ;
  assign n4667 = n4221 & n4666 ;
  assign n4670 = n4667 ^ n4661 ;
  assign n4671 = n4670 ^ x65 ;
  assign n4672 = ~n4265 & n4671 ;
  assign n4673 = n4672 ^ x65 ;
  assign n4668 = n4667 ^ n4666 ;
  assign n4669 = n4668 ^ n4661 ;
  assign n4674 = n4673 ^ n4669 ;
  assign n4675 = ~n4300 & n4674 ;
  assign n4678 = n4675 ^ n4669 ;
  assign n4679 = n4678 ^ x33 ;
  assign n4680 = ~n4343 & n4679 ;
  assign n4681 = n4680 ^ x33 ;
  assign n4676 = n4675 ^ n4674 ;
  assign n4677 = n4676 ^ n4669 ;
  assign n4682 = n4681 ^ n4677 ;
  assign n4683 = n4379 & n4682 ;
  assign n4686 = n4683 ^ n4677 ;
  assign n4687 = n4686 ^ x1 ;
  assign n4688 = ~n4425 & n4687 ;
  assign n4689 = n4688 ^ x1 ;
  assign n4684 = n4683 ^ n4682 ;
  assign n4685 = n4684 ^ n4677 ;
  assign n4690 = n4689 ^ n4685 ;
  assign n4691 = ~n4461 & n4690 ;
  assign n4692 = n4691 ^ n4690 ;
  assign n4693 = n4692 ^ n4685 ;
  assign n4694 = x482 ^ x450 ;
  assign n4695 = ~n3330 & n4694 ;
  assign n4698 = n4695 ^ x450 ;
  assign n4699 = n4698 ^ x418 ;
  assign n4700 = ~n3377 & n4699 ;
  assign n4701 = n4700 ^ x418 ;
  assign n4696 = n4695 ^ n4694 ;
  assign n4697 = n4696 ^ x450 ;
  assign n4702 = n4701 ^ n4697 ;
  assign n4703 = ~n3413 & n4702 ;
  assign n4706 = n4703 ^ n4697 ;
  assign n4707 = n4706 ^ x386 ;
  assign n4708 = ~n3457 & n4707 ;
  assign n4709 = n4708 ^ x386 ;
  assign n4704 = n4703 ^ n4702 ;
  assign n4705 = n4704 ^ n4697 ;
  assign n4710 = n4709 ^ n4705 ;
  assign n4711 = ~n3493 & n4710 ;
  assign n4714 = n4711 ^ n4705 ;
  assign n4715 = n4714 ^ x354 ;
  assign n4716 = ~n3537 & n4715 ;
  assign n4717 = n4716 ^ x354 ;
  assign n4712 = n4711 ^ n4710 ;
  assign n4713 = n4712 ^ n4705 ;
  assign n4718 = n4717 ^ n4713 ;
  assign n4719 = n3577 & n4718 ;
  assign n4722 = n4719 ^ n4713 ;
  assign n4723 = n4722 ^ x322 ;
  assign n4724 = ~n3620 & n4723 ;
  assign n4725 = n4724 ^ x322 ;
  assign n4720 = n4719 ^ n4718 ;
  assign n4721 = n4720 ^ n4713 ;
  assign n4726 = n4725 ^ n4721 ;
  assign n4727 = n3656 & n4726 ;
  assign n4730 = n4727 ^ n4721 ;
  assign n4731 = n4730 ^ x290 ;
  assign n4732 = ~n3700 & n4731 ;
  assign n4733 = n4732 ^ x290 ;
  assign n4728 = n4727 ^ n4726 ;
  assign n4729 = n4728 ^ n4721 ;
  assign n4734 = n4733 ^ n4729 ;
  assign n4735 = n3739 & n4734 ;
  assign n4738 = n4735 ^ n4729 ;
  assign n4739 = n4738 ^ x258 ;
  assign n4740 = ~n3783 & n4739 ;
  assign n4741 = n4740 ^ x258 ;
  assign n4736 = n4735 ^ n4734 ;
  assign n4737 = n4736 ^ n4729 ;
  assign n4742 = n4741 ^ n4737 ;
  assign n4743 = ~n3818 & n4742 ;
  assign n4746 = n4743 ^ n4737 ;
  assign n4747 = n4746 ^ x226 ;
  assign n4748 = ~n3861 & n4747 ;
  assign n4749 = n4748 ^ x226 ;
  assign n4744 = n4743 ^ n4742 ;
  assign n4745 = n4744 ^ n4737 ;
  assign n4750 = n4749 ^ n4745 ;
  assign n4751 = n3897 & n4750 ;
  assign n4754 = n4751 ^ n4745 ;
  assign n4755 = n4754 ^ x194 ;
  assign n4756 = ~n3941 & n4755 ;
  assign n4757 = n4756 ^ x194 ;
  assign n4752 = n4751 ^ n4750 ;
  assign n4753 = n4752 ^ n4745 ;
  assign n4758 = n4757 ^ n4753 ;
  assign n4759 = n3980 & n4758 ;
  assign n4762 = n4759 ^ n4753 ;
  assign n4763 = n4762 ^ x162 ;
  assign n4764 = ~n4024 & n4763 ;
  assign n4765 = n4764 ^ x162 ;
  assign n4760 = n4759 ^ n4758 ;
  assign n4761 = n4760 ^ n4753 ;
  assign n4766 = n4765 ^ n4761 ;
  assign n4767 = ~n4059 & n4766 ;
  assign n4770 = n4767 ^ n4761 ;
  assign n4771 = n4770 ^ x130 ;
  assign n4772 = ~n4102 & n4771 ;
  assign n4773 = n4772 ^ x130 ;
  assign n4768 = n4767 ^ n4766 ;
  assign n4769 = n4768 ^ n4761 ;
  assign n4774 = n4773 ^ n4769 ;
  assign n4775 = n4138 & n4774 ;
  assign n4778 = n4775 ^ n4769 ;
  assign n4779 = n4778 ^ x98 ;
  assign n4780 = ~n4182 & n4779 ;
  assign n4781 = n4780 ^ x98 ;
  assign n4776 = n4775 ^ n4774 ;
  assign n4777 = n4776 ^ n4769 ;
  assign n4782 = n4781 ^ n4777 ;
  assign n4783 = n4221 & n4782 ;
  assign n4786 = n4783 ^ n4777 ;
  assign n4787 = n4786 ^ x66 ;
  assign n4788 = ~n4265 & n4787 ;
  assign n4789 = n4788 ^ x66 ;
  assign n4784 = n4783 ^ n4782 ;
  assign n4785 = n4784 ^ n4777 ;
  assign n4790 = n4789 ^ n4785 ;
  assign n4791 = ~n4300 & n4790 ;
  assign n4794 = n4791 ^ n4785 ;
  assign n4795 = n4794 ^ x34 ;
  assign n4796 = ~n4343 & n4795 ;
  assign n4797 = n4796 ^ x34 ;
  assign n4792 = n4791 ^ n4790 ;
  assign n4793 = n4792 ^ n4785 ;
  assign n4798 = n4797 ^ n4793 ;
  assign n4799 = n4379 & n4798 ;
  assign n4802 = n4799 ^ n4793 ;
  assign n4803 = n4802 ^ x2 ;
  assign n4804 = ~n4425 & n4803 ;
  assign n4805 = n4804 ^ x2 ;
  assign n4800 = n4799 ^ n4798 ;
  assign n4801 = n4800 ^ n4793 ;
  assign n4806 = n4805 ^ n4801 ;
  assign n4807 = ~n4461 & n4806 ;
  assign n4808 = n4807 ^ n4806 ;
  assign n4809 = n4808 ^ n4801 ;
  assign n4810 = x483 ^ x451 ;
  assign n4811 = ~n3330 & n4810 ;
  assign n4814 = n4811 ^ x451 ;
  assign n4815 = n4814 ^ x419 ;
  assign n4816 = ~n3377 & n4815 ;
  assign n4817 = n4816 ^ x419 ;
  assign n4812 = n4811 ^ n4810 ;
  assign n4813 = n4812 ^ x451 ;
  assign n4818 = n4817 ^ n4813 ;
  assign n4819 = ~n3413 & n4818 ;
  assign n4822 = n4819 ^ n4813 ;
  assign n4823 = n4822 ^ x387 ;
  assign n4824 = ~n3457 & n4823 ;
  assign n4825 = n4824 ^ x387 ;
  assign n4820 = n4819 ^ n4818 ;
  assign n4821 = n4820 ^ n4813 ;
  assign n4826 = n4825 ^ n4821 ;
  assign n4827 = ~n3493 & n4826 ;
  assign n4830 = n4827 ^ n4821 ;
  assign n4831 = n4830 ^ x355 ;
  assign n4832 = ~n3537 & n4831 ;
  assign n4833 = n4832 ^ x355 ;
  assign n4828 = n4827 ^ n4826 ;
  assign n4829 = n4828 ^ n4821 ;
  assign n4834 = n4833 ^ n4829 ;
  assign n4835 = n3577 & n4834 ;
  assign n4838 = n4835 ^ n4829 ;
  assign n4839 = n4838 ^ x323 ;
  assign n4840 = ~n3620 & n4839 ;
  assign n4841 = n4840 ^ x323 ;
  assign n4836 = n4835 ^ n4834 ;
  assign n4837 = n4836 ^ n4829 ;
  assign n4842 = n4841 ^ n4837 ;
  assign n4843 = n3656 & n4842 ;
  assign n4846 = n4843 ^ n4837 ;
  assign n4847 = n4846 ^ x291 ;
  assign n4848 = ~n3700 & n4847 ;
  assign n4849 = n4848 ^ x291 ;
  assign n4844 = n4843 ^ n4842 ;
  assign n4845 = n4844 ^ n4837 ;
  assign n4850 = n4849 ^ n4845 ;
  assign n4851 = n3739 & n4850 ;
  assign n4854 = n4851 ^ n4845 ;
  assign n4855 = n4854 ^ x259 ;
  assign n4856 = ~n3783 & n4855 ;
  assign n4857 = n4856 ^ x259 ;
  assign n4852 = n4851 ^ n4850 ;
  assign n4853 = n4852 ^ n4845 ;
  assign n4858 = n4857 ^ n4853 ;
  assign n4859 = ~n3818 & n4858 ;
  assign n4862 = n4859 ^ n4853 ;
  assign n4863 = n4862 ^ x227 ;
  assign n4864 = ~n3861 & n4863 ;
  assign n4865 = n4864 ^ x227 ;
  assign n4860 = n4859 ^ n4858 ;
  assign n4861 = n4860 ^ n4853 ;
  assign n4866 = n4865 ^ n4861 ;
  assign n4867 = n3897 & n4866 ;
  assign n4870 = n4867 ^ n4861 ;
  assign n4871 = n4870 ^ x195 ;
  assign n4872 = ~n3941 & n4871 ;
  assign n4873 = n4872 ^ x195 ;
  assign n4868 = n4867 ^ n4866 ;
  assign n4869 = n4868 ^ n4861 ;
  assign n4874 = n4873 ^ n4869 ;
  assign n4875 = n3980 & n4874 ;
  assign n4878 = n4875 ^ n4869 ;
  assign n4879 = n4878 ^ x163 ;
  assign n4880 = ~n4024 & n4879 ;
  assign n4881 = n4880 ^ x163 ;
  assign n4876 = n4875 ^ n4874 ;
  assign n4877 = n4876 ^ n4869 ;
  assign n4882 = n4881 ^ n4877 ;
  assign n4883 = ~n4059 & n4882 ;
  assign n4886 = n4883 ^ n4877 ;
  assign n4887 = n4886 ^ x131 ;
  assign n4888 = ~n4102 & n4887 ;
  assign n4889 = n4888 ^ x131 ;
  assign n4884 = n4883 ^ n4882 ;
  assign n4885 = n4884 ^ n4877 ;
  assign n4890 = n4889 ^ n4885 ;
  assign n4891 = n4138 & n4890 ;
  assign n4894 = n4891 ^ n4885 ;
  assign n4895 = n4894 ^ x99 ;
  assign n4896 = ~n4182 & n4895 ;
  assign n4897 = n4896 ^ x99 ;
  assign n4892 = n4891 ^ n4890 ;
  assign n4893 = n4892 ^ n4885 ;
  assign n4898 = n4897 ^ n4893 ;
  assign n4899 = n4221 & n4898 ;
  assign n4902 = n4899 ^ n4893 ;
  assign n4903 = n4902 ^ x67 ;
  assign n4904 = ~n4265 & n4903 ;
  assign n4905 = n4904 ^ x67 ;
  assign n4900 = n4899 ^ n4898 ;
  assign n4901 = n4900 ^ n4893 ;
  assign n4906 = n4905 ^ n4901 ;
  assign n4907 = ~n4300 & n4906 ;
  assign n4910 = n4907 ^ n4901 ;
  assign n4911 = n4910 ^ x35 ;
  assign n4912 = ~n4343 & n4911 ;
  assign n4913 = n4912 ^ x35 ;
  assign n4908 = n4907 ^ n4906 ;
  assign n4909 = n4908 ^ n4901 ;
  assign n4914 = n4913 ^ n4909 ;
  assign n4915 = n4379 & n4914 ;
  assign n4918 = n4915 ^ n4909 ;
  assign n4919 = n4918 ^ x3 ;
  assign n4920 = ~n4425 & n4919 ;
  assign n4921 = n4920 ^ x3 ;
  assign n4916 = n4915 ^ n4914 ;
  assign n4917 = n4916 ^ n4909 ;
  assign n4922 = n4921 ^ n4917 ;
  assign n4923 = ~n4461 & n4922 ;
  assign n4924 = n4923 ^ n4922 ;
  assign n4925 = n4924 ^ n4917 ;
  assign n4926 = x484 ^ x452 ;
  assign n4927 = ~n3330 & n4926 ;
  assign n4930 = n4927 ^ x452 ;
  assign n4931 = n4930 ^ x420 ;
  assign n4932 = ~n3377 & n4931 ;
  assign n4933 = n4932 ^ x420 ;
  assign n4928 = n4927 ^ n4926 ;
  assign n4929 = n4928 ^ x452 ;
  assign n4934 = n4933 ^ n4929 ;
  assign n4935 = ~n3413 & n4934 ;
  assign n4938 = n4935 ^ n4929 ;
  assign n4939 = n4938 ^ x388 ;
  assign n4940 = ~n3457 & n4939 ;
  assign n4941 = n4940 ^ x388 ;
  assign n4936 = n4935 ^ n4934 ;
  assign n4937 = n4936 ^ n4929 ;
  assign n4942 = n4941 ^ n4937 ;
  assign n4943 = ~n3493 & n4942 ;
  assign n4946 = n4943 ^ n4937 ;
  assign n4947 = n4946 ^ x356 ;
  assign n4948 = ~n3537 & n4947 ;
  assign n4949 = n4948 ^ x356 ;
  assign n4944 = n4943 ^ n4942 ;
  assign n4945 = n4944 ^ n4937 ;
  assign n4950 = n4949 ^ n4945 ;
  assign n4951 = n3577 & n4950 ;
  assign n4954 = n4951 ^ n4945 ;
  assign n4955 = n4954 ^ x324 ;
  assign n4956 = ~n3620 & n4955 ;
  assign n4957 = n4956 ^ x324 ;
  assign n4952 = n4951 ^ n4950 ;
  assign n4953 = n4952 ^ n4945 ;
  assign n4958 = n4957 ^ n4953 ;
  assign n4959 = n3656 & n4958 ;
  assign n4962 = n4959 ^ n4953 ;
  assign n4963 = n4962 ^ x292 ;
  assign n4964 = ~n3700 & n4963 ;
  assign n4965 = n4964 ^ x292 ;
  assign n4960 = n4959 ^ n4958 ;
  assign n4961 = n4960 ^ n4953 ;
  assign n4966 = n4965 ^ n4961 ;
  assign n4967 = n3739 & n4966 ;
  assign n4970 = n4967 ^ n4961 ;
  assign n4971 = n4970 ^ x260 ;
  assign n4972 = ~n3783 & n4971 ;
  assign n4973 = n4972 ^ x260 ;
  assign n4968 = n4967 ^ n4966 ;
  assign n4969 = n4968 ^ n4961 ;
  assign n4974 = n4973 ^ n4969 ;
  assign n4975 = ~n3818 & n4974 ;
  assign n4978 = n4975 ^ n4969 ;
  assign n4979 = n4978 ^ x228 ;
  assign n4980 = ~n3861 & n4979 ;
  assign n4981 = n4980 ^ x228 ;
  assign n4976 = n4975 ^ n4974 ;
  assign n4977 = n4976 ^ n4969 ;
  assign n4982 = n4981 ^ n4977 ;
  assign n4983 = n3897 & n4982 ;
  assign n4986 = n4983 ^ n4977 ;
  assign n4987 = n4986 ^ x196 ;
  assign n4988 = ~n3941 & n4987 ;
  assign n4989 = n4988 ^ x196 ;
  assign n4984 = n4983 ^ n4982 ;
  assign n4985 = n4984 ^ n4977 ;
  assign n4990 = n4989 ^ n4985 ;
  assign n4991 = n3980 & n4990 ;
  assign n4994 = n4991 ^ n4985 ;
  assign n4995 = n4994 ^ x164 ;
  assign n4996 = ~n4024 & n4995 ;
  assign n4997 = n4996 ^ x164 ;
  assign n4992 = n4991 ^ n4990 ;
  assign n4993 = n4992 ^ n4985 ;
  assign n4998 = n4997 ^ n4993 ;
  assign n4999 = ~n4059 & n4998 ;
  assign n5002 = n4999 ^ n4993 ;
  assign n5003 = n5002 ^ x132 ;
  assign n5004 = ~n4102 & n5003 ;
  assign n5005 = n5004 ^ x132 ;
  assign n5000 = n4999 ^ n4998 ;
  assign n5001 = n5000 ^ n4993 ;
  assign n5006 = n5005 ^ n5001 ;
  assign n5007 = n4138 & n5006 ;
  assign n5010 = n5007 ^ n5001 ;
  assign n5011 = n5010 ^ x100 ;
  assign n5012 = ~n4182 & n5011 ;
  assign n5013 = n5012 ^ x100 ;
  assign n5008 = n5007 ^ n5006 ;
  assign n5009 = n5008 ^ n5001 ;
  assign n5014 = n5013 ^ n5009 ;
  assign n5015 = n4221 & n5014 ;
  assign n5018 = n5015 ^ n5009 ;
  assign n5019 = n5018 ^ x68 ;
  assign n5020 = ~n4265 & n5019 ;
  assign n5021 = n5020 ^ x68 ;
  assign n5016 = n5015 ^ n5014 ;
  assign n5017 = n5016 ^ n5009 ;
  assign n5022 = n5021 ^ n5017 ;
  assign n5023 = ~n4300 & n5022 ;
  assign n5026 = n5023 ^ n5017 ;
  assign n5027 = n5026 ^ x36 ;
  assign n5028 = ~n4343 & n5027 ;
  assign n5029 = n5028 ^ x36 ;
  assign n5024 = n5023 ^ n5022 ;
  assign n5025 = n5024 ^ n5017 ;
  assign n5030 = n5029 ^ n5025 ;
  assign n5031 = n4379 & n5030 ;
  assign n5034 = n5031 ^ n5025 ;
  assign n5035 = n5034 ^ x4 ;
  assign n5036 = ~n4425 & n5035 ;
  assign n5037 = n5036 ^ x4 ;
  assign n5032 = n5031 ^ n5030 ;
  assign n5033 = n5032 ^ n5025 ;
  assign n5038 = n5037 ^ n5033 ;
  assign n5039 = ~n4461 & n5038 ;
  assign n5040 = n5039 ^ n5038 ;
  assign n5041 = n5040 ^ n5033 ;
  assign n5042 = x485 ^ x453 ;
  assign n5043 = ~n3330 & n5042 ;
  assign n5046 = n5043 ^ x453 ;
  assign n5047 = n5046 ^ x421 ;
  assign n5048 = ~n3377 & n5047 ;
  assign n5049 = n5048 ^ x421 ;
  assign n5044 = n5043 ^ n5042 ;
  assign n5045 = n5044 ^ x453 ;
  assign n5050 = n5049 ^ n5045 ;
  assign n5051 = ~n3413 & n5050 ;
  assign n5054 = n5051 ^ n5045 ;
  assign n5055 = n5054 ^ x389 ;
  assign n5056 = ~n3457 & n5055 ;
  assign n5057 = n5056 ^ x389 ;
  assign n5052 = n5051 ^ n5050 ;
  assign n5053 = n5052 ^ n5045 ;
  assign n5058 = n5057 ^ n5053 ;
  assign n5059 = ~n3493 & n5058 ;
  assign n5062 = n5059 ^ n5053 ;
  assign n5063 = n5062 ^ x357 ;
  assign n5064 = ~n3537 & n5063 ;
  assign n5065 = n5064 ^ x357 ;
  assign n5060 = n5059 ^ n5058 ;
  assign n5061 = n5060 ^ n5053 ;
  assign n5066 = n5065 ^ n5061 ;
  assign n5067 = n3577 & n5066 ;
  assign n5070 = n5067 ^ n5061 ;
  assign n5071 = n5070 ^ x325 ;
  assign n5072 = ~n3620 & n5071 ;
  assign n5073 = n5072 ^ x325 ;
  assign n5068 = n5067 ^ n5066 ;
  assign n5069 = n5068 ^ n5061 ;
  assign n5074 = n5073 ^ n5069 ;
  assign n5075 = n3656 & n5074 ;
  assign n5078 = n5075 ^ n5069 ;
  assign n5079 = n5078 ^ x293 ;
  assign n5080 = ~n3700 & n5079 ;
  assign n5081 = n5080 ^ x293 ;
  assign n5076 = n5075 ^ n5074 ;
  assign n5077 = n5076 ^ n5069 ;
  assign n5082 = n5081 ^ n5077 ;
  assign n5083 = n3739 & n5082 ;
  assign n5086 = n5083 ^ n5077 ;
  assign n5087 = n5086 ^ x261 ;
  assign n5088 = ~n3783 & n5087 ;
  assign n5089 = n5088 ^ x261 ;
  assign n5084 = n5083 ^ n5082 ;
  assign n5085 = n5084 ^ n5077 ;
  assign n5090 = n5089 ^ n5085 ;
  assign n5091 = ~n3818 & n5090 ;
  assign n5094 = n5091 ^ n5085 ;
  assign n5095 = n5094 ^ x229 ;
  assign n5096 = ~n3861 & n5095 ;
  assign n5097 = n5096 ^ x229 ;
  assign n5092 = n5091 ^ n5090 ;
  assign n5093 = n5092 ^ n5085 ;
  assign n5098 = n5097 ^ n5093 ;
  assign n5099 = n3897 & n5098 ;
  assign n5102 = n5099 ^ n5093 ;
  assign n5103 = n5102 ^ x197 ;
  assign n5104 = ~n3941 & n5103 ;
  assign n5105 = n5104 ^ x197 ;
  assign n5100 = n5099 ^ n5098 ;
  assign n5101 = n5100 ^ n5093 ;
  assign n5106 = n5105 ^ n5101 ;
  assign n5107 = n3980 & n5106 ;
  assign n5110 = n5107 ^ n5101 ;
  assign n5111 = n5110 ^ x165 ;
  assign n5112 = ~n4024 & n5111 ;
  assign n5113 = n5112 ^ x165 ;
  assign n5108 = n5107 ^ n5106 ;
  assign n5109 = n5108 ^ n5101 ;
  assign n5114 = n5113 ^ n5109 ;
  assign n5115 = ~n4059 & n5114 ;
  assign n5118 = n5115 ^ n5109 ;
  assign n5119 = n5118 ^ x133 ;
  assign n5120 = ~n4102 & n5119 ;
  assign n5121 = n5120 ^ x133 ;
  assign n5116 = n5115 ^ n5114 ;
  assign n5117 = n5116 ^ n5109 ;
  assign n5122 = n5121 ^ n5117 ;
  assign n5123 = n4138 & n5122 ;
  assign n5126 = n5123 ^ n5117 ;
  assign n5127 = n5126 ^ x101 ;
  assign n5128 = ~n4182 & n5127 ;
  assign n5129 = n5128 ^ x101 ;
  assign n5124 = n5123 ^ n5122 ;
  assign n5125 = n5124 ^ n5117 ;
  assign n5130 = n5129 ^ n5125 ;
  assign n5131 = n4221 & n5130 ;
  assign n5134 = n5131 ^ n5125 ;
  assign n5135 = n5134 ^ x69 ;
  assign n5136 = ~n4265 & n5135 ;
  assign n5137 = n5136 ^ x69 ;
  assign n5132 = n5131 ^ n5130 ;
  assign n5133 = n5132 ^ n5125 ;
  assign n5138 = n5137 ^ n5133 ;
  assign n5139 = ~n4300 & n5138 ;
  assign n5142 = n5139 ^ n5133 ;
  assign n5143 = n5142 ^ x37 ;
  assign n5144 = ~n4343 & n5143 ;
  assign n5145 = n5144 ^ x37 ;
  assign n5140 = n5139 ^ n5138 ;
  assign n5141 = n5140 ^ n5133 ;
  assign n5146 = n5145 ^ n5141 ;
  assign n5147 = n4379 & n5146 ;
  assign n5150 = n5147 ^ n5141 ;
  assign n5151 = n5150 ^ x5 ;
  assign n5152 = ~n4425 & n5151 ;
  assign n5153 = n5152 ^ x5 ;
  assign n5148 = n5147 ^ n5146 ;
  assign n5149 = n5148 ^ n5141 ;
  assign n5154 = n5153 ^ n5149 ;
  assign n5155 = ~n4461 & n5154 ;
  assign n5156 = n5155 ^ n5154 ;
  assign n5157 = n5156 ^ n5149 ;
  assign n5158 = x486 ^ x454 ;
  assign n5159 = ~n3330 & n5158 ;
  assign n5162 = n5159 ^ x454 ;
  assign n5163 = n5162 ^ x422 ;
  assign n5164 = ~n3377 & n5163 ;
  assign n5165 = n5164 ^ x422 ;
  assign n5160 = n5159 ^ n5158 ;
  assign n5161 = n5160 ^ x454 ;
  assign n5166 = n5165 ^ n5161 ;
  assign n5167 = ~n3413 & n5166 ;
  assign n5170 = n5167 ^ n5161 ;
  assign n5171 = n5170 ^ x390 ;
  assign n5172 = ~n3457 & n5171 ;
  assign n5173 = n5172 ^ x390 ;
  assign n5168 = n5167 ^ n5166 ;
  assign n5169 = n5168 ^ n5161 ;
  assign n5174 = n5173 ^ n5169 ;
  assign n5175 = ~n3493 & n5174 ;
  assign n5178 = n5175 ^ n5169 ;
  assign n5179 = n5178 ^ x358 ;
  assign n5180 = ~n3537 & n5179 ;
  assign n5181 = n5180 ^ x358 ;
  assign n5176 = n5175 ^ n5174 ;
  assign n5177 = n5176 ^ n5169 ;
  assign n5182 = n5181 ^ n5177 ;
  assign n5183 = n3577 & n5182 ;
  assign n5186 = n5183 ^ n5177 ;
  assign n5187 = n5186 ^ x326 ;
  assign n5188 = ~n3620 & n5187 ;
  assign n5189 = n5188 ^ x326 ;
  assign n5184 = n5183 ^ n5182 ;
  assign n5185 = n5184 ^ n5177 ;
  assign n5190 = n5189 ^ n5185 ;
  assign n5191 = n3656 & n5190 ;
  assign n5194 = n5191 ^ n5185 ;
  assign n5195 = n5194 ^ x294 ;
  assign n5196 = ~n3700 & n5195 ;
  assign n5197 = n5196 ^ x294 ;
  assign n5192 = n5191 ^ n5190 ;
  assign n5193 = n5192 ^ n5185 ;
  assign n5198 = n5197 ^ n5193 ;
  assign n5199 = n3739 & n5198 ;
  assign n5202 = n5199 ^ n5193 ;
  assign n5203 = n5202 ^ x262 ;
  assign n5204 = ~n3783 & n5203 ;
  assign n5205 = n5204 ^ x262 ;
  assign n5200 = n5199 ^ n5198 ;
  assign n5201 = n5200 ^ n5193 ;
  assign n5206 = n5205 ^ n5201 ;
  assign n5207 = ~n3818 & n5206 ;
  assign n5210 = n5207 ^ n5201 ;
  assign n5211 = n5210 ^ x230 ;
  assign n5212 = ~n3861 & n5211 ;
  assign n5213 = n5212 ^ x230 ;
  assign n5208 = n5207 ^ n5206 ;
  assign n5209 = n5208 ^ n5201 ;
  assign n5214 = n5213 ^ n5209 ;
  assign n5215 = n3897 & n5214 ;
  assign n5218 = n5215 ^ n5209 ;
  assign n5219 = n5218 ^ x198 ;
  assign n5220 = ~n3941 & n5219 ;
  assign n5221 = n5220 ^ x198 ;
  assign n5216 = n5215 ^ n5214 ;
  assign n5217 = n5216 ^ n5209 ;
  assign n5222 = n5221 ^ n5217 ;
  assign n5223 = n3980 & n5222 ;
  assign n5226 = n5223 ^ n5217 ;
  assign n5227 = n5226 ^ x166 ;
  assign n5228 = ~n4024 & n5227 ;
  assign n5229 = n5228 ^ x166 ;
  assign n5224 = n5223 ^ n5222 ;
  assign n5225 = n5224 ^ n5217 ;
  assign n5230 = n5229 ^ n5225 ;
  assign n5231 = ~n4059 & n5230 ;
  assign n5234 = n5231 ^ n5225 ;
  assign n5235 = n5234 ^ x134 ;
  assign n5236 = ~n4102 & n5235 ;
  assign n5237 = n5236 ^ x134 ;
  assign n5232 = n5231 ^ n5230 ;
  assign n5233 = n5232 ^ n5225 ;
  assign n5238 = n5237 ^ n5233 ;
  assign n5239 = n4138 & n5238 ;
  assign n5242 = n5239 ^ n5233 ;
  assign n5243 = n5242 ^ x102 ;
  assign n5244 = ~n4182 & n5243 ;
  assign n5245 = n5244 ^ x102 ;
  assign n5240 = n5239 ^ n5238 ;
  assign n5241 = n5240 ^ n5233 ;
  assign n5246 = n5245 ^ n5241 ;
  assign n5247 = n4221 & n5246 ;
  assign n5250 = n5247 ^ n5241 ;
  assign n5251 = n5250 ^ x70 ;
  assign n5252 = ~n4265 & n5251 ;
  assign n5253 = n5252 ^ x70 ;
  assign n5248 = n5247 ^ n5246 ;
  assign n5249 = n5248 ^ n5241 ;
  assign n5254 = n5253 ^ n5249 ;
  assign n5255 = ~n4300 & n5254 ;
  assign n5258 = n5255 ^ n5249 ;
  assign n5259 = n5258 ^ x38 ;
  assign n5260 = ~n4343 & n5259 ;
  assign n5261 = n5260 ^ x38 ;
  assign n5256 = n5255 ^ n5254 ;
  assign n5257 = n5256 ^ n5249 ;
  assign n5262 = n5261 ^ n5257 ;
  assign n5263 = n4379 & n5262 ;
  assign n5266 = n5263 ^ n5257 ;
  assign n5267 = n5266 ^ x6 ;
  assign n5268 = ~n4425 & n5267 ;
  assign n5269 = n5268 ^ x6 ;
  assign n5264 = n5263 ^ n5262 ;
  assign n5265 = n5264 ^ n5257 ;
  assign n5270 = n5269 ^ n5265 ;
  assign n5271 = ~n4461 & n5270 ;
  assign n5272 = n5271 ^ n5270 ;
  assign n5273 = n5272 ^ n5265 ;
  assign n5274 = x487 ^ x455 ;
  assign n5275 = ~n3330 & n5274 ;
  assign n5278 = n5275 ^ x455 ;
  assign n5279 = n5278 ^ x423 ;
  assign n5280 = ~n3377 & n5279 ;
  assign n5281 = n5280 ^ x423 ;
  assign n5276 = n5275 ^ n5274 ;
  assign n5277 = n5276 ^ x455 ;
  assign n5282 = n5281 ^ n5277 ;
  assign n5283 = ~n3413 & n5282 ;
  assign n5286 = n5283 ^ n5277 ;
  assign n5287 = n5286 ^ x391 ;
  assign n5288 = ~n3457 & n5287 ;
  assign n5289 = n5288 ^ x391 ;
  assign n5284 = n5283 ^ n5282 ;
  assign n5285 = n5284 ^ n5277 ;
  assign n5290 = n5289 ^ n5285 ;
  assign n5291 = ~n3493 & n5290 ;
  assign n5294 = n5291 ^ n5285 ;
  assign n5295 = n5294 ^ x359 ;
  assign n5296 = ~n3537 & n5295 ;
  assign n5297 = n5296 ^ x359 ;
  assign n5292 = n5291 ^ n5290 ;
  assign n5293 = n5292 ^ n5285 ;
  assign n5298 = n5297 ^ n5293 ;
  assign n5299 = n3577 & n5298 ;
  assign n5302 = n5299 ^ n5293 ;
  assign n5303 = n5302 ^ x327 ;
  assign n5304 = ~n3620 & n5303 ;
  assign n5305 = n5304 ^ x327 ;
  assign n5300 = n5299 ^ n5298 ;
  assign n5301 = n5300 ^ n5293 ;
  assign n5306 = n5305 ^ n5301 ;
  assign n5307 = n3656 & n5306 ;
  assign n5310 = n5307 ^ n5301 ;
  assign n5311 = n5310 ^ x295 ;
  assign n5312 = ~n3700 & n5311 ;
  assign n5313 = n5312 ^ x295 ;
  assign n5308 = n5307 ^ n5306 ;
  assign n5309 = n5308 ^ n5301 ;
  assign n5314 = n5313 ^ n5309 ;
  assign n5315 = n3739 & n5314 ;
  assign n5318 = n5315 ^ n5309 ;
  assign n5319 = n5318 ^ x263 ;
  assign n5320 = ~n3783 & n5319 ;
  assign n5321 = n5320 ^ x263 ;
  assign n5316 = n5315 ^ n5314 ;
  assign n5317 = n5316 ^ n5309 ;
  assign n5322 = n5321 ^ n5317 ;
  assign n5323 = ~n3818 & n5322 ;
  assign n5326 = n5323 ^ n5317 ;
  assign n5327 = n5326 ^ x231 ;
  assign n5328 = ~n3861 & n5327 ;
  assign n5329 = n5328 ^ x231 ;
  assign n5324 = n5323 ^ n5322 ;
  assign n5325 = n5324 ^ n5317 ;
  assign n5330 = n5329 ^ n5325 ;
  assign n5331 = n3897 & n5330 ;
  assign n5334 = n5331 ^ n5325 ;
  assign n5335 = n5334 ^ x199 ;
  assign n5336 = ~n3941 & n5335 ;
  assign n5337 = n5336 ^ x199 ;
  assign n5332 = n5331 ^ n5330 ;
  assign n5333 = n5332 ^ n5325 ;
  assign n5338 = n5337 ^ n5333 ;
  assign n5339 = n3980 & n5338 ;
  assign n5342 = n5339 ^ n5333 ;
  assign n5343 = n5342 ^ x167 ;
  assign n5344 = ~n4024 & n5343 ;
  assign n5345 = n5344 ^ x167 ;
  assign n5340 = n5339 ^ n5338 ;
  assign n5341 = n5340 ^ n5333 ;
  assign n5346 = n5345 ^ n5341 ;
  assign n5347 = ~n4059 & n5346 ;
  assign n5350 = n5347 ^ n5341 ;
  assign n5351 = n5350 ^ x135 ;
  assign n5352 = ~n4102 & n5351 ;
  assign n5353 = n5352 ^ x135 ;
  assign n5348 = n5347 ^ n5346 ;
  assign n5349 = n5348 ^ n5341 ;
  assign n5354 = n5353 ^ n5349 ;
  assign n5355 = n4138 & n5354 ;
  assign n5358 = n5355 ^ n5349 ;
  assign n5359 = n5358 ^ x103 ;
  assign n5360 = ~n4182 & n5359 ;
  assign n5361 = n5360 ^ x103 ;
  assign n5356 = n5355 ^ n5354 ;
  assign n5357 = n5356 ^ n5349 ;
  assign n5362 = n5361 ^ n5357 ;
  assign n5363 = n4221 & n5362 ;
  assign n5366 = n5363 ^ n5357 ;
  assign n5367 = n5366 ^ x71 ;
  assign n5368 = ~n4265 & n5367 ;
  assign n5369 = n5368 ^ x71 ;
  assign n5364 = n5363 ^ n5362 ;
  assign n5365 = n5364 ^ n5357 ;
  assign n5370 = n5369 ^ n5365 ;
  assign n5371 = ~n4300 & n5370 ;
  assign n5374 = n5371 ^ n5365 ;
  assign n5375 = n5374 ^ x39 ;
  assign n5376 = ~n4343 & n5375 ;
  assign n5377 = n5376 ^ x39 ;
  assign n5372 = n5371 ^ n5370 ;
  assign n5373 = n5372 ^ n5365 ;
  assign n5378 = n5377 ^ n5373 ;
  assign n5379 = n4379 & n5378 ;
  assign n5382 = n5379 ^ n5373 ;
  assign n5383 = n5382 ^ x7 ;
  assign n5384 = ~n4425 & n5383 ;
  assign n5385 = n5384 ^ x7 ;
  assign n5380 = n5379 ^ n5378 ;
  assign n5381 = n5380 ^ n5373 ;
  assign n5386 = n5385 ^ n5381 ;
  assign n5387 = ~n4461 & n5386 ;
  assign n5388 = n5387 ^ n5386 ;
  assign n5389 = n5388 ^ n5381 ;
  assign n5390 = x488 ^ x456 ;
  assign n5391 = ~n3330 & n5390 ;
  assign n5394 = n5391 ^ x456 ;
  assign n5395 = n5394 ^ x424 ;
  assign n5396 = ~n3377 & n5395 ;
  assign n5397 = n5396 ^ x424 ;
  assign n5392 = n5391 ^ n5390 ;
  assign n5393 = n5392 ^ x456 ;
  assign n5398 = n5397 ^ n5393 ;
  assign n5399 = ~n3413 & n5398 ;
  assign n5402 = n5399 ^ n5393 ;
  assign n5403 = n5402 ^ x392 ;
  assign n5404 = ~n3457 & n5403 ;
  assign n5405 = n5404 ^ x392 ;
  assign n5400 = n5399 ^ n5398 ;
  assign n5401 = n5400 ^ n5393 ;
  assign n5406 = n5405 ^ n5401 ;
  assign n5407 = ~n3493 & n5406 ;
  assign n5410 = n5407 ^ n5401 ;
  assign n5411 = n5410 ^ x360 ;
  assign n5412 = ~n3537 & n5411 ;
  assign n5413 = n5412 ^ x360 ;
  assign n5408 = n5407 ^ n5406 ;
  assign n5409 = n5408 ^ n5401 ;
  assign n5414 = n5413 ^ n5409 ;
  assign n5415 = n3577 & n5414 ;
  assign n5418 = n5415 ^ n5409 ;
  assign n5419 = n5418 ^ x328 ;
  assign n5420 = ~n3620 & n5419 ;
  assign n5421 = n5420 ^ x328 ;
  assign n5416 = n5415 ^ n5414 ;
  assign n5417 = n5416 ^ n5409 ;
  assign n5422 = n5421 ^ n5417 ;
  assign n5423 = n3656 & n5422 ;
  assign n5426 = n5423 ^ n5417 ;
  assign n5427 = n5426 ^ x296 ;
  assign n5428 = ~n3700 & n5427 ;
  assign n5429 = n5428 ^ x296 ;
  assign n5424 = n5423 ^ n5422 ;
  assign n5425 = n5424 ^ n5417 ;
  assign n5430 = n5429 ^ n5425 ;
  assign n5431 = n3739 & n5430 ;
  assign n5434 = n5431 ^ n5425 ;
  assign n5435 = n5434 ^ x264 ;
  assign n5436 = ~n3783 & n5435 ;
  assign n5437 = n5436 ^ x264 ;
  assign n5432 = n5431 ^ n5430 ;
  assign n5433 = n5432 ^ n5425 ;
  assign n5438 = n5437 ^ n5433 ;
  assign n5439 = ~n3818 & n5438 ;
  assign n5442 = n5439 ^ n5433 ;
  assign n5443 = n5442 ^ x232 ;
  assign n5444 = ~n3861 & n5443 ;
  assign n5445 = n5444 ^ x232 ;
  assign n5440 = n5439 ^ n5438 ;
  assign n5441 = n5440 ^ n5433 ;
  assign n5446 = n5445 ^ n5441 ;
  assign n5447 = n3897 & n5446 ;
  assign n5450 = n5447 ^ n5441 ;
  assign n5451 = n5450 ^ x200 ;
  assign n5452 = ~n3941 & n5451 ;
  assign n5453 = n5452 ^ x200 ;
  assign n5448 = n5447 ^ n5446 ;
  assign n5449 = n5448 ^ n5441 ;
  assign n5454 = n5453 ^ n5449 ;
  assign n5455 = n3980 & n5454 ;
  assign n5458 = n5455 ^ n5449 ;
  assign n5459 = n5458 ^ x168 ;
  assign n5460 = ~n4024 & n5459 ;
  assign n5461 = n5460 ^ x168 ;
  assign n5456 = n5455 ^ n5454 ;
  assign n5457 = n5456 ^ n5449 ;
  assign n5462 = n5461 ^ n5457 ;
  assign n5463 = ~n4059 & n5462 ;
  assign n5466 = n5463 ^ n5457 ;
  assign n5467 = n5466 ^ x136 ;
  assign n5468 = ~n4102 & n5467 ;
  assign n5469 = n5468 ^ x136 ;
  assign n5464 = n5463 ^ n5462 ;
  assign n5465 = n5464 ^ n5457 ;
  assign n5470 = n5469 ^ n5465 ;
  assign n5471 = n4138 & n5470 ;
  assign n5474 = n5471 ^ n5465 ;
  assign n5475 = n5474 ^ x104 ;
  assign n5476 = ~n4182 & n5475 ;
  assign n5477 = n5476 ^ x104 ;
  assign n5472 = n5471 ^ n5470 ;
  assign n5473 = n5472 ^ n5465 ;
  assign n5478 = n5477 ^ n5473 ;
  assign n5479 = n4221 & n5478 ;
  assign n5482 = n5479 ^ n5473 ;
  assign n5483 = n5482 ^ x72 ;
  assign n5484 = ~n4265 & n5483 ;
  assign n5485 = n5484 ^ x72 ;
  assign n5480 = n5479 ^ n5478 ;
  assign n5481 = n5480 ^ n5473 ;
  assign n5486 = n5485 ^ n5481 ;
  assign n5487 = ~n4300 & n5486 ;
  assign n5490 = n5487 ^ n5481 ;
  assign n5491 = n5490 ^ x40 ;
  assign n5492 = ~n4343 & n5491 ;
  assign n5493 = n5492 ^ x40 ;
  assign n5488 = n5487 ^ n5486 ;
  assign n5489 = n5488 ^ n5481 ;
  assign n5494 = n5493 ^ n5489 ;
  assign n5495 = n4379 & n5494 ;
  assign n5498 = n5495 ^ n5489 ;
  assign n5499 = n5498 ^ x8 ;
  assign n5500 = ~n4425 & n5499 ;
  assign n5501 = n5500 ^ x8 ;
  assign n5496 = n5495 ^ n5494 ;
  assign n5497 = n5496 ^ n5489 ;
  assign n5502 = n5501 ^ n5497 ;
  assign n5503 = ~n4461 & n5502 ;
  assign n5504 = n5503 ^ n5502 ;
  assign n5505 = n5504 ^ n5497 ;
  assign n5506 = x489 ^ x457 ;
  assign n5507 = ~n3330 & n5506 ;
  assign n5510 = n5507 ^ x457 ;
  assign n5511 = n5510 ^ x425 ;
  assign n5512 = ~n3377 & n5511 ;
  assign n5513 = n5512 ^ x425 ;
  assign n5508 = n5507 ^ n5506 ;
  assign n5509 = n5508 ^ x457 ;
  assign n5514 = n5513 ^ n5509 ;
  assign n5515 = ~n3413 & n5514 ;
  assign n5518 = n5515 ^ n5509 ;
  assign n5519 = n5518 ^ x393 ;
  assign n5520 = ~n3457 & n5519 ;
  assign n5521 = n5520 ^ x393 ;
  assign n5516 = n5515 ^ n5514 ;
  assign n5517 = n5516 ^ n5509 ;
  assign n5522 = n5521 ^ n5517 ;
  assign n5523 = ~n3493 & n5522 ;
  assign n5526 = n5523 ^ n5517 ;
  assign n5527 = n5526 ^ x361 ;
  assign n5528 = ~n3537 & n5527 ;
  assign n5529 = n5528 ^ x361 ;
  assign n5524 = n5523 ^ n5522 ;
  assign n5525 = n5524 ^ n5517 ;
  assign n5530 = n5529 ^ n5525 ;
  assign n5531 = n3577 & n5530 ;
  assign n5534 = n5531 ^ n5525 ;
  assign n5535 = n5534 ^ x329 ;
  assign n5536 = ~n3620 & n5535 ;
  assign n5537 = n5536 ^ x329 ;
  assign n5532 = n5531 ^ n5530 ;
  assign n5533 = n5532 ^ n5525 ;
  assign n5538 = n5537 ^ n5533 ;
  assign n5539 = n3656 & n5538 ;
  assign n5542 = n5539 ^ n5533 ;
  assign n5543 = n5542 ^ x297 ;
  assign n5544 = ~n3700 & n5543 ;
  assign n5545 = n5544 ^ x297 ;
  assign n5540 = n5539 ^ n5538 ;
  assign n5541 = n5540 ^ n5533 ;
  assign n5546 = n5545 ^ n5541 ;
  assign n5547 = n3739 & n5546 ;
  assign n5550 = n5547 ^ n5541 ;
  assign n5551 = n5550 ^ x265 ;
  assign n5552 = ~n3783 & n5551 ;
  assign n5553 = n5552 ^ x265 ;
  assign n5548 = n5547 ^ n5546 ;
  assign n5549 = n5548 ^ n5541 ;
  assign n5554 = n5553 ^ n5549 ;
  assign n5555 = ~n3818 & n5554 ;
  assign n5558 = n5555 ^ n5549 ;
  assign n5559 = n5558 ^ x233 ;
  assign n5560 = ~n3861 & n5559 ;
  assign n5561 = n5560 ^ x233 ;
  assign n5556 = n5555 ^ n5554 ;
  assign n5557 = n5556 ^ n5549 ;
  assign n5562 = n5561 ^ n5557 ;
  assign n5563 = n3897 & n5562 ;
  assign n5566 = n5563 ^ n5557 ;
  assign n5567 = n5566 ^ x201 ;
  assign n5568 = ~n3941 & n5567 ;
  assign n5569 = n5568 ^ x201 ;
  assign n5564 = n5563 ^ n5562 ;
  assign n5565 = n5564 ^ n5557 ;
  assign n5570 = n5569 ^ n5565 ;
  assign n5571 = n3980 & n5570 ;
  assign n5574 = n5571 ^ n5565 ;
  assign n5575 = n5574 ^ x169 ;
  assign n5576 = ~n4024 & n5575 ;
  assign n5577 = n5576 ^ x169 ;
  assign n5572 = n5571 ^ n5570 ;
  assign n5573 = n5572 ^ n5565 ;
  assign n5578 = n5577 ^ n5573 ;
  assign n5579 = ~n4059 & n5578 ;
  assign n5582 = n5579 ^ n5573 ;
  assign n5583 = n5582 ^ x137 ;
  assign n5584 = ~n4102 & n5583 ;
  assign n5585 = n5584 ^ x137 ;
  assign n5580 = n5579 ^ n5578 ;
  assign n5581 = n5580 ^ n5573 ;
  assign n5586 = n5585 ^ n5581 ;
  assign n5587 = n4138 & n5586 ;
  assign n5590 = n5587 ^ n5581 ;
  assign n5591 = n5590 ^ x105 ;
  assign n5592 = ~n4182 & n5591 ;
  assign n5593 = n5592 ^ x105 ;
  assign n5588 = n5587 ^ n5586 ;
  assign n5589 = n5588 ^ n5581 ;
  assign n5594 = n5593 ^ n5589 ;
  assign n5595 = n4221 & n5594 ;
  assign n5598 = n5595 ^ n5589 ;
  assign n5599 = n5598 ^ x73 ;
  assign n5600 = ~n4265 & n5599 ;
  assign n5601 = n5600 ^ x73 ;
  assign n5596 = n5595 ^ n5594 ;
  assign n5597 = n5596 ^ n5589 ;
  assign n5602 = n5601 ^ n5597 ;
  assign n5603 = ~n4300 & n5602 ;
  assign n5606 = n5603 ^ n5597 ;
  assign n5607 = n5606 ^ x41 ;
  assign n5608 = ~n4343 & n5607 ;
  assign n5609 = n5608 ^ x41 ;
  assign n5604 = n5603 ^ n5602 ;
  assign n5605 = n5604 ^ n5597 ;
  assign n5610 = n5609 ^ n5605 ;
  assign n5611 = n4379 & n5610 ;
  assign n5614 = n5611 ^ n5605 ;
  assign n5615 = n5614 ^ x9 ;
  assign n5616 = ~n4425 & n5615 ;
  assign n5617 = n5616 ^ x9 ;
  assign n5612 = n5611 ^ n5610 ;
  assign n5613 = n5612 ^ n5605 ;
  assign n5618 = n5617 ^ n5613 ;
  assign n5619 = ~n4461 & n5618 ;
  assign n5620 = n5619 ^ n5618 ;
  assign n5621 = n5620 ^ n5613 ;
  assign n5622 = x490 ^ x458 ;
  assign n5623 = ~n3330 & n5622 ;
  assign n5626 = n5623 ^ x458 ;
  assign n5627 = n5626 ^ x426 ;
  assign n5628 = ~n3377 & n5627 ;
  assign n5629 = n5628 ^ x426 ;
  assign n5624 = n5623 ^ n5622 ;
  assign n5625 = n5624 ^ x458 ;
  assign n5630 = n5629 ^ n5625 ;
  assign n5631 = ~n3413 & n5630 ;
  assign n5634 = n5631 ^ n5625 ;
  assign n5635 = n5634 ^ x394 ;
  assign n5636 = ~n3457 & n5635 ;
  assign n5637 = n5636 ^ x394 ;
  assign n5632 = n5631 ^ n5630 ;
  assign n5633 = n5632 ^ n5625 ;
  assign n5638 = n5637 ^ n5633 ;
  assign n5639 = ~n3493 & n5638 ;
  assign n5642 = n5639 ^ n5633 ;
  assign n5643 = n5642 ^ x362 ;
  assign n5644 = ~n3537 & n5643 ;
  assign n5645 = n5644 ^ x362 ;
  assign n5640 = n5639 ^ n5638 ;
  assign n5641 = n5640 ^ n5633 ;
  assign n5646 = n5645 ^ n5641 ;
  assign n5647 = n3577 & n5646 ;
  assign n5650 = n5647 ^ n5641 ;
  assign n5651 = n5650 ^ x330 ;
  assign n5652 = ~n3620 & n5651 ;
  assign n5653 = n5652 ^ x330 ;
  assign n5648 = n5647 ^ n5646 ;
  assign n5649 = n5648 ^ n5641 ;
  assign n5654 = n5653 ^ n5649 ;
  assign n5655 = n3656 & n5654 ;
  assign n5658 = n5655 ^ n5649 ;
  assign n5659 = n5658 ^ x298 ;
  assign n5660 = ~n3700 & n5659 ;
  assign n5661 = n5660 ^ x298 ;
  assign n5656 = n5655 ^ n5654 ;
  assign n5657 = n5656 ^ n5649 ;
  assign n5662 = n5661 ^ n5657 ;
  assign n5663 = n3739 & n5662 ;
  assign n5666 = n5663 ^ n5657 ;
  assign n5667 = n5666 ^ x266 ;
  assign n5668 = ~n3783 & n5667 ;
  assign n5669 = n5668 ^ x266 ;
  assign n5664 = n5663 ^ n5662 ;
  assign n5665 = n5664 ^ n5657 ;
  assign n5670 = n5669 ^ n5665 ;
  assign n5671 = ~n3818 & n5670 ;
  assign n5674 = n5671 ^ n5665 ;
  assign n5675 = n5674 ^ x234 ;
  assign n5676 = ~n3861 & n5675 ;
  assign n5677 = n5676 ^ x234 ;
  assign n5672 = n5671 ^ n5670 ;
  assign n5673 = n5672 ^ n5665 ;
  assign n5678 = n5677 ^ n5673 ;
  assign n5679 = n3897 & n5678 ;
  assign n5682 = n5679 ^ n5673 ;
  assign n5683 = n5682 ^ x202 ;
  assign n5684 = ~n3941 & n5683 ;
  assign n5685 = n5684 ^ x202 ;
  assign n5680 = n5679 ^ n5678 ;
  assign n5681 = n5680 ^ n5673 ;
  assign n5686 = n5685 ^ n5681 ;
  assign n5687 = n3980 & n5686 ;
  assign n5690 = n5687 ^ n5681 ;
  assign n5691 = n5690 ^ x170 ;
  assign n5692 = ~n4024 & n5691 ;
  assign n5693 = n5692 ^ x170 ;
  assign n5688 = n5687 ^ n5686 ;
  assign n5689 = n5688 ^ n5681 ;
  assign n5694 = n5693 ^ n5689 ;
  assign n5695 = ~n4059 & n5694 ;
  assign n5698 = n5695 ^ n5689 ;
  assign n5699 = n5698 ^ x138 ;
  assign n5700 = ~n4102 & n5699 ;
  assign n5701 = n5700 ^ x138 ;
  assign n5696 = n5695 ^ n5694 ;
  assign n5697 = n5696 ^ n5689 ;
  assign n5702 = n5701 ^ n5697 ;
  assign n5703 = n4138 & n5702 ;
  assign n5706 = n5703 ^ n5697 ;
  assign n5707 = n5706 ^ x106 ;
  assign n5708 = ~n4182 & n5707 ;
  assign n5709 = n5708 ^ x106 ;
  assign n5704 = n5703 ^ n5702 ;
  assign n5705 = n5704 ^ n5697 ;
  assign n5710 = n5709 ^ n5705 ;
  assign n5711 = n4221 & n5710 ;
  assign n5714 = n5711 ^ n5705 ;
  assign n5715 = n5714 ^ x74 ;
  assign n5716 = ~n4265 & n5715 ;
  assign n5717 = n5716 ^ x74 ;
  assign n5712 = n5711 ^ n5710 ;
  assign n5713 = n5712 ^ n5705 ;
  assign n5718 = n5717 ^ n5713 ;
  assign n5719 = ~n4300 & n5718 ;
  assign n5722 = n5719 ^ n5713 ;
  assign n5723 = n5722 ^ x42 ;
  assign n5724 = ~n4343 & n5723 ;
  assign n5725 = n5724 ^ x42 ;
  assign n5720 = n5719 ^ n5718 ;
  assign n5721 = n5720 ^ n5713 ;
  assign n5726 = n5725 ^ n5721 ;
  assign n5727 = n4379 & n5726 ;
  assign n5730 = n5727 ^ n5721 ;
  assign n5731 = n5730 ^ x10 ;
  assign n5732 = ~n4425 & n5731 ;
  assign n5733 = n5732 ^ x10 ;
  assign n5728 = n5727 ^ n5726 ;
  assign n5729 = n5728 ^ n5721 ;
  assign n5734 = n5733 ^ n5729 ;
  assign n5735 = ~n4461 & n5734 ;
  assign n5736 = n5735 ^ n5734 ;
  assign n5737 = n5736 ^ n5729 ;
  assign n5738 = x491 ^ x459 ;
  assign n5739 = ~n3330 & n5738 ;
  assign n5742 = n5739 ^ x459 ;
  assign n5743 = n5742 ^ x427 ;
  assign n5744 = ~n3377 & n5743 ;
  assign n5745 = n5744 ^ x427 ;
  assign n5740 = n5739 ^ n5738 ;
  assign n5741 = n5740 ^ x459 ;
  assign n5746 = n5745 ^ n5741 ;
  assign n5747 = ~n3413 & n5746 ;
  assign n5750 = n5747 ^ n5741 ;
  assign n5751 = n5750 ^ x395 ;
  assign n5752 = ~n3457 & n5751 ;
  assign n5753 = n5752 ^ x395 ;
  assign n5748 = n5747 ^ n5746 ;
  assign n5749 = n5748 ^ n5741 ;
  assign n5754 = n5753 ^ n5749 ;
  assign n5755 = ~n3493 & n5754 ;
  assign n5758 = n5755 ^ n5749 ;
  assign n5759 = n5758 ^ x363 ;
  assign n5760 = ~n3537 & n5759 ;
  assign n5761 = n5760 ^ x363 ;
  assign n5756 = n5755 ^ n5754 ;
  assign n5757 = n5756 ^ n5749 ;
  assign n5762 = n5761 ^ n5757 ;
  assign n5763 = n3577 & n5762 ;
  assign n5766 = n5763 ^ n5757 ;
  assign n5767 = n5766 ^ x331 ;
  assign n5768 = ~n3620 & n5767 ;
  assign n5769 = n5768 ^ x331 ;
  assign n5764 = n5763 ^ n5762 ;
  assign n5765 = n5764 ^ n5757 ;
  assign n5770 = n5769 ^ n5765 ;
  assign n5771 = n3656 & n5770 ;
  assign n5774 = n5771 ^ n5765 ;
  assign n5775 = n5774 ^ x299 ;
  assign n5776 = ~n3700 & n5775 ;
  assign n5777 = n5776 ^ x299 ;
  assign n5772 = n5771 ^ n5770 ;
  assign n5773 = n5772 ^ n5765 ;
  assign n5778 = n5777 ^ n5773 ;
  assign n5779 = n3739 & n5778 ;
  assign n5782 = n5779 ^ n5773 ;
  assign n5783 = n5782 ^ x267 ;
  assign n5784 = ~n3783 & n5783 ;
  assign n5785 = n5784 ^ x267 ;
  assign n5780 = n5779 ^ n5778 ;
  assign n5781 = n5780 ^ n5773 ;
  assign n5786 = n5785 ^ n5781 ;
  assign n5787 = ~n3818 & n5786 ;
  assign n5790 = n5787 ^ n5781 ;
  assign n5791 = n5790 ^ x235 ;
  assign n5792 = ~n3861 & n5791 ;
  assign n5793 = n5792 ^ x235 ;
  assign n5788 = n5787 ^ n5786 ;
  assign n5789 = n5788 ^ n5781 ;
  assign n5794 = n5793 ^ n5789 ;
  assign n5795 = n3897 & n5794 ;
  assign n5798 = n5795 ^ n5789 ;
  assign n5799 = n5798 ^ x203 ;
  assign n5800 = ~n3941 & n5799 ;
  assign n5801 = n5800 ^ x203 ;
  assign n5796 = n5795 ^ n5794 ;
  assign n5797 = n5796 ^ n5789 ;
  assign n5802 = n5801 ^ n5797 ;
  assign n5803 = n3980 & n5802 ;
  assign n5806 = n5803 ^ n5797 ;
  assign n5807 = n5806 ^ x171 ;
  assign n5808 = ~n4024 & n5807 ;
  assign n5809 = n5808 ^ x171 ;
  assign n5804 = n5803 ^ n5802 ;
  assign n5805 = n5804 ^ n5797 ;
  assign n5810 = n5809 ^ n5805 ;
  assign n5811 = ~n4059 & n5810 ;
  assign n5814 = n5811 ^ n5805 ;
  assign n5815 = n5814 ^ x139 ;
  assign n5816 = ~n4102 & n5815 ;
  assign n5817 = n5816 ^ x139 ;
  assign n5812 = n5811 ^ n5810 ;
  assign n5813 = n5812 ^ n5805 ;
  assign n5818 = n5817 ^ n5813 ;
  assign n5819 = n4138 & n5818 ;
  assign n5822 = n5819 ^ n5813 ;
  assign n5823 = n5822 ^ x107 ;
  assign n5824 = ~n4182 & n5823 ;
  assign n5825 = n5824 ^ x107 ;
  assign n5820 = n5819 ^ n5818 ;
  assign n5821 = n5820 ^ n5813 ;
  assign n5826 = n5825 ^ n5821 ;
  assign n5827 = n4221 & n5826 ;
  assign n5830 = n5827 ^ n5821 ;
  assign n5831 = n5830 ^ x75 ;
  assign n5832 = ~n4265 & n5831 ;
  assign n5833 = n5832 ^ x75 ;
  assign n5828 = n5827 ^ n5826 ;
  assign n5829 = n5828 ^ n5821 ;
  assign n5834 = n5833 ^ n5829 ;
  assign n5835 = ~n4300 & n5834 ;
  assign n5838 = n5835 ^ n5829 ;
  assign n5839 = n5838 ^ x43 ;
  assign n5840 = ~n4343 & n5839 ;
  assign n5841 = n5840 ^ x43 ;
  assign n5836 = n5835 ^ n5834 ;
  assign n5837 = n5836 ^ n5829 ;
  assign n5842 = n5841 ^ n5837 ;
  assign n5843 = n4379 & n5842 ;
  assign n5846 = n5843 ^ n5837 ;
  assign n5847 = n5846 ^ x11 ;
  assign n5848 = ~n4425 & n5847 ;
  assign n5849 = n5848 ^ x11 ;
  assign n5844 = n5843 ^ n5842 ;
  assign n5845 = n5844 ^ n5837 ;
  assign n5850 = n5849 ^ n5845 ;
  assign n5851 = ~n4461 & n5850 ;
  assign n5852 = n5851 ^ n5850 ;
  assign n5853 = n5852 ^ n5845 ;
  assign n5854 = x492 ^ x460 ;
  assign n5855 = ~n3330 & n5854 ;
  assign n5858 = n5855 ^ x460 ;
  assign n5859 = n5858 ^ x428 ;
  assign n5860 = ~n3377 & n5859 ;
  assign n5861 = n5860 ^ x428 ;
  assign n5856 = n5855 ^ n5854 ;
  assign n5857 = n5856 ^ x460 ;
  assign n5862 = n5861 ^ n5857 ;
  assign n5863 = ~n3413 & n5862 ;
  assign n5866 = n5863 ^ n5857 ;
  assign n5867 = n5866 ^ x396 ;
  assign n5868 = ~n3457 & n5867 ;
  assign n5869 = n5868 ^ x396 ;
  assign n5864 = n5863 ^ n5862 ;
  assign n5865 = n5864 ^ n5857 ;
  assign n5870 = n5869 ^ n5865 ;
  assign n5871 = ~n3493 & n5870 ;
  assign n5874 = n5871 ^ n5865 ;
  assign n5875 = n5874 ^ x364 ;
  assign n5876 = ~n3537 & n5875 ;
  assign n5877 = n5876 ^ x364 ;
  assign n5872 = n5871 ^ n5870 ;
  assign n5873 = n5872 ^ n5865 ;
  assign n5878 = n5877 ^ n5873 ;
  assign n5879 = n3577 & n5878 ;
  assign n5882 = n5879 ^ n5873 ;
  assign n5883 = n5882 ^ x332 ;
  assign n5884 = ~n3620 & n5883 ;
  assign n5885 = n5884 ^ x332 ;
  assign n5880 = n5879 ^ n5878 ;
  assign n5881 = n5880 ^ n5873 ;
  assign n5886 = n5885 ^ n5881 ;
  assign n5887 = n3656 & n5886 ;
  assign n5890 = n5887 ^ n5881 ;
  assign n5891 = n5890 ^ x300 ;
  assign n5892 = ~n3700 & n5891 ;
  assign n5893 = n5892 ^ x300 ;
  assign n5888 = n5887 ^ n5886 ;
  assign n5889 = n5888 ^ n5881 ;
  assign n5894 = n5893 ^ n5889 ;
  assign n5895 = n3739 & n5894 ;
  assign n5898 = n5895 ^ n5889 ;
  assign n5899 = n5898 ^ x268 ;
  assign n5900 = ~n3783 & n5899 ;
  assign n5901 = n5900 ^ x268 ;
  assign n5896 = n5895 ^ n5894 ;
  assign n5897 = n5896 ^ n5889 ;
  assign n5902 = n5901 ^ n5897 ;
  assign n5903 = ~n3818 & n5902 ;
  assign n5906 = n5903 ^ n5897 ;
  assign n5907 = n5906 ^ x236 ;
  assign n5908 = ~n3861 & n5907 ;
  assign n5909 = n5908 ^ x236 ;
  assign n5904 = n5903 ^ n5902 ;
  assign n5905 = n5904 ^ n5897 ;
  assign n5910 = n5909 ^ n5905 ;
  assign n5911 = n3897 & n5910 ;
  assign n5914 = n5911 ^ n5905 ;
  assign n5915 = n5914 ^ x204 ;
  assign n5916 = ~n3941 & n5915 ;
  assign n5917 = n5916 ^ x204 ;
  assign n5912 = n5911 ^ n5910 ;
  assign n5913 = n5912 ^ n5905 ;
  assign n5918 = n5917 ^ n5913 ;
  assign n5919 = n3980 & n5918 ;
  assign n5922 = n5919 ^ n5913 ;
  assign n5923 = n5922 ^ x172 ;
  assign n5924 = ~n4024 & n5923 ;
  assign n5925 = n5924 ^ x172 ;
  assign n5920 = n5919 ^ n5918 ;
  assign n5921 = n5920 ^ n5913 ;
  assign n5926 = n5925 ^ n5921 ;
  assign n5927 = ~n4059 & n5926 ;
  assign n5930 = n5927 ^ n5921 ;
  assign n5931 = n5930 ^ x140 ;
  assign n5932 = ~n4102 & n5931 ;
  assign n5933 = n5932 ^ x140 ;
  assign n5928 = n5927 ^ n5926 ;
  assign n5929 = n5928 ^ n5921 ;
  assign n5934 = n5933 ^ n5929 ;
  assign n5935 = n4138 & n5934 ;
  assign n5938 = n5935 ^ n5929 ;
  assign n5939 = n5938 ^ x108 ;
  assign n5940 = ~n4182 & n5939 ;
  assign n5941 = n5940 ^ x108 ;
  assign n5936 = n5935 ^ n5934 ;
  assign n5937 = n5936 ^ n5929 ;
  assign n5942 = n5941 ^ n5937 ;
  assign n5943 = n4221 & n5942 ;
  assign n5946 = n5943 ^ n5937 ;
  assign n5947 = n5946 ^ x76 ;
  assign n5948 = ~n4265 & n5947 ;
  assign n5949 = n5948 ^ x76 ;
  assign n5944 = n5943 ^ n5942 ;
  assign n5945 = n5944 ^ n5937 ;
  assign n5950 = n5949 ^ n5945 ;
  assign n5951 = ~n4300 & n5950 ;
  assign n5954 = n5951 ^ n5945 ;
  assign n5955 = n5954 ^ x44 ;
  assign n5956 = ~n4343 & n5955 ;
  assign n5957 = n5956 ^ x44 ;
  assign n5952 = n5951 ^ n5950 ;
  assign n5953 = n5952 ^ n5945 ;
  assign n5958 = n5957 ^ n5953 ;
  assign n5959 = n4379 & n5958 ;
  assign n5962 = n5959 ^ n5953 ;
  assign n5963 = n5962 ^ x12 ;
  assign n5964 = ~n4425 & n5963 ;
  assign n5965 = n5964 ^ x12 ;
  assign n5960 = n5959 ^ n5958 ;
  assign n5961 = n5960 ^ n5953 ;
  assign n5966 = n5965 ^ n5961 ;
  assign n5967 = ~n4461 & n5966 ;
  assign n5968 = n5967 ^ n5966 ;
  assign n5969 = n5968 ^ n5961 ;
  assign n5970 = x493 ^ x461 ;
  assign n5971 = ~n3330 & n5970 ;
  assign n5974 = n5971 ^ x461 ;
  assign n5975 = n5974 ^ x429 ;
  assign n5976 = ~n3377 & n5975 ;
  assign n5977 = n5976 ^ x429 ;
  assign n5972 = n5971 ^ n5970 ;
  assign n5973 = n5972 ^ x461 ;
  assign n5978 = n5977 ^ n5973 ;
  assign n5979 = ~n3413 & n5978 ;
  assign n5982 = n5979 ^ n5973 ;
  assign n5983 = n5982 ^ x397 ;
  assign n5984 = ~n3457 & n5983 ;
  assign n5985 = n5984 ^ x397 ;
  assign n5980 = n5979 ^ n5978 ;
  assign n5981 = n5980 ^ n5973 ;
  assign n5986 = n5985 ^ n5981 ;
  assign n5987 = ~n3493 & n5986 ;
  assign n5990 = n5987 ^ n5981 ;
  assign n5991 = n5990 ^ x365 ;
  assign n5992 = ~n3537 & n5991 ;
  assign n5993 = n5992 ^ x365 ;
  assign n5988 = n5987 ^ n5986 ;
  assign n5989 = n5988 ^ n5981 ;
  assign n5994 = n5993 ^ n5989 ;
  assign n5995 = n3577 & n5994 ;
  assign n5998 = n5995 ^ n5989 ;
  assign n5999 = n5998 ^ x333 ;
  assign n6000 = ~n3620 & n5999 ;
  assign n6001 = n6000 ^ x333 ;
  assign n5996 = n5995 ^ n5994 ;
  assign n5997 = n5996 ^ n5989 ;
  assign n6002 = n6001 ^ n5997 ;
  assign n6003 = n3656 & n6002 ;
  assign n6006 = n6003 ^ n5997 ;
  assign n6007 = n6006 ^ x301 ;
  assign n6008 = ~n3700 & n6007 ;
  assign n6009 = n6008 ^ x301 ;
  assign n6004 = n6003 ^ n6002 ;
  assign n6005 = n6004 ^ n5997 ;
  assign n6010 = n6009 ^ n6005 ;
  assign n6011 = n3739 & n6010 ;
  assign n6014 = n6011 ^ n6005 ;
  assign n6015 = n6014 ^ x269 ;
  assign n6016 = ~n3783 & n6015 ;
  assign n6017 = n6016 ^ x269 ;
  assign n6012 = n6011 ^ n6010 ;
  assign n6013 = n6012 ^ n6005 ;
  assign n6018 = n6017 ^ n6013 ;
  assign n6019 = ~n3818 & n6018 ;
  assign n6022 = n6019 ^ n6013 ;
  assign n6023 = n6022 ^ x237 ;
  assign n6024 = ~n3861 & n6023 ;
  assign n6025 = n6024 ^ x237 ;
  assign n6020 = n6019 ^ n6018 ;
  assign n6021 = n6020 ^ n6013 ;
  assign n6026 = n6025 ^ n6021 ;
  assign n6027 = n3897 & n6026 ;
  assign n6030 = n6027 ^ n6021 ;
  assign n6031 = n6030 ^ x205 ;
  assign n6032 = ~n3941 & n6031 ;
  assign n6033 = n6032 ^ x205 ;
  assign n6028 = n6027 ^ n6026 ;
  assign n6029 = n6028 ^ n6021 ;
  assign n6034 = n6033 ^ n6029 ;
  assign n6035 = n3980 & n6034 ;
  assign n6038 = n6035 ^ n6029 ;
  assign n6039 = n6038 ^ x173 ;
  assign n6040 = ~n4024 & n6039 ;
  assign n6041 = n6040 ^ x173 ;
  assign n6036 = n6035 ^ n6034 ;
  assign n6037 = n6036 ^ n6029 ;
  assign n6042 = n6041 ^ n6037 ;
  assign n6043 = ~n4059 & n6042 ;
  assign n6046 = n6043 ^ n6037 ;
  assign n6047 = n6046 ^ x141 ;
  assign n6048 = ~n4102 & n6047 ;
  assign n6049 = n6048 ^ x141 ;
  assign n6044 = n6043 ^ n6042 ;
  assign n6045 = n6044 ^ n6037 ;
  assign n6050 = n6049 ^ n6045 ;
  assign n6051 = n4138 & n6050 ;
  assign n6054 = n6051 ^ n6045 ;
  assign n6055 = n6054 ^ x109 ;
  assign n6056 = ~n4182 & n6055 ;
  assign n6057 = n6056 ^ x109 ;
  assign n6052 = n6051 ^ n6050 ;
  assign n6053 = n6052 ^ n6045 ;
  assign n6058 = n6057 ^ n6053 ;
  assign n6059 = n4221 & n6058 ;
  assign n6062 = n6059 ^ n6053 ;
  assign n6063 = n6062 ^ x77 ;
  assign n6064 = ~n4265 & n6063 ;
  assign n6065 = n6064 ^ x77 ;
  assign n6060 = n6059 ^ n6058 ;
  assign n6061 = n6060 ^ n6053 ;
  assign n6066 = n6065 ^ n6061 ;
  assign n6067 = ~n4300 & n6066 ;
  assign n6070 = n6067 ^ n6061 ;
  assign n6071 = n6070 ^ x45 ;
  assign n6072 = ~n4343 & n6071 ;
  assign n6073 = n6072 ^ x45 ;
  assign n6068 = n6067 ^ n6066 ;
  assign n6069 = n6068 ^ n6061 ;
  assign n6074 = n6073 ^ n6069 ;
  assign n6075 = n4379 & n6074 ;
  assign n6078 = n6075 ^ n6069 ;
  assign n6079 = n6078 ^ x13 ;
  assign n6080 = ~n4425 & n6079 ;
  assign n6081 = n6080 ^ x13 ;
  assign n6076 = n6075 ^ n6074 ;
  assign n6077 = n6076 ^ n6069 ;
  assign n6082 = n6081 ^ n6077 ;
  assign n6083 = ~n4461 & n6082 ;
  assign n6084 = n6083 ^ n6082 ;
  assign n6085 = n6084 ^ n6077 ;
  assign n6086 = x494 ^ x462 ;
  assign n6087 = ~n3330 & n6086 ;
  assign n6090 = n6087 ^ x462 ;
  assign n6091 = n6090 ^ x430 ;
  assign n6092 = ~n3377 & n6091 ;
  assign n6093 = n6092 ^ x430 ;
  assign n6088 = n6087 ^ n6086 ;
  assign n6089 = n6088 ^ x462 ;
  assign n6094 = n6093 ^ n6089 ;
  assign n6095 = ~n3413 & n6094 ;
  assign n6098 = n6095 ^ n6089 ;
  assign n6099 = n6098 ^ x398 ;
  assign n6100 = ~n3457 & n6099 ;
  assign n6101 = n6100 ^ x398 ;
  assign n6096 = n6095 ^ n6094 ;
  assign n6097 = n6096 ^ n6089 ;
  assign n6102 = n6101 ^ n6097 ;
  assign n6103 = ~n3493 & n6102 ;
  assign n6106 = n6103 ^ n6097 ;
  assign n6107 = n6106 ^ x366 ;
  assign n6108 = ~n3537 & n6107 ;
  assign n6109 = n6108 ^ x366 ;
  assign n6104 = n6103 ^ n6102 ;
  assign n6105 = n6104 ^ n6097 ;
  assign n6110 = n6109 ^ n6105 ;
  assign n6111 = n3577 & n6110 ;
  assign n6114 = n6111 ^ n6105 ;
  assign n6115 = n6114 ^ x334 ;
  assign n6116 = ~n3620 & n6115 ;
  assign n6117 = n6116 ^ x334 ;
  assign n6112 = n6111 ^ n6110 ;
  assign n6113 = n6112 ^ n6105 ;
  assign n6118 = n6117 ^ n6113 ;
  assign n6119 = n3656 & n6118 ;
  assign n6122 = n6119 ^ n6113 ;
  assign n6123 = n6122 ^ x302 ;
  assign n6124 = ~n3700 & n6123 ;
  assign n6125 = n6124 ^ x302 ;
  assign n6120 = n6119 ^ n6118 ;
  assign n6121 = n6120 ^ n6113 ;
  assign n6126 = n6125 ^ n6121 ;
  assign n6127 = n3739 & n6126 ;
  assign n6130 = n6127 ^ n6121 ;
  assign n6131 = n6130 ^ x270 ;
  assign n6132 = ~n3783 & n6131 ;
  assign n6133 = n6132 ^ x270 ;
  assign n6128 = n6127 ^ n6126 ;
  assign n6129 = n6128 ^ n6121 ;
  assign n6134 = n6133 ^ n6129 ;
  assign n6135 = ~n3818 & n6134 ;
  assign n6138 = n6135 ^ n6129 ;
  assign n6139 = n6138 ^ x238 ;
  assign n6140 = ~n3861 & n6139 ;
  assign n6141 = n6140 ^ x238 ;
  assign n6136 = n6135 ^ n6134 ;
  assign n6137 = n6136 ^ n6129 ;
  assign n6142 = n6141 ^ n6137 ;
  assign n6143 = n3897 & n6142 ;
  assign n6146 = n6143 ^ n6137 ;
  assign n6147 = n6146 ^ x206 ;
  assign n6148 = ~n3941 & n6147 ;
  assign n6149 = n6148 ^ x206 ;
  assign n6144 = n6143 ^ n6142 ;
  assign n6145 = n6144 ^ n6137 ;
  assign n6150 = n6149 ^ n6145 ;
  assign n6151 = n3980 & n6150 ;
  assign n6154 = n6151 ^ n6145 ;
  assign n6155 = n6154 ^ x174 ;
  assign n6156 = ~n4024 & n6155 ;
  assign n6157 = n6156 ^ x174 ;
  assign n6152 = n6151 ^ n6150 ;
  assign n6153 = n6152 ^ n6145 ;
  assign n6158 = n6157 ^ n6153 ;
  assign n6159 = ~n4059 & n6158 ;
  assign n6162 = n6159 ^ n6153 ;
  assign n6163 = n6162 ^ x142 ;
  assign n6164 = ~n4102 & n6163 ;
  assign n6165 = n6164 ^ x142 ;
  assign n6160 = n6159 ^ n6158 ;
  assign n6161 = n6160 ^ n6153 ;
  assign n6166 = n6165 ^ n6161 ;
  assign n6167 = n4138 & n6166 ;
  assign n6170 = n6167 ^ n6161 ;
  assign n6171 = n6170 ^ x110 ;
  assign n6172 = ~n4182 & n6171 ;
  assign n6173 = n6172 ^ x110 ;
  assign n6168 = n6167 ^ n6166 ;
  assign n6169 = n6168 ^ n6161 ;
  assign n6174 = n6173 ^ n6169 ;
  assign n6175 = n4221 & n6174 ;
  assign n6178 = n6175 ^ n6169 ;
  assign n6179 = n6178 ^ x78 ;
  assign n6180 = ~n4265 & n6179 ;
  assign n6181 = n6180 ^ x78 ;
  assign n6176 = n6175 ^ n6174 ;
  assign n6177 = n6176 ^ n6169 ;
  assign n6182 = n6181 ^ n6177 ;
  assign n6183 = ~n4300 & n6182 ;
  assign n6186 = n6183 ^ n6177 ;
  assign n6187 = n6186 ^ x46 ;
  assign n6188 = ~n4343 & n6187 ;
  assign n6189 = n6188 ^ x46 ;
  assign n6184 = n6183 ^ n6182 ;
  assign n6185 = n6184 ^ n6177 ;
  assign n6190 = n6189 ^ n6185 ;
  assign n6191 = n4379 & n6190 ;
  assign n6194 = n6191 ^ n6185 ;
  assign n6195 = n6194 ^ x14 ;
  assign n6196 = ~n4425 & n6195 ;
  assign n6197 = n6196 ^ x14 ;
  assign n6192 = n6191 ^ n6190 ;
  assign n6193 = n6192 ^ n6185 ;
  assign n6198 = n6197 ^ n6193 ;
  assign n6199 = ~n4461 & n6198 ;
  assign n6200 = n6199 ^ n6198 ;
  assign n6201 = n6200 ^ n6193 ;
  assign n6202 = x495 ^ x463 ;
  assign n6203 = ~n3330 & n6202 ;
  assign n6206 = n6203 ^ x463 ;
  assign n6207 = n6206 ^ x431 ;
  assign n6208 = ~n3377 & n6207 ;
  assign n6209 = n6208 ^ x431 ;
  assign n6204 = n6203 ^ n6202 ;
  assign n6205 = n6204 ^ x463 ;
  assign n6210 = n6209 ^ n6205 ;
  assign n6211 = ~n3413 & n6210 ;
  assign n6214 = n6211 ^ n6205 ;
  assign n6215 = n6214 ^ x399 ;
  assign n6216 = ~n3457 & n6215 ;
  assign n6217 = n6216 ^ x399 ;
  assign n6212 = n6211 ^ n6210 ;
  assign n6213 = n6212 ^ n6205 ;
  assign n6218 = n6217 ^ n6213 ;
  assign n6219 = ~n3493 & n6218 ;
  assign n6222 = n6219 ^ n6213 ;
  assign n6223 = n6222 ^ x367 ;
  assign n6224 = ~n3537 & n6223 ;
  assign n6225 = n6224 ^ x367 ;
  assign n6220 = n6219 ^ n6218 ;
  assign n6221 = n6220 ^ n6213 ;
  assign n6226 = n6225 ^ n6221 ;
  assign n6227 = n3577 & n6226 ;
  assign n6230 = n6227 ^ n6221 ;
  assign n6231 = n6230 ^ x335 ;
  assign n6232 = ~n3620 & n6231 ;
  assign n6233 = n6232 ^ x335 ;
  assign n6228 = n6227 ^ n6226 ;
  assign n6229 = n6228 ^ n6221 ;
  assign n6234 = n6233 ^ n6229 ;
  assign n6235 = n3656 & n6234 ;
  assign n6238 = n6235 ^ n6229 ;
  assign n6239 = n6238 ^ x303 ;
  assign n6240 = ~n3700 & n6239 ;
  assign n6241 = n6240 ^ x303 ;
  assign n6236 = n6235 ^ n6234 ;
  assign n6237 = n6236 ^ n6229 ;
  assign n6242 = n6241 ^ n6237 ;
  assign n6243 = n3739 & n6242 ;
  assign n6246 = n6243 ^ n6237 ;
  assign n6247 = n6246 ^ x271 ;
  assign n6248 = ~n3783 & n6247 ;
  assign n6249 = n6248 ^ x271 ;
  assign n6244 = n6243 ^ n6242 ;
  assign n6245 = n6244 ^ n6237 ;
  assign n6250 = n6249 ^ n6245 ;
  assign n6251 = ~n3818 & n6250 ;
  assign n6254 = n6251 ^ n6245 ;
  assign n6255 = n6254 ^ x239 ;
  assign n6256 = ~n3861 & n6255 ;
  assign n6257 = n6256 ^ x239 ;
  assign n6252 = n6251 ^ n6250 ;
  assign n6253 = n6252 ^ n6245 ;
  assign n6258 = n6257 ^ n6253 ;
  assign n6259 = n3897 & n6258 ;
  assign n6262 = n6259 ^ n6253 ;
  assign n6263 = n6262 ^ x207 ;
  assign n6264 = ~n3941 & n6263 ;
  assign n6265 = n6264 ^ x207 ;
  assign n6260 = n6259 ^ n6258 ;
  assign n6261 = n6260 ^ n6253 ;
  assign n6266 = n6265 ^ n6261 ;
  assign n6267 = n3980 & n6266 ;
  assign n6270 = n6267 ^ n6261 ;
  assign n6271 = n6270 ^ x175 ;
  assign n6272 = ~n4024 & n6271 ;
  assign n6273 = n6272 ^ x175 ;
  assign n6268 = n6267 ^ n6266 ;
  assign n6269 = n6268 ^ n6261 ;
  assign n6274 = n6273 ^ n6269 ;
  assign n6275 = ~n4059 & n6274 ;
  assign n6278 = n6275 ^ n6269 ;
  assign n6279 = n6278 ^ x143 ;
  assign n6280 = ~n4102 & n6279 ;
  assign n6281 = n6280 ^ x143 ;
  assign n6276 = n6275 ^ n6274 ;
  assign n6277 = n6276 ^ n6269 ;
  assign n6282 = n6281 ^ n6277 ;
  assign n6283 = n4138 & n6282 ;
  assign n6286 = n6283 ^ n6277 ;
  assign n6287 = n6286 ^ x111 ;
  assign n6288 = ~n4182 & n6287 ;
  assign n6289 = n6288 ^ x111 ;
  assign n6284 = n6283 ^ n6282 ;
  assign n6285 = n6284 ^ n6277 ;
  assign n6290 = n6289 ^ n6285 ;
  assign n6291 = n4221 & n6290 ;
  assign n6294 = n6291 ^ n6285 ;
  assign n6295 = n6294 ^ x79 ;
  assign n6296 = ~n4265 & n6295 ;
  assign n6297 = n6296 ^ x79 ;
  assign n6292 = n6291 ^ n6290 ;
  assign n6293 = n6292 ^ n6285 ;
  assign n6298 = n6297 ^ n6293 ;
  assign n6299 = ~n4300 & n6298 ;
  assign n6302 = n6299 ^ n6293 ;
  assign n6303 = n6302 ^ x47 ;
  assign n6304 = ~n4343 & n6303 ;
  assign n6305 = n6304 ^ x47 ;
  assign n6300 = n6299 ^ n6298 ;
  assign n6301 = n6300 ^ n6293 ;
  assign n6306 = n6305 ^ n6301 ;
  assign n6307 = n4379 & n6306 ;
  assign n6310 = n6307 ^ n6301 ;
  assign n6311 = n6310 ^ x15 ;
  assign n6312 = ~n4425 & n6311 ;
  assign n6313 = n6312 ^ x15 ;
  assign n6308 = n6307 ^ n6306 ;
  assign n6309 = n6308 ^ n6301 ;
  assign n6314 = n6313 ^ n6309 ;
  assign n6315 = ~n4461 & n6314 ;
  assign n6316 = n6315 ^ n6314 ;
  assign n6317 = n6316 ^ n6309 ;
  assign n6318 = x496 ^ x464 ;
  assign n6319 = ~n3330 & n6318 ;
  assign n6322 = n6319 ^ x464 ;
  assign n6323 = n6322 ^ x432 ;
  assign n6324 = ~n3377 & n6323 ;
  assign n6325 = n6324 ^ x432 ;
  assign n6320 = n6319 ^ n6318 ;
  assign n6321 = n6320 ^ x464 ;
  assign n6326 = n6325 ^ n6321 ;
  assign n6327 = ~n3413 & n6326 ;
  assign n6330 = n6327 ^ n6321 ;
  assign n6331 = n6330 ^ x400 ;
  assign n6332 = ~n3457 & n6331 ;
  assign n6333 = n6332 ^ x400 ;
  assign n6328 = n6327 ^ n6326 ;
  assign n6329 = n6328 ^ n6321 ;
  assign n6334 = n6333 ^ n6329 ;
  assign n6335 = ~n3493 & n6334 ;
  assign n6338 = n6335 ^ n6329 ;
  assign n6339 = n6338 ^ x368 ;
  assign n6340 = ~n3537 & n6339 ;
  assign n6341 = n6340 ^ x368 ;
  assign n6336 = n6335 ^ n6334 ;
  assign n6337 = n6336 ^ n6329 ;
  assign n6342 = n6341 ^ n6337 ;
  assign n6343 = n3577 & n6342 ;
  assign n6346 = n6343 ^ n6337 ;
  assign n6347 = n6346 ^ x336 ;
  assign n6348 = ~n3620 & n6347 ;
  assign n6349 = n6348 ^ x336 ;
  assign n6344 = n6343 ^ n6342 ;
  assign n6345 = n6344 ^ n6337 ;
  assign n6350 = n6349 ^ n6345 ;
  assign n6351 = n3656 & n6350 ;
  assign n6354 = n6351 ^ n6345 ;
  assign n6355 = n6354 ^ x304 ;
  assign n6356 = ~n3700 & n6355 ;
  assign n6357 = n6356 ^ x304 ;
  assign n6352 = n6351 ^ n6350 ;
  assign n6353 = n6352 ^ n6345 ;
  assign n6358 = n6357 ^ n6353 ;
  assign n6359 = n3739 & n6358 ;
  assign n6362 = n6359 ^ n6353 ;
  assign n6363 = n6362 ^ x272 ;
  assign n6364 = ~n3783 & n6363 ;
  assign n6365 = n6364 ^ x272 ;
  assign n6360 = n6359 ^ n6358 ;
  assign n6361 = n6360 ^ n6353 ;
  assign n6366 = n6365 ^ n6361 ;
  assign n6367 = ~n3818 & n6366 ;
  assign n6370 = n6367 ^ n6361 ;
  assign n6371 = n6370 ^ x240 ;
  assign n6372 = ~n3861 & n6371 ;
  assign n6373 = n6372 ^ x240 ;
  assign n6368 = n6367 ^ n6366 ;
  assign n6369 = n6368 ^ n6361 ;
  assign n6374 = n6373 ^ n6369 ;
  assign n6375 = n3897 & n6374 ;
  assign n6378 = n6375 ^ n6369 ;
  assign n6379 = n6378 ^ x208 ;
  assign n6380 = ~n3941 & n6379 ;
  assign n6381 = n6380 ^ x208 ;
  assign n6376 = n6375 ^ n6374 ;
  assign n6377 = n6376 ^ n6369 ;
  assign n6382 = n6381 ^ n6377 ;
  assign n6383 = n3980 & n6382 ;
  assign n6386 = n6383 ^ n6377 ;
  assign n6387 = n6386 ^ x176 ;
  assign n6388 = ~n4024 & n6387 ;
  assign n6389 = n6388 ^ x176 ;
  assign n6384 = n6383 ^ n6382 ;
  assign n6385 = n6384 ^ n6377 ;
  assign n6390 = n6389 ^ n6385 ;
  assign n6391 = ~n4059 & n6390 ;
  assign n6394 = n6391 ^ n6385 ;
  assign n6395 = n6394 ^ x144 ;
  assign n6396 = ~n4102 & n6395 ;
  assign n6397 = n6396 ^ x144 ;
  assign n6392 = n6391 ^ n6390 ;
  assign n6393 = n6392 ^ n6385 ;
  assign n6398 = n6397 ^ n6393 ;
  assign n6399 = n4138 & n6398 ;
  assign n6402 = n6399 ^ n6393 ;
  assign n6403 = n6402 ^ x112 ;
  assign n6404 = ~n4182 & n6403 ;
  assign n6405 = n6404 ^ x112 ;
  assign n6400 = n6399 ^ n6398 ;
  assign n6401 = n6400 ^ n6393 ;
  assign n6406 = n6405 ^ n6401 ;
  assign n6407 = n4221 & n6406 ;
  assign n6410 = n6407 ^ n6401 ;
  assign n6411 = n6410 ^ x80 ;
  assign n6412 = ~n4265 & n6411 ;
  assign n6413 = n6412 ^ x80 ;
  assign n6408 = n6407 ^ n6406 ;
  assign n6409 = n6408 ^ n6401 ;
  assign n6414 = n6413 ^ n6409 ;
  assign n6415 = ~n4300 & n6414 ;
  assign n6418 = n6415 ^ n6409 ;
  assign n6419 = n6418 ^ x48 ;
  assign n6420 = ~n4343 & n6419 ;
  assign n6421 = n6420 ^ x48 ;
  assign n6416 = n6415 ^ n6414 ;
  assign n6417 = n6416 ^ n6409 ;
  assign n6422 = n6421 ^ n6417 ;
  assign n6423 = n4379 & n6422 ;
  assign n6426 = n6423 ^ n6417 ;
  assign n6427 = n6426 ^ x16 ;
  assign n6428 = ~n4425 & n6427 ;
  assign n6429 = n6428 ^ x16 ;
  assign n6424 = n6423 ^ n6422 ;
  assign n6425 = n6424 ^ n6417 ;
  assign n6430 = n6429 ^ n6425 ;
  assign n6431 = ~n4461 & n6430 ;
  assign n6432 = n6431 ^ n6430 ;
  assign n6433 = n6432 ^ n6425 ;
  assign n6434 = x497 ^ x465 ;
  assign n6435 = ~n3330 & n6434 ;
  assign n6438 = n6435 ^ x465 ;
  assign n6439 = n6438 ^ x433 ;
  assign n6440 = ~n3377 & n6439 ;
  assign n6441 = n6440 ^ x433 ;
  assign n6436 = n6435 ^ n6434 ;
  assign n6437 = n6436 ^ x465 ;
  assign n6442 = n6441 ^ n6437 ;
  assign n6443 = ~n3413 & n6442 ;
  assign n6446 = n6443 ^ n6437 ;
  assign n6447 = n6446 ^ x401 ;
  assign n6448 = ~n3457 & n6447 ;
  assign n6449 = n6448 ^ x401 ;
  assign n6444 = n6443 ^ n6442 ;
  assign n6445 = n6444 ^ n6437 ;
  assign n6450 = n6449 ^ n6445 ;
  assign n6451 = ~n3493 & n6450 ;
  assign n6454 = n6451 ^ n6445 ;
  assign n6455 = n6454 ^ x369 ;
  assign n6456 = ~n3537 & n6455 ;
  assign n6457 = n6456 ^ x369 ;
  assign n6452 = n6451 ^ n6450 ;
  assign n6453 = n6452 ^ n6445 ;
  assign n6458 = n6457 ^ n6453 ;
  assign n6459 = n3577 & n6458 ;
  assign n6462 = n6459 ^ n6453 ;
  assign n6463 = n6462 ^ x337 ;
  assign n6464 = ~n3620 & n6463 ;
  assign n6465 = n6464 ^ x337 ;
  assign n6460 = n6459 ^ n6458 ;
  assign n6461 = n6460 ^ n6453 ;
  assign n6466 = n6465 ^ n6461 ;
  assign n6467 = n3656 & n6466 ;
  assign n6470 = n6467 ^ n6461 ;
  assign n6471 = n6470 ^ x305 ;
  assign n6472 = ~n3700 & n6471 ;
  assign n6473 = n6472 ^ x305 ;
  assign n6468 = n6467 ^ n6466 ;
  assign n6469 = n6468 ^ n6461 ;
  assign n6474 = n6473 ^ n6469 ;
  assign n6475 = n3739 & n6474 ;
  assign n6478 = n6475 ^ n6469 ;
  assign n6479 = n6478 ^ x273 ;
  assign n6480 = ~n3783 & n6479 ;
  assign n6481 = n6480 ^ x273 ;
  assign n6476 = n6475 ^ n6474 ;
  assign n6477 = n6476 ^ n6469 ;
  assign n6482 = n6481 ^ n6477 ;
  assign n6483 = ~n3818 & n6482 ;
  assign n6486 = n6483 ^ n6477 ;
  assign n6487 = n6486 ^ x241 ;
  assign n6488 = ~n3861 & n6487 ;
  assign n6489 = n6488 ^ x241 ;
  assign n6484 = n6483 ^ n6482 ;
  assign n6485 = n6484 ^ n6477 ;
  assign n6490 = n6489 ^ n6485 ;
  assign n6491 = n3897 & n6490 ;
  assign n6494 = n6491 ^ n6485 ;
  assign n6495 = n6494 ^ x209 ;
  assign n6496 = ~n3941 & n6495 ;
  assign n6497 = n6496 ^ x209 ;
  assign n6492 = n6491 ^ n6490 ;
  assign n6493 = n6492 ^ n6485 ;
  assign n6498 = n6497 ^ n6493 ;
  assign n6499 = n3980 & n6498 ;
  assign n6502 = n6499 ^ n6493 ;
  assign n6503 = n6502 ^ x177 ;
  assign n6504 = ~n4024 & n6503 ;
  assign n6505 = n6504 ^ x177 ;
  assign n6500 = n6499 ^ n6498 ;
  assign n6501 = n6500 ^ n6493 ;
  assign n6506 = n6505 ^ n6501 ;
  assign n6507 = ~n4059 & n6506 ;
  assign n6510 = n6507 ^ n6501 ;
  assign n6511 = n6510 ^ x145 ;
  assign n6512 = ~n4102 & n6511 ;
  assign n6513 = n6512 ^ x145 ;
  assign n6508 = n6507 ^ n6506 ;
  assign n6509 = n6508 ^ n6501 ;
  assign n6514 = n6513 ^ n6509 ;
  assign n6515 = n4138 & n6514 ;
  assign n6518 = n6515 ^ n6509 ;
  assign n6519 = n6518 ^ x113 ;
  assign n6520 = ~n4182 & n6519 ;
  assign n6521 = n6520 ^ x113 ;
  assign n6516 = n6515 ^ n6514 ;
  assign n6517 = n6516 ^ n6509 ;
  assign n6522 = n6521 ^ n6517 ;
  assign n6523 = n4221 & n6522 ;
  assign n6526 = n6523 ^ n6517 ;
  assign n6527 = n6526 ^ x81 ;
  assign n6528 = ~n4265 & n6527 ;
  assign n6529 = n6528 ^ x81 ;
  assign n6524 = n6523 ^ n6522 ;
  assign n6525 = n6524 ^ n6517 ;
  assign n6530 = n6529 ^ n6525 ;
  assign n6531 = ~n4300 & n6530 ;
  assign n6534 = n6531 ^ n6525 ;
  assign n6535 = n6534 ^ x49 ;
  assign n6536 = ~n4343 & n6535 ;
  assign n6537 = n6536 ^ x49 ;
  assign n6532 = n6531 ^ n6530 ;
  assign n6533 = n6532 ^ n6525 ;
  assign n6538 = n6537 ^ n6533 ;
  assign n6539 = n4379 & n6538 ;
  assign n6542 = n6539 ^ n6533 ;
  assign n6543 = n6542 ^ x17 ;
  assign n6544 = ~n4425 & n6543 ;
  assign n6545 = n6544 ^ x17 ;
  assign n6540 = n6539 ^ n6538 ;
  assign n6541 = n6540 ^ n6533 ;
  assign n6546 = n6545 ^ n6541 ;
  assign n6547 = ~n4461 & n6546 ;
  assign n6548 = n6547 ^ n6546 ;
  assign n6549 = n6548 ^ n6541 ;
  assign n6550 = x498 ^ x466 ;
  assign n6551 = ~n3330 & n6550 ;
  assign n6554 = n6551 ^ x466 ;
  assign n6555 = n6554 ^ x434 ;
  assign n6556 = ~n3377 & n6555 ;
  assign n6557 = n6556 ^ x434 ;
  assign n6552 = n6551 ^ n6550 ;
  assign n6553 = n6552 ^ x466 ;
  assign n6558 = n6557 ^ n6553 ;
  assign n6559 = ~n3413 & n6558 ;
  assign n6562 = n6559 ^ n6553 ;
  assign n6563 = n6562 ^ x402 ;
  assign n6564 = ~n3457 & n6563 ;
  assign n6565 = n6564 ^ x402 ;
  assign n6560 = n6559 ^ n6558 ;
  assign n6561 = n6560 ^ n6553 ;
  assign n6566 = n6565 ^ n6561 ;
  assign n6567 = ~n3493 & n6566 ;
  assign n6570 = n6567 ^ n6561 ;
  assign n6571 = n6570 ^ x370 ;
  assign n6572 = ~n3537 & n6571 ;
  assign n6573 = n6572 ^ x370 ;
  assign n6568 = n6567 ^ n6566 ;
  assign n6569 = n6568 ^ n6561 ;
  assign n6574 = n6573 ^ n6569 ;
  assign n6575 = n3577 & n6574 ;
  assign n6578 = n6575 ^ n6569 ;
  assign n6579 = n6578 ^ x338 ;
  assign n6580 = ~n3620 & n6579 ;
  assign n6581 = n6580 ^ x338 ;
  assign n6576 = n6575 ^ n6574 ;
  assign n6577 = n6576 ^ n6569 ;
  assign n6582 = n6581 ^ n6577 ;
  assign n6583 = n3656 & n6582 ;
  assign n6586 = n6583 ^ n6577 ;
  assign n6587 = n6586 ^ x306 ;
  assign n6588 = ~n3700 & n6587 ;
  assign n6589 = n6588 ^ x306 ;
  assign n6584 = n6583 ^ n6582 ;
  assign n6585 = n6584 ^ n6577 ;
  assign n6590 = n6589 ^ n6585 ;
  assign n6591 = n3739 & n6590 ;
  assign n6594 = n6591 ^ n6585 ;
  assign n6595 = n6594 ^ x274 ;
  assign n6596 = ~n3783 & n6595 ;
  assign n6597 = n6596 ^ x274 ;
  assign n6592 = n6591 ^ n6590 ;
  assign n6593 = n6592 ^ n6585 ;
  assign n6598 = n6597 ^ n6593 ;
  assign n6599 = ~n3818 & n6598 ;
  assign n6602 = n6599 ^ n6593 ;
  assign n6603 = n6602 ^ x242 ;
  assign n6604 = ~n3861 & n6603 ;
  assign n6605 = n6604 ^ x242 ;
  assign n6600 = n6599 ^ n6598 ;
  assign n6601 = n6600 ^ n6593 ;
  assign n6606 = n6605 ^ n6601 ;
  assign n6607 = n3897 & n6606 ;
  assign n6610 = n6607 ^ n6601 ;
  assign n6611 = n6610 ^ x210 ;
  assign n6612 = ~n3941 & n6611 ;
  assign n6613 = n6612 ^ x210 ;
  assign n6608 = n6607 ^ n6606 ;
  assign n6609 = n6608 ^ n6601 ;
  assign n6614 = n6613 ^ n6609 ;
  assign n6615 = n3980 & n6614 ;
  assign n6618 = n6615 ^ n6609 ;
  assign n6619 = n6618 ^ x178 ;
  assign n6620 = ~n4024 & n6619 ;
  assign n6621 = n6620 ^ x178 ;
  assign n6616 = n6615 ^ n6614 ;
  assign n6617 = n6616 ^ n6609 ;
  assign n6622 = n6621 ^ n6617 ;
  assign n6623 = ~n4059 & n6622 ;
  assign n6626 = n6623 ^ n6617 ;
  assign n6627 = n6626 ^ x146 ;
  assign n6628 = ~n4102 & n6627 ;
  assign n6629 = n6628 ^ x146 ;
  assign n6624 = n6623 ^ n6622 ;
  assign n6625 = n6624 ^ n6617 ;
  assign n6630 = n6629 ^ n6625 ;
  assign n6631 = n4138 & n6630 ;
  assign n6634 = n6631 ^ n6625 ;
  assign n6635 = n6634 ^ x114 ;
  assign n6636 = ~n4182 & n6635 ;
  assign n6637 = n6636 ^ x114 ;
  assign n6632 = n6631 ^ n6630 ;
  assign n6633 = n6632 ^ n6625 ;
  assign n6638 = n6637 ^ n6633 ;
  assign n6639 = n4221 & n6638 ;
  assign n6642 = n6639 ^ n6633 ;
  assign n6643 = n6642 ^ x82 ;
  assign n6644 = ~n4265 & n6643 ;
  assign n6645 = n6644 ^ x82 ;
  assign n6640 = n6639 ^ n6638 ;
  assign n6641 = n6640 ^ n6633 ;
  assign n6646 = n6645 ^ n6641 ;
  assign n6647 = ~n4300 & n6646 ;
  assign n6650 = n6647 ^ n6641 ;
  assign n6651 = n6650 ^ x50 ;
  assign n6652 = ~n4343 & n6651 ;
  assign n6653 = n6652 ^ x50 ;
  assign n6648 = n6647 ^ n6646 ;
  assign n6649 = n6648 ^ n6641 ;
  assign n6654 = n6653 ^ n6649 ;
  assign n6655 = n4379 & n6654 ;
  assign n6658 = n6655 ^ n6649 ;
  assign n6659 = n6658 ^ x18 ;
  assign n6660 = ~n4425 & n6659 ;
  assign n6661 = n6660 ^ x18 ;
  assign n6656 = n6655 ^ n6654 ;
  assign n6657 = n6656 ^ n6649 ;
  assign n6662 = n6661 ^ n6657 ;
  assign n6663 = ~n4461 & n6662 ;
  assign n6664 = n6663 ^ n6662 ;
  assign n6665 = n6664 ^ n6657 ;
  assign n6666 = x499 ^ x467 ;
  assign n6667 = ~n3330 & n6666 ;
  assign n6670 = n6667 ^ x467 ;
  assign n6671 = n6670 ^ x435 ;
  assign n6672 = ~n3377 & n6671 ;
  assign n6673 = n6672 ^ x435 ;
  assign n6668 = n6667 ^ n6666 ;
  assign n6669 = n6668 ^ x467 ;
  assign n6674 = n6673 ^ n6669 ;
  assign n6675 = ~n3413 & n6674 ;
  assign n6678 = n6675 ^ n6669 ;
  assign n6679 = n6678 ^ x403 ;
  assign n6680 = ~n3457 & n6679 ;
  assign n6681 = n6680 ^ x403 ;
  assign n6676 = n6675 ^ n6674 ;
  assign n6677 = n6676 ^ n6669 ;
  assign n6682 = n6681 ^ n6677 ;
  assign n6683 = ~n3493 & n6682 ;
  assign n6686 = n6683 ^ n6677 ;
  assign n6687 = n6686 ^ x371 ;
  assign n6688 = ~n3537 & n6687 ;
  assign n6689 = n6688 ^ x371 ;
  assign n6684 = n6683 ^ n6682 ;
  assign n6685 = n6684 ^ n6677 ;
  assign n6690 = n6689 ^ n6685 ;
  assign n6691 = n3577 & n6690 ;
  assign n6694 = n6691 ^ n6685 ;
  assign n6695 = n6694 ^ x339 ;
  assign n6696 = ~n3620 & n6695 ;
  assign n6697 = n6696 ^ x339 ;
  assign n6692 = n6691 ^ n6690 ;
  assign n6693 = n6692 ^ n6685 ;
  assign n6698 = n6697 ^ n6693 ;
  assign n6699 = n3656 & n6698 ;
  assign n6702 = n6699 ^ n6693 ;
  assign n6703 = n6702 ^ x307 ;
  assign n6704 = ~n3700 & n6703 ;
  assign n6705 = n6704 ^ x307 ;
  assign n6700 = n6699 ^ n6698 ;
  assign n6701 = n6700 ^ n6693 ;
  assign n6706 = n6705 ^ n6701 ;
  assign n6707 = n3739 & n6706 ;
  assign n6710 = n6707 ^ n6701 ;
  assign n6711 = n6710 ^ x275 ;
  assign n6712 = ~n3783 & n6711 ;
  assign n6713 = n6712 ^ x275 ;
  assign n6708 = n6707 ^ n6706 ;
  assign n6709 = n6708 ^ n6701 ;
  assign n6714 = n6713 ^ n6709 ;
  assign n6715 = ~n3818 & n6714 ;
  assign n6718 = n6715 ^ n6709 ;
  assign n6719 = n6718 ^ x243 ;
  assign n6720 = ~n3861 & n6719 ;
  assign n6721 = n6720 ^ x243 ;
  assign n6716 = n6715 ^ n6714 ;
  assign n6717 = n6716 ^ n6709 ;
  assign n6722 = n6721 ^ n6717 ;
  assign n6723 = n3897 & n6722 ;
  assign n6726 = n6723 ^ n6717 ;
  assign n6727 = n6726 ^ x211 ;
  assign n6728 = ~n3941 & n6727 ;
  assign n6729 = n6728 ^ x211 ;
  assign n6724 = n6723 ^ n6722 ;
  assign n6725 = n6724 ^ n6717 ;
  assign n6730 = n6729 ^ n6725 ;
  assign n6731 = n3980 & n6730 ;
  assign n6734 = n6731 ^ n6725 ;
  assign n6735 = n6734 ^ x179 ;
  assign n6736 = ~n4024 & n6735 ;
  assign n6737 = n6736 ^ x179 ;
  assign n6732 = n6731 ^ n6730 ;
  assign n6733 = n6732 ^ n6725 ;
  assign n6738 = n6737 ^ n6733 ;
  assign n6739 = ~n4059 & n6738 ;
  assign n6742 = n6739 ^ n6733 ;
  assign n6743 = n6742 ^ x147 ;
  assign n6744 = ~n4102 & n6743 ;
  assign n6745 = n6744 ^ x147 ;
  assign n6740 = n6739 ^ n6738 ;
  assign n6741 = n6740 ^ n6733 ;
  assign n6746 = n6745 ^ n6741 ;
  assign n6747 = n4138 & n6746 ;
  assign n6750 = n6747 ^ n6741 ;
  assign n6751 = n6750 ^ x115 ;
  assign n6752 = ~n4182 & n6751 ;
  assign n6753 = n6752 ^ x115 ;
  assign n6748 = n6747 ^ n6746 ;
  assign n6749 = n6748 ^ n6741 ;
  assign n6754 = n6753 ^ n6749 ;
  assign n6755 = n4221 & n6754 ;
  assign n6758 = n6755 ^ n6749 ;
  assign n6759 = n6758 ^ x83 ;
  assign n6760 = ~n4265 & n6759 ;
  assign n6761 = n6760 ^ x83 ;
  assign n6756 = n6755 ^ n6754 ;
  assign n6757 = n6756 ^ n6749 ;
  assign n6762 = n6761 ^ n6757 ;
  assign n6763 = ~n4300 & n6762 ;
  assign n6766 = n6763 ^ n6757 ;
  assign n6767 = n6766 ^ x51 ;
  assign n6768 = ~n4343 & n6767 ;
  assign n6769 = n6768 ^ x51 ;
  assign n6764 = n6763 ^ n6762 ;
  assign n6765 = n6764 ^ n6757 ;
  assign n6770 = n6769 ^ n6765 ;
  assign n6771 = n4379 & n6770 ;
  assign n6774 = n6771 ^ n6765 ;
  assign n6775 = n6774 ^ x19 ;
  assign n6776 = ~n4425 & n6775 ;
  assign n6777 = n6776 ^ x19 ;
  assign n6772 = n6771 ^ n6770 ;
  assign n6773 = n6772 ^ n6765 ;
  assign n6778 = n6777 ^ n6773 ;
  assign n6779 = ~n4461 & n6778 ;
  assign n6780 = n6779 ^ n6778 ;
  assign n6781 = n6780 ^ n6773 ;
  assign n6782 = x500 ^ x468 ;
  assign n6783 = ~n3330 & n6782 ;
  assign n6786 = n6783 ^ x468 ;
  assign n6787 = n6786 ^ x436 ;
  assign n6788 = ~n3377 & n6787 ;
  assign n6789 = n6788 ^ x436 ;
  assign n6784 = n6783 ^ n6782 ;
  assign n6785 = n6784 ^ x468 ;
  assign n6790 = n6789 ^ n6785 ;
  assign n6791 = ~n3413 & n6790 ;
  assign n6794 = n6791 ^ n6785 ;
  assign n6795 = n6794 ^ x404 ;
  assign n6796 = ~n3457 & n6795 ;
  assign n6797 = n6796 ^ x404 ;
  assign n6792 = n6791 ^ n6790 ;
  assign n6793 = n6792 ^ n6785 ;
  assign n6798 = n6797 ^ n6793 ;
  assign n6799 = ~n3493 & n6798 ;
  assign n6802 = n6799 ^ n6793 ;
  assign n6803 = n6802 ^ x372 ;
  assign n6804 = ~n3537 & n6803 ;
  assign n6805 = n6804 ^ x372 ;
  assign n6800 = n6799 ^ n6798 ;
  assign n6801 = n6800 ^ n6793 ;
  assign n6806 = n6805 ^ n6801 ;
  assign n6807 = n3577 & n6806 ;
  assign n6810 = n6807 ^ n6801 ;
  assign n6811 = n6810 ^ x340 ;
  assign n6812 = ~n3620 & n6811 ;
  assign n6813 = n6812 ^ x340 ;
  assign n6808 = n6807 ^ n6806 ;
  assign n6809 = n6808 ^ n6801 ;
  assign n6814 = n6813 ^ n6809 ;
  assign n6815 = n3656 & n6814 ;
  assign n6818 = n6815 ^ n6809 ;
  assign n6819 = n6818 ^ x308 ;
  assign n6820 = ~n3700 & n6819 ;
  assign n6821 = n6820 ^ x308 ;
  assign n6816 = n6815 ^ n6814 ;
  assign n6817 = n6816 ^ n6809 ;
  assign n6822 = n6821 ^ n6817 ;
  assign n6823 = n3739 & n6822 ;
  assign n6826 = n6823 ^ n6817 ;
  assign n6827 = n6826 ^ x276 ;
  assign n6828 = ~n3783 & n6827 ;
  assign n6829 = n6828 ^ x276 ;
  assign n6824 = n6823 ^ n6822 ;
  assign n6825 = n6824 ^ n6817 ;
  assign n6830 = n6829 ^ n6825 ;
  assign n6831 = ~n3818 & n6830 ;
  assign n6834 = n6831 ^ n6825 ;
  assign n6835 = n6834 ^ x244 ;
  assign n6836 = ~n3861 & n6835 ;
  assign n6837 = n6836 ^ x244 ;
  assign n6832 = n6831 ^ n6830 ;
  assign n6833 = n6832 ^ n6825 ;
  assign n6838 = n6837 ^ n6833 ;
  assign n6839 = n3897 & n6838 ;
  assign n6842 = n6839 ^ n6833 ;
  assign n6843 = n6842 ^ x212 ;
  assign n6844 = ~n3941 & n6843 ;
  assign n6845 = n6844 ^ x212 ;
  assign n6840 = n6839 ^ n6838 ;
  assign n6841 = n6840 ^ n6833 ;
  assign n6846 = n6845 ^ n6841 ;
  assign n6847 = n3980 & n6846 ;
  assign n6850 = n6847 ^ n6841 ;
  assign n6851 = n6850 ^ x180 ;
  assign n6852 = ~n4024 & n6851 ;
  assign n6853 = n6852 ^ x180 ;
  assign n6848 = n6847 ^ n6846 ;
  assign n6849 = n6848 ^ n6841 ;
  assign n6854 = n6853 ^ n6849 ;
  assign n6855 = ~n4059 & n6854 ;
  assign n6858 = n6855 ^ n6849 ;
  assign n6859 = n6858 ^ x148 ;
  assign n6860 = ~n4102 & n6859 ;
  assign n6861 = n6860 ^ x148 ;
  assign n6856 = n6855 ^ n6854 ;
  assign n6857 = n6856 ^ n6849 ;
  assign n6862 = n6861 ^ n6857 ;
  assign n6863 = n4138 & n6862 ;
  assign n6866 = n6863 ^ n6857 ;
  assign n6867 = n6866 ^ x116 ;
  assign n6868 = ~n4182 & n6867 ;
  assign n6869 = n6868 ^ x116 ;
  assign n6864 = n6863 ^ n6862 ;
  assign n6865 = n6864 ^ n6857 ;
  assign n6870 = n6869 ^ n6865 ;
  assign n6871 = n4221 & n6870 ;
  assign n6874 = n6871 ^ n6865 ;
  assign n6875 = n6874 ^ x84 ;
  assign n6876 = ~n4265 & n6875 ;
  assign n6877 = n6876 ^ x84 ;
  assign n6872 = n6871 ^ n6870 ;
  assign n6873 = n6872 ^ n6865 ;
  assign n6878 = n6877 ^ n6873 ;
  assign n6879 = ~n4300 & n6878 ;
  assign n6882 = n6879 ^ n6873 ;
  assign n6883 = n6882 ^ x52 ;
  assign n6884 = ~n4343 & n6883 ;
  assign n6885 = n6884 ^ x52 ;
  assign n6880 = n6879 ^ n6878 ;
  assign n6881 = n6880 ^ n6873 ;
  assign n6886 = n6885 ^ n6881 ;
  assign n6887 = n4379 & n6886 ;
  assign n6890 = n6887 ^ n6881 ;
  assign n6891 = n6890 ^ x20 ;
  assign n6892 = ~n4425 & n6891 ;
  assign n6893 = n6892 ^ x20 ;
  assign n6888 = n6887 ^ n6886 ;
  assign n6889 = n6888 ^ n6881 ;
  assign n6894 = n6893 ^ n6889 ;
  assign n6895 = ~n4461 & n6894 ;
  assign n6896 = n6895 ^ n6894 ;
  assign n6897 = n6896 ^ n6889 ;
  assign n6898 = x501 ^ x469 ;
  assign n6899 = ~n3330 & n6898 ;
  assign n6902 = n6899 ^ x469 ;
  assign n6903 = n6902 ^ x437 ;
  assign n6904 = ~n3377 & n6903 ;
  assign n6905 = n6904 ^ x437 ;
  assign n6900 = n6899 ^ n6898 ;
  assign n6901 = n6900 ^ x469 ;
  assign n6906 = n6905 ^ n6901 ;
  assign n6907 = ~n3413 & n6906 ;
  assign n6910 = n6907 ^ n6901 ;
  assign n6911 = n6910 ^ x405 ;
  assign n6912 = ~n3457 & n6911 ;
  assign n6913 = n6912 ^ x405 ;
  assign n6908 = n6907 ^ n6906 ;
  assign n6909 = n6908 ^ n6901 ;
  assign n6914 = n6913 ^ n6909 ;
  assign n6915 = ~n3493 & n6914 ;
  assign n6918 = n6915 ^ n6909 ;
  assign n6919 = n6918 ^ x373 ;
  assign n6920 = ~n3537 & n6919 ;
  assign n6921 = n6920 ^ x373 ;
  assign n6916 = n6915 ^ n6914 ;
  assign n6917 = n6916 ^ n6909 ;
  assign n6922 = n6921 ^ n6917 ;
  assign n6923 = n3577 & n6922 ;
  assign n6926 = n6923 ^ n6917 ;
  assign n6927 = n6926 ^ x341 ;
  assign n6928 = ~n3620 & n6927 ;
  assign n6929 = n6928 ^ x341 ;
  assign n6924 = n6923 ^ n6922 ;
  assign n6925 = n6924 ^ n6917 ;
  assign n6930 = n6929 ^ n6925 ;
  assign n6931 = n3656 & n6930 ;
  assign n6934 = n6931 ^ n6925 ;
  assign n6935 = n6934 ^ x309 ;
  assign n6936 = ~n3700 & n6935 ;
  assign n6937 = n6936 ^ x309 ;
  assign n6932 = n6931 ^ n6930 ;
  assign n6933 = n6932 ^ n6925 ;
  assign n6938 = n6937 ^ n6933 ;
  assign n6939 = n3739 & n6938 ;
  assign n6942 = n6939 ^ n6933 ;
  assign n6943 = n6942 ^ x277 ;
  assign n6944 = ~n3783 & n6943 ;
  assign n6945 = n6944 ^ x277 ;
  assign n6940 = n6939 ^ n6938 ;
  assign n6941 = n6940 ^ n6933 ;
  assign n6946 = n6945 ^ n6941 ;
  assign n6947 = ~n3818 & n6946 ;
  assign n6950 = n6947 ^ n6941 ;
  assign n6951 = n6950 ^ x245 ;
  assign n6952 = ~n3861 & n6951 ;
  assign n6953 = n6952 ^ x245 ;
  assign n6948 = n6947 ^ n6946 ;
  assign n6949 = n6948 ^ n6941 ;
  assign n6954 = n6953 ^ n6949 ;
  assign n6955 = n3897 & n6954 ;
  assign n6958 = n6955 ^ n6949 ;
  assign n6959 = n6958 ^ x213 ;
  assign n6960 = ~n3941 & n6959 ;
  assign n6961 = n6960 ^ x213 ;
  assign n6956 = n6955 ^ n6954 ;
  assign n6957 = n6956 ^ n6949 ;
  assign n6962 = n6961 ^ n6957 ;
  assign n6963 = n3980 & n6962 ;
  assign n6966 = n6963 ^ n6957 ;
  assign n6967 = n6966 ^ x181 ;
  assign n6968 = ~n4024 & n6967 ;
  assign n6969 = n6968 ^ x181 ;
  assign n6964 = n6963 ^ n6962 ;
  assign n6965 = n6964 ^ n6957 ;
  assign n6970 = n6969 ^ n6965 ;
  assign n6971 = ~n4059 & n6970 ;
  assign n6974 = n6971 ^ n6965 ;
  assign n6975 = n6974 ^ x149 ;
  assign n6976 = ~n4102 & n6975 ;
  assign n6977 = n6976 ^ x149 ;
  assign n6972 = n6971 ^ n6970 ;
  assign n6973 = n6972 ^ n6965 ;
  assign n6978 = n6977 ^ n6973 ;
  assign n6979 = n4138 & n6978 ;
  assign n6982 = n6979 ^ n6973 ;
  assign n6983 = n6982 ^ x117 ;
  assign n6984 = ~n4182 & n6983 ;
  assign n6985 = n6984 ^ x117 ;
  assign n6980 = n6979 ^ n6978 ;
  assign n6981 = n6980 ^ n6973 ;
  assign n6986 = n6985 ^ n6981 ;
  assign n6987 = n4221 & n6986 ;
  assign n6990 = n6987 ^ n6981 ;
  assign n6991 = n6990 ^ x85 ;
  assign n6992 = ~n4265 & n6991 ;
  assign n6993 = n6992 ^ x85 ;
  assign n6988 = n6987 ^ n6986 ;
  assign n6989 = n6988 ^ n6981 ;
  assign n6994 = n6993 ^ n6989 ;
  assign n6995 = ~n4300 & n6994 ;
  assign n6998 = n6995 ^ n6989 ;
  assign n6999 = n6998 ^ x53 ;
  assign n7000 = ~n4343 & n6999 ;
  assign n7001 = n7000 ^ x53 ;
  assign n6996 = n6995 ^ n6994 ;
  assign n6997 = n6996 ^ n6989 ;
  assign n7002 = n7001 ^ n6997 ;
  assign n7003 = n4379 & n7002 ;
  assign n7006 = n7003 ^ n6997 ;
  assign n7007 = n7006 ^ x21 ;
  assign n7008 = ~n4425 & n7007 ;
  assign n7009 = n7008 ^ x21 ;
  assign n7004 = n7003 ^ n7002 ;
  assign n7005 = n7004 ^ n6997 ;
  assign n7010 = n7009 ^ n7005 ;
  assign n7011 = ~n4461 & n7010 ;
  assign n7012 = n7011 ^ n7010 ;
  assign n7013 = n7012 ^ n7005 ;
  assign n7014 = x502 ^ x470 ;
  assign n7015 = ~n3330 & n7014 ;
  assign n7018 = n7015 ^ x470 ;
  assign n7019 = n7018 ^ x438 ;
  assign n7020 = ~n3377 & n7019 ;
  assign n7021 = n7020 ^ x438 ;
  assign n7016 = n7015 ^ n7014 ;
  assign n7017 = n7016 ^ x470 ;
  assign n7022 = n7021 ^ n7017 ;
  assign n7023 = ~n3413 & n7022 ;
  assign n7026 = n7023 ^ n7017 ;
  assign n7027 = n7026 ^ x406 ;
  assign n7028 = ~n3457 & n7027 ;
  assign n7029 = n7028 ^ x406 ;
  assign n7024 = n7023 ^ n7022 ;
  assign n7025 = n7024 ^ n7017 ;
  assign n7030 = n7029 ^ n7025 ;
  assign n7031 = ~n3493 & n7030 ;
  assign n7034 = n7031 ^ n7025 ;
  assign n7035 = n7034 ^ x374 ;
  assign n7036 = ~n3537 & n7035 ;
  assign n7037 = n7036 ^ x374 ;
  assign n7032 = n7031 ^ n7030 ;
  assign n7033 = n7032 ^ n7025 ;
  assign n7038 = n7037 ^ n7033 ;
  assign n7039 = n3577 & n7038 ;
  assign n7042 = n7039 ^ n7033 ;
  assign n7043 = n7042 ^ x342 ;
  assign n7044 = ~n3620 & n7043 ;
  assign n7045 = n7044 ^ x342 ;
  assign n7040 = n7039 ^ n7038 ;
  assign n7041 = n7040 ^ n7033 ;
  assign n7046 = n7045 ^ n7041 ;
  assign n7047 = n3656 & n7046 ;
  assign n7050 = n7047 ^ n7041 ;
  assign n7051 = n7050 ^ x310 ;
  assign n7052 = ~n3700 & n7051 ;
  assign n7053 = n7052 ^ x310 ;
  assign n7048 = n7047 ^ n7046 ;
  assign n7049 = n7048 ^ n7041 ;
  assign n7054 = n7053 ^ n7049 ;
  assign n7055 = n3739 & n7054 ;
  assign n7058 = n7055 ^ n7049 ;
  assign n7059 = n7058 ^ x278 ;
  assign n7060 = ~n3783 & n7059 ;
  assign n7061 = n7060 ^ x278 ;
  assign n7056 = n7055 ^ n7054 ;
  assign n7057 = n7056 ^ n7049 ;
  assign n7062 = n7061 ^ n7057 ;
  assign n7063 = ~n3818 & n7062 ;
  assign n7066 = n7063 ^ n7057 ;
  assign n7067 = n7066 ^ x246 ;
  assign n7068 = ~n3861 & n7067 ;
  assign n7069 = n7068 ^ x246 ;
  assign n7064 = n7063 ^ n7062 ;
  assign n7065 = n7064 ^ n7057 ;
  assign n7070 = n7069 ^ n7065 ;
  assign n7071 = n3897 & n7070 ;
  assign n7074 = n7071 ^ n7065 ;
  assign n7075 = n7074 ^ x214 ;
  assign n7076 = ~n3941 & n7075 ;
  assign n7077 = n7076 ^ x214 ;
  assign n7072 = n7071 ^ n7070 ;
  assign n7073 = n7072 ^ n7065 ;
  assign n7078 = n7077 ^ n7073 ;
  assign n7079 = n3980 & n7078 ;
  assign n7082 = n7079 ^ n7073 ;
  assign n7083 = n7082 ^ x182 ;
  assign n7084 = ~n4024 & n7083 ;
  assign n7085 = n7084 ^ x182 ;
  assign n7080 = n7079 ^ n7078 ;
  assign n7081 = n7080 ^ n7073 ;
  assign n7086 = n7085 ^ n7081 ;
  assign n7087 = ~n4059 & n7086 ;
  assign n7090 = n7087 ^ n7081 ;
  assign n7091 = n7090 ^ x150 ;
  assign n7092 = ~n4102 & n7091 ;
  assign n7093 = n7092 ^ x150 ;
  assign n7088 = n7087 ^ n7086 ;
  assign n7089 = n7088 ^ n7081 ;
  assign n7094 = n7093 ^ n7089 ;
  assign n7095 = n4138 & n7094 ;
  assign n7098 = n7095 ^ n7089 ;
  assign n7099 = n7098 ^ x118 ;
  assign n7100 = ~n4182 & n7099 ;
  assign n7101 = n7100 ^ x118 ;
  assign n7096 = n7095 ^ n7094 ;
  assign n7097 = n7096 ^ n7089 ;
  assign n7102 = n7101 ^ n7097 ;
  assign n7103 = n4221 & n7102 ;
  assign n7106 = n7103 ^ n7097 ;
  assign n7107 = n7106 ^ x86 ;
  assign n7108 = ~n4265 & n7107 ;
  assign n7109 = n7108 ^ x86 ;
  assign n7104 = n7103 ^ n7102 ;
  assign n7105 = n7104 ^ n7097 ;
  assign n7110 = n7109 ^ n7105 ;
  assign n7111 = ~n4300 & n7110 ;
  assign n7114 = n7111 ^ n7105 ;
  assign n7115 = n7114 ^ x54 ;
  assign n7116 = ~n4343 & n7115 ;
  assign n7117 = n7116 ^ x54 ;
  assign n7112 = n7111 ^ n7110 ;
  assign n7113 = n7112 ^ n7105 ;
  assign n7118 = n7117 ^ n7113 ;
  assign n7119 = n4379 & n7118 ;
  assign n7122 = n7119 ^ n7113 ;
  assign n7123 = n7122 ^ x22 ;
  assign n7124 = ~n4425 & n7123 ;
  assign n7125 = n7124 ^ x22 ;
  assign n7120 = n7119 ^ n7118 ;
  assign n7121 = n7120 ^ n7113 ;
  assign n7126 = n7125 ^ n7121 ;
  assign n7127 = ~n4461 & n7126 ;
  assign n7128 = n7127 ^ n7126 ;
  assign n7129 = n7128 ^ n7121 ;
  assign n7130 = x503 ^ x471 ;
  assign n7131 = ~n3330 & n7130 ;
  assign n7134 = n7131 ^ x471 ;
  assign n7135 = n7134 ^ x439 ;
  assign n7136 = ~n3377 & n7135 ;
  assign n7137 = n7136 ^ x439 ;
  assign n7132 = n7131 ^ n7130 ;
  assign n7133 = n7132 ^ x471 ;
  assign n7138 = n7137 ^ n7133 ;
  assign n7139 = ~n3413 & n7138 ;
  assign n7142 = n7139 ^ n7133 ;
  assign n7143 = n7142 ^ x407 ;
  assign n7144 = ~n3457 & n7143 ;
  assign n7145 = n7144 ^ x407 ;
  assign n7140 = n7139 ^ n7138 ;
  assign n7141 = n7140 ^ n7133 ;
  assign n7146 = n7145 ^ n7141 ;
  assign n7147 = ~n3493 & n7146 ;
  assign n7150 = n7147 ^ n7141 ;
  assign n7151 = n7150 ^ x375 ;
  assign n7152 = ~n3537 & n7151 ;
  assign n7153 = n7152 ^ x375 ;
  assign n7148 = n7147 ^ n7146 ;
  assign n7149 = n7148 ^ n7141 ;
  assign n7154 = n7153 ^ n7149 ;
  assign n7155 = n3577 & n7154 ;
  assign n7158 = n7155 ^ n7149 ;
  assign n7159 = n7158 ^ x343 ;
  assign n7160 = ~n3620 & n7159 ;
  assign n7161 = n7160 ^ x343 ;
  assign n7156 = n7155 ^ n7154 ;
  assign n7157 = n7156 ^ n7149 ;
  assign n7162 = n7161 ^ n7157 ;
  assign n7163 = n3656 & n7162 ;
  assign n7166 = n7163 ^ n7157 ;
  assign n7167 = n7166 ^ x311 ;
  assign n7168 = ~n3700 & n7167 ;
  assign n7169 = n7168 ^ x311 ;
  assign n7164 = n7163 ^ n7162 ;
  assign n7165 = n7164 ^ n7157 ;
  assign n7170 = n7169 ^ n7165 ;
  assign n7171 = n3739 & n7170 ;
  assign n7174 = n7171 ^ n7165 ;
  assign n7175 = n7174 ^ x279 ;
  assign n7176 = ~n3783 & n7175 ;
  assign n7177 = n7176 ^ x279 ;
  assign n7172 = n7171 ^ n7170 ;
  assign n7173 = n7172 ^ n7165 ;
  assign n7178 = n7177 ^ n7173 ;
  assign n7179 = ~n3818 & n7178 ;
  assign n7182 = n7179 ^ n7173 ;
  assign n7183 = n7182 ^ x247 ;
  assign n7184 = ~n3861 & n7183 ;
  assign n7185 = n7184 ^ x247 ;
  assign n7180 = n7179 ^ n7178 ;
  assign n7181 = n7180 ^ n7173 ;
  assign n7186 = n7185 ^ n7181 ;
  assign n7187 = n3897 & n7186 ;
  assign n7190 = n7187 ^ n7181 ;
  assign n7191 = n7190 ^ x215 ;
  assign n7192 = ~n3941 & n7191 ;
  assign n7193 = n7192 ^ x215 ;
  assign n7188 = n7187 ^ n7186 ;
  assign n7189 = n7188 ^ n7181 ;
  assign n7194 = n7193 ^ n7189 ;
  assign n7195 = n3980 & n7194 ;
  assign n7198 = n7195 ^ n7189 ;
  assign n7199 = n7198 ^ x183 ;
  assign n7200 = ~n4024 & n7199 ;
  assign n7201 = n7200 ^ x183 ;
  assign n7196 = n7195 ^ n7194 ;
  assign n7197 = n7196 ^ n7189 ;
  assign n7202 = n7201 ^ n7197 ;
  assign n7203 = ~n4059 & n7202 ;
  assign n7206 = n7203 ^ n7197 ;
  assign n7207 = n7206 ^ x151 ;
  assign n7208 = ~n4102 & n7207 ;
  assign n7209 = n7208 ^ x151 ;
  assign n7204 = n7203 ^ n7202 ;
  assign n7205 = n7204 ^ n7197 ;
  assign n7210 = n7209 ^ n7205 ;
  assign n7211 = n4138 & n7210 ;
  assign n7214 = n7211 ^ n7205 ;
  assign n7215 = n7214 ^ x119 ;
  assign n7216 = ~n4182 & n7215 ;
  assign n7217 = n7216 ^ x119 ;
  assign n7212 = n7211 ^ n7210 ;
  assign n7213 = n7212 ^ n7205 ;
  assign n7218 = n7217 ^ n7213 ;
  assign n7219 = n4221 & n7218 ;
  assign n7222 = n7219 ^ n7213 ;
  assign n7223 = n7222 ^ x87 ;
  assign n7224 = ~n4265 & n7223 ;
  assign n7225 = n7224 ^ x87 ;
  assign n7220 = n7219 ^ n7218 ;
  assign n7221 = n7220 ^ n7213 ;
  assign n7226 = n7225 ^ n7221 ;
  assign n7227 = ~n4300 & n7226 ;
  assign n7230 = n7227 ^ n7221 ;
  assign n7231 = n7230 ^ x55 ;
  assign n7232 = ~n4343 & n7231 ;
  assign n7233 = n7232 ^ x55 ;
  assign n7228 = n7227 ^ n7226 ;
  assign n7229 = n7228 ^ n7221 ;
  assign n7234 = n7233 ^ n7229 ;
  assign n7235 = n4379 & n7234 ;
  assign n7238 = n7235 ^ n7229 ;
  assign n7239 = n7238 ^ x23 ;
  assign n7240 = ~n4425 & n7239 ;
  assign n7241 = n7240 ^ x23 ;
  assign n7236 = n7235 ^ n7234 ;
  assign n7237 = n7236 ^ n7229 ;
  assign n7242 = n7241 ^ n7237 ;
  assign n7243 = ~n4461 & n7242 ;
  assign n7244 = n7243 ^ n7242 ;
  assign n7245 = n7244 ^ n7237 ;
  assign n7246 = x504 ^ x472 ;
  assign n7247 = ~n3330 & n7246 ;
  assign n7250 = n7247 ^ x472 ;
  assign n7251 = n7250 ^ x440 ;
  assign n7252 = ~n3377 & n7251 ;
  assign n7253 = n7252 ^ x440 ;
  assign n7248 = n7247 ^ n7246 ;
  assign n7249 = n7248 ^ x472 ;
  assign n7254 = n7253 ^ n7249 ;
  assign n7255 = ~n3413 & n7254 ;
  assign n7258 = n7255 ^ n7249 ;
  assign n7259 = n7258 ^ x408 ;
  assign n7260 = ~n3457 & n7259 ;
  assign n7261 = n7260 ^ x408 ;
  assign n7256 = n7255 ^ n7254 ;
  assign n7257 = n7256 ^ n7249 ;
  assign n7262 = n7261 ^ n7257 ;
  assign n7263 = ~n3493 & n7262 ;
  assign n7266 = n7263 ^ n7257 ;
  assign n7267 = n7266 ^ x376 ;
  assign n7268 = ~n3537 & n7267 ;
  assign n7269 = n7268 ^ x376 ;
  assign n7264 = n7263 ^ n7262 ;
  assign n7265 = n7264 ^ n7257 ;
  assign n7270 = n7269 ^ n7265 ;
  assign n7271 = n3577 & n7270 ;
  assign n7274 = n7271 ^ n7265 ;
  assign n7275 = n7274 ^ x344 ;
  assign n7276 = ~n3620 & n7275 ;
  assign n7277 = n7276 ^ x344 ;
  assign n7272 = n7271 ^ n7270 ;
  assign n7273 = n7272 ^ n7265 ;
  assign n7278 = n7277 ^ n7273 ;
  assign n7279 = n3656 & n7278 ;
  assign n7282 = n7279 ^ n7273 ;
  assign n7283 = n7282 ^ x312 ;
  assign n7284 = ~n3700 & n7283 ;
  assign n7285 = n7284 ^ x312 ;
  assign n7280 = n7279 ^ n7278 ;
  assign n7281 = n7280 ^ n7273 ;
  assign n7286 = n7285 ^ n7281 ;
  assign n7287 = n3739 & n7286 ;
  assign n7290 = n7287 ^ n7281 ;
  assign n7291 = n7290 ^ x280 ;
  assign n7292 = ~n3783 & n7291 ;
  assign n7293 = n7292 ^ x280 ;
  assign n7288 = n7287 ^ n7286 ;
  assign n7289 = n7288 ^ n7281 ;
  assign n7294 = n7293 ^ n7289 ;
  assign n7295 = ~n3818 & n7294 ;
  assign n7298 = n7295 ^ n7289 ;
  assign n7299 = n7298 ^ x248 ;
  assign n7300 = ~n3861 & n7299 ;
  assign n7301 = n7300 ^ x248 ;
  assign n7296 = n7295 ^ n7294 ;
  assign n7297 = n7296 ^ n7289 ;
  assign n7302 = n7301 ^ n7297 ;
  assign n7303 = n3897 & n7302 ;
  assign n7306 = n7303 ^ n7297 ;
  assign n7307 = n7306 ^ x216 ;
  assign n7308 = ~n3941 & n7307 ;
  assign n7309 = n7308 ^ x216 ;
  assign n7304 = n7303 ^ n7302 ;
  assign n7305 = n7304 ^ n7297 ;
  assign n7310 = n7309 ^ n7305 ;
  assign n7311 = n3980 & n7310 ;
  assign n7314 = n7311 ^ n7305 ;
  assign n7315 = n7314 ^ x184 ;
  assign n7316 = ~n4024 & n7315 ;
  assign n7317 = n7316 ^ x184 ;
  assign n7312 = n7311 ^ n7310 ;
  assign n7313 = n7312 ^ n7305 ;
  assign n7318 = n7317 ^ n7313 ;
  assign n7319 = ~n4059 & n7318 ;
  assign n7322 = n7319 ^ n7313 ;
  assign n7323 = n7322 ^ x152 ;
  assign n7324 = ~n4102 & n7323 ;
  assign n7325 = n7324 ^ x152 ;
  assign n7320 = n7319 ^ n7318 ;
  assign n7321 = n7320 ^ n7313 ;
  assign n7326 = n7325 ^ n7321 ;
  assign n7327 = n4138 & n7326 ;
  assign n7330 = n7327 ^ n7321 ;
  assign n7331 = n7330 ^ x120 ;
  assign n7332 = ~n4182 & n7331 ;
  assign n7333 = n7332 ^ x120 ;
  assign n7328 = n7327 ^ n7326 ;
  assign n7329 = n7328 ^ n7321 ;
  assign n7334 = n7333 ^ n7329 ;
  assign n7335 = n4221 & n7334 ;
  assign n7338 = n7335 ^ n7329 ;
  assign n7339 = n7338 ^ x88 ;
  assign n7340 = ~n4265 & n7339 ;
  assign n7341 = n7340 ^ x88 ;
  assign n7336 = n7335 ^ n7334 ;
  assign n7337 = n7336 ^ n7329 ;
  assign n7342 = n7341 ^ n7337 ;
  assign n7343 = ~n4300 & n7342 ;
  assign n7346 = n7343 ^ n7337 ;
  assign n7347 = n7346 ^ x56 ;
  assign n7348 = ~n4343 & n7347 ;
  assign n7349 = n7348 ^ x56 ;
  assign n7344 = n7343 ^ n7342 ;
  assign n7345 = n7344 ^ n7337 ;
  assign n7350 = n7349 ^ n7345 ;
  assign n7351 = n4379 & n7350 ;
  assign n7354 = n7351 ^ n7345 ;
  assign n7355 = n7354 ^ x24 ;
  assign n7356 = ~n4425 & n7355 ;
  assign n7357 = n7356 ^ x24 ;
  assign n7352 = n7351 ^ n7350 ;
  assign n7353 = n7352 ^ n7345 ;
  assign n7358 = n7357 ^ n7353 ;
  assign n7359 = ~n4461 & n7358 ;
  assign n7360 = n7359 ^ n7358 ;
  assign n7361 = n7360 ^ n7353 ;
  assign n7362 = x505 ^ x473 ;
  assign n7363 = ~n3330 & n7362 ;
  assign n7366 = n7363 ^ x473 ;
  assign n7367 = n7366 ^ x441 ;
  assign n7368 = ~n3377 & n7367 ;
  assign n7369 = n7368 ^ x441 ;
  assign n7364 = n7363 ^ n7362 ;
  assign n7365 = n7364 ^ x473 ;
  assign n7370 = n7369 ^ n7365 ;
  assign n7371 = ~n3413 & n7370 ;
  assign n7374 = n7371 ^ n7365 ;
  assign n7375 = n7374 ^ x409 ;
  assign n7376 = ~n3457 & n7375 ;
  assign n7377 = n7376 ^ x409 ;
  assign n7372 = n7371 ^ n7370 ;
  assign n7373 = n7372 ^ n7365 ;
  assign n7378 = n7377 ^ n7373 ;
  assign n7379 = ~n3493 & n7378 ;
  assign n7382 = n7379 ^ n7373 ;
  assign n7383 = n7382 ^ x377 ;
  assign n7384 = ~n3537 & n7383 ;
  assign n7385 = n7384 ^ x377 ;
  assign n7380 = n7379 ^ n7378 ;
  assign n7381 = n7380 ^ n7373 ;
  assign n7386 = n7385 ^ n7381 ;
  assign n7387 = n3577 & n7386 ;
  assign n7390 = n7387 ^ n7381 ;
  assign n7391 = n7390 ^ x345 ;
  assign n7392 = ~n3620 & n7391 ;
  assign n7393 = n7392 ^ x345 ;
  assign n7388 = n7387 ^ n7386 ;
  assign n7389 = n7388 ^ n7381 ;
  assign n7394 = n7393 ^ n7389 ;
  assign n7395 = n3656 & n7394 ;
  assign n7398 = n7395 ^ n7389 ;
  assign n7399 = n7398 ^ x313 ;
  assign n7400 = ~n3700 & n7399 ;
  assign n7401 = n7400 ^ x313 ;
  assign n7396 = n7395 ^ n7394 ;
  assign n7397 = n7396 ^ n7389 ;
  assign n7402 = n7401 ^ n7397 ;
  assign n7403 = n3739 & n7402 ;
  assign n7406 = n7403 ^ n7397 ;
  assign n7407 = n7406 ^ x281 ;
  assign n7408 = ~n3783 & n7407 ;
  assign n7409 = n7408 ^ x281 ;
  assign n7404 = n7403 ^ n7402 ;
  assign n7405 = n7404 ^ n7397 ;
  assign n7410 = n7409 ^ n7405 ;
  assign n7411 = ~n3818 & n7410 ;
  assign n7414 = n7411 ^ n7405 ;
  assign n7415 = n7414 ^ x249 ;
  assign n7416 = ~n3861 & n7415 ;
  assign n7417 = n7416 ^ x249 ;
  assign n7412 = n7411 ^ n7410 ;
  assign n7413 = n7412 ^ n7405 ;
  assign n7418 = n7417 ^ n7413 ;
  assign n7419 = n3897 & n7418 ;
  assign n7422 = n7419 ^ n7413 ;
  assign n7423 = n7422 ^ x217 ;
  assign n7424 = ~n3941 & n7423 ;
  assign n7425 = n7424 ^ x217 ;
  assign n7420 = n7419 ^ n7418 ;
  assign n7421 = n7420 ^ n7413 ;
  assign n7426 = n7425 ^ n7421 ;
  assign n7427 = n3980 & n7426 ;
  assign n7430 = n7427 ^ n7421 ;
  assign n7431 = n7430 ^ x185 ;
  assign n7432 = ~n4024 & n7431 ;
  assign n7433 = n7432 ^ x185 ;
  assign n7428 = n7427 ^ n7426 ;
  assign n7429 = n7428 ^ n7421 ;
  assign n7434 = n7433 ^ n7429 ;
  assign n7435 = ~n4059 & n7434 ;
  assign n7438 = n7435 ^ n7429 ;
  assign n7439 = n7438 ^ x153 ;
  assign n7440 = ~n4102 & n7439 ;
  assign n7441 = n7440 ^ x153 ;
  assign n7436 = n7435 ^ n7434 ;
  assign n7437 = n7436 ^ n7429 ;
  assign n7442 = n7441 ^ n7437 ;
  assign n7443 = n4138 & n7442 ;
  assign n7446 = n7443 ^ n7437 ;
  assign n7447 = n7446 ^ x121 ;
  assign n7448 = ~n4182 & n7447 ;
  assign n7449 = n7448 ^ x121 ;
  assign n7444 = n7443 ^ n7442 ;
  assign n7445 = n7444 ^ n7437 ;
  assign n7450 = n7449 ^ n7445 ;
  assign n7451 = n4221 & n7450 ;
  assign n7454 = n7451 ^ n7445 ;
  assign n7455 = n7454 ^ x89 ;
  assign n7456 = ~n4265 & n7455 ;
  assign n7457 = n7456 ^ x89 ;
  assign n7452 = n7451 ^ n7450 ;
  assign n7453 = n7452 ^ n7445 ;
  assign n7458 = n7457 ^ n7453 ;
  assign n7459 = ~n4300 & n7458 ;
  assign n7462 = n7459 ^ n7453 ;
  assign n7463 = n7462 ^ x57 ;
  assign n7464 = ~n4343 & n7463 ;
  assign n7465 = n7464 ^ x57 ;
  assign n7460 = n7459 ^ n7458 ;
  assign n7461 = n7460 ^ n7453 ;
  assign n7466 = n7465 ^ n7461 ;
  assign n7467 = n4379 & n7466 ;
  assign n7470 = n7467 ^ n7461 ;
  assign n7471 = n7470 ^ x25 ;
  assign n7472 = ~n4425 & n7471 ;
  assign n7473 = n7472 ^ x25 ;
  assign n7468 = n7467 ^ n7466 ;
  assign n7469 = n7468 ^ n7461 ;
  assign n7474 = n7473 ^ n7469 ;
  assign n7475 = ~n4461 & n7474 ;
  assign n7476 = n7475 ^ n7474 ;
  assign n7477 = n7476 ^ n7469 ;
  assign n7478 = x506 ^ x474 ;
  assign n7479 = ~n3330 & n7478 ;
  assign n7482 = n7479 ^ x474 ;
  assign n7483 = n7482 ^ x442 ;
  assign n7484 = ~n3377 & n7483 ;
  assign n7485 = n7484 ^ x442 ;
  assign n7480 = n7479 ^ n7478 ;
  assign n7481 = n7480 ^ x474 ;
  assign n7486 = n7485 ^ n7481 ;
  assign n7487 = ~n3413 & n7486 ;
  assign n7490 = n7487 ^ n7481 ;
  assign n7491 = n7490 ^ x410 ;
  assign n7492 = ~n3457 & n7491 ;
  assign n7493 = n7492 ^ x410 ;
  assign n7488 = n7487 ^ n7486 ;
  assign n7489 = n7488 ^ n7481 ;
  assign n7494 = n7493 ^ n7489 ;
  assign n7495 = ~n3493 & n7494 ;
  assign n7498 = n7495 ^ n7489 ;
  assign n7499 = n7498 ^ x378 ;
  assign n7500 = ~n3537 & n7499 ;
  assign n7501 = n7500 ^ x378 ;
  assign n7496 = n7495 ^ n7494 ;
  assign n7497 = n7496 ^ n7489 ;
  assign n7502 = n7501 ^ n7497 ;
  assign n7503 = n3577 & n7502 ;
  assign n7506 = n7503 ^ n7497 ;
  assign n7507 = n7506 ^ x346 ;
  assign n7508 = ~n3620 & n7507 ;
  assign n7509 = n7508 ^ x346 ;
  assign n7504 = n7503 ^ n7502 ;
  assign n7505 = n7504 ^ n7497 ;
  assign n7510 = n7509 ^ n7505 ;
  assign n7511 = n3656 & n7510 ;
  assign n7514 = n7511 ^ n7505 ;
  assign n7515 = n7514 ^ x314 ;
  assign n7516 = ~n3700 & n7515 ;
  assign n7517 = n7516 ^ x314 ;
  assign n7512 = n7511 ^ n7510 ;
  assign n7513 = n7512 ^ n7505 ;
  assign n7518 = n7517 ^ n7513 ;
  assign n7519 = n3739 & n7518 ;
  assign n7522 = n7519 ^ n7513 ;
  assign n7523 = n7522 ^ x282 ;
  assign n7524 = ~n3783 & n7523 ;
  assign n7525 = n7524 ^ x282 ;
  assign n7520 = n7519 ^ n7518 ;
  assign n7521 = n7520 ^ n7513 ;
  assign n7526 = n7525 ^ n7521 ;
  assign n7527 = ~n3818 & n7526 ;
  assign n7530 = n7527 ^ n7521 ;
  assign n7531 = n7530 ^ x250 ;
  assign n7532 = ~n3861 & n7531 ;
  assign n7533 = n7532 ^ x250 ;
  assign n7528 = n7527 ^ n7526 ;
  assign n7529 = n7528 ^ n7521 ;
  assign n7534 = n7533 ^ n7529 ;
  assign n7535 = n3897 & n7534 ;
  assign n7538 = n7535 ^ n7529 ;
  assign n7539 = n7538 ^ x218 ;
  assign n7540 = ~n3941 & n7539 ;
  assign n7541 = n7540 ^ x218 ;
  assign n7536 = n7535 ^ n7534 ;
  assign n7537 = n7536 ^ n7529 ;
  assign n7542 = n7541 ^ n7537 ;
  assign n7543 = n3980 & n7542 ;
  assign n7546 = n7543 ^ n7537 ;
  assign n7547 = n7546 ^ x186 ;
  assign n7548 = ~n4024 & n7547 ;
  assign n7549 = n7548 ^ x186 ;
  assign n7544 = n7543 ^ n7542 ;
  assign n7545 = n7544 ^ n7537 ;
  assign n7550 = n7549 ^ n7545 ;
  assign n7551 = ~n4059 & n7550 ;
  assign n7554 = n7551 ^ n7545 ;
  assign n7555 = n7554 ^ x154 ;
  assign n7556 = ~n4102 & n7555 ;
  assign n7557 = n7556 ^ x154 ;
  assign n7552 = n7551 ^ n7550 ;
  assign n7553 = n7552 ^ n7545 ;
  assign n7558 = n7557 ^ n7553 ;
  assign n7559 = n4138 & n7558 ;
  assign n7562 = n7559 ^ n7553 ;
  assign n7563 = n7562 ^ x122 ;
  assign n7564 = ~n4182 & n7563 ;
  assign n7565 = n7564 ^ x122 ;
  assign n7560 = n7559 ^ n7558 ;
  assign n7561 = n7560 ^ n7553 ;
  assign n7566 = n7565 ^ n7561 ;
  assign n7567 = n4221 & n7566 ;
  assign n7570 = n7567 ^ n7561 ;
  assign n7571 = n7570 ^ x90 ;
  assign n7572 = ~n4265 & n7571 ;
  assign n7573 = n7572 ^ x90 ;
  assign n7568 = n7567 ^ n7566 ;
  assign n7569 = n7568 ^ n7561 ;
  assign n7574 = n7573 ^ n7569 ;
  assign n7575 = ~n4300 & n7574 ;
  assign n7578 = n7575 ^ n7569 ;
  assign n7579 = n7578 ^ x58 ;
  assign n7580 = ~n4343 & n7579 ;
  assign n7581 = n7580 ^ x58 ;
  assign n7576 = n7575 ^ n7574 ;
  assign n7577 = n7576 ^ n7569 ;
  assign n7582 = n7581 ^ n7577 ;
  assign n7583 = n4379 & n7582 ;
  assign n7586 = n7583 ^ n7577 ;
  assign n7587 = n7586 ^ x26 ;
  assign n7588 = ~n4425 & n7587 ;
  assign n7589 = n7588 ^ x26 ;
  assign n7584 = n7583 ^ n7582 ;
  assign n7585 = n7584 ^ n7577 ;
  assign n7590 = n7589 ^ n7585 ;
  assign n7591 = ~n4461 & n7590 ;
  assign n7592 = n7591 ^ n7590 ;
  assign n7593 = n7592 ^ n7585 ;
  assign n7594 = x507 ^ x475 ;
  assign n7595 = ~n3330 & n7594 ;
  assign n7598 = n7595 ^ x475 ;
  assign n7599 = n7598 ^ x443 ;
  assign n7600 = ~n3377 & n7599 ;
  assign n7601 = n7600 ^ x443 ;
  assign n7596 = n7595 ^ n7594 ;
  assign n7597 = n7596 ^ x475 ;
  assign n7602 = n7601 ^ n7597 ;
  assign n7603 = ~n3413 & n7602 ;
  assign n7606 = n7603 ^ n7597 ;
  assign n7607 = n7606 ^ x411 ;
  assign n7608 = ~n3457 & n7607 ;
  assign n7609 = n7608 ^ x411 ;
  assign n7604 = n7603 ^ n7602 ;
  assign n7605 = n7604 ^ n7597 ;
  assign n7610 = n7609 ^ n7605 ;
  assign n7611 = ~n3493 & n7610 ;
  assign n7614 = n7611 ^ n7605 ;
  assign n7615 = n7614 ^ x379 ;
  assign n7616 = ~n3537 & n7615 ;
  assign n7617 = n7616 ^ x379 ;
  assign n7612 = n7611 ^ n7610 ;
  assign n7613 = n7612 ^ n7605 ;
  assign n7618 = n7617 ^ n7613 ;
  assign n7619 = n3577 & n7618 ;
  assign n7622 = n7619 ^ n7613 ;
  assign n7623 = n7622 ^ x347 ;
  assign n7624 = ~n3620 & n7623 ;
  assign n7625 = n7624 ^ x347 ;
  assign n7620 = n7619 ^ n7618 ;
  assign n7621 = n7620 ^ n7613 ;
  assign n7626 = n7625 ^ n7621 ;
  assign n7627 = n3656 & n7626 ;
  assign n7630 = n7627 ^ n7621 ;
  assign n7631 = n7630 ^ x315 ;
  assign n7632 = ~n3700 & n7631 ;
  assign n7633 = n7632 ^ x315 ;
  assign n7628 = n7627 ^ n7626 ;
  assign n7629 = n7628 ^ n7621 ;
  assign n7634 = n7633 ^ n7629 ;
  assign n7635 = n3739 & n7634 ;
  assign n7638 = n7635 ^ n7629 ;
  assign n7639 = n7638 ^ x283 ;
  assign n7640 = ~n3783 & n7639 ;
  assign n7641 = n7640 ^ x283 ;
  assign n7636 = n7635 ^ n7634 ;
  assign n7637 = n7636 ^ n7629 ;
  assign n7642 = n7641 ^ n7637 ;
  assign n7643 = ~n3818 & n7642 ;
  assign n7646 = n7643 ^ n7637 ;
  assign n7647 = n7646 ^ x251 ;
  assign n7648 = ~n3861 & n7647 ;
  assign n7649 = n7648 ^ x251 ;
  assign n7644 = n7643 ^ n7642 ;
  assign n7645 = n7644 ^ n7637 ;
  assign n7650 = n7649 ^ n7645 ;
  assign n7651 = n3897 & n7650 ;
  assign n7654 = n7651 ^ n7645 ;
  assign n7655 = n7654 ^ x219 ;
  assign n7656 = ~n3941 & n7655 ;
  assign n7657 = n7656 ^ x219 ;
  assign n7652 = n7651 ^ n7650 ;
  assign n7653 = n7652 ^ n7645 ;
  assign n7658 = n7657 ^ n7653 ;
  assign n7659 = n3980 & n7658 ;
  assign n7662 = n7659 ^ n7653 ;
  assign n7663 = n7662 ^ x187 ;
  assign n7664 = ~n4024 & n7663 ;
  assign n7665 = n7664 ^ x187 ;
  assign n7660 = n7659 ^ n7658 ;
  assign n7661 = n7660 ^ n7653 ;
  assign n7666 = n7665 ^ n7661 ;
  assign n7667 = ~n4059 & n7666 ;
  assign n7670 = n7667 ^ n7661 ;
  assign n7671 = n7670 ^ x155 ;
  assign n7672 = ~n4102 & n7671 ;
  assign n7673 = n7672 ^ x155 ;
  assign n7668 = n7667 ^ n7666 ;
  assign n7669 = n7668 ^ n7661 ;
  assign n7674 = n7673 ^ n7669 ;
  assign n7675 = n4138 & n7674 ;
  assign n7678 = n7675 ^ n7669 ;
  assign n7679 = n7678 ^ x123 ;
  assign n7680 = ~n4182 & n7679 ;
  assign n7681 = n7680 ^ x123 ;
  assign n7676 = n7675 ^ n7674 ;
  assign n7677 = n7676 ^ n7669 ;
  assign n7682 = n7681 ^ n7677 ;
  assign n7683 = n4221 & n7682 ;
  assign n7686 = n7683 ^ n7677 ;
  assign n7687 = n7686 ^ x91 ;
  assign n7688 = ~n4265 & n7687 ;
  assign n7689 = n7688 ^ x91 ;
  assign n7684 = n7683 ^ n7682 ;
  assign n7685 = n7684 ^ n7677 ;
  assign n7690 = n7689 ^ n7685 ;
  assign n7691 = ~n4300 & n7690 ;
  assign n7694 = n7691 ^ n7685 ;
  assign n7695 = n7694 ^ x59 ;
  assign n7696 = ~n4343 & n7695 ;
  assign n7697 = n7696 ^ x59 ;
  assign n7692 = n7691 ^ n7690 ;
  assign n7693 = n7692 ^ n7685 ;
  assign n7698 = n7697 ^ n7693 ;
  assign n7699 = n4379 & n7698 ;
  assign n7702 = n7699 ^ n7693 ;
  assign n7703 = n7702 ^ x27 ;
  assign n7704 = ~n4425 & n7703 ;
  assign n7705 = n7704 ^ x27 ;
  assign n7700 = n7699 ^ n7698 ;
  assign n7701 = n7700 ^ n7693 ;
  assign n7706 = n7705 ^ n7701 ;
  assign n7707 = ~n4461 & n7706 ;
  assign n7708 = n7707 ^ n7706 ;
  assign n7709 = n7708 ^ n7701 ;
  assign n7710 = x508 ^ x476 ;
  assign n7711 = ~n3330 & n7710 ;
  assign n7714 = n7711 ^ x476 ;
  assign n7715 = n7714 ^ x444 ;
  assign n7716 = ~n3377 & n7715 ;
  assign n7717 = n7716 ^ x444 ;
  assign n7712 = n7711 ^ n7710 ;
  assign n7713 = n7712 ^ x476 ;
  assign n7718 = n7717 ^ n7713 ;
  assign n7719 = ~n3413 & n7718 ;
  assign n7722 = n7719 ^ n7713 ;
  assign n7723 = n7722 ^ x412 ;
  assign n7724 = ~n3457 & n7723 ;
  assign n7725 = n7724 ^ x412 ;
  assign n7720 = n7719 ^ n7718 ;
  assign n7721 = n7720 ^ n7713 ;
  assign n7726 = n7725 ^ n7721 ;
  assign n7727 = ~n3493 & n7726 ;
  assign n7730 = n7727 ^ n7721 ;
  assign n7731 = n7730 ^ x380 ;
  assign n7732 = ~n3537 & n7731 ;
  assign n7733 = n7732 ^ x380 ;
  assign n7728 = n7727 ^ n7726 ;
  assign n7729 = n7728 ^ n7721 ;
  assign n7734 = n7733 ^ n7729 ;
  assign n7735 = n3577 & n7734 ;
  assign n7738 = n7735 ^ n7729 ;
  assign n7739 = n7738 ^ x348 ;
  assign n7740 = ~n3620 & n7739 ;
  assign n7741 = n7740 ^ x348 ;
  assign n7736 = n7735 ^ n7734 ;
  assign n7737 = n7736 ^ n7729 ;
  assign n7742 = n7741 ^ n7737 ;
  assign n7743 = n3656 & n7742 ;
  assign n7746 = n7743 ^ n7737 ;
  assign n7747 = n7746 ^ x316 ;
  assign n7748 = ~n3700 & n7747 ;
  assign n7749 = n7748 ^ x316 ;
  assign n7744 = n7743 ^ n7742 ;
  assign n7745 = n7744 ^ n7737 ;
  assign n7750 = n7749 ^ n7745 ;
  assign n7751 = n3739 & n7750 ;
  assign n7754 = n7751 ^ n7745 ;
  assign n7755 = n7754 ^ x284 ;
  assign n7756 = ~n3783 & n7755 ;
  assign n7757 = n7756 ^ x284 ;
  assign n7752 = n7751 ^ n7750 ;
  assign n7753 = n7752 ^ n7745 ;
  assign n7758 = n7757 ^ n7753 ;
  assign n7759 = ~n3818 & n7758 ;
  assign n7762 = n7759 ^ n7753 ;
  assign n7763 = n7762 ^ x252 ;
  assign n7764 = ~n3861 & n7763 ;
  assign n7765 = n7764 ^ x252 ;
  assign n7760 = n7759 ^ n7758 ;
  assign n7761 = n7760 ^ n7753 ;
  assign n7766 = n7765 ^ n7761 ;
  assign n7767 = n3897 & n7766 ;
  assign n7770 = n7767 ^ n7761 ;
  assign n7771 = n7770 ^ x220 ;
  assign n7772 = ~n3941 & n7771 ;
  assign n7773 = n7772 ^ x220 ;
  assign n7768 = n7767 ^ n7766 ;
  assign n7769 = n7768 ^ n7761 ;
  assign n7774 = n7773 ^ n7769 ;
  assign n7775 = n3980 & n7774 ;
  assign n7778 = n7775 ^ n7769 ;
  assign n7779 = n7778 ^ x188 ;
  assign n7780 = ~n4024 & n7779 ;
  assign n7781 = n7780 ^ x188 ;
  assign n7776 = n7775 ^ n7774 ;
  assign n7777 = n7776 ^ n7769 ;
  assign n7782 = n7781 ^ n7777 ;
  assign n7783 = ~n4059 & n7782 ;
  assign n7786 = n7783 ^ n7777 ;
  assign n7787 = n7786 ^ x156 ;
  assign n7788 = ~n4102 & n7787 ;
  assign n7789 = n7788 ^ x156 ;
  assign n7784 = n7783 ^ n7782 ;
  assign n7785 = n7784 ^ n7777 ;
  assign n7790 = n7789 ^ n7785 ;
  assign n7791 = n4138 & n7790 ;
  assign n7794 = n7791 ^ n7785 ;
  assign n7795 = n7794 ^ x124 ;
  assign n7796 = ~n4182 & n7795 ;
  assign n7797 = n7796 ^ x124 ;
  assign n7792 = n7791 ^ n7790 ;
  assign n7793 = n7792 ^ n7785 ;
  assign n7798 = n7797 ^ n7793 ;
  assign n7799 = n4221 & n7798 ;
  assign n7802 = n7799 ^ n7793 ;
  assign n7803 = n7802 ^ x92 ;
  assign n7804 = ~n4265 & n7803 ;
  assign n7805 = n7804 ^ x92 ;
  assign n7800 = n7799 ^ n7798 ;
  assign n7801 = n7800 ^ n7793 ;
  assign n7806 = n7805 ^ n7801 ;
  assign n7807 = ~n4300 & n7806 ;
  assign n7810 = n7807 ^ n7801 ;
  assign n7811 = n7810 ^ x60 ;
  assign n7812 = ~n4343 & n7811 ;
  assign n7813 = n7812 ^ x60 ;
  assign n7808 = n7807 ^ n7806 ;
  assign n7809 = n7808 ^ n7801 ;
  assign n7814 = n7813 ^ n7809 ;
  assign n7815 = n4379 & n7814 ;
  assign n7818 = n7815 ^ n7809 ;
  assign n7819 = n7818 ^ x28 ;
  assign n7820 = ~n4425 & n7819 ;
  assign n7821 = n7820 ^ x28 ;
  assign n7816 = n7815 ^ n7814 ;
  assign n7817 = n7816 ^ n7809 ;
  assign n7822 = n7821 ^ n7817 ;
  assign n7823 = ~n4461 & n7822 ;
  assign n7824 = n7823 ^ n7822 ;
  assign n7825 = n7824 ^ n7817 ;
  assign n7826 = x509 ^ x477 ;
  assign n7827 = ~n3330 & n7826 ;
  assign n7830 = n7827 ^ x477 ;
  assign n7831 = n7830 ^ x445 ;
  assign n7832 = ~n3377 & n7831 ;
  assign n7833 = n7832 ^ x445 ;
  assign n7828 = n7827 ^ n7826 ;
  assign n7829 = n7828 ^ x477 ;
  assign n7834 = n7833 ^ n7829 ;
  assign n7835 = ~n3413 & n7834 ;
  assign n7838 = n7835 ^ n7829 ;
  assign n7839 = n7838 ^ x413 ;
  assign n7840 = ~n3457 & n7839 ;
  assign n7841 = n7840 ^ x413 ;
  assign n7836 = n7835 ^ n7834 ;
  assign n7837 = n7836 ^ n7829 ;
  assign n7842 = n7841 ^ n7837 ;
  assign n7843 = ~n3493 & n7842 ;
  assign n7846 = n7843 ^ n7837 ;
  assign n7847 = n7846 ^ x381 ;
  assign n7848 = ~n3537 & n7847 ;
  assign n7849 = n7848 ^ x381 ;
  assign n7844 = n7843 ^ n7842 ;
  assign n7845 = n7844 ^ n7837 ;
  assign n7850 = n7849 ^ n7845 ;
  assign n7851 = n3577 & n7850 ;
  assign n7854 = n7851 ^ n7845 ;
  assign n7855 = n7854 ^ x349 ;
  assign n7856 = ~n3620 & n7855 ;
  assign n7857 = n7856 ^ x349 ;
  assign n7852 = n7851 ^ n7850 ;
  assign n7853 = n7852 ^ n7845 ;
  assign n7858 = n7857 ^ n7853 ;
  assign n7859 = n3656 & n7858 ;
  assign n7862 = n7859 ^ n7853 ;
  assign n7863 = n7862 ^ x317 ;
  assign n7864 = ~n3700 & n7863 ;
  assign n7865 = n7864 ^ x317 ;
  assign n7860 = n7859 ^ n7858 ;
  assign n7861 = n7860 ^ n7853 ;
  assign n7866 = n7865 ^ n7861 ;
  assign n7867 = n3739 & n7866 ;
  assign n7870 = n7867 ^ n7861 ;
  assign n7871 = n7870 ^ x285 ;
  assign n7872 = ~n3783 & n7871 ;
  assign n7873 = n7872 ^ x285 ;
  assign n7868 = n7867 ^ n7866 ;
  assign n7869 = n7868 ^ n7861 ;
  assign n7874 = n7873 ^ n7869 ;
  assign n7875 = ~n3818 & n7874 ;
  assign n7878 = n7875 ^ n7869 ;
  assign n7879 = n7878 ^ x253 ;
  assign n7880 = ~n3861 & n7879 ;
  assign n7881 = n7880 ^ x253 ;
  assign n7876 = n7875 ^ n7874 ;
  assign n7877 = n7876 ^ n7869 ;
  assign n7882 = n7881 ^ n7877 ;
  assign n7883 = n3897 & n7882 ;
  assign n7886 = n7883 ^ n7877 ;
  assign n7887 = n7886 ^ x221 ;
  assign n7888 = ~n3941 & n7887 ;
  assign n7889 = n7888 ^ x221 ;
  assign n7884 = n7883 ^ n7882 ;
  assign n7885 = n7884 ^ n7877 ;
  assign n7890 = n7889 ^ n7885 ;
  assign n7891 = n3980 & n7890 ;
  assign n7894 = n7891 ^ n7885 ;
  assign n7895 = n7894 ^ x189 ;
  assign n7896 = ~n4024 & n7895 ;
  assign n7897 = n7896 ^ x189 ;
  assign n7892 = n7891 ^ n7890 ;
  assign n7893 = n7892 ^ n7885 ;
  assign n7898 = n7897 ^ n7893 ;
  assign n7899 = ~n4059 & n7898 ;
  assign n7902 = n7899 ^ n7893 ;
  assign n7903 = n7902 ^ x157 ;
  assign n7904 = ~n4102 & n7903 ;
  assign n7905 = n7904 ^ x157 ;
  assign n7900 = n7899 ^ n7898 ;
  assign n7901 = n7900 ^ n7893 ;
  assign n7906 = n7905 ^ n7901 ;
  assign n7907 = n4138 & n7906 ;
  assign n7910 = n7907 ^ n7901 ;
  assign n7911 = n7910 ^ x125 ;
  assign n7912 = ~n4182 & n7911 ;
  assign n7913 = n7912 ^ x125 ;
  assign n7908 = n7907 ^ n7906 ;
  assign n7909 = n7908 ^ n7901 ;
  assign n7914 = n7913 ^ n7909 ;
  assign n7915 = n4221 & n7914 ;
  assign n7918 = n7915 ^ n7909 ;
  assign n7919 = n7918 ^ x93 ;
  assign n7920 = ~n4265 & n7919 ;
  assign n7921 = n7920 ^ x93 ;
  assign n7916 = n7915 ^ n7914 ;
  assign n7917 = n7916 ^ n7909 ;
  assign n7922 = n7921 ^ n7917 ;
  assign n7923 = ~n4300 & n7922 ;
  assign n7926 = n7923 ^ n7917 ;
  assign n7927 = n7926 ^ x61 ;
  assign n7928 = ~n4343 & n7927 ;
  assign n7929 = n7928 ^ x61 ;
  assign n7924 = n7923 ^ n7922 ;
  assign n7925 = n7924 ^ n7917 ;
  assign n7930 = n7929 ^ n7925 ;
  assign n7931 = n4379 & n7930 ;
  assign n7934 = n7931 ^ n7925 ;
  assign n7935 = n7934 ^ x29 ;
  assign n7936 = ~n4425 & n7935 ;
  assign n7937 = n7936 ^ x29 ;
  assign n7932 = n7931 ^ n7930 ;
  assign n7933 = n7932 ^ n7925 ;
  assign n7938 = n7937 ^ n7933 ;
  assign n7939 = ~n4461 & n7938 ;
  assign n7940 = n7939 ^ n7938 ;
  assign n7941 = n7940 ^ n7933 ;
  assign n7942 = x510 ^ x478 ;
  assign n7943 = ~n3330 & n7942 ;
  assign n7946 = n7943 ^ x478 ;
  assign n7947 = n7946 ^ x446 ;
  assign n7948 = ~n3377 & n7947 ;
  assign n7949 = n7948 ^ x446 ;
  assign n7944 = n7943 ^ n7942 ;
  assign n7945 = n7944 ^ x478 ;
  assign n7950 = n7949 ^ n7945 ;
  assign n7951 = ~n3413 & n7950 ;
  assign n7954 = n7951 ^ n7945 ;
  assign n7955 = n7954 ^ x414 ;
  assign n7956 = ~n3457 & n7955 ;
  assign n7957 = n7956 ^ x414 ;
  assign n7952 = n7951 ^ n7950 ;
  assign n7953 = n7952 ^ n7945 ;
  assign n7958 = n7957 ^ n7953 ;
  assign n7959 = ~n3493 & n7958 ;
  assign n7962 = n7959 ^ n7953 ;
  assign n7963 = n7962 ^ x382 ;
  assign n7964 = ~n3537 & n7963 ;
  assign n7965 = n7964 ^ x382 ;
  assign n7960 = n7959 ^ n7958 ;
  assign n7961 = n7960 ^ n7953 ;
  assign n7966 = n7965 ^ n7961 ;
  assign n7967 = n3577 & n7966 ;
  assign n7970 = n7967 ^ n7961 ;
  assign n7971 = n7970 ^ x350 ;
  assign n7972 = ~n3620 & n7971 ;
  assign n7973 = n7972 ^ x350 ;
  assign n7968 = n7967 ^ n7966 ;
  assign n7969 = n7968 ^ n7961 ;
  assign n7974 = n7973 ^ n7969 ;
  assign n7975 = n3656 & n7974 ;
  assign n7978 = n7975 ^ n7969 ;
  assign n7979 = n7978 ^ x318 ;
  assign n7980 = ~n3700 & n7979 ;
  assign n7981 = n7980 ^ x318 ;
  assign n7976 = n7975 ^ n7974 ;
  assign n7977 = n7976 ^ n7969 ;
  assign n7982 = n7981 ^ n7977 ;
  assign n7983 = n3739 & n7982 ;
  assign n7986 = n7983 ^ n7977 ;
  assign n7987 = n7986 ^ x286 ;
  assign n7988 = ~n3783 & n7987 ;
  assign n7989 = n7988 ^ x286 ;
  assign n7984 = n7983 ^ n7982 ;
  assign n7985 = n7984 ^ n7977 ;
  assign n7990 = n7989 ^ n7985 ;
  assign n7991 = ~n3818 & n7990 ;
  assign n7994 = n7991 ^ n7985 ;
  assign n7995 = n7994 ^ x254 ;
  assign n7996 = ~n3861 & n7995 ;
  assign n7997 = n7996 ^ x254 ;
  assign n7992 = n7991 ^ n7990 ;
  assign n7993 = n7992 ^ n7985 ;
  assign n7998 = n7997 ^ n7993 ;
  assign n7999 = n3897 & n7998 ;
  assign n8002 = n7999 ^ n7993 ;
  assign n8003 = n8002 ^ x222 ;
  assign n8004 = ~n3941 & n8003 ;
  assign n8005 = n8004 ^ x222 ;
  assign n8000 = n7999 ^ n7998 ;
  assign n8001 = n8000 ^ n7993 ;
  assign n8006 = n8005 ^ n8001 ;
  assign n8007 = n3980 & n8006 ;
  assign n8010 = n8007 ^ n8001 ;
  assign n8011 = n8010 ^ x190 ;
  assign n8012 = ~n4024 & n8011 ;
  assign n8013 = n8012 ^ x190 ;
  assign n8008 = n8007 ^ n8006 ;
  assign n8009 = n8008 ^ n8001 ;
  assign n8014 = n8013 ^ n8009 ;
  assign n8015 = ~n4059 & n8014 ;
  assign n8018 = n8015 ^ n8009 ;
  assign n8019 = n8018 ^ x158 ;
  assign n8020 = ~n4102 & n8019 ;
  assign n8021 = n8020 ^ x158 ;
  assign n8016 = n8015 ^ n8014 ;
  assign n8017 = n8016 ^ n8009 ;
  assign n8022 = n8021 ^ n8017 ;
  assign n8023 = n4138 & n8022 ;
  assign n8026 = n8023 ^ n8017 ;
  assign n8027 = n8026 ^ x126 ;
  assign n8028 = ~n4182 & n8027 ;
  assign n8029 = n8028 ^ x126 ;
  assign n8024 = n8023 ^ n8022 ;
  assign n8025 = n8024 ^ n8017 ;
  assign n8030 = n8029 ^ n8025 ;
  assign n8031 = n4221 & n8030 ;
  assign n8034 = n8031 ^ n8025 ;
  assign n8035 = n8034 ^ x94 ;
  assign n8036 = ~n4265 & n8035 ;
  assign n8037 = n8036 ^ x94 ;
  assign n8032 = n8031 ^ n8030 ;
  assign n8033 = n8032 ^ n8025 ;
  assign n8038 = n8037 ^ n8033 ;
  assign n8039 = ~n4300 & n8038 ;
  assign n8042 = n8039 ^ n8033 ;
  assign n8043 = n8042 ^ x62 ;
  assign n8044 = ~n4343 & n8043 ;
  assign n8045 = n8044 ^ x62 ;
  assign n8040 = n8039 ^ n8038 ;
  assign n8041 = n8040 ^ n8033 ;
  assign n8046 = n8045 ^ n8041 ;
  assign n8047 = n4379 & n8046 ;
  assign n8050 = n8047 ^ n8041 ;
  assign n8051 = n8050 ^ x30 ;
  assign n8052 = ~n4425 & n8051 ;
  assign n8053 = n8052 ^ x30 ;
  assign n8048 = n8047 ^ n8046 ;
  assign n8049 = n8048 ^ n8041 ;
  assign n8054 = n8053 ^ n8049 ;
  assign n8055 = ~n4461 & n8054 ;
  assign n8056 = n8055 ^ n8054 ;
  assign n8057 = n8056 ^ n8049 ;
  assign n8058 = x511 ^ x479 ;
  assign n8059 = ~n3330 & n8058 ;
  assign n8062 = n8059 ^ x479 ;
  assign n8063 = n8062 ^ x447 ;
  assign n8064 = ~n3377 & n8063 ;
  assign n8065 = n8064 ^ x447 ;
  assign n8060 = n8059 ^ n8058 ;
  assign n8061 = n8060 ^ x479 ;
  assign n8066 = n8065 ^ n8061 ;
  assign n8067 = ~n3413 & n8066 ;
  assign n8070 = n8067 ^ n8061 ;
  assign n8071 = n8070 ^ x415 ;
  assign n8072 = ~n3457 & n8071 ;
  assign n8073 = n8072 ^ x415 ;
  assign n8068 = n8067 ^ n8066 ;
  assign n8069 = n8068 ^ n8061 ;
  assign n8074 = n8073 ^ n8069 ;
  assign n8075 = ~n3493 & n8074 ;
  assign n8078 = n8075 ^ n8069 ;
  assign n8079 = n8078 ^ x383 ;
  assign n8080 = ~n3537 & n8079 ;
  assign n8081 = n8080 ^ x383 ;
  assign n8076 = n8075 ^ n8074 ;
  assign n8077 = n8076 ^ n8069 ;
  assign n8082 = n8081 ^ n8077 ;
  assign n8083 = n3577 & n8082 ;
  assign n8086 = n8083 ^ n8077 ;
  assign n8087 = n8086 ^ x351 ;
  assign n8088 = ~n3620 & n8087 ;
  assign n8089 = n8088 ^ x351 ;
  assign n8084 = n8083 ^ n8082 ;
  assign n8085 = n8084 ^ n8077 ;
  assign n8090 = n8089 ^ n8085 ;
  assign n8091 = n3656 & n8090 ;
  assign n8094 = n8091 ^ n8085 ;
  assign n8095 = n8094 ^ x319 ;
  assign n8096 = ~n3700 & n8095 ;
  assign n8097 = n8096 ^ x319 ;
  assign n8092 = n8091 ^ n8090 ;
  assign n8093 = n8092 ^ n8085 ;
  assign n8098 = n8097 ^ n8093 ;
  assign n8099 = n3739 & n8098 ;
  assign n8102 = n8099 ^ n8093 ;
  assign n8103 = n8102 ^ x287 ;
  assign n8104 = ~n3783 & n8103 ;
  assign n8105 = n8104 ^ x287 ;
  assign n8100 = n8099 ^ n8098 ;
  assign n8101 = n8100 ^ n8093 ;
  assign n8106 = n8105 ^ n8101 ;
  assign n8107 = ~n3818 & n8106 ;
  assign n8110 = n8107 ^ n8101 ;
  assign n8111 = n8110 ^ x255 ;
  assign n8112 = ~n3861 & n8111 ;
  assign n8113 = n8112 ^ x255 ;
  assign n8108 = n8107 ^ n8106 ;
  assign n8109 = n8108 ^ n8101 ;
  assign n8114 = n8113 ^ n8109 ;
  assign n8115 = n3897 & n8114 ;
  assign n8118 = n8115 ^ n8109 ;
  assign n8119 = n8118 ^ x223 ;
  assign n8120 = ~n3941 & n8119 ;
  assign n8121 = n8120 ^ x223 ;
  assign n8116 = n8115 ^ n8114 ;
  assign n8117 = n8116 ^ n8109 ;
  assign n8122 = n8121 ^ n8117 ;
  assign n8123 = n3980 & n8122 ;
  assign n8126 = n8123 ^ n8117 ;
  assign n8127 = n8126 ^ x191 ;
  assign n8128 = ~n4024 & n8127 ;
  assign n8129 = n8128 ^ x191 ;
  assign n8124 = n8123 ^ n8122 ;
  assign n8125 = n8124 ^ n8117 ;
  assign n8130 = n8129 ^ n8125 ;
  assign n8131 = ~n4059 & n8130 ;
  assign n8134 = n8131 ^ n8125 ;
  assign n8135 = n8134 ^ x159 ;
  assign n8136 = ~n4102 & n8135 ;
  assign n8137 = n8136 ^ x159 ;
  assign n8132 = n8131 ^ n8130 ;
  assign n8133 = n8132 ^ n8125 ;
  assign n8138 = n8137 ^ n8133 ;
  assign n8139 = n4138 & n8138 ;
  assign n8142 = n8139 ^ n8133 ;
  assign n8143 = n8142 ^ x127 ;
  assign n8144 = ~n4182 & n8143 ;
  assign n8145 = n8144 ^ x127 ;
  assign n8140 = n8139 ^ n8138 ;
  assign n8141 = n8140 ^ n8133 ;
  assign n8146 = n8145 ^ n8141 ;
  assign n8147 = n4221 & n8146 ;
  assign n8150 = n8147 ^ n8141 ;
  assign n8151 = n8150 ^ x95 ;
  assign n8152 = ~n4265 & n8151 ;
  assign n8153 = n8152 ^ x95 ;
  assign n8148 = n8147 ^ n8146 ;
  assign n8149 = n8148 ^ n8141 ;
  assign n8154 = n8153 ^ n8149 ;
  assign n8155 = ~n4300 & n8154 ;
  assign n8158 = n8155 ^ n8149 ;
  assign n8159 = n8158 ^ x63 ;
  assign n8160 = ~n4343 & n8159 ;
  assign n8161 = n8160 ^ x63 ;
  assign n8156 = n8155 ^ n8154 ;
  assign n8157 = n8156 ^ n8149 ;
  assign n8162 = n8161 ^ n8157 ;
  assign n8163 = n4379 & n8162 ;
  assign n8166 = n8163 ^ n8157 ;
  assign n8167 = n8166 ^ x31 ;
  assign n8168 = ~n4425 & n8167 ;
  assign n8169 = n8168 ^ x31 ;
  assign n8164 = n8163 ^ n8162 ;
  assign n8165 = n8164 ^ n8157 ;
  assign n8170 = n8169 ^ n8165 ;
  assign n8171 = ~n4461 & n8170 ;
  assign n8172 = n8171 ^ n8170 ;
  assign n8173 = n8172 ^ n8165 ;
  assign n8174 = n4575 ^ n4569 ;
  assign n8175 = n4691 ^ n4685 ;
  assign n8176 = n4807 ^ n4801 ;
  assign n8177 = n4923 ^ n4917 ;
  assign n8178 = n5039 ^ n5033 ;
  assign n8179 = n5155 ^ n5149 ;
  assign n8180 = n5271 ^ n5265 ;
  assign n8181 = n5387 ^ n5381 ;
  assign n8182 = n5503 ^ n5497 ;
  assign n8183 = n5619 ^ n5613 ;
  assign n8184 = n5735 ^ n5729 ;
  assign n8185 = n5851 ^ n5845 ;
  assign n8186 = n5967 ^ n5961 ;
  assign n8187 = n6083 ^ n6077 ;
  assign n8188 = n6199 ^ n6193 ;
  assign n8189 = n6315 ^ n6309 ;
  assign n8190 = n6431 ^ n6425 ;
  assign n8191 = n6547 ^ n6541 ;
  assign n8192 = n6663 ^ n6657 ;
  assign n8193 = n6779 ^ n6773 ;
  assign n8194 = n6895 ^ n6889 ;
  assign n8195 = n7011 ^ n7005 ;
  assign n8196 = n7127 ^ n7121 ;
  assign n8197 = n7243 ^ n7237 ;
  assign n8198 = n7359 ^ n7353 ;
  assign n8199 = n7475 ^ n7469 ;
  assign n8200 = n7591 ^ n7585 ;
  assign n8201 = n7707 ^ n7701 ;
  assign n8202 = n7823 ^ n7817 ;
  assign n8203 = n7939 ^ n7933 ;
  assign n8204 = n8055 ^ n8049 ;
  assign n8205 = n8171 ^ n8165 ;
  assign y0 = n4577 ;
  assign y1 = n4693 ;
  assign y2 = n4809 ;
  assign y3 = n4925 ;
  assign y4 = n5041 ;
  assign y5 = n5157 ;
  assign y6 = n5273 ;
  assign y7 = n5389 ;
  assign y8 = n5505 ;
  assign y9 = n5621 ;
  assign y10 = n5737 ;
  assign y11 = n5853 ;
  assign y12 = n5969 ;
  assign y13 = n6085 ;
  assign y14 = n6201 ;
  assign y15 = n6317 ;
  assign y16 = n6433 ;
  assign y17 = n6549 ;
  assign y18 = n6665 ;
  assign y19 = n6781 ;
  assign y20 = n6897 ;
  assign y21 = n7013 ;
  assign y22 = n7129 ;
  assign y23 = n7245 ;
  assign y24 = n7361 ;
  assign y25 = n7477 ;
  assign y26 = n7593 ;
  assign y27 = n7709 ;
  assign y28 = n7825 ;
  assign y29 = n7941 ;
  assign y30 = n8057 ;
  assign y31 = n8173 ;
  assign y32 = n8174 ;
  assign y33 = n8175 ;
  assign y34 = n8176 ;
  assign y35 = n8177 ;
  assign y36 = n8178 ;
  assign y37 = n8179 ;
  assign y38 = n8180 ;
  assign y39 = n8181 ;
  assign y40 = n8182 ;
  assign y41 = n8183 ;
  assign y42 = n8184 ;
  assign y43 = n8185 ;
  assign y44 = n8186 ;
  assign y45 = n8187 ;
  assign y46 = n8188 ;
  assign y47 = n8189 ;
  assign y48 = n8190 ;
  assign y49 = n8191 ;
  assign y50 = n8192 ;
  assign y51 = n8193 ;
  assign y52 = n8194 ;
  assign y53 = n8195 ;
  assign y54 = n8196 ;
  assign y55 = n8197 ;
  assign y56 = n8198 ;
  assign y57 = n8199 ;
  assign y58 = n8200 ;
  assign y59 = n8201 ;
  assign y60 = n8202 ;
  assign y61 = n8203 ;
  assign y62 = n8204 ;
  assign y63 = n8205 ;
endmodule
