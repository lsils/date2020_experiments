module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336;
  assign n25 = x2 ^ x1;
  assign n62 = x19 & ~x22;
  assign n27 = ~x0 & x1;
  assign n28 = n27 ^ x0;
  assign n29 = ~n25 & ~n28;
  assign n30 = ~x3 & n29;
  assign n31 = ~x4 & n30;
  assign n32 = ~x5 & n31;
  assign n33 = ~x6 & ~x7;
  assign n34 = n32 & n33;
  assign n35 = ~x8 & n34;
  assign n36 = ~x9 & n35;
  assign n37 = ~x10 & n36;
  assign n38 = ~x11 & n37;
  assign n39 = ~x12 & ~x13;
  assign n40 = ~x14 & n39;
  assign n41 = n38 & n40;
  assign n45 = ~x15 & n41;
  assign n86 = n45 ^ x18;
  assign n87 = n86 ^ x22;
  assign n88 = x17 ^ x16;
  assign n89 = ~n45 & ~n88;
  assign n47 = ~x16 & x17;
  assign n48 = n47 ^ x16;
  assign n90 = n89 ^ n48;
  assign n91 = n90 ^ n86;
  assign n92 = n87 & n91;
  assign n93 = n92 ^ n89;
  assign n94 = n93 ^ n48;
  assign n95 = n94 ^ x22;
  assign n96 = ~n86 & n95;
  assign n97 = n96 ^ n86;
  assign n49 = x18 & ~x19;
  assign n50 = n49 ^ x18;
  assign n135 = ~n48 & n50;
  assign n136 = n97 & ~n135;
  assign n137 = ~n62 & ~n136;
  assign n26 = x22 ^ x21;
  assign n46 = ~x22 & ~n45;
  assign n51 = n50 ^ x19;
  assign n52 = n51 ^ x18;
  assign n53 = ~n48 & ~n52;
  assign n54 = ~n46 & n53;
  assign n55 = ~x22 & ~n54;
  assign n56 = n55 ^ x20;
  assign n57 = ~n26 & n56;
  assign n147 = n57 ^ n56;
  assign n42 = ~x22 & ~n41;
  assign n43 = n42 ^ x15;
  assign n74 = n43 & ~n56;
  assign n75 = n74 ^ n43;
  assign n58 = ~n43 & ~n57;
  assign n59 = n58 ^ n43;
  assign n60 = n59 ^ n57;
  assign n76 = n75 ^ n60;
  assign n203 = n147 ^ n76;
  assign n237 = n137 & ~n203;
  assign n68 = n48 ^ x17;
  assign n121 = n62 ^ x22;
  assign n81 = x22 & n49;
  assign n120 = n81 ^ n49;
  assign n122 = n121 ^ n120;
  assign n149 = n122 ^ n52;
  assign n158 = n68 & n149;
  assign n65 = n62 ^ x19;
  assign n63 = ~x18 & n62;
  assign n64 = n63 ^ n51;
  assign n66 = n65 ^ n64;
  assign n67 = n66 ^ n50;
  assign n77 = n45 ^ x16;
  assign n78 = ~x17 & ~n77;
  assign n79 = n78 ^ n77;
  assign n157 = n67 & ~n79;
  assign n159 = n158 ^ n157;
  assign n104 = x21 ^ x20;
  assign n105 = n55 ^ x21;
  assign n106 = n104 & n105;
  assign n44 = ~n26 & n43;
  assign n61 = n60 ^ n44;
  assign n183 = n106 ^ n61;
  assign n236 = n159 & ~n183;
  assign n238 = n237 ^ n236;
  assign n69 = n68 ^ x16;
  assign n168 = n64 & n69;
  assign n167 = n78 & n120;
  assign n169 = n168 ^ n167;
  assign n117 = n26 & ~n104;
  assign n118 = ~n43 & n117;
  assign n241 = n118 ^ n75;
  assign n242 = n169 & n241;
  assign n239 = n118 & n169;
  assign n190 = n57 & n169;
  assign n171 = ~n43 & n169;
  assign n170 = n58 & n169;
  assign n172 = n171 ^ n170;
  assign n191 = n190 ^ n172;
  assign n240 = n239 ^ n191;
  assign n243 = n242 ^ n240;
  assign n127 = n66 & n68;
  assign n126 = ~n79 & ~n122;
  assign n128 = n127 ^ n126;
  assign n195 = n106 & n128;
  assign n175 = ~n61 & n128;
  assign n196 = n195 ^ n175;
  assign n244 = n243 ^ n196;
  assign n245 = ~n238 & ~n244;
  assign n70 = ~n45 & n69;
  assign n71 = n67 & n70;
  assign n72 = n71 ^ n54;
  assign n247 = n72 ^ n61;
  assign n73 = n61 & ~n72;
  assign n248 = n247 ^ n73;
  assign n246 = n128 & ~n203;
  assign n249 = n248 ^ n246;
  assign n119 = n118 ^ n117;
  assign n153 = n47 & n149;
  assign n130 = n90 ^ n77;
  assign n152 = n67 & ~n130;
  assign n154 = n153 ^ n152;
  assign n251 = n119 & n154;
  assign n82 = n68 & n81;
  assign n80 = n63 & ~n79;
  assign n83 = n82 ^ n80;
  assign n250 = n83 & ~n203;
  assign n252 = n251 ^ n250;
  assign n253 = ~n249 & ~n252;
  assign n254 = n245 & n253;
  assign n225 = n69 & n81;
  assign n224 = n63 & n78;
  assign n226 = n225 ^ n224;
  assign n99 = ~n48 & n81;
  assign n98 = x19 & ~n97;
  assign n100 = n99 ^ n98;
  assign n261 = n226 ^ n100;
  assign n262 = n57 & n261;
  assign n256 = ~n46 & n51;
  assign n257 = ~n48 & n256;
  assign n255 = n70 & n120;
  assign n258 = n257 ^ n255;
  assign n214 = n64 & n68;
  assign n213 = ~n79 & n120;
  assign n215 = n214 ^ n213;
  assign n259 = n258 ^ n215;
  assign n260 = n106 & n259;
  assign n263 = n262 ^ n260;
  assign n270 = n57 & n128;
  assign n267 = n169 & ~n183;
  assign n266 = n239 ^ n170;
  assign n268 = n267 ^ n266;
  assign n264 = n117 & n159;
  assign n265 = n264 ^ n72;
  assign n269 = n268 ^ n265;
  assign n271 = n270 ^ n269;
  assign n272 = ~n263 & ~n271;
  assign n207 = n47 & n81;
  assign n206 = n63 & ~n130;
  assign n208 = n207 ^ n206;
  assign n280 = n76 & ~n208;
  assign n279 = n208 ^ n76;
  assign n281 = n280 ^ n279;
  assign n150 = n69 & n149;
  assign n148 = n67 & n78;
  assign n151 = n150 ^ n148;
  assign n277 = n118 & n151;
  assign n276 = n117 & n151;
  assign n278 = n277 ^ n276;
  assign n282 = n281 ^ n278;
  assign n124 = n66 & n69;
  assign n123 = n78 & ~n122;
  assign n125 = n124 ^ n123;
  assign n274 = ~n61 & n125;
  assign n273 = ~n60 & n208;
  assign n275 = n274 ^ n273;
  assign n283 = n282 ^ n275;
  assign n284 = n272 & ~n283;
  assign n132 = n47 & n66;
  assign n131 = ~n122 & ~n130;
  assign n133 = n132 ^ n131;
  assign n287 = ~n59 & n133;
  assign n285 = ~n61 & n159;
  assign n286 = n285 ^ n277;
  assign n288 = n287 ^ n286;
  assign n293 = ~n76 & n137;
  assign n290 = n118 & n154;
  assign n289 = n100 & n118;
  assign n291 = n290 ^ n289;
  assign n218 = n57 & n215;
  assign n216 = ~n43 & n215;
  assign n217 = n57 & n216;
  assign n219 = n218 ^ n217;
  assign n292 = n291 ^ n219;
  assign n294 = n293 ^ n292;
  assign n295 = ~n288 & ~n294;
  assign n296 = n284 & n295;
  assign n297 = n254 & n296;
  assign n101 = n76 & ~n100;
  assign n84 = ~n76 & n83;
  assign n85 = n84 ^ n83;
  assign n102 = n101 ^ n85;
  assign n103 = ~n73 & ~n102;
  assign n110 = ~n59 & n72;
  assign n109 = ~n60 & n72;
  assign n111 = n110 ^ n109;
  assign n112 = n75 ^ n56;
  assign n113 = n72 & n112;
  assign n114 = ~n111 & ~n113;
  assign n115 = n114 ^ n111;
  assign n107 = n100 ^ n83;
  assign n108 = n106 & n107;
  assign n116 = n115 ^ n108;
  assign n129 = n128 ^ n125;
  assign n134 = n133 ^ n129;
  assign n142 = n118 & ~n134;
  assign n143 = n142 ^ n118;
  assign n138 = n137 ^ n133;
  assign n139 = n43 & n138;
  assign n140 = ~n134 & ~n139;
  assign n141 = n119 & ~n140;
  assign n144 = n143 ^ n141;
  assign n145 = n116 & ~n144;
  assign n146 = ~n103 & n145;
  assign n164 = n47 & n64;
  assign n163 = n120 & ~n130;
  assign n165 = n164 ^ n163;
  assign n166 = ~n59 & n165;
  assign n173 = n172 ^ n166;
  assign n179 = n57 & n151;
  assign n177 = ~n60 & n165;
  assign n174 = ~n61 & n137;
  assign n176 = n175 ^ n174;
  assign n178 = n177 ^ n176;
  assign n180 = n179 ^ n178;
  assign n181 = ~n173 & ~n180;
  assign n298 = ~n59 & n159;
  assign n194 = n137 & ~n183;
  assign n299 = n298 ^ n194;
  assign n307 = ~n118 & ~n226;
  assign n309 = n76 & n307;
  assign n308 = n307 ^ n76;
  assign n310 = n309 ^ n308;
  assign n186 = ~n76 & n125;
  assign n311 = n310 ^ n186;
  assign n303 = ~n43 & n208;
  assign n304 = n147 & n303;
  assign n301 = ~n59 & n226;
  assign n300 = n112 & n226;
  assign n302 = n301 ^ n300;
  assign n305 = n304 ^ n302;
  assign n306 = n305 ^ n84;
  assign n312 = n311 ^ n306;
  assign n313 = ~n299 & n312;
  assign n314 = n181 & n313;
  assign n315 = n146 & n314;
  assign n316 = n297 & n315;
  assign n184 = n183 ^ n76;
  assign n185 = n125 & n184;
  assign n187 = n186 ^ n185;
  assign n182 = ~n57 & ~n133;
  assign n188 = n187 ^ n182;
  assign n189 = ~n106 & ~n137;
  assign n192 = n191 ^ n189;
  assign n193 = ~n188 & ~n192;
  assign n197 = n196 ^ n194;
  assign n198 = ~n193 & ~n197;
  assign n199 = n181 & n198;
  assign n419 = ~n61 & n208;
  assign n544 = n226 ^ n169;
  assign n545 = n544 ^ n165;
  assign n546 = n106 & n545;
  assign n547 = ~n419 & ~n546;
  assign n548 = ~n263 & n547;
  assign n549 = n274 ^ n57;
  assign n550 = n548 & ~n549;
  assign n551 = n199 & n550;
  assign n552 = ~x22 & ~n38;
  assign n751 = n552 ^ x12;
  assign n752 = ~x22 & ~n37;
  assign n753 = n752 ^ x11;
  assign n1954 = n751 & n753;
  assign n754 = n753 ^ n751;
  assign n1955 = n1954 ^ n754;
  assign n553 = x12 & ~x22;
  assign n554 = ~n552 & ~n553;
  assign n581 = x13 & ~x22;
  assign n582 = n554 & ~n581;
  assign n583 = n582 ^ x14;
  assign n555 = n554 ^ x13;
  assign n584 = n583 ^ n555;
  assign n1956 = n1955 ^ n584;
  assign n1957 = ~n551 & ~n1956;
  assign n557 = n106 & n551;
  assign n204 = n125 & ~n203;
  assign n200 = n169 ^ n128;
  assign n201 = n200 ^ n139;
  assign n202 = n147 & n201;
  assign n205 = n204 ^ n202;
  assign n565 = ~n76 & n165;
  assign n566 = n565 ^ n186;
  assign n561 = n159 ^ n72;
  assign n155 = n154 ^ n151;
  assign n562 = n561 ^ n155;
  assign n563 = ~n183 & n562;
  assign n363 = ~n61 & n133;
  assign n559 = n363 ^ n133;
  assign n445 = n203 ^ n61;
  assign n558 = n133 & ~n445;
  assign n560 = n559 ^ n558;
  assign n564 = n563 ^ n560;
  assign n567 = n566 ^ n564;
  assign n568 = ~n237 & ~n567;
  assign n569 = ~n205 & n568;
  assign n570 = ~n557 & n569;
  assign n1958 = n570 & ~n583;
  assign n1959 = n1958 ^ n583;
  assign n1960 = ~n1957 & n1959;
  assign n348 = ~n60 & n128;
  assign n347 = n75 & n128;
  assign n349 = n348 ^ n347;
  assign n342 = n83 & n118;
  assign n334 = ~n83 & ~n119;
  assign n333 = n119 ^ n83;
  assign n335 = n334 ^ n333;
  assign n343 = n342 ^ n335;
  assign n340 = n183 ^ n118;
  assign n341 = n83 & ~n340;
  assign n344 = n343 ^ n341;
  assign n337 = n106 & n151;
  assign n336 = ~n61 & n151;
  assign n338 = n337 ^ n336;
  assign n339 = n338 ^ n335;
  assign n345 = n344 ^ n339;
  assign n346 = n345 ^ n194;
  assign n350 = n349 ^ n346;
  assign n446 = ~n43 & ~n165;
  assign n447 = n165 ^ n83;
  assign n448 = ~n446 & n447;
  assign n449 = n445 & n448;
  assign n450 = n133 & ~n183;
  assign n319 = n118 & n258;
  assign n451 = n450 ^ n319;
  assign n452 = ~n449 & ~n451;
  assign n689 = ~n350 & n452;
  assign n676 = n147 & n216;
  assign n666 = n57 & n125;
  assign n428 = ~n60 & n125;
  assign n667 = n666 ^ n428;
  assign n690 = n676 ^ n667;
  assign n373 = n119 & n165;
  assign n691 = n690 ^ n373;
  assign n692 = n100 ^ n76;
  assign n693 = n692 ^ n101;
  assign n370 = n112 & n258;
  assign n317 = n118 ^ n59;
  assign n318 = n258 & ~n317;
  assign n320 = n319 ^ n318;
  assign n371 = n370 ^ n320;
  assign n694 = n693 ^ n371;
  assign n695 = ~n691 & ~n694;
  assign n696 = n689 & n695;
  assign n700 = ~n61 & n169;
  assign n701 = n700 ^ n320;
  assign n383 = ~n61 & n100;
  assign n702 = n701 ^ n383;
  assign n574 = n118 & n137;
  assign n697 = n574 ^ n186;
  assign n698 = n697 ^ n273;
  assign n699 = n698 ^ n336;
  assign n703 = n702 ^ n699;
  assign n704 = n696 & ~n703;
  assign n456 = n363 ^ n173;
  assign n453 = n57 & n303;
  assign n454 = n453 ^ n217;
  assign n412 = ~n76 & n133;
  assign n413 = n412 ^ n250;
  assign n455 = n454 ^ n413;
  assign n457 = n456 ^ n455;
  assign n639 = ~n57 & ~n208;
  assign n705 = n307 ^ n117;
  assign n670 = n117 & n226;
  assign n706 = n705 ^ n670;
  assign n707 = n706 ^ n219;
  assign n708 = ~n639 & ~n707;
  assign n683 = n348 ^ n270;
  assign n709 = n683 ^ n560;
  assign n481 = n226 ^ n60;
  assign n479 = n44 & n226;
  assign n227 = ~n61 & n226;
  assign n480 = n479 ^ n227;
  assign n482 = n481 ^ n480;
  assign n484 = n119 & n133;
  assign n483 = n133 ^ n119;
  assign n485 = n484 ^ n483;
  assign n486 = ~n482 & n485;
  assign n710 = n709 ^ n486;
  assign n711 = ~n708 & ~n710;
  assign n712 = ~n457 & n711;
  assign n656 = n75 & n258;
  assign n713 = n656 ^ n115;
  assign n714 = n560 ^ n174;
  assign n461 = n100 & ~n203;
  assign n715 = n714 ^ n461;
  assign n716 = n713 & ~n715;
  assign n426 = n226 ^ n118;
  assign n427 = n426 ^ n307;
  assign n717 = n427 ^ n204;
  assign n718 = n717 ^ n277;
  assign n719 = n716 & n718;
  assign n720 = n712 & n719;
  assign n721 = n704 & n720;
  assign n522 = n57 & n83;
  assign n430 = n118 & n208;
  assign n722 = n522 ^ n430;
  assign n723 = n722 ^ n251;
  assign n492 = n119 & n169;
  assign n352 = n119 & n125;
  assign n351 = n117 & n125;
  assign n353 = n352 ^ n351;
  assign n724 = n492 ^ n353;
  assign n725 = ~n723 & ~n724;
  assign n355 = ~n76 & n151;
  assign n726 = n355 ^ n352;
  assign n727 = n726 ^ n278;
  assign n731 = n428 ^ n191;
  assign n732 = n731 ^ n177;
  assign n733 = n732 ^ n287;
  assign n728 = n303 ^ n128;
  assign n729 = n106 & n728;
  assign n730 = n729 ^ n290;
  assign n734 = n733 ^ n730;
  assign n735 = ~n727 & ~n734;
  assign n736 = n725 & n735;
  assign n374 = ~n76 & n215;
  assign n738 = n374 ^ n348;
  assign n737 = ~n59 & n137;
  assign n739 = n738 ^ n737;
  assign n743 = n383 ^ n267;
  assign n380 = ~n100 & ~n106;
  assign n379 = n106 ^ n100;
  assign n381 = n380 ^ n379;
  assign n744 = n743 ^ n381;
  assign n740 = n72 & ~n76;
  assign n532 = n137 ^ n59;
  assign n530 = n60 & ~n137;
  assign n531 = n530 ^ n57;
  assign n533 = n532 ^ n531;
  assign n741 = n740 ^ n533;
  assign n742 = n741 ^ n239;
  assign n745 = n744 ^ n742;
  assign n746 = ~n739 & n745;
  assign n747 = n736 & n746;
  assign n748 = n721 & n747;
  assign n365 = ~n60 & n159;
  assign n589 = n449 ^ n365;
  assign n590 = n589 ^ n183;
  assign n591 = n446 ^ n303;
  assign n592 = ~n590 & ~n591;
  assign n415 = n75 & n159;
  assign n416 = n415 ^ n365;
  assign n593 = n416 ^ n251;
  assign n436 = ~n119 & ~n137;
  assign n435 = n137 ^ n119;
  assign n437 = n436 ^ n435;
  assign n525 = n437 ^ n338;
  assign n594 = n558 ^ n525;
  assign n595 = ~n593 & n594;
  assign n596 = ~n592 & n595;
  assign n597 = n203 & n596;
  assign n598 = n109 ^ n72;
  assign n599 = n598 ^ n482;
  assign n600 = ~n597 & ~n599;
  assign n601 = n133 ^ n100;
  assign n602 = n106 & n562;
  assign n603 = n602 ^ n106;
  assign n604 = n603 ^ n142;
  assign n605 = ~n601 & ~n604;
  assign n606 = n83 ^ n59;
  assign n223 = ~n60 & n83;
  assign n523 = n522 ^ n223;
  assign n607 = n606 ^ n523;
  assign n608 = ~n605 & ~n607;
  assign n609 = n226 ^ n133;
  assign n610 = n183 & ~n609;
  assign n405 = n119 & n208;
  assign n611 = n405 ^ n208;
  assign n612 = n611 ^ n334;
  assign n613 = ~n610 & ~n612;
  assign n402 = ~n60 & n154;
  assign n614 = n402 ^ n191;
  assign n212 = ~n60 & n100;
  assign n615 = n614 ^ n212;
  assign n616 = ~n613 & ~n615;
  assign n617 = ~n60 & n151;
  assign n618 = n617 ^ n179;
  assign n619 = n618 ^ n173;
  assign n620 = n616 & ~n619;
  assign n621 = ~n608 & n620;
  assign n622 = ~n600 & n621;
  assign n625 = n319 ^ n310;
  assign n623 = n165 & ~n203;
  assign n624 = n623 ^ n428;
  assign n626 = n625 ^ n624;
  assign n627 = n622 & n626;
  assign n629 = n335 ^ n248;
  assign n628 = n370 ^ n298;
  assign n630 = n629 ^ n628;
  assign n631 = n525 ^ n289;
  assign n632 = n631 ^ n383;
  assign n633 = n630 & n632;
  assign n634 = n258 ^ n119;
  assign n575 = n119 & n258;
  assign n635 = n634 ^ n575;
  assign n636 = ~n72 & ~n635;
  assign n637 = ~n101 & ~n636;
  assign n322 = n118 & n128;
  assign n466 = n353 ^ n322;
  assign n467 = n466 ^ n143;
  assign n638 = n467 ^ n303;
  assign n642 = n215 ^ n208;
  assign n640 = n215 ^ n57;
  assign n641 = n640 ^ n218;
  assign n643 = n642 ^ n641;
  assign n644 = n643 ^ n639;
  assign n645 = ~n638 & n644;
  assign n646 = ~n637 & n645;
  assign n650 = n301 ^ n110;
  assign n651 = n650 ^ n523;
  assign n647 = n226 ^ n72;
  assign n648 = n57 & n647;
  assign n649 = n648 ^ n374;
  assign n652 = n651 ^ n649;
  assign n653 = n646 & ~n652;
  assign n654 = n633 & n653;
  assign n655 = n627 & n654;
  assign n498 = ~n76 & n258;
  assign n657 = n656 ^ n498;
  assign n658 = n657 ^ n301;
  assign n659 = n658 ^ n427;
  assign n464 = n336 ^ n84;
  assign n660 = n659 ^ n464;
  assign n661 = n72 ^ n59;
  assign n662 = n661 ^ n110;
  assign n663 = ~n189 & ~n662;
  assign n664 = n663 ^ n322;
  assign n665 = n660 & ~n664;
  assign n671 = n670 ^ n427;
  assign n672 = n671 ^ n172;
  assign n515 = n226 ^ n208;
  assign n668 = ~n76 & n515;
  assign n669 = n668 ^ n667;
  assign n673 = n672 ^ n669;
  assign n489 = n43 & n154;
  assign n490 = n106 & n489;
  assign n677 = n676 ^ n490;
  assign n678 = n677 ^ n348;
  assign n674 = n187 ^ n110;
  assign n675 = n674 ^ n533;
  assign n679 = n678 ^ n675;
  assign n680 = n673 & ~n679;
  assign n681 = n145 & n680;
  assign n682 = n665 & n681;
  assign n401 = n57 & n154;
  assign n403 = n402 ^ n401;
  assign n400 = n154 & ~n183;
  assign n404 = n403 ^ n400;
  assign n406 = n405 ^ n404;
  assign n408 = n274 ^ n236;
  assign n409 = n408 ^ n352;
  assign n407 = n223 ^ n177;
  assign n410 = n409 ^ n407;
  assign n411 = ~n406 & ~n410;
  assign n684 = n683 ^ n285;
  assign n685 = n684 ^ n617;
  assign n686 = n411 & ~n685;
  assign n687 = n682 & n686;
  assign n688 = n655 & n687;
  assign n758 = n748 ^ n688;
  assign n571 = n215 ^ n169;
  assign n572 = n571 ^ n165;
  assign n573 = n117 & n572;
  assign n576 = n575 ^ n574;
  assign n577 = ~n573 & ~n576;
  assign n578 = n146 & n577;
  assign n579 = n570 & n578;
  assign n759 = n688 ^ n579;
  assign n760 = n688 ^ n583;
  assign n761 = n759 & n760;
  assign n762 = n761 ^ n688;
  assign n763 = ~n758 & ~n762;
  assign n764 = n763 ^ n579;
  assign n749 = ~n688 & ~n748;
  assign n750 = ~n579 & ~n749;
  assign n755 = ~n551 & n754;
  assign n756 = ~n750 & ~n755;
  assign n782 = n555 & ~n756;
  assign n556 = ~n551 & n555;
  assign n580 = ~n147 & n579;
  assign n585 = n570 & n584;
  assign n586 = n585 ^ n555;
  assign n587 = ~n580 & ~n586;
  assign n588 = ~n556 & ~n587;
  assign n765 = ~n551 & ~n751;
  assign n766 = n580 & ~n765;
  assign n767 = n556 ^ n555;
  assign n768 = n767 ^ n751;
  assign n769 = n570 & ~n768;
  assign n770 = n769 ^ n751;
  assign n771 = ~n766 & n770;
  assign n781 = n588 & ~n771;
  assign n783 = n782 ^ n781;
  assign n784 = n764 & n783;
  assign n785 = n784 ^ n781;
  assign n786 = ~n551 & n785;
  assign n775 = n588 & ~n756;
  assign n757 = n756 ^ n588;
  assign n772 = n764 & ~n771;
  assign n773 = ~n757 & n772;
  assign n1952 = n775 ^ n773;
  assign n1953 = ~n786 & ~n1952;
  assign n1961 = n1960 ^ n1953;
  assign n2300 = ~n555 & ~n1955;
  assign n2301 = n2300 ^ n1955;
  assign n2302 = ~n583 & n2301;
  assign n2303 = ~n551 & n2302;
  assign n2304 = n1959 & ~n2303;
  assign n2306 = n2300 ^ n555;
  assign n2307 = ~n551 & ~n2306;
  assign n2350 = n2304 & ~n2307;
  assign n793 = ~x22 & ~n35;
  assign n794 = n793 ^ x9;
  assign n791 = ~x22 & ~n36;
  assign n792 = n791 ^ x10;
  assign n795 = n794 ^ n792;
  assign n360 = ~n61 & n258;
  assign n359 = n106 & n258;
  assign n361 = n360 ^ n359;
  assign n834 = n560 ^ n361;
  assign n378 = n100 & n119;
  assign n382 = n381 ^ n378;
  assign n384 = n383 ^ n382;
  assign n835 = n834 ^ n384;
  assign n836 = n335 ^ n186;
  assign n837 = n835 & n836;
  assign n838 = ~n280 & n635;
  assign n839 = n838 ^ n322;
  assign n840 = n118 & n215;
  assign n841 = n840 ^ n250;
  assign n842 = n841 ^ n618;
  assign n843 = ~n839 & ~n842;
  assign n844 = n837 & n843;
  assign n418 = n106 & n208;
  assign n420 = n419 ^ n418;
  assign n845 = n420 ^ n194;
  assign n325 = n165 & ~n183;
  assign n846 = n845 ^ n325;
  assign n847 = n846 ^ n659;
  assign n848 = n844 & n847;
  assign n854 = n352 ^ n243;
  assign n855 = n854 ^ n479;
  assign n850 = ~n118 & ~n147;
  assign n849 = n147 ^ n118;
  assign n851 = n850 ^ n849;
  assign n326 = ~n43 & ~n151;
  assign n327 = ~n147 & n326;
  assign n328 = n327 ^ n326;
  assign n329 = n328 ^ n203;
  assign n852 = n851 ^ n329;
  assign n853 = n852 ^ n239;
  assign n856 = n855 ^ n853;
  assign n857 = n119 ^ n59;
  assign n858 = n561 & ~n857;
  assign n395 = n118 & n165;
  assign n859 = n574 ^ n395;
  assign n860 = n859 ^ n246;
  assign n861 = ~n858 & ~n860;
  assign n862 = n617 ^ n461;
  assign n863 = n861 & ~n862;
  assign n864 = ~n856 & n863;
  assign n865 = n236 ^ n175;
  assign n866 = n865 ^ n490;
  assign n867 = n866 ^ n133;
  assign n868 = n106 & n867;
  assign n870 = ~n59 & n100;
  assign n871 = n870 ^ n298;
  assign n872 = n871 ^ n109;
  assign n869 = n250 ^ n212;
  assign n873 = n872 ^ n869;
  assign n874 = n873 ^ n282;
  assign n875 = ~n868 & ~n874;
  assign n876 = n864 & n875;
  assign n877 = n848 & n876;
  assign n878 = n676 ^ n304;
  assign n879 = n878 ^ n484;
  assign n880 = ~n318 & ~n879;
  assign n881 = ~n416 & n880;
  assign n882 = n251 ^ n103;
  assign n809 = n226 ^ n137;
  assign n810 = n809 ^ n154;
  assign n811 = ~n76 & n810;
  assign n883 = n811 ^ n217;
  assign n884 = ~n882 & ~n883;
  assign n885 = n881 & n884;
  assign n510 = ~n61 & n215;
  assign n886 = n700 ^ n510;
  assign n887 = n886 ^ n623;
  assign n536 = n118 & n159;
  assign n817 = n536 ^ n264;
  assign n888 = n817 ^ n467;
  assign n889 = ~n887 & ~n888;
  assign n890 = n885 & n889;
  assign n891 = n877 & n890;
  assign n796 = n215 ^ n151;
  assign n797 = ~n445 & ~n796;
  assign n798 = n530 ^ n329;
  assign n799 = ~n797 & n798;
  assign n424 = n119 & n215;
  assign n801 = n424 ^ n363;
  assign n800 = n739 ^ n196;
  assign n802 = n801 ^ n800;
  assign n803 = ~n799 & ~n802;
  assign n804 = n467 ^ n177;
  assign n805 = ~n697 & ~n804;
  assign n478 = n325 ^ n204;
  assign n806 = n478 ^ n404;
  assign n807 = n805 & ~n806;
  assign n808 = n803 & n807;
  assign n491 = n490 ^ n335;
  assign n812 = n491 ^ n395;
  assign n813 = ~n286 & n812;
  assign n814 = n536 ^ n413;
  assign n815 = n813 & ~n814;
  assign n816 = ~n811 & n815;
  assign n460 = n154 & ~n203;
  assign n818 = n817 ^ n460;
  assign n819 = n818 ^ n741;
  assign n820 = n683 ^ n360;
  assign n821 = n820 ^ n510;
  assign n423 = n106 & n216;
  assign n493 = n492 ^ n423;
  assign n822 = n821 ^ n493;
  assign n823 = ~n819 & ~n822;
  assign n825 = n450 ^ n246;
  assign n433 = n119 & n128;
  assign n824 = n433 ^ n278;
  assign n826 = n825 ^ n824;
  assign n827 = n666 ^ n175;
  assign n828 = n827 ^ n693;
  assign n829 = ~n826 & ~n828;
  assign n830 = n823 & n829;
  assign n831 = n816 & n830;
  assign n832 = n808 & n831;
  assign n833 = n627 & n832;
  assign n893 = n891 ^ n833;
  assign n892 = n833 & n891;
  assign n894 = n893 ^ n892;
  assign n896 = n748 & ~n894;
  assign n895 = n894 ^ n748;
  assign n897 = n896 ^ n895;
  assign n898 = n897 ^ n792;
  assign n899 = n795 & n898;
  assign n900 = n899 ^ n794;
  assign n905 = n900 ^ n753;
  assign n906 = ~n551 & n905;
  assign n901 = n771 ^ n764;
  assign n907 = n906 ^ n901;
  assign n915 = n580 ^ n570;
  assign n916 = n751 & n915;
  assign n917 = n570 ^ n551;
  assign n918 = n753 & n917;
  assign n919 = n918 ^ n551;
  assign n920 = ~n916 & n919;
  assign n908 = n579 ^ n555;
  assign n909 = n748 ^ n579;
  assign n910 = n759 & n909;
  assign n911 = n908 & n910;
  assign n912 = n583 ^ n579;
  assign n913 = n758 & n912;
  assign n914 = ~n911 & ~n913;
  assign n921 = n920 ^ n914;
  assign n926 = n758 & n908;
  assign n924 = n751 ^ n579;
  assign n925 = n910 & ~n924;
  assign n927 = n926 ^ n925;
  assign n922 = ~n551 & ~n794;
  assign n923 = n922 ^ n551;
  assign n928 = n927 ^ n923;
  assign n929 = n833 ^ n748;
  assign n930 = n833 ^ n583;
  assign n931 = n929 & n930;
  assign n932 = n931 ^ n833;
  assign n933 = ~n893 & ~n932;
  assign n934 = n933 ^ n748;
  assign n935 = n934 ^ n923;
  assign n936 = n928 & n935;
  assign n937 = n936 ^ n927;
  assign n938 = n937 ^ n914;
  assign n939 = ~n921 & ~n938;
  assign n940 = n939 ^ n937;
  assign n941 = n940 ^ n907;
  assign n942 = n941 ^ n753;
  assign n943 = n942 ^ n905;
  assign n944 = n907 & ~n943;
  assign n902 = n900 & ~n901;
  assign n903 = n551 & n902;
  assign n904 = n903 ^ n900;
  assign n945 = n944 ^ n904;
  assign n774 = n551 & n757;
  assign n776 = n775 ^ n757;
  assign n777 = ~n753 & n776;
  assign n778 = ~n774 & ~n777;
  assign n779 = n771 & ~n778;
  assign n780 = ~n773 & ~n779;
  assign n787 = ~n774 & ~n775;
  assign n788 = ~n764 & ~n787;
  assign n789 = ~n786 & ~n788;
  assign n790 = n780 & n789;
  assign n946 = n945 ^ n790;
  assign n1082 = n748 ^ n555;
  assign n1109 = n893 & n1082;
  assign n1083 = ~n748 & n892;
  assign n1084 = n1083 ^ n896;
  assign n1107 = n751 ^ n748;
  assign n1108 = n1084 & ~n1107;
  assign n1110 = n1109 ^ n1108;
  assign n956 = ~x22 & ~n32;
  assign n957 = x6 & ~x22;
  assign n958 = ~n956 & ~n957;
  assign n959 = n958 ^ x7;
  assign n1106 = ~n551 & ~n959;
  assign n1111 = n1110 ^ n1106;
  assign n1008 = n700 ^ n243;
  assign n1009 = n1008 ^ n268;
  assign n1010 = n1009 ^ n450;
  assign n1013 = ~n76 & n154;
  assign n1014 = n1013 ^ n817;
  assign n1015 = n1014 ^ n186;
  assign n1011 = n322 ^ n277;
  assign n1012 = n1011 ^ n194;
  assign n1016 = n1015 ^ n1012;
  assign n1017 = ~n1010 & ~n1016;
  assign n1019 = n437 ^ n236;
  assign n1018 = n460 ^ n341;
  assign n1020 = n1019 ^ n1018;
  assign n1021 = n1017 & n1020;
  assign n1022 = n183 & n1021;
  assign n1023 = n436 ^ n378;
  assign n1024 = n1023 ^ n384;
  assign n1025 = ~n1022 & n1024;
  assign n1026 = n165 ^ n133;
  assign n1027 = n60 & ~n1026;
  assign n1028 = ~n73 & ~n1027;
  assign n971 = n840 ^ n400;
  assign n972 = n971 ^ n575;
  assign n973 = ~n204 & ~n972;
  assign n1029 = ~n727 & n973;
  assign n229 = ~n183 & n226;
  assign n1031 = n617 ^ n216;
  assign n1030 = n348 ^ n250;
  assign n1032 = n1031 ^ n1030;
  assign n1033 = ~n229 & ~n1032;
  assign n1035 = n359 ^ n177;
  assign n1034 = n623 ^ n480;
  assign n1036 = n1035 ^ n1034;
  assign n1037 = n353 ^ n277;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = n1033 & n1038;
  assign n1040 = n1029 & n1039;
  assign n1041 = ~n1028 & n1040;
  assign n1042 = ~n1025 & n1041;
  assign n1043 = n574 ^ n267;
  assign n1044 = n1043 ^ n416;
  assign n519 = n72 & n119;
  assign n1046 = n519 ^ n298;
  assign n1045 = n574 ^ n325;
  assign n1047 = n1046 ^ n1045;
  assign n1048 = ~n1044 & ~n1047;
  assign n1050 = n237 ^ n174;
  assign n1049 = n673 ^ n492;
  assign n1051 = n1050 ^ n1049;
  assign n1052 = n1048 & n1051;
  assign n228 = n227 ^ n223;
  assign n502 = n258 ^ n151;
  assign n503 = ~n203 & n502;
  assign n504 = n503 ^ n419;
  assign n505 = ~n228 & ~n504;
  assign n506 = n402 ^ n287;
  assign n507 = n506 ^ n185;
  assign n508 = n505 & ~n507;
  assign n1053 = n427 ^ n251;
  assign n1054 = ~n249 & n1053;
  assign n1055 = ~n709 & n1054;
  assign n1056 = n508 & n1055;
  assign n1057 = n1052 & n1056;
  assign n1058 = n169 ^ n100;
  assign n1059 = n1058 ^ n154;
  assign n1060 = n290 ^ n61;
  assign n1061 = n1059 & ~n1060;
  assign n1062 = ~n275 & ~n1061;
  assign n362 = ~n60 & n133;
  assign n1063 = n362 ^ n212;
  assign n1064 = n1063 ^ n319;
  assign n414 = n159 & ~n203;
  assign n1065 = n693 ^ n414;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = n1062 & n1066;
  assign n509 = n72 & n118;
  assign n511 = n510 ^ n509;
  assign n1068 = n536 ^ n511;
  assign n1069 = n484 ^ n428;
  assign n1070 = n1069 ^ n268;
  assign n1071 = ~n1068 & ~n1070;
  assign n1072 = n1067 & n1071;
  assign n1073 = n1057 & n1072;
  assign n1074 = n1042 & n1073;
  assign n961 = n428 ^ n196;
  assign n962 = n871 ^ n657;
  assign n963 = ~n961 & ~n962;
  assign n964 = n450 ^ n424;
  assign n965 = n964 ^ n275;
  assign n966 = n403 ^ n236;
  assign n967 = n966 ^ n740;
  assign n968 = n967 ^ n246;
  assign n969 = ~n965 & ~n968;
  assign n970 = n963 & n969;
  assign n974 = n533 ^ n318;
  assign n975 = n973 & ~n974;
  assign n976 = n737 ^ n667;
  assign n977 = n976 ^ n287;
  assign n978 = n977 ^ n347;
  assign n979 = n978 ^ n427;
  assign n980 = n975 & n979;
  assign n981 = n970 & n980;
  assign n982 = n676 ^ n454;
  assign n983 = n353 ^ n115;
  assign n984 = n983 ^ n423;
  assign n985 = ~n982 & n984;
  assign n986 = n616 & n985;
  assign n987 = n383 ^ n281;
  assign n988 = n987 ^ n170;
  assign n989 = n986 & ~n988;
  assign n991 = n395 ^ n363;
  assign n990 = n248 ^ n229;
  assign n992 = n991 ^ n990;
  assign n995 = n361 ^ n329;
  assign n993 = n373 ^ n352;
  assign n994 = n993 ^ n683;
  assign n996 = n995 ^ n994;
  assign n997 = ~n992 & n996;
  assign n1001 = ~n76 & n571;
  assign n1002 = n1001 ^ n846;
  assign n1003 = n1002 ^ n362;
  assign n998 = ~n203 & n261;
  assign n999 = n998 ^ n355;
  assign n1000 = n999 ^ n336;
  assign n1004 = n1003 ^ n1000;
  assign n1005 = n997 & ~n1004;
  assign n1006 = n989 & n1005;
  assign n1007 = n981 & n1006;
  assign n1112 = n1074 ^ n1007;
  assign n1113 = n1007 ^ n891;
  assign n1114 = n1007 ^ n583;
  assign n1115 = n1113 & n1114;
  assign n1116 = n1115 ^ n1007;
  assign n1117 = ~n1112 & ~n1116;
  assign n1118 = n1117 ^ n891;
  assign n1119 = n1118 ^ n1110;
  assign n1120 = ~n1111 & n1119;
  assign n1121 = n1120 ^ n1106;
  assign n954 = ~x22 & ~n34;
  assign n955 = n954 ^ x8;
  assign n960 = n959 ^ n955;
  assign n1104 = ~n551 & ~n960;
  assign n1075 = ~n1007 & ~n1074;
  assign n1076 = ~n891 & ~n1075;
  assign n1105 = n1104 ^ n1076;
  assign n1122 = n1121 ^ n1105;
  assign n1221 = ~n551 & ~n955;
  assign n1222 = n580 & ~n1221;
  assign n1223 = n922 ^ n794;
  assign n1224 = n1223 ^ n955;
  assign n1225 = n570 & n1224;
  assign n1226 = n1225 ^ n955;
  assign n1227 = ~n1222 & n1226;
  assign n1123 = ~n147 & ~n592;
  assign n1124 = n165 ^ n100;
  assign n1125 = ~n112 & n1124;
  assign n1126 = n1125 ^ n169;
  assign n1127 = ~n1123 & n1126;
  assign n1128 = ~n484 & ~n1127;
  assign n1129 = n602 ^ n203;
  assign n1130 = n154 & ~n1129;
  assign n1132 = n310 ^ n109;
  assign n1131 = n575 ^ n519;
  assign n1133 = n1132 ^ n1131;
  assign n1134 = ~n348 & n1133;
  assign n1135 = ~n1130 & n1134;
  assign n1136 = n453 ^ n424;
  assign n1137 = n1136 ^ n489;
  assign n1138 = ~n194 & ~n1137;
  assign n1139 = n725 & n1138;
  assign n1140 = n1054 & n1139;
  assign n1141 = n1135 & n1140;
  assign n1142 = n1128 & n1141;
  assign n417 = n416 ^ n414;
  assign n421 = n420 ^ n417;
  assign n422 = ~n413 & ~n421;
  assign n1143 = n422 & ~n691;
  assign n1144 = n963 & n1143;
  assign n1145 = n533 ^ n322;
  assign n1146 = ~n990 & ~n1145;
  assign n1147 = n450 ^ n338;
  assign n1148 = n1147 ^ n290;
  assign n1149 = n1148 ^ n186;
  assign n1150 = n1146 & ~n1149;
  assign n1151 = n1144 & n1150;
  assign n494 = n493 ^ n381;
  assign n495 = n491 & n494;
  assign n496 = n479 ^ n137;
  assign n497 = n56 & n496;
  assign n499 = n498 ^ n281;
  assign n500 = ~n497 & ~n499;
  assign n501 = n495 & n500;
  assign n1153 = n151 ^ n133;
  assign n1154 = n1153 ^ n259;
  assign n1155 = ~n61 & n1154;
  assign n1156 = n1155 ^ n289;
  assign n1152 = n618 ^ n212;
  assign n1157 = n1156 ^ n1152;
  assign n1158 = ~n511 & ~n1157;
  assign n1159 = n501 & n1158;
  assign n1160 = n1151 & n1159;
  assign n1161 = n1142 & n1160;
  assign n1162 = n1074 & n1161;
  assign n1163 = n956 ^ x6;
  assign n1164 = ~n551 & n1163;
  assign n1165 = ~n1162 & ~n1164;
  assign n1166 = n433 ^ n166;
  assign n1167 = ~n658 & ~n1064;
  assign n1168 = ~n1166 & n1167;
  assign n1169 = n666 ^ n228;
  assign n1170 = n1169 ^ n287;
  assign n1172 = n374 ^ n329;
  assign n321 = n72 & ~n183;
  assign n1171 = n342 ^ n321;
  assign n1173 = n1172 ^ n1171;
  assign n1174 = ~n1170 & n1173;
  assign n1175 = n1168 & n1174;
  assign n1176 = n424 ^ n285;
  assign n1177 = n1176 ^ n289;
  assign n1179 = n428 ^ n273;
  assign n1180 = n1179 ^ n533;
  assign n1178 = n510 ^ n490;
  assign n1181 = n1180 ^ n1178;
  assign n1182 = ~n1177 & ~n1181;
  assign n1183 = n1175 & n1182;
  assign n1184 = n1128 & n1183;
  assign n1185 = ~n183 & n642;
  assign n1186 = n1185 ^ n817;
  assign n366 = n365 ^ n109;
  assign n1187 = n1186 ^ n366;
  assign n1188 = ~n674 & ~n1187;
  assign n1189 = ~n1043 & n1188;
  assign n1190 = n1058 ^ n647;
  assign n1191 = n61 & ~n1190;
  assign n1192 = n334 & ~n1058;
  assign n1193 = n74 & ~n1192;
  assign n1194 = ~n1191 & n1193;
  assign n1196 = n359 ^ n195;
  assign n1197 = n1196 ^ n427;
  assign n1195 = n536 ^ n509;
  assign n1198 = n1197 ^ n1195;
  assign n1199 = ~n991 & n1198;
  assign n1200 = ~n1194 & n1199;
  assign n1201 = n1189 & n1200;
  assign n390 = n137 ^ n128;
  assign n1202 = n390 ^ n311;
  assign n1203 = ~n850 & ~n1202;
  assign n1204 = n1201 & ~n1203;
  assign n462 = n461 ^ n460;
  assign n459 = n302 ^ n115;
  assign n463 = n462 ^ n459;
  assign n465 = n464 ^ n463;
  assign n1205 = ~n59 & ~n1192;
  assign n1206 = n1205 ^ n617;
  assign n1207 = n623 ^ n560;
  assign n1208 = n1207 ^ n414;
  assign n1209 = n1208 ^ n454;
  assign n1210 = ~n1206 & ~n1209;
  assign n1211 = n465 & n1210;
  assign n1212 = n1204 & n1211;
  assign n1213 = n1184 & n1212;
  assign n1218 = ~n1074 & n1213;
  assign n1215 = ~n1161 & ~n1213;
  assign n1214 = n1213 ^ n1161;
  assign n1216 = n1215 ^ n1214;
  assign n1217 = ~n1074 & ~n1216;
  assign n1219 = n1218 ^ n1217;
  assign n1220 = ~n1165 & ~n1219;
  assign n1228 = n1227 ^ n1220;
  assign n1094 = n753 ^ n579;
  assign n1231 = n758 & ~n1094;
  assign n1229 = n792 ^ n579;
  assign n1230 = n910 & ~n1229;
  assign n1232 = n1231 ^ n1230;
  assign n1233 = n1232 ^ n1220;
  assign n1234 = ~n1228 & n1233;
  assign n1235 = n1234 ^ n1232;
  assign n1236 = n1235 ^ n1121;
  assign n1237 = ~n1122 & ~n1236;
  assign n1238 = n1237 ^ n1235;
  assign n1102 = n934 ^ n928;
  assign n1089 = n570 & n795;
  assign n1090 = n1089 ^ n794;
  assign n1091 = ~n580 & n1090;
  assign n1092 = ~n922 & ~n1091;
  assign n1085 = n1082 & n1084;
  assign n1086 = n748 ^ n583;
  assign n1087 = n893 & n1086;
  assign n1088 = ~n1085 & ~n1087;
  assign n1093 = n1092 ^ n1088;
  assign n1096 = n758 & ~n924;
  assign n1095 = n910 & ~n1094;
  assign n1097 = n1096 ^ n1095;
  assign n1098 = n1097 ^ n1088;
  assign n1099 = ~n1093 & ~n1098;
  assign n1100 = n1099 ^ n1097;
  assign n1077 = n1076 ^ n959;
  assign n1078 = ~n960 & n1077;
  assign n1079 = n1078 ^ n959;
  assign n1080 = ~n551 & ~n1079;
  assign n947 = n551 & n580;
  assign n948 = n551 & n570;
  assign n949 = ~n753 & n948;
  assign n950 = ~n947 & ~n949;
  assign n951 = n792 & ~n915;
  assign n952 = n951 ^ n570;
  assign n953 = n950 & n952;
  assign n1081 = n1080 ^ n953;
  assign n1101 = n1100 ^ n1081;
  assign n1103 = n1102 ^ n1101;
  assign n1239 = n1238 ^ n1103;
  assign n1240 = n1235 ^ n1122;
  assign n1269 = n893 & ~n1107;
  assign n1267 = n753 ^ n748;
  assign n1268 = n1084 & ~n1267;
  assign n1270 = n1269 ^ n1268;
  assign n1273 = n1270 ^ n1164;
  assign n1282 = ~x22 & ~n31;
  assign n1283 = n1282 ^ x5;
  assign n1285 = n551 & ~n1283;
  assign n1284 = n1283 ^ n551;
  assign n1286 = n1285 ^ n1284;
  assign n1276 = n1219 ^ n1162;
  assign n1274 = n1161 ^ n1074;
  assign n1275 = n1274 ^ n1215;
  assign n1277 = n1276 ^ n1275;
  assign n1278 = n1277 ^ n1216;
  assign n1279 = ~n583 & n1278;
  assign n1287 = ~n1276 & ~n1279;
  assign n1288 = n1286 & n1287;
  assign n1280 = ~n1161 & n1279;
  assign n1281 = n1280 ^ n1219;
  assign n1289 = n1288 ^ n1281;
  assign n1290 = n1289 ^ n1219;
  assign n1291 = n1290 ^ n1270;
  assign n1292 = ~n1273 & n1291;
  assign n1272 = n1220 ^ n1165;
  assign n1293 = n1292 ^ n1272;
  assign n1271 = ~n1162 & n1270;
  assign n1294 = n1293 ^ n1271;
  assign n1252 = n891 ^ n555;
  assign n1253 = n1074 ^ n891;
  assign n1254 = n1252 & n1253;
  assign n1251 = n891 ^ n583;
  assign n1255 = n1254 ^ n1251;
  assign n1256 = ~n1112 & n1255;
  assign n1257 = n1256 ^ n1251;
  assign n1248 = n959 ^ n551;
  assign n1245 = n570 & ~n955;
  assign n1246 = n1245 ^ n959;
  assign n1247 = ~n917 & n1246;
  assign n1249 = n1248 ^ n1247;
  assign n1250 = ~n947 & n1249;
  assign n1258 = n1257 ^ n1250;
  assign n1261 = n758 & ~n1229;
  assign n1259 = n794 ^ n579;
  assign n1260 = n910 & ~n1259;
  assign n1262 = n1261 ^ n1260;
  assign n1263 = n1262 ^ n1257;
  assign n1264 = ~n1258 & n1263;
  assign n1265 = n1264 ^ n1262;
  assign n1242 = n1118 ^ n1106;
  assign n1243 = n1242 ^ n1110;
  assign n1241 = n1232 ^ n1228;
  assign n1244 = n1243 ^ n1241;
  assign n1266 = n1265 ^ n1244;
  assign n1295 = n1294 ^ n1266;
  assign n1304 = n1112 & n1252;
  assign n1301 = ~n1112 & n1253;
  assign n1302 = n891 ^ n751;
  assign n1303 = n1301 & ~n1302;
  assign n1305 = n1304 ^ n1303;
  assign n1299 = n893 & ~n1267;
  assign n1297 = n792 ^ n748;
  assign n1298 = n1084 & ~n1297;
  assign n1300 = n1299 ^ n1298;
  assign n1306 = n1305 ^ n1300;
  assign n1309 = n758 & ~n1259;
  assign n1307 = n955 ^ n579;
  assign n1308 = n910 & ~n1307;
  assign n1310 = n1309 ^ n1308;
  assign n1311 = n1310 ^ n1300;
  assign n1312 = ~n1306 & n1311;
  assign n1313 = n1312 ^ n1310;
  assign n1296 = n1262 ^ n1258;
  assign n1314 = n1313 ^ n1296;
  assign n1325 = n1112 & ~n1302;
  assign n1323 = n891 ^ n753;
  assign n1324 = n1301 & ~n1323;
  assign n1326 = n1325 ^ n1324;
  assign n1321 = n893 & ~n1297;
  assign n1319 = n794 ^ n748;
  assign n1320 = n1084 & ~n1319;
  assign n1322 = n1321 ^ n1320;
  assign n1327 = n1326 ^ n1322;
  assign n1330 = n758 & ~n1307;
  assign n1328 = n959 ^ n579;
  assign n1329 = n910 & n1328;
  assign n1331 = n1330 ^ n1329;
  assign n1332 = n1331 ^ n1322;
  assign n1333 = ~n1327 & n1332;
  assign n1334 = n1333 ^ n1331;
  assign n1315 = n915 & ~n959;
  assign n1316 = n917 & n1163;
  assign n1317 = n1316 ^ n551;
  assign n1318 = ~n1315 & n1317;
  assign n1335 = n1334 ^ n1318;
  assign n1340 = ~n555 & n1278;
  assign n1344 = n1274 ^ n583;
  assign n1341 = n1218 ^ n1074;
  assign n1342 = n1341 ^ n583;
  assign n1343 = ~n1214 & n1342;
  assign n1345 = n1344 ^ n1343;
  assign n1346 = ~n1340 & ~n1345;
  assign n1336 = ~x22 & ~n30;
  assign n1337 = n1336 ^ x4;
  assign n1338 = ~n551 & ~n1337;
  assign n1339 = n1338 ^ n551;
  assign n1347 = n1346 ^ n1339;
  assign n1348 = n1339 ^ n1161;
  assign n1349 = ~n1213 & n1348;
  assign n1350 = n1349 ^ n1161;
  assign n1351 = n1347 & ~n1350;
  assign n1352 = ~n555 & ~n1277;
  assign n1353 = n1339 & ~n1352;
  assign n1354 = n555 & n1218;
  assign n1355 = n1161 & ~n1354;
  assign n1356 = ~n1353 & ~n1355;
  assign n1357 = ~n1351 & ~n1356;
  assign n1358 = n1357 ^ n1318;
  assign n1359 = ~n1335 & ~n1358;
  assign n1360 = n1359 ^ n1334;
  assign n1361 = n1360 ^ n1313;
  assign n1362 = ~n1314 & n1361;
  assign n1363 = n1362 ^ n1360;
  assign n1364 = n1363 ^ n1294;
  assign n1365 = n1295 & ~n1364;
  assign n1366 = n1365 ^ n1363;
  assign n1367 = n1366 ^ n1240;
  assign n1368 = ~n1240 & ~n1367;
  assign n1369 = n1368 ^ n1367;
  assign n1370 = n1239 & n1369;
  assign n1373 = n1287 ^ n1286;
  assign n1372 = n1310 ^ n1306;
  assign n1374 = n1373 ^ n1372;
  assign n1385 = x22 ^ x2;
  assign n1386 = x1 & ~x2;
  assign n1387 = n1386 ^ n25;
  assign n1388 = n1385 & ~n1387;
  assign n1391 = n1388 ^ x22;
  assign n1389 = n28 & n1388;
  assign n1390 = n1389 ^ n29;
  assign n1392 = n1391 ^ n1390;
  assign n1393 = n1392 ^ x3;
  assign n1394 = ~n551 & ~n1393;
  assign n1379 = n1277 ^ n1217;
  assign n1380 = n1074 ^ n751;
  assign n1381 = ~n1379 & ~n1380;
  assign n1382 = n1074 ^ n555;
  assign n1383 = n1214 & n1382;
  assign n1384 = ~n1381 & ~n1383;
  assign n1395 = n1394 ^ n1384;
  assign n323 = n322 ^ n321;
  assign n324 = ~n320 & ~n323;
  assign n330 = n329 ^ n325;
  assign n331 = n330 ^ n273;
  assign n332 = n324 & n331;
  assign n354 = n353 ^ n196;
  assign n356 = n355 ^ n354;
  assign n357 = ~n350 & ~n356;
  assign n358 = n332 & n357;
  assign n364 = n363 ^ n362;
  assign n367 = n366 ^ n364;
  assign n368 = ~n361 & ~n367;
  assign n369 = n358 & n368;
  assign n1396 = n369 & ~n536;
  assign n394 = n267 ^ n186;
  assign n1399 = n394 ^ n223;
  assign n1397 = n290 ^ n285;
  assign n1398 = n1397 ^ n1178;
  assign n1400 = n1399 ^ n1398;
  assign n1401 = n718 & ~n1400;
  assign n1402 = n119 & n809;
  assign n1403 = n1402 ^ n676;
  assign n1404 = ~n623 & ~n1403;
  assign n1406 = n336 ^ n73;
  assign n1405 = n72 & n850;
  assign n1407 = n1406 ^ n1405;
  assign n1408 = n1407 ^ n61;
  assign n1409 = n1404 & ~n1408;
  assign n1410 = n1401 & n1409;
  assign n1411 = n137 ^ n83;
  assign n1412 = ~n43 & n1411;
  assign n1413 = ~n117 & ~n1412;
  assign n1414 = ~n58 & n1411;
  assign n1415 = n1414 ^ n100;
  assign n1416 = ~n1413 & n1415;
  assign n1417 = n693 ^ n84;
  assign n1418 = n1417 ^ n467;
  assign n1419 = ~n1416 & ~n1418;
  assign n1420 = n181 & n1419;
  assign n1421 = n1410 & n1420;
  assign n1422 = n1396 & n1421;
  assign n1423 = ~n583 & n1422;
  assign n1424 = ~n1161 & ~n1423;
  assign n1425 = n1424 ^ n1384;
  assign n1426 = ~n1395 & n1425;
  assign n1427 = n1426 ^ n1394;
  assign n1375 = n915 & n1163;
  assign n1376 = n917 & n1283;
  assign n1377 = n1376 ^ n551;
  assign n1378 = ~n1375 & n1377;
  assign n1428 = n1427 ^ n1378;
  assign n1435 = n1112 & ~n1323;
  assign n1433 = n891 ^ n792;
  assign n1434 = n1301 & ~n1433;
  assign n1436 = n1435 ^ n1434;
  assign n1431 = n893 & ~n1319;
  assign n1429 = n955 ^ n748;
  assign n1430 = n1084 & ~n1429;
  assign n1432 = n1431 ^ n1430;
  assign n1437 = n1436 ^ n1432;
  assign n1440 = n758 & n1328;
  assign n1438 = n1163 ^ n579;
  assign n1439 = n910 & ~n1438;
  assign n1441 = n1440 ^ n1439;
  assign n1442 = n1441 ^ n1432;
  assign n1443 = ~n1437 & n1442;
  assign n1444 = n1443 ^ n1441;
  assign n1445 = n1444 ^ n1378;
  assign n1446 = ~n1428 & n1445;
  assign n1447 = n1446 ^ n1427;
  assign n1448 = n1447 ^ n1372;
  assign n1449 = ~n1374 & n1448;
  assign n1450 = n1449 ^ n1447;
  assign n1371 = n1363 ^ n1295;
  assign n1451 = n1450 ^ n1371;
  assign n1452 = n1290 ^ n1162;
  assign n1453 = n1452 ^ n1273;
  assign n1454 = n1453 ^ n1450;
  assign n1456 = n1357 ^ n1335;
  assign n1455 = n1447 ^ n1374;
  assign n1457 = n1456 ^ n1455;
  assign n1458 = n1331 ^ n1327;
  assign n1459 = n1458 ^ n1347;
  assign n1466 = n580 & ~n1338;
  assign n1467 = n1337 ^ n1285;
  assign n1468 = n570 & ~n1467;
  assign n1469 = n1468 ^ n1337;
  assign n1470 = ~n1466 & n1469;
  assign n1461 = n1161 ^ n583;
  assign n1460 = n555 & ~n1161;
  assign n1462 = n1461 ^ n1460;
  assign n1463 = n1422 & n1462;
  assign n1464 = n1463 ^ n1461;
  assign n1465 = ~n551 & n1464;
  assign n1471 = n1470 ^ n1465;
  assign n1478 = n1112 & ~n1433;
  assign n1476 = n891 ^ n794;
  assign n1477 = n1301 & ~n1476;
  assign n1479 = n1478 ^ n1477;
  assign n1474 = n893 & ~n1429;
  assign n1472 = n959 ^ n748;
  assign n1473 = n1084 & n1472;
  assign n1475 = n1474 ^ n1473;
  assign n1480 = n1479 ^ n1475;
  assign n1483 = n758 & ~n1438;
  assign n1481 = n1283 ^ n579;
  assign n1482 = n910 & ~n1481;
  assign n1484 = n1483 ^ n1482;
  assign n1485 = n1484 ^ n1475;
  assign n1486 = ~n1480 & n1485;
  assign n1487 = n1486 ^ n1484;
  assign n1488 = n1487 ^ n1465;
  assign n1489 = ~n1471 & n1488;
  assign n1490 = n1489 ^ n1487;
  assign n1491 = n1490 ^ n1458;
  assign n1492 = n1459 & n1491;
  assign n1493 = n1492 ^ n1490;
  assign n1494 = n1493 ^ n1455;
  assign n1495 = ~n1457 & n1494;
  assign n1496 = n1495 ^ n1493;
  assign n1497 = n1496 ^ n1450;
  assign n1498 = n1454 & n1497;
  assign n1499 = n1498 ^ n1454;
  assign n1500 = ~n1451 & n1499;
  assign n1501 = n1500 ^ n1371;
  assign n1502 = n1360 ^ n1314;
  assign n1504 = n1490 ^ n1459;
  assign n1503 = n1493 ^ n1457;
  assign n1505 = n1504 ^ n1503;
  assign n1506 = n1444 ^ n1428;
  assign n1507 = n1506 ^ n1504;
  assign n1527 = n1441 ^ n1437;
  assign n1513 = n1393 ^ n551;
  assign n1512 = n570 & n1337;
  assign n1514 = n1513 ^ n1512;
  assign n1515 = ~n917 & n1514;
  assign n1516 = n1515 ^ n1513;
  assign n1517 = ~n947 & n1516;
  assign n1511 = n1464 ^ n551;
  assign n1518 = n1517 ^ n1511;
  assign n1521 = n1214 & ~n1380;
  assign n1519 = n1074 ^ n753;
  assign n1520 = ~n1379 & ~n1519;
  assign n1522 = n1521 ^ n1520;
  assign n1523 = n1522 ^ n1511;
  assign n1524 = n1518 & ~n1523;
  assign n1525 = n1524 ^ n1522;
  assign n1509 = n1424 ^ n1394;
  assign n1510 = n1509 ^ n1384;
  assign n1526 = n1525 ^ n1510;
  assign n1528 = n1527 ^ n1526;
  assign n1508 = n1487 ^ n1471;
  assign n1529 = n1528 ^ n1508;
  assign n1537 = n1112 & ~n1476;
  assign n1535 = n955 ^ n891;
  assign n1536 = n1301 & ~n1535;
  assign n1538 = n1537 ^ n1536;
  assign n1533 = n893 & n1472;
  assign n1531 = n1163 ^ n748;
  assign n1532 = n1084 & ~n1531;
  assign n1534 = n1533 ^ n1532;
  assign n1539 = n1538 ^ n1534;
  assign n1540 = n758 & ~n1393;
  assign n1541 = n750 & ~n1540;
  assign n1543 = n1161 ^ n751;
  assign n1542 = ~n753 & ~n1161;
  assign n1544 = n1543 ^ n1542;
  assign n1545 = n1422 & ~n1544;
  assign n1546 = n1545 ^ n1543;
  assign n1547 = n1541 & ~n1546;
  assign n1548 = n1547 ^ n1538;
  assign n1549 = n1539 & ~n1548;
  assign n1550 = n1549 ^ n1534;
  assign n1530 = n1484 ^ n1480;
  assign n1551 = n1550 ^ n1530;
  assign n1559 = n1214 & ~n1519;
  assign n1557 = n1074 ^ n792;
  assign n1558 = ~n1379 & ~n1557;
  assign n1560 = n1559 ^ n1558;
  assign n1553 = n1161 ^ n555;
  assign n1552 = ~n751 & ~n1161;
  assign n1554 = n1553 ^ n1552;
  assign n1555 = n1422 & n1554;
  assign n1556 = n1555 ^ n1553;
  assign n1561 = n1560 ^ n1556;
  assign n1564 = n758 & ~n1481;
  assign n1562 = n1337 ^ n579;
  assign n1563 = n910 & ~n1562;
  assign n1565 = n1564 ^ n1563;
  assign n1566 = n1565 ^ n1560;
  assign n1567 = ~n1561 & n1566;
  assign n1568 = n1567 ^ n1565;
  assign n1569 = n1568 ^ n1530;
  assign n1570 = n1551 & ~n1569;
  assign n1571 = n1570 ^ n1550;
  assign n1572 = n1571 ^ n1508;
  assign n1573 = n1529 & n1572;
  assign n1574 = n1573 ^ n1571;
  assign n1575 = n1574 ^ n1504;
  assign n1576 = ~n1507 & n1575;
  assign n1577 = ~n1505 & n1576;
  assign n1578 = n1577 ^ n1503;
  assign n1590 = n1163 ^ n891;
  assign n1618 = n1112 & ~n1590;
  assign n1616 = n1283 ^ n891;
  assign n1617 = n1301 & ~n1616;
  assign n1619 = n1618 ^ n1617;
  assign n1584 = n1074 ^ n955;
  assign n1614 = n1214 & ~n1584;
  assign n1612 = n1074 ^ n959;
  assign n1613 = ~n1379 & n1612;
  assign n1615 = n1614 ^ n1613;
  assign n1620 = n1619 ^ n1615;
  assign n1622 = n1084 & ~n1393;
  assign n1605 = n1337 ^ n748;
  assign n1621 = n893 & ~n1605;
  assign n1623 = n1622 ^ n1621;
  assign n1624 = n1623 ^ n1083;
  assign n1625 = n1624 ^ n1615;
  assign n1626 = n1620 & ~n1625;
  assign n1627 = n1626 ^ n1619;
  assign n1607 = n1283 ^ n748;
  assign n1608 = n893 & ~n1607;
  assign n1606 = n1084 & ~n1605;
  assign n1609 = n1608 ^ n1606;
  assign n1610 = n1609 ^ n1540;
  assign n1596 = n897 & n1393;
  assign n1597 = ~n1083 & ~n1596;
  assign n1599 = n1161 ^ n792;
  assign n1598 = ~n794 & ~n1161;
  assign n1600 = n1599 ^ n1598;
  assign n1601 = n1422 & ~n1600;
  assign n1602 = n1601 ^ n1599;
  assign n1603 = ~n1597 & ~n1602;
  assign n1592 = n959 ^ n891;
  assign n1593 = n1112 & n1592;
  assign n1591 = n1301 & ~n1590;
  assign n1594 = n1593 ^ n1591;
  assign n1586 = n1074 ^ n794;
  assign n1587 = n1214 & ~n1586;
  assign n1585 = ~n1379 & ~n1584;
  assign n1588 = n1587 ^ n1585;
  assign n1580 = n1161 ^ n753;
  assign n1579 = ~n792 & ~n1161;
  assign n1581 = n1580 ^ n1579;
  assign n1582 = n1422 & ~n1581;
  assign n1583 = n1582 ^ n1580;
  assign n1589 = n1588 ^ n1583;
  assign n1595 = n1594 ^ n1589;
  assign n1604 = n1603 ^ n1595;
  assign n1611 = n1610 ^ n1604;
  assign n1628 = n1627 ^ n1611;
  assign n1635 = n1214 & n1612;
  assign n1633 = n1163 ^ n1074;
  assign n1634 = ~n1379 & ~n1633;
  assign n1636 = n1635 ^ n1634;
  assign n1631 = n1112 & ~n1616;
  assign n1629 = n1337 ^ n891;
  assign n1630 = n1301 & ~n1629;
  assign n1632 = n1631 ^ n1630;
  assign n1637 = n1636 ^ n1632;
  assign n1639 = n1161 ^ n794;
  assign n1638 = ~n955 & ~n1161;
  assign n1640 = n1639 ^ n1638;
  assign n1641 = n1422 & ~n1640;
  assign n1642 = n1641 ^ n1639;
  assign n1643 = n1642 ^ n1632;
  assign n1644 = n1637 & n1643;
  assign n1645 = n1644 ^ n1636;
  assign n1653 = n1214 & ~n1633;
  assign n1651 = n1283 ^ n1074;
  assign n1652 = ~n1379 & ~n1651;
  assign n1654 = n1653 ^ n1652;
  assign n1647 = n1161 ^ n955;
  assign n1646 = n959 & ~n1161;
  assign n1648 = n1647 ^ n1646;
  assign n1649 = n1422 & ~n1648;
  assign n1650 = n1649 ^ n1647;
  assign n1655 = n1654 ^ n1650;
  assign n1657 = n1393 ^ n1075;
  assign n1658 = n1301 & n1657;
  assign n1656 = n1112 & ~n1629;
  assign n1659 = n1658 ^ n1656;
  assign n1660 = n1112 & ~n1393;
  assign n1661 = n1076 & ~n1660;
  assign n1662 = ~n1659 & ~n1661;
  assign n1663 = n1662 ^ n1650;
  assign n1664 = ~n1655 & ~n1663;
  assign n1665 = n1664 ^ n1654;
  assign n1666 = n893 & ~n1393;
  assign n1667 = n1661 ^ n1659;
  assign n1668 = n1667 ^ n1662;
  assign n1670 = n1666 ^ n1665;
  assign n1669 = ~n1650 & n1654;
  assign n1671 = n1670 ^ n1669;
  assign n1672 = n1668 & ~n1671;
  assign n1673 = n1672 ^ n1669;
  assign n1674 = ~n1666 & ~n1673;
  assign n1675 = n1665 & ~n1674;
  assign n1677 = n1645 & n1675;
  assign n1676 = n1675 ^ n1645;
  assign n1678 = n1677 ^ n1676;
  assign n1679 = ~n1628 & n1678;
  assign n1680 = n1642 ^ n1637;
  assign n1681 = n1680 ^ n1673;
  assign n1689 = n1214 & ~n1651;
  assign n1687 = n1337 ^ n1074;
  assign n1688 = ~n1379 & ~n1687;
  assign n1690 = n1689 ^ n1688;
  assign n1683 = n1161 ^ n959;
  assign n1682 = ~n1161 & ~n1163;
  assign n1684 = n1683 ^ n1682;
  assign n1685 = n1422 & n1684;
  assign n1686 = n1685 ^ n1683;
  assign n1691 = n1690 ^ n1686;
  assign n1692 = n1393 ^ n1213;
  assign n1693 = n1214 & n1692;
  assign n1694 = n1693 ^ n1213;
  assign n1695 = ~n1074 & n1694;
  assign n1696 = ~n1660 & ~n1695;
  assign n1697 = n1691 & ~n1696;
  assign n1701 = n1163 ^ n1161;
  assign n1698 = ~n1161 & n1283;
  assign n1699 = n1698 ^ n1163;
  assign n1700 = n1422 & n1699;
  assign n1702 = n1701 ^ n1700;
  assign n1703 = ~n1697 & n1702;
  assign n1705 = ~n1379 & ~n1393;
  assign n1706 = n1705 ^ n1217;
  assign n1704 = n1214 & ~n1687;
  assign n1707 = n1706 ^ n1704;
  assign n1709 = n1691 & n1707;
  assign n1708 = n1707 ^ n1691;
  assign n1710 = n1709 ^ n1708;
  assign n1711 = ~n1695 & ~n1710;
  assign n1712 = ~n1703 & ~n1711;
  assign n1713 = ~n1660 & ~n1709;
  assign n1714 = n1712 & ~n1713;
  assign n1716 = n1283 & ~n1422;
  assign n1715 = ~n1213 & ~n1393;
  assign n1717 = n1716 ^ n1715;
  assign n1718 = n1422 ^ n1393;
  assign n1719 = n1422 ^ n1161;
  assign n1720 = ~n1422 & n1719;
  assign n1721 = n1720 ^ n1422;
  assign n1722 = n1718 & ~n1721;
  assign n1723 = n1722 ^ n1720;
  assign n1724 = n1723 ^ n1422;
  assign n1725 = n1724 ^ n1161;
  assign n1726 = n1337 & n1725;
  assign n1728 = n1726 ^ n1161;
  assign n1727 = n1716 & ~n1726;
  assign n1729 = n1728 ^ n1727;
  assign n1730 = ~n1717 & ~n1729;
  assign n1731 = ~n1714 & ~n1730;
  assign n1732 = n1710 & ~n1713;
  assign n1733 = n1702 & ~n1732;
  assign n1734 = n1667 ^ n1655;
  assign n1735 = n1734 ^ n1696;
  assign n1736 = n1734 ^ n1686;
  assign n1737 = n1734 ^ n1691;
  assign n1738 = n1734 & ~n1737;
  assign n1739 = n1738 ^ n1734;
  assign n1740 = ~n1736 & n1739;
  assign n1741 = n1740 ^ n1738;
  assign n1742 = n1741 ^ n1734;
  assign n1743 = n1742 ^ n1691;
  assign n1744 = n1735 & ~n1743;
  assign n1745 = n1744 ^ n1734;
  assign n1746 = ~n1733 & ~n1745;
  assign n1747 = ~n1731 & n1746;
  assign n1748 = n1747 ^ n1680;
  assign n1749 = n1748 ^ n1680;
  assign n1750 = n1695 & ~n1702;
  assign n1751 = n1750 ^ n1686;
  assign n1752 = n1691 & ~n1751;
  assign n1753 = n1752 ^ n1690;
  assign n1754 = ~n1734 & n1753;
  assign n1755 = n1754 ^ n1680;
  assign n1756 = n1755 ^ n1680;
  assign n1757 = ~n1749 & ~n1756;
  assign n1758 = n1757 ^ n1680;
  assign n1759 = n1681 & ~n1758;
  assign n1760 = n1759 ^ n1673;
  assign n1761 = ~n1679 & n1760;
  assign n1762 = n1628 & ~n1677;
  assign n1763 = n1602 ^ n1597;
  assign n1764 = n1624 ^ n1620;
  assign n1766 = n1763 & n1764;
  assign n1765 = n1764 ^ n1763;
  assign n1767 = n1766 ^ n1765;
  assign n1768 = ~n1762 & n1767;
  assign n1769 = ~n1761 & n1768;
  assign n1770 = n1766 ^ n1628;
  assign n1771 = n1760 ^ n1645;
  assign n1772 = n1676 & n1771;
  assign n1773 = n1772 ^ n1675;
  assign n1774 = n1773 ^ n1766;
  assign n1775 = ~n1770 & ~n1774;
  assign n1776 = n1775 ^ n1628;
  assign n1777 = ~n1769 & n1776;
  assign n1786 = n893 & ~n1531;
  assign n1785 = n1084 & ~n1607;
  assign n1787 = n1786 ^ n1785;
  assign n1782 = n1214 & ~n1557;
  assign n1781 = ~n1379 & ~n1586;
  assign n1783 = n1782 ^ n1781;
  assign n1779 = n1112 & ~n1535;
  assign n1778 = n1301 & n1592;
  assign n1780 = n1779 ^ n1778;
  assign n1784 = n1783 ^ n1780;
  assign n1788 = n1787 ^ n1784;
  assign n1789 = n1777 & ~n1788;
  assign n1808 = n1787 ^ n1780;
  assign n1809 = ~n1784 & n1808;
  assign n1810 = n1809 ^ n1787;
  assign n1806 = n915 & ~n1393;
  assign n1805 = n1547 ^ n1539;
  assign n1807 = n1806 ^ n1805;
  assign n1811 = n1810 ^ n1807;
  assign n1795 = n1393 ^ n579;
  assign n1796 = n910 & n1795;
  assign n1794 = n758 & ~n1562;
  assign n1797 = n1796 ^ n1794;
  assign n1793 = n1546 ^ n1541;
  assign n1798 = n1797 ^ n1793;
  assign n1790 = n1594 ^ n1583;
  assign n1791 = ~n1589 & n1790;
  assign n1792 = n1791 ^ n1588;
  assign n1801 = n1797 ^ n1792;
  assign n1802 = n1798 & n1801;
  assign n1803 = n1802 ^ n1792;
  assign n1800 = n1565 ^ n1561;
  assign n1804 = n1803 ^ n1800;
  assign n1812 = n1811 ^ n1804;
  assign n1799 = n1798 ^ n1792;
  assign n1813 = n1812 ^ n1799;
  assign n1814 = n1540 & n1609;
  assign n1817 = n1814 ^ n1610;
  assign n1818 = ~n1603 & ~n1817;
  assign n1815 = n1603 & n1814;
  assign n1816 = n1815 ^ n1610;
  assign n1819 = n1818 ^ n1816;
  assign n1820 = n1819 ^ n1603;
  assign n1823 = n1627 ^ n1595;
  assign n1821 = ~n1595 & n1627;
  assign n1824 = n1823 ^ n1821;
  assign n1827 = n1820 & n1824;
  assign n1828 = n1818 & ~n1821;
  assign n1829 = ~n1827 & ~n1828;
  assign n1822 = ~n1820 & n1821;
  assign n1825 = n1815 & ~n1824;
  assign n1826 = ~n1822 & ~n1825;
  assign n1830 = n1829 ^ n1826;
  assign n1831 = ~n1812 & n1830;
  assign n1832 = n1831 ^ n1829;
  assign n1833 = ~n1813 & n1832;
  assign n1834 = n1833 ^ n1799;
  assign n1835 = ~n1789 & ~n1834;
  assign n1836 = ~n1799 & n1829;
  assign n1837 = n1826 & ~n1836;
  assign n1838 = n1837 ^ n1812;
  assign n1839 = n1788 ^ n1777;
  assign n1840 = n1839 ^ n1789;
  assign n1841 = n1840 ^ n1837;
  assign n1842 = ~n1838 & n1841;
  assign n1843 = n1842 ^ n1812;
  assign n1844 = ~n1835 & ~n1843;
  assign n1845 = n1571 ^ n1529;
  assign n1846 = n1522 ^ n1518;
  assign n1847 = n1811 ^ n1800;
  assign n1848 = n1804 & ~n1847;
  assign n1849 = n1848 ^ n1803;
  assign n1851 = ~n1846 & n1849;
  assign n1850 = n1849 ^ n1846;
  assign n1852 = n1851 ^ n1850;
  assign n1853 = ~n1845 & ~n1852;
  assign n1854 = n1844 & ~n1853;
  assign n1855 = n1845 & ~n1851;
  assign n1856 = n1568 ^ n1551;
  assign n1857 = n1810 ^ n1806;
  assign n1858 = n1807 & ~n1857;
  assign n1859 = n1858 ^ n1805;
  assign n1861 = n1856 & n1859;
  assign n1860 = n1859 ^ n1856;
  assign n1862 = n1861 ^ n1860;
  assign n1863 = ~n1855 & n1862;
  assign n1864 = ~n1854 & n1863;
  assign n1865 = n1861 ^ n1845;
  assign n1866 = n1849 ^ n1844;
  assign n1867 = n1850 & n1866;
  assign n1868 = n1867 ^ n1850;
  assign n1869 = n1868 ^ n1844;
  assign n1870 = n1869 ^ n1845;
  assign n1871 = ~n1865 & n1870;
  assign n1872 = n1871 ^ n1845;
  assign n1873 = ~n1864 & n1872;
  assign n1874 = n1527 ^ n1510;
  assign n1875 = ~n1526 & n1874;
  assign n1876 = n1875 ^ n1525;
  assign n1878 = n1873 & ~n1876;
  assign n1877 = n1876 ^ n1873;
  assign n1879 = n1878 ^ n1877;
  assign n1880 = ~n1578 & ~n1879;
  assign n1881 = n1576 ^ n1507;
  assign n1882 = n1881 ^ n1574;
  assign n1883 = n1882 ^ n1878;
  assign n1884 = n1882 ^ n1503;
  assign n1885 = n1883 & ~n1884;
  assign n1886 = n1885 ^ n1882;
  assign n1887 = ~n1880 & ~n1886;
  assign n1889 = ~n1502 & ~n1887;
  assign n1888 = n1887 ^ n1502;
  assign n1890 = n1889 ^ n1888;
  assign n1891 = n1501 & n1890;
  assign n1892 = n1498 ^ n1496;
  assign n1893 = n1892 ^ n1889;
  assign n1894 = n1892 ^ n1371;
  assign n1895 = ~n1893 & ~n1894;
  assign n1896 = n1895 ^ n1892;
  assign n1897 = ~n1891 & n1896;
  assign n1898 = ~n1370 & n1897;
  assign n1899 = ~n1239 & ~n1368;
  assign n1900 = n1097 ^ n1093;
  assign n1901 = n1265 ^ n1243;
  assign n1902 = n1244 & ~n1901;
  assign n1903 = n1902 ^ n1241;
  assign n1905 = ~n1900 & ~n1903;
  assign n1904 = n1903 ^ n1900;
  assign n1906 = n1905 ^ n1904;
  assign n1907 = ~n1899 & n1906;
  assign n1908 = ~n1898 & n1907;
  assign n1909 = n1905 ^ n1239;
  assign n1910 = n1897 ^ n1366;
  assign n1911 = n1367 & ~n1910;
  assign n1912 = n1911 ^ n1240;
  assign n1913 = n1912 ^ n1239;
  assign n1914 = n1909 & n1913;
  assign n1915 = n1914 ^ n1905;
  assign n1916 = ~n1908 & ~n1915;
  assign n1917 = n1238 ^ n1101;
  assign n1918 = n1103 & n1917;
  assign n1919 = n1918 ^ n1238;
  assign n1920 = n937 ^ n921;
  assign n1921 = n1100 ^ n1080;
  assign n1922 = ~n1081 & n1921;
  assign n1923 = n1922 ^ n1100;
  assign n1924 = n1923 ^ n1920;
  assign n1925 = ~n551 & n795;
  assign n1926 = n1925 ^ n897;
  assign n1927 = n1926 ^ n1923;
  assign n1928 = n1924 & n1927;
  assign n1929 = n1928 ^ n1927;
  assign n1930 = n1920 & n1929;
  assign n1932 = ~n1919 & ~n1930;
  assign n1931 = n1930 ^ n1919;
  assign n1933 = n1932 ^ n1931;
  assign n1934 = ~n941 & n1933;
  assign n1940 = n1930 ^ n1929;
  assign n1941 = ~n1919 & n1940;
  assign n1942 = n1941 ^ n1933;
  assign n1937 = n1928 ^ n1920;
  assign n1938 = ~n1932 & n1937;
  assign n1935 = n1926 ^ n1924;
  assign n1936 = n1935 ^ n1919;
  assign n1939 = n1938 ^ n1936;
  assign n1943 = n1942 ^ n1939;
  assign n1944 = ~n1934 & ~n1943;
  assign n1945 = ~n1916 & ~n1944;
  assign n1946 = n941 & ~n1941;
  assign n1947 = ~n1938 & ~n1946;
  assign n1948 = ~n1945 & ~n1947;
  assign n1949 = n1948 ^ n945;
  assign n1950 = n946 & n1949;
  assign n1951 = n1950 ^ n1948;
  assign n2351 = n2350 ^ n1951;
  assign n2352 = n1961 & n2351;
  assign n458 = n133 & n457;
  assign n468 = n467 ^ n378;
  assign n469 = n468 ^ n424;
  assign n470 = n469 ^ n267;
  assign n471 = n395 ^ n177;
  assign n472 = n471 ^ n353;
  assign n473 = n472 ^ n400;
  assign n474 = ~n470 & ~n473;
  assign n475 = n465 & n474;
  assign n476 = ~n458 & n475;
  assign n477 = n452 & n476;
  assign n487 = n486 ^ n478;
  assign n488 = n477 & ~n487;
  assign n512 = n511 ^ n403;
  assign n513 = n508 & ~n512;
  assign n514 = n501 & n513;
  assign n516 = n515 ^ n83;
  assign n517 = ~n183 & n516;
  assign n518 = ~n274 & ~n517;
  assign n520 = n519 ^ n166;
  assign n521 = n518 & ~n520;
  assign n524 = n523 ^ n219;
  assign n526 = n525 ^ n524;
  assign n527 = n521 & n526;
  assign n534 = n533 ^ n414;
  assign n528 = ~n59 & n502;
  assign n529 = n528 ^ n360;
  assign n535 = n534 ^ n529;
  assign n537 = n536 ^ n361;
  assign n538 = n537 ^ n342;
  assign n539 = n538 ^ n239;
  assign n540 = ~n535 & ~n539;
  assign n541 = n527 & n540;
  assign n542 = n514 & n541;
  assign n543 = n488 & n542;
  assign n1963 = n523 ^ n293;
  assign n1964 = n1963 ^ n114;
  assign n1965 = ~n882 & n1964;
  assign n1966 = n838 ^ n671;
  assign n1967 = n977 ^ n421;
  assign n1968 = n1966 & ~n1967;
  assign n1969 = n1965 & n1968;
  assign n1970 = n430 ^ n349;
  assign n1971 = n834 ^ n363;
  assign n1972 = n1971 ^ n84;
  assign n1973 = ~n1970 & ~n1972;
  assign n1974 = n1969 & n1973;
  assign n1975 = n657 ^ n403;
  assign n1976 = n1975 ^ n310;
  assign n1977 = n353 ^ n229;
  assign n1978 = n1977 ^ n384;
  assign n1979 = n1976 & n1978;
  assign n1980 = n1021 & n1979;
  assign n1981 = n1974 & n1980;
  assign n1982 = n374 ^ n174;
  assign n1983 = ~n1397 & ~n1982;
  assign n1985 = n453 ^ n204;
  assign n1986 = n1985 ^ n302;
  assign n425 = n424 ^ n423;
  assign n1984 = n425 ^ n250;
  assign n1987 = n1986 ^ n1984;
  assign n1988 = n1983 & ~n1987;
  assign n1989 = n617 ^ n219;
  assign n1990 = n1989 ^ n575;
  assign n1991 = n1990 ^ n820;
  assign n1992 = n419 ^ n173;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = ~n856 & n1993;
  assign n1995 = n1988 & n1994;
  assign n1996 = n1981 & n1995;
  assign n1962 = n1961 ^ n1951;
  assign n1997 = n1996 ^ n1962;
  assign n2005 = n1013 ^ n175;
  assign n2006 = n2005 ^ n1990;
  assign n2004 = n355 ^ n274;
  assign n2007 = n2006 ^ n2004;
  assign n2008 = n452 & ~n2007;
  assign n2009 = n1972 ^ n223;
  assign n2010 = n2009 ^ n344;
  assign n2011 = n2008 & n2010;
  assign n2013 = n1069 ^ n403;
  assign n2012 = n674 ^ n490;
  assign n2014 = n2013 ^ n2012;
  assign n2015 = n2011 & ~n2014;
  assign n2016 = n486 ^ n402;
  assign n2017 = n430 ^ n360;
  assign n2018 = n2017 ^ n304;
  assign n2019 = ~n2016 & ~n2018;
  assign n2020 = n840 ^ n281;
  assign n2021 = n2020 ^ n227;
  assign n2022 = n2019 & ~n2021;
  assign n2023 = ~n141 & ~n664;
  assign n2024 = n2022 & n2023;
  assign n2025 = ~n703 & n2024;
  assign n2026 = n694 ^ n510;
  assign n2027 = n817 ^ n191;
  assign n2028 = ~n2026 & ~n2027;
  assign n2029 = ~n691 & n2028;
  assign n2030 = n254 & ~n652;
  assign n2031 = n2029 & n2030;
  assign n2032 = n2025 & n2031;
  assign n2033 = n2015 & n2032;
  assign n1999 = n1943 ^ n1938;
  assign n2000 = ~n1916 & n1999;
  assign n2001 = n2000 ^ n1938;
  assign n2002 = n1942 & ~n2001;
  assign n2003 = n2002 ^ n941;
  assign n2034 = n2033 ^ n2003;
  assign n2036 = n492 ^ n378;
  assign n2037 = n2036 ^ n172;
  assign n2038 = n2015 & ~n2037;
  assign n2039 = n427 ^ n243;
  assign n2040 = n2039 ^ n61;
  assign n2041 = n544 & n2040;
  assign n2042 = ~n871 & ~n2041;
  assign n2044 = n331 ^ n278;
  assign n2045 = n2044 ^ n337;
  assign n2043 = n511 ^ n348;
  assign n2046 = n2045 ^ n2043;
  assign n2047 = n2042 & n2046;
  assign n2048 = n159 ^ n100;
  assign n2049 = ~n43 & n2048;
  assign n2050 = n2049 ^ n728;
  assign n2051 = n289 ^ n147;
  assign n2052 = n2050 & n2051;
  assign n2053 = ~n267 & ~n2052;
  assign n2054 = n1154 ^ n76;
  assign n2055 = ~n59 & n2054;
  assign n2056 = n2055 ^ n76;
  assign n2057 = ~n532 & n2056;
  assign n2058 = n2057 ^ n137;
  assign n2059 = ~n351 & ~n2058;
  assign n2060 = n2053 & n2059;
  assign n2061 = n1988 & n2060;
  assign n2062 = n2047 & n2061;
  assign n2063 = n2038 & n2062;
  assign n2035 = n1936 ^ n1916;
  assign n2064 = n2063 ^ n2035;
  assign n2095 = n1904 ^ n1367;
  assign n2096 = n1904 ^ n1897;
  assign n2097 = n2095 & ~n2096;
  assign n2094 = n1906 ^ n1368;
  assign n2098 = n2097 ^ n2094;
  assign n2099 = n2098 ^ n1239;
  assign n2065 = n1028 ^ n471;
  assign n2066 = ~n1177 & ~n2065;
  assign n2067 = n454 ^ n243;
  assign n2068 = n2067 ^ n204;
  assign n2069 = n324 & ~n2068;
  assign n2070 = n2066 & n2069;
  assign n2071 = ~n1025 & n2070;
  assign n2072 = n510 ^ n242;
  assign n2073 = n2072 ^ n300;
  assign n2074 = n623 ^ n355;
  assign n2075 = n2074 ^ n740;
  assign n2076 = ~n2073 & ~n2075;
  assign n2077 = n258 ^ n137;
  assign n2078 = n59 & ~n2077;
  assign n2079 = ~n101 & ~n2078;
  assign n2080 = n467 ^ n342;
  assign n2081 = n2080 ^ n349;
  assign n2082 = n2081 ^ n840;
  assign n2083 = ~n2079 & ~n2082;
  assign n2084 = n617 ^ n403;
  assign n2085 = n2084 ^ n365;
  assign n2086 = n2083 & ~n2085;
  assign n2087 = n2076 & n2086;
  assign n2088 = n74 & n447;
  assign n2089 = n2088 ^ n412;
  assign n2090 = n2089 ^ n657;
  assign n2091 = n2087 & ~n2090;
  assign n2092 = n1057 & n2091;
  assign n2093 = n2071 & n2092;
  assign n2100 = n2099 ^ n2093;
  assign n2114 = n2095 ^ n1897;
  assign n375 = n374 ^ n373;
  assign n372 = n371 ^ n342;
  assign n376 = n375 ^ n372;
  assign n377 = n237 ^ n229;
  assign n385 = n384 ^ n377;
  assign n386 = ~n376 & n385;
  assign n387 = n335 ^ n217;
  assign n388 = n387 ^ n281;
  assign n389 = n386 & n388;
  assign n2101 = n817 ^ n519;
  assign n2102 = n2101 ^ n321;
  assign n2103 = ~n306 & ~n2102;
  assign n2104 = n973 & n2103;
  assign n2105 = n389 & n2104;
  assign n2106 = n301 ^ n172;
  assign n2107 = n2106 ^ n228;
  assign n2108 = n2107 ^ n693;
  assign n2109 = n1038 & ~n2108;
  assign n2110 = ~n978 & n2109;
  assign n2111 = n2105 & n2110;
  assign n2112 = n596 & n970;
  assign n2113 = n2111 & n2112;
  assign n2115 = n2114 ^ n2113;
  assign n2123 = ~n383 & n518;
  assign n2124 = n2123 ^ n618;
  assign n2121 = n365 ^ n278;
  assign n2122 = n2121 ^ n676;
  assign n2125 = n2124 ^ n2122;
  assign n2126 = n492 ^ n349;
  assign n2127 = n2126 ^ n430;
  assign n2128 = n2125 & ~n2127;
  assign n2129 = n1055 & n2128;
  assign n2130 = n565 ^ n454;
  assign n2131 = n484 ^ n187;
  assign n2132 = n2131 ^ n290;
  assign n2133 = n227 ^ n196;
  assign n2134 = ~n2132 & ~n2133;
  assign n2135 = ~n2130 & n2134;
  assign n2136 = n666 ^ n223;
  assign n2137 = n2136 ^ n1009;
  assign n2138 = ~n839 & ~n2137;
  assign n2139 = n2135 & n2138;
  assign n2140 = n2129 & n2139;
  assign n2141 = n488 & n2140;
  assign n2116 = n1892 ^ n1502;
  assign n2117 = n2116 ^ n1499;
  assign n2118 = ~n1888 & ~n2117;
  assign n2119 = n2118 ^ n1499;
  assign n2120 = n2119 ^ n1371;
  assign n2142 = n2141 ^ n2120;
  assign n2145 = n425 ^ n249;
  assign n2146 = ~n2021 & ~n2145;
  assign n2148 = n870 ^ n301;
  assign n2149 = n2148 ^ n372;
  assign n2147 = n732 ^ n273;
  assign n2150 = n2149 ^ n2147;
  assign n2151 = n2146 & ~n2150;
  assign n2152 = ~n814 & ~n2127;
  assign n2153 = n241 & n502;
  assign n2154 = n2153 ^ n360;
  assign n2155 = n2152 & ~n2154;
  assign n2157 = n336 ^ n274;
  assign n2156 = n693 ^ n565;
  assign n2158 = n2157 ^ n2156;
  assign n2159 = n2158 ^ n353;
  assign n2160 = n183 ^ n72;
  assign n2161 = n607 ^ n100;
  assign n2162 = n2161 ^ n870;
  assign n2163 = ~n2160 & ~n2162;
  assign n2164 = n2163 ^ n498;
  assign n2165 = ~n2159 & ~n2164;
  assign n2168 = n977 ^ n467;
  assign n2166 = n74 & n137;
  assign n2167 = n2166 ^ n450;
  assign n2169 = n2168 ^ n2167;
  assign n2170 = n2165 & ~n2169;
  assign n2171 = n2155 & n2170;
  assign n2172 = n2151 & n2171;
  assign n2173 = n890 & n2172;
  assign n2143 = n1496 ^ n1454;
  assign n2144 = n2143 ^ n1888;
  assign n2174 = n2173 ^ n2144;
  assign n2182 = n348 ^ n84;
  assign n2183 = n400 ^ n187;
  assign n2184 = n2183 ^ n405;
  assign n2185 = ~n2182 & ~n2184;
  assign n2186 = ~n327 & ~n380;
  assign n2187 = n43 & ~n159;
  assign n2188 = n2186 & ~n2187;
  assign n2189 = ~n670 & ~n2188;
  assign n2190 = n2185 & n2189;
  assign n2191 = n2017 ^ n1985;
  assign n2192 = n2191 ^ n190;
  assign n2193 = n2190 & ~n2192;
  assign n2194 = n320 ^ n236;
  assign n2195 = ~n2126 & ~n2194;
  assign n2197 = n524 ^ n484;
  assign n2196 = n840 ^ n459;
  assign n2198 = n2197 ^ n2196;
  assign n2199 = n2195 & n2198;
  assign n2200 = n165 ^ n125;
  assign n2201 = ~n61 & n2200;
  assign n2202 = n2201 ^ n510;
  assign n2203 = n2202 ^ n565;
  assign n2204 = ~n826 & ~n2203;
  assign n2205 = n2199 & n2204;
  assign n2206 = n2193 & n2205;
  assign n2207 = n389 & n2206;
  assign n2180 = n1574 ^ n1507;
  assign n2181 = n2180 ^ n1877;
  assign n2208 = n2207 ^ n2181;
  assign n2209 = n1869 ^ n1859;
  assign n2210 = n2209 ^ n1867;
  assign n2211 = ~n1860 & n2210;
  assign n2212 = n2211 ^ n1867;
  assign n2213 = n2212 ^ n1845;
  assign n2214 = n445 & ~n1142;
  assign n2216 = n100 & n117;
  assign n2215 = n337 ^ n195;
  assign n2217 = n2216 ^ n2215;
  assign n2218 = ~n267 & ~n2217;
  assign n2219 = ~n865 & n2218;
  assign n2220 = n1145 ^ n677;
  assign n2221 = n2219 & ~n2220;
  assign n2222 = n889 & ~n1047;
  assign n2223 = n2221 & n2222;
  assign n2224 = n2151 & n2223;
  assign n2225 = n1974 & n2224;
  assign n2226 = ~n2214 & n2225;
  assign n2227 = n2213 & n2226;
  assign n2228 = n2227 ^ n2207;
  assign n2229 = ~n2208 & ~n2228;
  assign n2230 = n2229 ^ n2181;
  assign n2175 = n1882 ^ n1876;
  assign n2176 = n2175 ^ n1576;
  assign n2177 = n1877 & n2176;
  assign n2178 = n2177 ^ n1576;
  assign n2179 = n2178 ^ n1503;
  assign n2231 = n2230 ^ n2179;
  assign n2232 = n625 ^ n267;
  assign n2233 = n361 ^ n251;
  assign n2234 = n2233 ^ n320;
  assign n2235 = n2234 ^ n109;
  assign n2236 = n2232 & ~n2235;
  assign n2237 = n423 ^ n175;
  assign n2238 = n963 & ~n2237;
  assign n2239 = n2236 & n2238;
  assign n2240 = n2165 & n2239;
  assign n2241 = n513 & n712;
  assign n2242 = n2240 & n2241;
  assign n2243 = n993 ^ n278;
  assign n2244 = n2243 ^ n322;
  assign n2245 = ~n462 & ~n2244;
  assign n2246 = n2126 ^ n2039;
  assign n2247 = n2245 & n2246;
  assign n2248 = n433 ^ n237;
  assign n2249 = n414 ^ n291;
  assign n2250 = ~n2248 & ~n2249;
  assign n2251 = n2247 & n2250;
  assign n2252 = ~n469 & n2104;
  assign n2253 = n2251 & n2252;
  assign n2254 = n2242 & n2253;
  assign n2255 = n2254 ^ n2230;
  assign n2256 = n2231 & n2255;
  assign n2257 = n2256 ^ n2179;
  assign n2258 = n2257 ^ n2144;
  assign n2259 = n2174 & n2258;
  assign n2260 = n2259 ^ n2257;
  assign n2261 = n2260 ^ n2141;
  assign n2262 = n2142 & n2261;
  assign n2263 = n2262 ^ n2120;
  assign n2264 = n2263 ^ n2114;
  assign n2265 = ~n2115 & n2264;
  assign n2266 = n2265 ^ n2263;
  assign n2267 = n2266 ^ n2099;
  assign n2268 = n2100 & ~n2267;
  assign n2269 = n2268 ^ n2266;
  assign n2270 = n2269 ^ n2035;
  assign n2271 = n2064 & ~n2270;
  assign n2272 = n2271 ^ n2269;
  assign n2273 = n2272 ^ n2003;
  assign n2274 = ~n2034 & n2273;
  assign n2275 = n2274 ^ n2272;
  assign n1998 = n1948 ^ n946;
  assign n2276 = n2275 ^ n1998;
  assign n2277 = n419 ^ n278;
  assign n2278 = n2277 ^ n115;
  assign n2279 = n506 ^ n285;
  assign n2280 = n2278 & ~n2279;
  assign n2282 = n484 ^ n239;
  assign n2283 = n2282 ^ n674;
  assign n2281 = n137 & ~n850;
  assign n2284 = n2283 ^ n2281;
  assign n2285 = n2280 & ~n2284;
  assign n2286 = n818 ^ n709;
  assign n2287 = ~n887 & ~n2286;
  assign n2288 = n646 & n2287;
  assign n2289 = n2285 & n2288;
  assign n2290 = n1151 & n2289;
  assign n2291 = ~n348 & ~n1004;
  assign n2292 = n2290 & n2291;
  assign n2293 = n2292 ^ n1998;
  assign n2294 = ~n2276 & n2293;
  assign n2295 = n2294 ^ n2275;
  assign n2296 = n2295 ^ n1962;
  assign n2297 = ~n1997 & n2296;
  assign n2298 = n2297 ^ n2295;
  assign n2353 = n543 & n2298;
  assign n2299 = n2298 ^ n543;
  assign n2381 = n2353 ^ n2299;
  assign n2382 = ~n2352 & ~n2381;
  assign n2354 = n2352 & n2353;
  assign n2406 = n2382 ^ n2354;
  assign n2305 = n1953 & ~n2304;
  assign n2308 = n1958 & n2307;
  assign n2309 = ~n2305 & ~n2308;
  assign n2310 = n1951 & ~n2309;
  assign n2311 = n2310 ^ n543;
  assign n2312 = n2299 & ~n2311;
  assign n2313 = n2312 ^ n2298;
  assign n2407 = n2406 ^ n2313;
  assign n2355 = n2295 ^ n1997;
  assign n2356 = n2292 ^ n2276;
  assign n2357 = n2272 ^ n2034;
  assign n2358 = n2269 ^ n2064;
  assign n2359 = n2266 ^ n2100;
  assign n2360 = n2263 ^ n2115;
  assign n2361 = n2260 ^ n2142;
  assign n2362 = n2257 ^ n2174;
  assign n2363 = n2254 ^ n2179;
  assign n2364 = n2363 ^ n2230;
  assign n2368 = n2227 ^ n2208;
  assign n2408 = ~n2364 & n2368;
  assign n2409 = n2362 & ~n2408;
  assign n2410 = n2361 & ~n2409;
  assign n2411 = n2360 & ~n2410;
  assign n2412 = n2359 & ~n2411;
  assign n2413 = ~n2358 & ~n2412;
  assign n2414 = ~n2357 & ~n2413;
  assign n2415 = ~n2356 & ~n2414;
  assign n2416 = ~n2355 & ~n2415;
  assign n2417 = ~n2407 & ~n2416;
  assign n2418 = n2417 ^ n2313;
  assign n2317 = n1013 ^ n523;
  assign n2318 = n2317 ^ n419;
  assign n2319 = n274 ^ n248;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = n2182 ^ n1166;
  assign n2322 = n1970 ^ n486;
  assign n2323 = ~n2321 & ~n2322;
  assign n2324 = n273 ^ n191;
  assign n2325 = n2324 ^ n174;
  assign n2326 = n2323 & ~n2325;
  assign n2327 = n2320 & n2326;
  assign n2328 = n848 & n2327;
  assign n2329 = n437 ^ n414;
  assign n2330 = n2329 ^ n110;
  assign n2331 = n2080 ^ n243;
  assign n2332 = n2331 ^ n450;
  assign n2333 = n2332 ^ n321;
  assign n2334 = n2330 & ~n2333;
  assign n2335 = n258 ^ n154;
  assign n2336 = ~n1129 & n2335;
  assign n2337 = n2334 & ~n2336;
  assign n2339 = ~n61 & n1124;
  assign n2340 = n2339 ^ n365;
  assign n2338 = n667 ^ n268;
  assign n2341 = n2340 ^ n2338;
  assign n2342 = ~n1991 & ~n2341;
  assign n2343 = n2337 & n2342;
  assign n2344 = n881 & n2343;
  assign n2345 = n2328 & n2344;
  assign n2419 = n2417 ^ n2345;
  assign n156 = n155 ^ n100;
  assign n391 = n390 ^ n156;
  assign n392 = ~n59 & n391;
  assign n396 = n395 ^ n394;
  assign n393 = n219 ^ n191;
  assign n397 = n396 ^ n393;
  assign n398 = ~n392 & ~n397;
  assign n399 = n389 & n398;
  assign n431 = n430 ^ n268;
  assign n429 = n428 ^ n427;
  assign n432 = n431 ^ n429;
  assign n434 = n433 ^ n197;
  assign n438 = n437 ^ n434;
  assign n439 = n432 & n438;
  assign n440 = ~n425 & n439;
  assign n441 = n422 & n440;
  assign n442 = n411 & n441;
  assign n443 = n399 & n442;
  assign n444 = n369 & n443;
  assign n2420 = n2345 ^ n444;
  assign n2421 = n2419 & n2420;
  assign n2422 = ~n2418 & n2421;
  assign n2423 = n2422 ^ n2345;
  assign n2424 = ~n316 & ~n2423;
  assign n2315 = ~n444 & ~n2313;
  assign n2314 = n2313 ^ n444;
  assign n2316 = n2315 ^ n2314;
  assign n2347 = n2316 & ~n2345;
  assign n2365 = n2226 ^ n2213;
  assign n2366 = ~n2208 & n2365;
  assign n2367 = n2366 ^ n2365;
  assign n2369 = n2368 ^ n2367;
  assign n2370 = n2364 & ~n2369;
  assign n2371 = ~n2362 & ~n2370;
  assign n2372 = ~n2361 & ~n2371;
  assign n2373 = ~n2360 & ~n2372;
  assign n2374 = ~n2359 & ~n2373;
  assign n2375 = n2358 & ~n2374;
  assign n2376 = n2357 & ~n2375;
  assign n2377 = n2356 & ~n2376;
  assign n2378 = n2355 & ~n2377;
  assign n2383 = ~n2378 & n2382;
  assign n2384 = n2383 ^ n2313;
  assign n2379 = n2313 & n2378;
  assign n2380 = ~n2354 & ~n2379;
  assign n2385 = n2384 ^ n2380;
  assign n2386 = n444 & n2385;
  assign n2387 = n2386 ^ n2380;
  assign n2388 = n2347 & n2387;
  assign n2389 = n316 & ~n2388;
  assign n3258 = n2424 ^ n2389;
  assign n3259 = n25 & n3258;
  assign n3260 = n3259 ^ x1;
  assign n2346 = n2345 ^ n2316;
  assign n2348 = n2347 ^ n2346;
  assign n2349 = n316 & n2348;
  assign n160 = n159 ^ n156;
  assign n161 = n147 & n160;
  assign n162 = n146 & ~n161;
  assign n209 = n208 ^ n107;
  assign n210 = n106 ^ n59;
  assign n211 = n209 & ~n210;
  assign n220 = n219 ^ n212;
  assign n221 = ~n211 & ~n220;
  assign n230 = n229 ^ n228;
  assign n222 = n138 & ~n203;
  assign n231 = n230 ^ n222;
  assign n232 = n221 & ~n231;
  assign n233 = ~n205 & n232;
  assign n234 = n199 & n233;
  assign n235 = n162 & n234;
  assign n2447 = n2349 ^ n235;
  assign n3257 = n2447 ^ x22;
  assign n3261 = n3260 ^ n3257;
  assign n3225 = n2348 ^ n316;
  assign n3255 = n3225 ^ n1385;
  assign n3256 = x1 & n3255;
  assign n3262 = n3261 ^ n3256;
  assign n3263 = n3262 ^ n3261;
  assign n3264 = n1387 & ~n2346;
  assign n3265 = ~n3263 & ~n3264;
  assign n3266 = n3265 ^ n3261;
  assign n3267 = ~x0 & ~n3266;
  assign n3268 = n3267 ^ n3261;
  assign n2936 = n2416 ^ n2385;
  assign n2937 = n2936 ^ n2417;
  assign n2938 = n2937 ^ n2416;
  assign n2471 = x22 & n27;
  assign n2472 = n2471 ^ n25;
  assign n2466 = n25 & n27;
  assign n2467 = n2466 ^ n25;
  assign n2465 = n29 ^ n28;
  assign n2468 = n2467 ^ n2465;
  assign n2453 = x0 & ~x22;
  assign n2454 = n2453 ^ x0;
  assign n2461 = n2454 ^ x1;
  assign n2462 = n2461 ^ n27;
  assign n2459 = n2453 ^ x2;
  assign n2456 = ~x2 & ~n2453;
  assign n2460 = n2459 ^ n2456;
  assign n2463 = n2462 ^ n2460;
  assign n2464 = ~n1390 & ~n2463;
  assign n2469 = n2468 ^ n2464;
  assign n2470 = n2469 ^ n1390;
  assign n2473 = n2472 ^ n2470;
  assign n2455 = x2 & ~n2454;
  assign n2457 = n2456 ^ n2455;
  assign n2458 = n2457 ^ n1389;
  assign n2474 = n2473 ^ n2458;
  assign n2475 = n2474 ^ n2464;
  assign n2476 = n2475 ^ n29;
  assign n2942 = n2476 ^ n1393;
  assign n3193 = n2314 ^ n1337;
  assign n3194 = ~n2942 & n3193;
  assign n3195 = n2938 & n3194;
  assign n2957 = ~n1393 & ~n2476;
  assign n2958 = n2957 ^ n2476;
  assign n2959 = ~n1337 & ~n2958;
  assign n3196 = n2355 & n2959;
  assign n3197 = n3196 ^ n2958;
  assign n3198 = n1337 & n2407;
  assign n2947 = n1283 & ~n1337;
  assign n3199 = n3198 ^ n2947;
  assign n3200 = ~n3197 & n3199;
  assign n2995 = ~n1283 & n2959;
  assign n2991 = n2959 ^ n1283;
  assign n2961 = n2959 ^ n2958;
  assign n2943 = ~n1337 & ~n2942;
  assign n2956 = n2943 ^ n1337;
  assign n2960 = n2959 ^ n2956;
  assign n2962 = n2961 ^ n2960;
  assign n2990 = n2962 ^ n2942;
  assign n2992 = n2991 ^ n2990;
  assign n2988 = n1283 & ~n2962;
  assign n2969 = n1283 & n2942;
  assign n2989 = n2988 ^ n2969;
  assign n2993 = n2992 ^ n2989;
  assign n2994 = n2993 ^ n2959;
  assign n2996 = n2995 ^ n2994;
  assign n3202 = ~n2355 & n2996;
  assign n3201 = n2407 & ~n2960;
  assign n3203 = n3202 ^ n3201;
  assign n3204 = ~n3200 & ~n3203;
  assign n3206 = ~n1283 & n3204;
  assign n3205 = n3204 ^ n1283;
  assign n3207 = n3206 ^ n3205;
  assign n3208 = ~n3195 & ~n3207;
  assign n2970 = n2969 ^ n1283;
  assign n2939 = n2406 ^ n444;
  assign n2940 = ~n2938 & ~n2939;
  assign n3209 = n2940 ^ n2417;
  assign n3210 = n3209 ^ n2938;
  assign n3211 = n2970 & ~n3210;
  assign n3212 = n3208 & ~n3211;
  assign n3213 = ~n2942 & ~n3209;
  assign n3214 = n3206 & ~n3213;
  assign n3215 = n3212 & ~n3214;
  assign n2674 = n754 & ~n2365;
  assign n2482 = n794 & n955;
  assign n2478 = n955 ^ n794;
  assign n2483 = n2482 ^ n2478;
  assign n2675 = n792 & ~n2365;
  assign n2676 = ~n2483 & ~n2675;
  assign n2677 = n2482 ^ n2365;
  assign n2678 = n2208 ^ n792;
  assign n2679 = n2482 & n2678;
  assign n2680 = n2679 ^ n2208;
  assign n2681 = n2677 & n2680;
  assign n2682 = n2681 ^ n2365;
  assign n2683 = ~n2676 & ~n2682;
  assign n2684 = n753 & n2683;
  assign n2685 = n2684 ^ n753;
  assign n2689 = n792 ^ n753;
  assign n2690 = n2367 & n2689;
  assign n2691 = n2690 ^ n2364;
  assign n2692 = n2478 & ~n2691;
  assign n2479 = n792 & n2478;
  assign n2489 = ~n753 & n2479;
  assign n2486 = n2483 ^ n753;
  assign n2487 = n2483 ^ n792;
  assign n2488 = n2486 & ~n2487;
  assign n2490 = n2489 ^ n2488;
  assign n2687 = ~n2365 & n2490;
  assign n2480 = n2479 ^ n2478;
  assign n2481 = n2480 ^ n792;
  assign n2484 = n2483 ^ n2481;
  assign n2686 = n2368 & n2484;
  assign n2688 = n2687 ^ n2686;
  assign n2693 = n2692 ^ n2688;
  assign n2694 = n2685 & ~n2693;
  assign n2695 = ~n2674 & ~n2694;
  assign n2696 = ~n2364 & n2484;
  assign n2697 = n2368 & n2490;
  assign n2698 = ~n2696 & ~n2697;
  assign n2507 = n2408 ^ n2370;
  assign n2699 = ~n2507 & n2689;
  assign n2700 = n2699 ^ n2362;
  assign n2701 = n2478 & ~n2700;
  assign n2702 = n2698 & ~n2701;
  assign n2703 = n2702 ^ n753;
  assign n2704 = ~n2695 & ~n2703;
  assign n2668 = n751 & ~n2365;
  assign n2669 = n2668 ^ n2368;
  assign n2670 = ~n754 & n2669;
  assign n2671 = n2670 ^ n2368;
  assign n2524 = ~n555 & ~n2365;
  assign n2672 = n2671 ^ n2524;
  assign n2550 = n2409 ^ n2371;
  assign n2651 = n2361 & n2478;
  assign n2652 = n2550 & n2651;
  assign n2653 = ~n2362 & n2484;
  assign n2654 = ~n2364 & n2490;
  assign n2655 = ~n2653 & ~n2654;
  assign n2656 = ~n2652 & n2655;
  assign n2657 = ~n753 & ~n2656;
  assign n2658 = n2478 & ~n2550;
  assign n2660 = n2361 ^ n792;
  assign n2659 = n753 & n2655;
  assign n2661 = n2660 ^ n2659;
  assign n2662 = n2661 ^ n2660;
  assign n2663 = ~n2651 & n2662;
  assign n2664 = n2663 ^ n2660;
  assign n2665 = ~n2658 & n2664;
  assign n2666 = n2665 ^ n2660;
  assign n2667 = ~n2657 & ~n2666;
  assign n2673 = n2672 ^ n2667;
  assign n2807 = n2704 ^ n2673;
  assign n2493 = n2413 ^ n2375;
  assign n2578 = n2493 ^ n2374;
  assign n2719 = n1283 ^ n1163;
  assign n2798 = n2578 & n2719;
  assign n2722 = n1163 & n1283;
  assign n2736 = ~n955 & n2722;
  assign n2737 = n2736 ^ n959;
  assign n2723 = n2722 ^ n2719;
  assign n2732 = ~n955 & ~n2723;
  assign n2733 = n2732 ^ n2723;
  assign n2726 = ~n955 & n959;
  assign n2727 = n2723 & ~n2726;
  assign n2728 = n2727 ^ n2726;
  assign n2734 = n2733 ^ n2728;
  assign n2720 = n959 & n2719;
  assign n2721 = n2720 ^ n959;
  assign n2724 = n2723 ^ n2721;
  assign n2730 = n955 & ~n2724;
  assign n2731 = n2730 ^ n2724;
  assign n2735 = n2734 ^ n2731;
  assign n2738 = n2737 ^ n2735;
  assign n2725 = ~n959 & n2724;
  assign n2729 = n2728 ^ n2725;
  assign n2739 = n2738 ^ n2729;
  assign n2795 = ~n2360 & ~n2739;
  assign n2794 = n2359 & ~n2724;
  assign n2796 = n2795 ^ n2794;
  assign n2576 = n2412 ^ n2374;
  assign n2793 = ~n2576 & n2719;
  assign n2797 = n2796 ^ n2793;
  assign n2799 = n2798 ^ n2797;
  assign n2800 = ~n955 & n2799;
  assign n2801 = n955 & ~n2796;
  assign n2802 = ~n2798 & n2801;
  assign n2803 = n2358 ^ n959;
  assign n2804 = n2793 & ~n2803;
  assign n2805 = ~n2802 & ~n2804;
  assign n2806 = ~n2800 & n2805;
  assign n2808 = n2807 ^ n2806;
  assign n2827 = n2703 ^ n2674;
  assign n2828 = n2827 ^ n2694;
  assign n2829 = n2694 & n2703;
  assign n2830 = n2828 & ~n2829;
  assign n2594 = n2411 ^ n2373;
  assign n2818 = n2594 ^ n2361;
  assign n2819 = n2739 & ~n2818;
  assign n2820 = n2819 ^ n2361;
  assign n2821 = n2820 ^ n2360;
  assign n2817 = n959 & ~n2594;
  assign n2822 = n2821 ^ n2817;
  assign n2823 = n2822 ^ n2820;
  assign n2824 = n2724 & n2823;
  assign n2825 = n2824 ^ n2821;
  assign n2602 = n2576 ^ n2373;
  assign n2810 = n2602 ^ n955;
  assign n2606 = n2594 ^ n2359;
  assign n2607 = n2606 ^ n2602;
  assign n2608 = n2607 ^ n2359;
  assign n2811 = n2810 ^ n2608;
  assign n2812 = n2811 ^ n2724;
  assign n2813 = ~n2594 & n2724;
  assign n2814 = n2812 & n2813;
  assign n2815 = n2814 ^ n2812;
  assign n2809 = n2359 & n2719;
  assign n2816 = n2815 ^ n2809;
  assign n2826 = n2825 ^ n2816;
  assign n2831 = n2830 ^ n2826;
  assign n2865 = n794 & ~n2365;
  assign n2866 = n2865 ^ n2368;
  assign n2867 = ~n2478 & n2866;
  assign n2868 = n2867 ^ n2368;
  assign n2869 = n2868 ^ n2675;
  assign n2840 = n2507 ^ n2368;
  assign n2841 = n2739 & ~n2840;
  assign n2842 = n2841 ^ n2368;
  assign n2834 = ~n2507 & n2724;
  assign n2839 = n959 & n2834;
  assign n2843 = n2842 ^ n2839;
  assign n2838 = ~n2364 & ~n2724;
  assign n2844 = n2843 ^ n2838;
  assign n2835 = n2507 ^ n955;
  assign n2836 = ~n2834 & ~n2835;
  assign n2833 = ~n2362 & n2719;
  assign n2837 = n2836 ^ n2833;
  assign n2845 = n2844 ^ n2837;
  assign n2846 = ~n960 & n2367;
  assign n2847 = n2846 ^ n2364;
  assign n2848 = n2719 & ~n2847;
  assign n2850 = ~n2365 & ~n2739;
  assign n2849 = n2368 & ~n2724;
  assign n2851 = n2850 ^ n2849;
  assign n2852 = ~n2848 & ~n2851;
  assign n2853 = n2722 ^ n2721;
  assign n2854 = n2368 & n2719;
  assign n2855 = n2365 & ~n2854;
  assign n2856 = ~n2853 & ~n2855;
  assign n2857 = n955 & n2856;
  assign n2858 = n2857 ^ n955;
  assign n2859 = n2852 & n2858;
  assign n2860 = ~n2365 & n2478;
  assign n2862 = n2859 & n2860;
  assign n2861 = n2860 ^ n2859;
  assign n2863 = n2862 ^ n2861;
  assign n2864 = n2845 & n2863;
  assign n2870 = n2869 ^ n2864;
  assign n2878 = ~n2364 & ~n2739;
  assign n2877 = ~n2362 & ~n2724;
  assign n2879 = n2878 ^ n2877;
  assign n2875 = ~n2550 & n2720;
  assign n2871 = ~n955 & ~n2550;
  assign n2872 = n2871 ^ n2361;
  assign n2873 = n2719 & n2872;
  assign n2874 = n2873 ^ n955;
  assign n2876 = n2875 ^ n2874;
  assign n2880 = n2879 ^ n2876;
  assign n2881 = n2880 ^ n2869;
  assign n2882 = n2870 & ~n2881;
  assign n2883 = n2882 ^ n2864;
  assign n2832 = n2693 ^ n2684;
  assign n2884 = n2883 ^ n2832;
  assign n2563 = n2410 ^ n2372;
  assign n2895 = n2563 ^ n2362;
  assign n2896 = n2739 & n2895;
  assign n2897 = n2896 ^ n2362;
  assign n2898 = n2897 ^ n2361;
  assign n2894 = ~n959 & ~n2563;
  assign n2899 = n2898 ^ n2894;
  assign n2900 = n2899 ^ n2897;
  assign n2901 = n2724 & ~n2900;
  assign n2902 = n2901 ^ n2898;
  assign n2888 = n2594 ^ n2410;
  assign n2633 = n2594 ^ n2372;
  assign n2886 = n2633 ^ n955;
  assign n2887 = n2886 ^ n2724;
  assign n2889 = n2888 ^ n2887;
  assign n2890 = ~n2563 & n2724;
  assign n2891 = ~n2889 & n2890;
  assign n2892 = n2891 ^ n2889;
  assign n2885 = ~n2360 & n2719;
  assign n2893 = n2892 ^ n2885;
  assign n2903 = n2902 ^ n2893;
  assign n2904 = n2903 ^ n2832;
  assign n2905 = ~n2884 & n2904;
  assign n2906 = n2905 ^ n2903;
  assign n2907 = n2906 ^ n2826;
  assign n2908 = n2831 & n2907;
  assign n2909 = n2908 ^ n2906;
  assign n2910 = n2909 ^ n2806;
  assign n2911 = ~n2808 & ~n2910;
  assign n2912 = n2911 ^ n2909;
  assign n2787 = n2493 ^ n2359;
  assign n2788 = ~n2739 & ~n2787;
  assign n2780 = ~n2493 & n2724;
  assign n2785 = n959 & n2780;
  assign n2786 = n2785 ^ n2724;
  assign n2789 = n2788 ^ n2786;
  assign n2784 = n2358 & ~n2724;
  assign n2790 = n2789 ^ n2784;
  assign n2782 = ~n2357 & n2719;
  assign n2756 = n2724 ^ n955;
  assign n2781 = n2756 & ~n2780;
  assign n2783 = n2782 ^ n2781;
  assign n2791 = n2790 ^ n2783;
  assign n2705 = n2704 ^ n2672;
  assign n2706 = ~n2673 & ~n2705;
  assign n2707 = n2706 ^ n2667;
  assign n2525 = n583 & ~n1955;
  assign n2526 = n2525 ^ n1955;
  assign n2527 = ~n2524 & ~n2526;
  assign n2528 = ~n2366 & ~n2527;
  assign n2529 = n555 & n1954;
  assign n2530 = ~n2365 & n2529;
  assign n2531 = n2530 ^ n1954;
  assign n2532 = n2528 & ~n2531;
  assign n2648 = ~n583 & n2532;
  assign n2533 = n584 & n2367;
  assign n2534 = n2533 ^ n2364;
  assign n2535 = n754 & ~n2534;
  assign n2536 = n2529 ^ n2300;
  assign n2537 = n2368 & n2536;
  assign n2538 = ~n583 & n1954;
  assign n2539 = n2538 ^ n1954;
  assign n2540 = n2539 ^ n2526;
  assign n2541 = n584 & ~n2540;
  assign n2542 = ~n2365 & n2541;
  assign n2543 = ~n2537 & ~n2542;
  assign n2544 = ~n2535 & n2543;
  assign n2649 = n2648 ^ n2544;
  assign n2622 = ~n792 & ~n2563;
  assign n2623 = ~n2360 & ~n2622;
  assign n2624 = n2361 & n2484;
  assign n2625 = ~n2362 & n2490;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = ~n2563 & n2626;
  assign n2628 = n2627 ^ n2478;
  assign n2629 = ~n753 & n2628;
  assign n2630 = n2629 ^ n2478;
  assign n2631 = n2623 & n2630;
  assign n2632 = n2626 ^ n753;
  assign n2634 = n2478 & n2633;
  assign n2635 = n2634 ^ n753;
  assign n2636 = n2360 & n2480;
  assign n2637 = ~n2563 & n2636;
  assign n2638 = n2637 ^ n753;
  assign n2639 = ~n753 & n2638;
  assign n2640 = n2639 ^ n753;
  assign n2641 = ~n2635 & ~n2640;
  assign n2642 = n2641 ^ n2639;
  assign n2643 = n2642 ^ n753;
  assign n2644 = n2643 ^ n2637;
  assign n2645 = n2632 & n2644;
  assign n2646 = n2645 ^ n2637;
  assign n2647 = ~n2631 & ~n2646;
  assign n2650 = n2649 ^ n2647;
  assign n2779 = n2707 ^ n2650;
  assign n2792 = n2791 ^ n2779;
  assign n3011 = n2912 ^ n2792;
  assign n2740 = n2416 ^ n2378;
  assign n2946 = n1337 ^ n1283;
  assign n2948 = n2947 ^ n2946;
  assign n2949 = n2948 ^ n2947;
  assign n2983 = ~n2740 & n2949;
  assign n2984 = n2983 ^ n1283;
  assign n2985 = n2984 ^ n2407;
  assign n2986 = ~n2942 & ~n2985;
  assign n2998 = n2988 ^ n1283;
  assign n2971 = n2970 ^ n2942;
  assign n2987 = n2971 ^ n1283;
  assign n2997 = n2996 ^ n2987;
  assign n2999 = n2998 ^ n2997;
  assign n3000 = ~n2355 & n2999;
  assign n3001 = n3000 ^ n2997;
  assign n3002 = n2996 ^ n2959;
  assign n3003 = ~n2356 & n3002;
  assign n3004 = n3003 ^ n2959;
  assign n3005 = n3001 ^ n2995;
  assign n3006 = n3004 & ~n3005;
  assign n3007 = n3006 ^ n2995;
  assign n3008 = ~n3001 & n3007;
  assign n3009 = n3008 ^ n3001;
  assign n3010 = ~n2986 & ~n3009;
  assign n3012 = n3011 ^ n3010;
  assign n3014 = n1283 & ~n2357;
  assign n3015 = n3014 ^ n2356;
  assign n3016 = ~n1337 & n3015;
  assign n3017 = n3016 ^ n2356;
  assign n3018 = ~n2958 & n3017;
  assign n3020 = ~n2357 & n2996;
  assign n3019 = n2356 & ~n2960;
  assign n3021 = n3020 ^ n3019;
  assign n3022 = ~n3018 & ~n3021;
  assign n3023 = n3022 ^ n1283;
  assign n2741 = n2740 ^ n2377;
  assign n3024 = ~n2741 & ~n2971;
  assign n3025 = n2355 ^ n1337;
  assign n2743 = n2415 ^ n2414;
  assign n2744 = n2743 ^ n2377;
  assign n2495 = n2414 ^ n2376;
  assign n2745 = n2744 ^ n2495;
  assign n2746 = n2745 ^ n2376;
  assign n3026 = ~n2746 & ~n2942;
  assign n3027 = ~n3025 & n3026;
  assign n3028 = ~n3024 & ~n3027;
  assign n2747 = n2746 ^ n2741;
  assign n3029 = n2747 & n2970;
  assign n3030 = n3028 & ~n3029;
  assign n3031 = ~n3023 & n3030;
  assign n3032 = n3031 ^ n3028;
  assign n3013 = n2909 ^ n2808;
  assign n3033 = n3032 ^ n3013;
  assign n3049 = n2906 ^ n2831;
  assign n3034 = ~n2744 & n2970;
  assign n3036 = n2358 & n2993;
  assign n3035 = ~n2357 & n2962;
  assign n3037 = n3036 ^ n3035;
  assign n3039 = ~n1283 & ~n3037;
  assign n3038 = n3037 ^ n1283;
  assign n3040 = n3039 ^ n3038;
  assign n3041 = ~n3034 & n3040;
  assign n3042 = n2356 ^ n1337;
  assign n3043 = ~n2495 & ~n2942;
  assign n3044 = ~n3042 & n3043;
  assign n3045 = n3041 & ~n3044;
  assign n3046 = n2745 & ~n2942;
  assign n3047 = n3039 & ~n3046;
  assign n3048 = n3045 & ~n3047;
  assign n3050 = n3049 ^ n3048;
  assign n3067 = n2903 ^ n2884;
  assign n2496 = n2495 ^ n2413;
  assign n3051 = n2496 & ~n2942;
  assign n3053 = n2359 & n2993;
  assign n3052 = n2358 & n2962;
  assign n3054 = n3053 ^ n3052;
  assign n3056 = ~n1283 & n3054;
  assign n3055 = n3054 ^ n1283;
  assign n3057 = n3056 ^ n3055;
  assign n3058 = ~n3051 & n3057;
  assign n3059 = ~n2493 & ~n2942;
  assign n3060 = n2357 ^ n1337;
  assign n3061 = n3059 & ~n3060;
  assign n3062 = ~n3058 & ~n3061;
  assign n3063 = n2495 ^ n2375;
  assign n3064 = ~n2971 & ~n3063;
  assign n3065 = ~n3056 & ~n3064;
  assign n3066 = n3062 & n3065;
  assign n3068 = n3067 ^ n3066;
  assign n3088 = n2880 ^ n2870;
  assign n3069 = ~n2576 & ~n2942;
  assign n3070 = n2358 ^ n1337;
  assign n3071 = n3069 & ~n3070;
  assign n3073 = ~n2360 & n2993;
  assign n3072 = n2359 & n2962;
  assign n3074 = n3073 ^ n3072;
  assign n3075 = n3074 ^ n1283;
  assign n3076 = n2578 & ~n2942;
  assign n3077 = n3076 ^ n3074;
  assign n3078 = n2493 ^ n2412;
  assign n3079 = n2970 & ~n3078;
  assign n3080 = n3079 ^ n3076;
  assign n3081 = ~n3077 & n3080;
  assign n3082 = n3081 ^ n3079;
  assign n3083 = n3082 ^ n3076;
  assign n3084 = n3083 ^ n3079;
  assign n3085 = ~n3075 & ~n3084;
  assign n3086 = n3085 ^ n3079;
  assign n3087 = ~n3071 & ~n3086;
  assign n3089 = n3088 ^ n3087;
  assign n3107 = n2863 ^ n2845;
  assign n3108 = ~n2862 & ~n3107;
  assign n3090 = n1337 & ~n2594;
  assign n3091 = n2359 & ~n3090;
  assign n3093 = n2361 & n2993;
  assign n3092 = ~n2360 & n2962;
  assign n3094 = n3093 ^ n3092;
  assign n3095 = ~n2594 & ~n3094;
  assign n3096 = n3095 ^ n2942;
  assign n3097 = n1283 & ~n3096;
  assign n3098 = n3097 ^ n2942;
  assign n3099 = n3091 & ~n3098;
  assign n3100 = n3094 ^ n1283;
  assign n2944 = n2943 ^ n2942;
  assign n3101 = n2607 & ~n2944;
  assign n3102 = n2608 & n2970;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = n3100 & n3103;
  assign n3105 = n3104 ^ n3101;
  assign n3106 = ~n3099 & ~n3105;
  assign n3109 = n3108 ^ n3106;
  assign n3125 = n2857 ^ n2852;
  assign n3110 = ~n2888 & ~n2971;
  assign n3112 = ~n2362 & n2993;
  assign n3111 = n2361 & n2962;
  assign n3113 = n3112 ^ n3111;
  assign n3115 = n1283 & ~n3113;
  assign n3114 = n3113 ^ n1283;
  assign n3116 = n3115 ^ n3114;
  assign n3117 = ~n3110 & ~n3116;
  assign n3118 = n2360 ^ n1337;
  assign n3119 = ~n2563 & ~n2942;
  assign n3120 = ~n3118 & n3119;
  assign n3121 = n3117 & ~n3120;
  assign n3122 = n2633 & ~n2942;
  assign n3123 = n3115 & ~n3122;
  assign n3124 = n3121 & ~n3123;
  assign n3126 = n3125 ^ n3124;
  assign n3132 = ~n2507 & n2949;
  assign n3133 = n3132 ^ n2362;
  assign n3134 = ~n2942 & ~n3133;
  assign n3136 = n2368 & n2993;
  assign n3135 = ~n2364 & n2962;
  assign n3137 = n3136 ^ n3135;
  assign n3138 = ~n3134 & ~n3137;
  assign n3139 = ~n2366 & ~n2990;
  assign n3140 = n1283 & ~n3139;
  assign n3146 = n1393 ^ n1337;
  assign n3147 = n2368 & ~n3146;
  assign n3143 = ~n1393 & n2949;
  assign n3144 = n3143 ^ n2947;
  assign n3145 = ~n2365 & n3144;
  assign n3148 = n3147 ^ n3145;
  assign n3141 = n2367 & n2949;
  assign n3142 = n3141 ^ n2364;
  assign n3149 = n3148 ^ n3142;
  assign n3150 = n2942 & ~n3149;
  assign n3151 = n3150 ^ n3142;
  assign n3152 = n3140 & n3151;
  assign n3153 = n3138 & ~n3152;
  assign n3130 = ~n2365 & n2719;
  assign n3154 = n3138 ^ n3130;
  assign n3155 = ~n3153 & n3154;
  assign n3131 = n1283 & n3130;
  assign n3156 = n3155 ^ n3131;
  assign n3127 = n2722 ^ n959;
  assign n3128 = ~n2365 & ~n3127;
  assign n3129 = n3128 ^ n2854;
  assign n3157 = n3156 ^ n3129;
  assign n3162 = ~n2364 & n3144;
  assign n3161 = ~n2362 & ~n3146;
  assign n3163 = n3162 ^ n3161;
  assign n3164 = n3163 ^ n1283;
  assign n3158 = ~n2550 & n2949;
  assign n3159 = n3158 ^ n1283;
  assign n3160 = n3159 ^ n2361;
  assign n3165 = n3164 ^ n3160;
  assign n3166 = n2942 & n3165;
  assign n3167 = n3166 ^ n3160;
  assign n3168 = n3167 ^ n3129;
  assign n3169 = n3157 & ~n3168;
  assign n3170 = n3169 ^ n3156;
  assign n3171 = n3170 ^ n3125;
  assign n3172 = n3126 & n3171;
  assign n3173 = n3172 ^ n3124;
  assign n3174 = n3173 ^ n3108;
  assign n3175 = n3109 & ~n3174;
  assign n3176 = n3175 ^ n3106;
  assign n3177 = n3176 ^ n3088;
  assign n3178 = n3089 & n3177;
  assign n3179 = n3178 ^ n3087;
  assign n3180 = n3179 ^ n3067;
  assign n3181 = ~n3068 & ~n3180;
  assign n3182 = n3181 ^ n3066;
  assign n3183 = n3182 ^ n3049;
  assign n3184 = ~n3050 & ~n3183;
  assign n3185 = n3184 ^ n3048;
  assign n3186 = n3185 ^ n3032;
  assign n3187 = n3033 & ~n3186;
  assign n3188 = n3187 ^ n3185;
  assign n3189 = n3188 ^ n3011;
  assign n3190 = n3012 & ~n3189;
  assign n3191 = n3190 ^ n3010;
  assign n2913 = n2912 ^ n2779;
  assign n2914 = n2792 & ~n2913;
  assign n2915 = n2914 ^ n2791;
  assign n2773 = n959 & ~n2495;
  assign n2774 = n2773 ^ n2414;
  assign n2775 = n2724 & n2774;
  assign n2776 = n2775 ^ n2414;
  assign n2767 = n2495 ^ n2358;
  assign n2768 = n2739 ^ n2495;
  assign n2764 = ~n2495 & n2724;
  assign n2769 = n2768 ^ n2764;
  assign n2770 = ~n2767 & n2769;
  assign n2765 = ~n955 & n2764;
  assign n2766 = n2765 ^ n955;
  assign n2771 = n2770 ^ n2766;
  assign n2763 = n2356 & n2719;
  assign n2772 = n2771 ^ n2763;
  assign n2777 = n2776 ^ n2772;
  assign n2708 = n2707 ^ n2649;
  assign n2709 = ~n2650 & ~n2708;
  assign n2710 = n2709 ^ n2647;
  assign n2545 = ~n2532 & n2544;
  assign n2615 = n2545 ^ n2365;
  assign n2508 = n584 & ~n2507;
  assign n2509 = n2508 ^ n2362;
  assign n2510 = n754 & n2509;
  assign n2511 = n555 & ~n583;
  assign n2514 = n2511 ^ n584;
  assign n2515 = n2368 & n2514;
  assign n2516 = n1954 & ~n2515;
  assign n2512 = n2368 & n2511;
  assign n2513 = ~n1955 & ~n2512;
  assign n2517 = n2516 ^ n2513;
  assign n2518 = n2516 ^ n555;
  assign n2519 = n2364 & ~n2518;
  assign n2520 = n2519 ^ n555;
  assign n2521 = n2517 & ~n2520;
  assign n2522 = n2521 ^ n2513;
  assign n2523 = ~n2510 & ~n2522;
  assign n2616 = n2523 ^ n583;
  assign n2617 = n2545 & n2616;
  assign n2618 = n2617 ^ n583;
  assign n2619 = n2615 & ~n2618;
  assign n2620 = n2619 ^ n2523;
  assign n2595 = n2478 & ~n2594;
  assign n2596 = n2359 ^ n792;
  assign n2597 = n2595 & ~n2596;
  assign n2598 = ~n2360 & n2484;
  assign n2599 = n2361 & n2490;
  assign n2600 = ~n2598 & ~n2599;
  assign n2601 = n2600 ^ n753;
  assign n2609 = n2478 & n2608;
  assign n2610 = ~n753 & n2609;
  assign n2603 = n753 & ~n2478;
  assign n2604 = n2603 ^ n753;
  assign n2605 = ~n2602 & n2604;
  assign n2611 = n2610 ^ n2605;
  assign n2612 = n2601 & ~n2611;
  assign n2613 = n2612 ^ n2605;
  assign n2614 = ~n2597 & ~n2613;
  assign n2621 = n2620 ^ n2614;
  assign n2762 = n2710 ^ n2621;
  assign n2778 = n2777 ^ n2762;
  assign n2982 = n2915 ^ n2778;
  assign n3192 = n3191 ^ n2982;
  assign n3254 = n3215 ^ n3192;
  assign n3269 = n3268 ^ n3254;
  assign n3274 = n1387 & ~n2314;
  assign n3273 = x1 & n2346;
  assign n3275 = n3274 ^ n3273;
  assign n2972 = n2423 ^ n2388;
  assign n3271 = n25 & ~n2972;
  assign n3272 = n3271 ^ n3225;
  assign n3276 = n3275 ^ n3272;
  assign n3277 = ~x0 & ~n3276;
  assign n3278 = n3277 ^ n3272;
  assign n3279 = n3278 ^ n2476;
  assign n3270 = n3188 ^ n3012;
  assign n3281 = n3279 ^ n3270;
  assign n3280 = n3270 & ~n3279;
  assign n3282 = n3281 ^ n3280;
  assign n3300 = n2476 ^ n2314;
  assign n3299 = n25 & n2938;
  assign n3301 = n3300 ^ n3299;
  assign n3297 = n2407 ^ n1385;
  assign n3298 = x1 & ~n3297;
  assign n3302 = n3301 ^ n3298;
  assign n3303 = n3302 ^ n3301;
  assign n3304 = n1387 & n2355;
  assign n3305 = ~n3303 & ~n3304;
  assign n3306 = n3305 ^ n3301;
  assign n3307 = ~x0 & n3306;
  assign n3308 = n3307 ^ n3301;
  assign n3296 = n3182 ^ n3050;
  assign n3309 = n3308 ^ n3296;
  assign n3319 = n3179 ^ n3068;
  assign n3313 = n1387 & n2356;
  assign n3312 = x1 & ~n2355;
  assign n3314 = n3313 ^ n3312;
  assign n3310 = n25 & ~n2740;
  assign n3311 = n3310 ^ n2407;
  assign n3315 = n3314 ^ n3311;
  assign n3316 = ~x0 & n3315;
  assign n3317 = n3316 ^ n3311;
  assign n3318 = n3317 ^ n2476;
  assign n3320 = n3319 ^ n3318;
  assign n3329 = n3176 ^ n3089;
  assign n3325 = ~n2357 & ~n2465;
  assign n3324 = n27 & n2356;
  assign n3326 = n3325 ^ n3324;
  assign n3322 = ~n2468 & ~n2746;
  assign n3321 = x0 & ~n2355;
  assign n3323 = n3322 ^ n3321;
  assign n3327 = n3326 ^ n3323;
  assign n3328 = n3327 ^ n2476;
  assign n3330 = n3329 ^ n3328;
  assign n3334 = x1 & n2358;
  assign n3333 = n1387 & n2359;
  assign n3335 = n3334 ^ n3333;
  assign n3331 = n25 & ~n2493;
  assign n3332 = n3331 ^ n2357;
  assign n3336 = n3335 ^ n3332;
  assign n3337 = ~x0 & ~n3336;
  assign n3338 = n3337 ^ n3332;
  assign n3339 = n3338 ^ n2476;
  assign n3340 = n3173 ^ n3109;
  assign n3341 = n25 & ~n2495;
  assign n3342 = n3341 ^ n2356;
  assign n3343 = x0 & n3342;
  assign n3345 = n2358 & ~n2465;
  assign n3344 = n27 & ~n2357;
  assign n3346 = n3345 ^ n3344;
  assign n3347 = ~n3343 & ~n3346;
  assign n3348 = n3347 ^ n3338;
  assign n3349 = ~n3340 & n3348;
  assign n3350 = n3339 & n3349;
  assign n3351 = n3350 ^ n3339;
  assign n3352 = n3170 ^ n3126;
  assign n3361 = n3167 ^ n3157;
  assign n3353 = n25 & ~n2576;
  assign n3354 = n3353 ^ n2358;
  assign n3355 = x0 & n3354;
  assign n3357 = ~n2360 & ~n2465;
  assign n3356 = n27 & n2359;
  assign n3358 = n3357 ^ n3356;
  assign n3359 = ~n3355 & ~n3358;
  assign n3360 = n3359 ^ n2476;
  assign n3362 = n3361 ^ n3360;
  assign n3375 = ~n2468 & ~n2606;
  assign n3371 = n2361 & ~n2465;
  assign n3239 = n2468 ^ x0;
  assign n3370 = n2359 & ~n3239;
  assign n3372 = n3371 ^ n3370;
  assign n3369 = n27 & ~n2360;
  assign n3373 = n3372 ^ n3369;
  assign n3374 = n3373 ^ n2476;
  assign n3376 = n3375 ^ n3374;
  assign n3364 = n3152 ^ n1283;
  assign n3365 = n3364 ^ n3138;
  assign n3363 = n3153 ^ n1163;
  assign n3366 = n3365 ^ n3363;
  assign n3367 = n2365 & n3366;
  assign n3368 = n3367 ^ n3363;
  assign n3377 = n3376 ^ n3368;
  assign n3398 = ~n1337 & ~n2476;
  assign n3402 = n3398 ^ n2476;
  assign n3400 = n2958 ^ n1337;
  assign n3399 = n3398 ^ n1393;
  assign n3401 = n3400 ^ n3399;
  assign n3403 = n3402 ^ n3401;
  assign n3404 = ~n2365 & ~n3403;
  assign n3378 = n2368 & ~n2942;
  assign n3405 = n3404 ^ n3378;
  assign n3382 = n25 & ~n2507;
  assign n3383 = n3382 ^ n2362;
  assign n3384 = x0 & ~n3383;
  assign n3386 = n2368 & ~n2465;
  assign n3385 = n27 & ~n2364;
  assign n3387 = n3386 ^ n3385;
  assign n3388 = ~n3384 & ~n3387;
  assign n3394 = ~n2365 & n2957;
  assign n3389 = ~n2208 & n2364;
  assign n3390 = n3389 ^ n1393;
  assign n3391 = n2365 & n3390;
  assign n3392 = n3391 ^ n1393;
  assign n3393 = n2476 & n3392;
  assign n3395 = n3394 ^ n3393;
  assign n3396 = ~n3388 & n3395;
  assign n3397 = n3396 ^ n3393;
  assign n3406 = n3405 ^ n3397;
  assign n3412 = n2361 & ~n3239;
  assign n3413 = n3412 ^ x0;
  assign n3410 = n2364 & ~n2465;
  assign n3409 = n27 & n2362;
  assign n3411 = n3410 ^ n3409;
  assign n3414 = n3413 ^ n3411;
  assign n3415 = n3414 ^ n2475;
  assign n3407 = n2550 ^ n2361;
  assign n3408 = ~n2468 & ~n3407;
  assign n3416 = n3415 ^ n3408;
  assign n3417 = n3416 ^ n3405;
  assign n3418 = n3406 & n3417;
  assign n3419 = n3418 ^ n3397;
  assign n3379 = n2365 & ~n3378;
  assign n3380 = n2989 & ~n3379;
  assign n3381 = n3380 ^ n3151;
  assign n3420 = n3419 ^ n3381;
  assign n3425 = ~n2362 & ~n2465;
  assign n3424 = ~n2360 & ~n3239;
  assign n3426 = n3425 ^ n3424;
  assign n3423 = n27 & n2361;
  assign n3427 = n3426 ^ n3423;
  assign n3428 = n3427 ^ n2476;
  assign n3421 = n2563 ^ n2360;
  assign n3422 = ~n2468 & n3421;
  assign n3429 = n3428 ^ n3422;
  assign n3430 = n3429 ^ n3381;
  assign n3431 = ~n3420 & n3430;
  assign n3432 = n3431 ^ n3419;
  assign n3433 = n3432 ^ n3368;
  assign n3434 = ~n3377 & n3433;
  assign n3435 = n3434 ^ n3376;
  assign n3436 = n3435 ^ n3361;
  assign n3437 = ~n3362 & ~n3436;
  assign n3438 = n3437 ^ n3360;
  assign n3440 = ~n3352 & n3438;
  assign n3439 = n3438 ^ n3352;
  assign n3441 = n3440 ^ n3439;
  assign n3442 = n3351 & ~n3441;
  assign n3443 = n3347 ^ n2476;
  assign n3444 = n3443 ^ n3340;
  assign n3445 = n3443 ^ n3440;
  assign n3446 = n3444 & ~n3445;
  assign n3447 = n3446 ^ n3340;
  assign n3448 = ~n3442 & ~n3447;
  assign n3449 = n3448 ^ n3329;
  assign n3450 = ~n3330 & n3449;
  assign n3451 = n3450 ^ n3328;
  assign n3452 = n3451 ^ n3319;
  assign n3453 = ~n3320 & n3452;
  assign n3454 = n3453 ^ n3318;
  assign n3455 = n3454 ^ n3296;
  assign n3456 = ~n3309 & ~n3455;
  assign n3457 = n3456 ^ n3308;
  assign n3292 = ~x0 & n2346;
  assign n2941 = n2940 ^ n2346;
  assign n3290 = n2941 ^ n2469;
  assign n3291 = n2940 & n3290;
  assign n3293 = n3292 ^ n3291;
  assign n3288 = n27 & ~n2314;
  assign n3286 = n2941 ^ n2464;
  assign n3287 = ~n2940 & n3286;
  assign n3289 = n3288 ^ n3287;
  assign n3294 = n3293 ^ n3289;
  assign n3283 = ~n28 & n2407;
  assign n3284 = ~n29 & ~n3283;
  assign n3285 = n3284 ^ n2474;
  assign n3295 = n3294 ^ n3285;
  assign n3458 = n3457 ^ n3295;
  assign n3459 = n3185 ^ n3033;
  assign n3460 = n3459 ^ n3295;
  assign n3461 = n3458 & ~n3460;
  assign n3462 = n3461 ^ n3457;
  assign n3514 = n683 ^ n229;
  assign n3515 = n3514 ^ n427;
  assign n3516 = n2278 & n3515;
  assign n3517 = n2076 & n3516;
  assign n3518 = n676 ^ n433;
  assign n3519 = n3517 & ~n3518;
  assign n3520 = ~n110 & n3519;
  assign n3521 = n281 ^ n166;
  assign n3522 = n3521 ^ n400;
  assign n3523 = n44 & n155;
  assign n3524 = n3523 ^ n2126;
  assign n3525 = ~n3522 & ~n3524;
  assign n3526 = n2135 & n3525;
  assign n3527 = n525 ^ n194;
  assign n3528 = n2232 & n3527;
  assign n3529 = n3526 & n3528;
  assign n3530 = n480 ^ n362;
  assign n3531 = ~n535 & ~n3530;
  assign n3532 = n815 & n3531;
  assign n3533 = n3529 & n3532;
  assign n3534 = n3520 & n3533;
  assign n3535 = ~n3462 & ~n3534;
  assign n3536 = n352 ^ n61;
  assign n3537 = n3536 ^ n378;
  assign n3538 = n352 ^ n125;
  assign n3539 = n3538 ^ n334;
  assign n3540 = ~n3537 & ~n3539;
  assign n3541 = n1182 & ~n3540;
  assign n3474 = n623 ^ n310;
  assign n3475 = n3474 ^ n290;
  assign n3542 = n840 ^ n416;
  assign n3543 = n3475 & ~n3542;
  assign n3544 = ~n473 & n3543;
  assign n3545 = n3541 & n3544;
  assign n3546 = n826 ^ n498;
  assign n3547 = n3546 ^ n196;
  assign n3548 = n3545 & ~n3547;
  assign n3549 = n412 ^ n236;
  assign n3550 = n2329 & ~n3549;
  assign n3551 = ~n990 & n3550;
  assign n3552 = ~n309 & ~n530;
  assign n3553 = n3552 ^ n871;
  assign n3554 = n3551 & ~n3553;
  assign n3555 = ~n2192 & n3554;
  assign n3556 = n467 ^ n166;
  assign n3557 = n363 ^ n227;
  assign n3558 = n3557 ^ n217;
  assign n3559 = ~n3556 & ~n3558;
  assign n3560 = n2237 ^ n715;
  assign n3561 = n3559 & ~n3560;
  assign n3562 = n817 ^ n371;
  assign n3563 = n671 ^ n492;
  assign n3564 = n3563 ^ n304;
  assign n3565 = ~n3562 & n3564;
  assign n3566 = n3561 & n3565;
  assign n3567 = n3555 & n3566;
  assign n3568 = n3548 & n3567;
  assign n3570 = ~n3535 & n3568;
  assign n3569 = n3568 ^ n3535;
  assign n3571 = n3570 ^ n3569;
  assign n3572 = n3571 ^ n3462;
  assign n3573 = ~n3281 & ~n3572;
  assign n3574 = n3573 ^ n3571;
  assign n3575 = ~n3282 & n3574;
  assign n3576 = n3575 ^ n3280;
  assign n3577 = n3269 & ~n3576;
  assign n3578 = ~n3280 & n3568;
  assign n3579 = ~n3269 & ~n3578;
  assign n3580 = n3282 & ~n3535;
  assign n3581 = n3579 & ~n3580;
  assign n3463 = ~n3280 & n3462;
  assign n3582 = n3463 & n3534;
  assign n3583 = n3581 & ~n3582;
  assign n3584 = ~n3577 & ~n3583;
  assign n3585 = ~n3281 & ~n3534;
  assign n3586 = n3570 & ~n3585;
  assign n3587 = ~n3584 & ~n3586;
  assign n3484 = n72 & ~n2071;
  assign n3486 = n565 ^ n175;
  assign n3485 = n657 ^ n191;
  assign n3487 = n3486 ^ n3485;
  assign n3488 = ~n964 & ~n3487;
  assign n3489 = n119 & n156;
  assign n3490 = n3489 ^ n617;
  assign n3491 = n44 & n83;
  assign n3492 = n3491 ^ n484;
  assign n3493 = n3492 ^ n273;
  assign n3494 = ~n3490 & ~n3493;
  assign n3495 = n2074 ^ n299;
  assign n3496 = n3494 & ~n3495;
  assign n3497 = n3488 & n3496;
  assign n3498 = n836 & n3497;
  assign n3499 = ~n3484 & n3498;
  assign n3500 = ~n237 & n712;
  assign n3501 = n618 ^ n174;
  assign n3502 = n3501 ^ n700;
  assign n3503 = n3502 ^ n246;
  assign n3504 = ~n2341 & ~n3503;
  assign n3505 = n746 & n3504;
  assign n3506 = ~n537 & ~n2318;
  assign n3507 = n804 ^ n287;
  assign n3508 = ~n408 & ~n3507;
  assign n3509 = ~n2026 & n3508;
  assign n3510 = n3506 & n3509;
  assign n3511 = n3505 & n3510;
  assign n3512 = n3500 & n3511;
  assign n3513 = n3499 & n3512;
  assign n3588 = n3587 ^ n3513;
  assign n3464 = ~n3282 & ~n3463;
  assign n3465 = n3464 ^ n3254;
  assign n3466 = n3269 & ~n3465;
  assign n3467 = n3466 ^ n3268;
  assign n3216 = n3215 ^ n3191;
  assign n3217 = ~n3192 & n3216;
  assign n3218 = n3217 ^ n3215;
  assign n2916 = n2915 ^ n2762;
  assign n2917 = n2778 & ~n2916;
  assign n2918 = n2917 ^ n2777;
  assign n2758 = ~n2355 & n2719;
  assign n2751 = n2724 & ~n2746;
  assign n2757 = ~n2751 & n2756;
  assign n2759 = n2758 ^ n2757;
  assign n2752 = n959 & n2751;
  assign n2753 = n2752 ^ n2724;
  assign n2750 = n2356 & ~n2724;
  assign n2754 = n2753 ^ n2750;
  assign n2742 = n2741 ^ n2357;
  assign n2748 = n2747 ^ n2742;
  assign n2749 = ~n2739 & n2748;
  assign n2755 = n2754 ^ n2749;
  assign n2760 = n2759 ^ n2755;
  assign n2711 = n2710 ^ n2620;
  assign n2712 = n2621 & ~n2711;
  assign n2713 = n2712 ^ n2614;
  assign n2546 = ~n583 & ~n2365;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = ~n2523 & ~n2547;
  assign n2549 = n2548 ^ n2368;
  assign n2589 = ~n2548 & ~n2549;
  assign n2590 = n583 & n2589;
  assign n2591 = n2590 ^ n2549;
  assign n2551 = n584 & ~n2550;
  assign n2552 = n2551 ^ n2361;
  assign n2553 = n754 & n2552;
  assign n2554 = ~n2362 & n2536;
  assign n2555 = ~n2364 & n2541;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = ~n2553 & n2556;
  assign n2592 = n2591 ^ n2557;
  assign n2573 = n2359 & n2484;
  assign n2574 = ~n2360 & n2490;
  assign n2575 = ~n2573 & ~n2574;
  assign n2579 = n2478 & n2578;
  assign n2577 = n2478 & ~n2576;
  assign n2580 = n2579 ^ n2577;
  assign n2581 = n2575 & ~n2580;
  assign n2582 = ~n753 & ~n2581;
  assign n2583 = n753 & n2575;
  assign n2584 = ~n2579 & n2583;
  assign n2585 = n2358 ^ n792;
  assign n2586 = n2577 & n2585;
  assign n2587 = ~n2584 & ~n2586;
  assign n2588 = ~n2582 & n2587;
  assign n2593 = n2592 ^ n2588;
  assign n2718 = n2713 ^ n2593;
  assign n2761 = n2760 ^ n2718;
  assign n2980 = n2918 ^ n2761;
  assign n2950 = ~n2346 & ~n2949;
  assign n2951 = n2950 ^ n1283;
  assign n2952 = ~n2942 & n2951;
  assign n2945 = n2940 & ~n2944;
  assign n2953 = n2952 ^ n2945;
  assign n2954 = ~n2941 & n2953;
  assign n2955 = n2954 ^ n2952;
  assign n2973 = n2972 ^ n2387;
  assign n2974 = n2973 ^ n2407;
  assign n2975 = ~n2971 & ~n2974;
  assign n2965 = n2407 & ~n2962;
  assign n2966 = n2962 ^ n1283;
  assign n2967 = n2966 ^ n2407;
  assign n2968 = ~n2965 & n2967;
  assign n2976 = n2975 ^ n2968;
  assign n2964 = n2407 & ~n2959;
  assign n2977 = n2976 ^ n2964;
  assign n2963 = n2314 & n2962;
  assign n2978 = n2977 ^ n2963;
  assign n2979 = ~n2955 & n2978;
  assign n2981 = n2980 ^ n2979;
  assign n3252 = n3218 ^ n2981;
  assign n3248 = n2465 ^ n2457;
  assign n3247 = n27 & ~n2447;
  assign n3249 = n3248 ^ n3247;
  assign n2425 = n235 & ~n2349;
  assign n2426 = ~n2424 & n2425;
  assign n2390 = n2389 ^ n2349;
  assign n2391 = n235 & ~n2390;
  assign n2392 = n2391 ^ n2389;
  assign n3243 = n2426 ^ n2392;
  assign n2393 = n162 & ~n250;
  assign n2394 = n502 ^ n83;
  assign n2395 = n57 & n2394;
  assign n2396 = ~n273 & ~n2395;
  assign n2397 = ~n420 & n2396;
  assign n2398 = n448 ^ n259;
  assign n2399 = n2398 ^ n515;
  assign n2400 = n147 & n2399;
  assign n2401 = ~n2130 & ~n2400;
  assign n2402 = n2397 & n2401;
  assign n2403 = n548 & n2402;
  assign n2404 = n2393 & n2403;
  assign n2427 = n2425 ^ n235;
  assign n2428 = ~n2404 & ~n2427;
  assign n3244 = n3243 ^ n2428;
  assign n3245 = ~n2468 & ~n3244;
  assign n3246 = n3245 ^ n2470;
  assign n3250 = n3249 ^ n3246;
  assign n3240 = n2428 & ~n3239;
  assign n3241 = n3240 ^ n2473;
  assign n3238 = ~n2465 & n3225;
  assign n3242 = n3241 ^ n3238;
  assign n3251 = n3250 ^ n3242;
  assign n3253 = n3252 ^ n3251;
  assign n3589 = n3467 ^ n3253;
  assign n3590 = n3589 ^ n3513;
  assign n3591 = ~n3588 & ~n3590;
  assign n3592 = n3591 ^ n3590;
  assign n3472 = n2237 ^ n450;
  assign n3473 = ~n252 & ~n3472;
  assign n3476 = n3475 ^ n519;
  assign n3477 = n3473 & n3476;
  assign n3478 = n2044 & n2320;
  assign n3479 = n3477 & n3478;
  assign n3480 = n680 & n3479;
  assign n3481 = n2071 & n3480;
  assign n3482 = n622 & n3481;
  assign n3468 = n3467 ^ n3251;
  assign n3469 = n3253 & n3468;
  assign n3470 = n3469 ^ n3467;
  assign n3223 = n2949 & ~n2972;
  assign n3224 = n3223 ^ n1283;
  assign n3226 = n3225 ^ n3224;
  assign n3227 = ~n2942 & n3226;
  assign n3228 = n2314 & n2995;
  assign n3229 = n3228 ^ n2314;
  assign n3230 = n3002 & n3229;
  assign n3231 = n3230 ^ n2959;
  assign n3232 = n2346 & n2999;
  assign n3233 = n3232 ^ n2997;
  assign n3234 = ~n3231 & ~n3233;
  assign n3235 = ~n3227 & n3234;
  assign n3219 = n3218 ^ n2979;
  assign n3220 = n2981 & n3219;
  assign n3221 = n3220 ^ n3218;
  assign n2930 = n2740 ^ n2356;
  assign n2931 = ~n2739 & ~n2930;
  assign n2923 = n2724 & n2740;
  assign n2929 = ~n2725 & ~n2923;
  assign n2932 = n2931 ^ n2929;
  assign n2928 = ~n2355 & ~n2724;
  assign n2933 = n2932 ^ n2928;
  assign n2926 = n2407 & n2719;
  assign n2924 = ~n955 & n2923;
  assign n2925 = n2924 ^ n2730;
  assign n2927 = n2926 ^ n2925;
  assign n2934 = n2933 ^ n2927;
  assign n2919 = n2918 ^ n2760;
  assign n2920 = n2761 & n2919;
  assign n2921 = n2920 ^ n2918;
  assign n2714 = n2713 ^ n2592;
  assign n2715 = ~n2593 & ~n2714;
  assign n2716 = n2715 ^ n2588;
  assign n2564 = n584 & ~n2563;
  assign n2565 = n2564 ^ n2360;
  assign n2566 = n754 & ~n2565;
  assign n2567 = n2361 & n2536;
  assign n2568 = ~n2362 & n2541;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = ~n2566 & n2569;
  assign n2558 = n2557 ^ n2548;
  assign n2559 = n2549 & ~n2558;
  assign n2560 = n2559 ^ n2368;
  assign n2561 = n2560 ^ n2364;
  assign n2562 = ~n583 & n2561;
  assign n2571 = n2570 ^ n2562;
  assign n2485 = n2358 & n2484;
  assign n2491 = n2359 & n2490;
  assign n2492 = ~n2485 & ~n2491;
  assign n2497 = n2478 & n2496;
  assign n2494 = n2478 & ~n2493;
  assign n2498 = n2497 ^ n2494;
  assign n2499 = n2492 & ~n2498;
  assign n2500 = ~n753 & ~n2499;
  assign n2501 = n753 & n2492;
  assign n2502 = ~n2497 & n2501;
  assign n2503 = n2357 ^ n792;
  assign n2504 = n2494 & ~n2503;
  assign n2505 = ~n2502 & ~n2504;
  assign n2506 = ~n2500 & n2505;
  assign n2572 = n2571 ^ n2506;
  assign n2717 = n2716 ^ n2572;
  assign n2922 = n2921 ^ n2717;
  assign n2935 = n2934 ^ n2922;
  assign n3222 = n3221 ^ n2935;
  assign n3236 = n3235 ^ n3222;
  assign n2448 = n1387 & ~n2447;
  assign n2446 = x1 & n2428;
  assign n2449 = n2448 ^ n2446;
  assign n2432 = n809 ^ n642;
  assign n2433 = ~n61 & n2432;
  assign n2434 = n276 ^ n251;
  assign n2435 = n2434 ^ n373;
  assign n2436 = ~n2433 & ~n2435;
  assign n2437 = n840 ^ n325;
  assign n2438 = n2436 & ~n2437;
  assign n2439 = n117 & n2399;
  assign n2440 = n604 ^ n401;
  assign n2441 = n2440 ^ n298;
  assign n2442 = ~n2439 & ~n2441;
  assign n2443 = n2438 & n2442;
  assign n2444 = n1201 & n2443;
  assign n2429 = ~n2426 & n2428;
  assign n2405 = n2392 & n2404;
  assign n2430 = n2429 ^ n2405;
  assign n2431 = n25 & ~n2430;
  assign n2445 = n2444 ^ n2431;
  assign n2450 = n2449 ^ n2445;
  assign n2451 = ~x0 & ~n2450;
  assign n2452 = n2451 ^ n2445;
  assign n2477 = n2476 ^ n2452;
  assign n3237 = n3236 ^ n2477;
  assign n3471 = n3470 ^ n3237;
  assign n3483 = n3482 ^ n3471;
  assign n3593 = n3592 ^ n3483;
  assign n3747 = x23 ^ x22;
  assign n3743 = ~n3589 & ~n3592;
  assign n3753 = n3747 ^ n3743;
  assign n3754 = n3743 ^ n3483;
  assign n3755 = ~n3753 & ~n3754;
  assign n3751 = n3471 & n3482;
  assign n3752 = n3751 ^ n3483;
  assign n3756 = n3755 ^ n3752;
  assign n3744 = n3743 ^ n3592;
  assign n3748 = ~n3744 & n3747;
  assign n3745 = n3483 & n3744;
  assign n3746 = n3745 ^ n3483;
  assign n3749 = n3748 ^ n3746;
  assign n3722 = n533 ^ n362;
  assign n3723 = n3722 ^ n383;
  assign n3721 = n840 ^ n693;
  assign n3724 = n3723 ^ n3721;
  assign n3725 = ~n2318 & ~n3724;
  assign n3727 = n3514 ^ n342;
  assign n3726 = ~n61 & n2335;
  assign n3728 = n3727 ^ n3726;
  assign n3729 = n3725 & ~n3728;
  assign n3730 = n2060 & n3729;
  assign n3731 = ~n674 & ~n838;
  assign n3732 = n412 ^ n301;
  assign n3733 = n3731 & ~n3732;
  assign n3734 = n3730 & n3733;
  assign n3735 = n3497 & n3734;
  assign n3598 = n281 ^ n268;
  assign n3599 = n3598 ^ n329;
  assign n3736 = n3599 ^ n220;
  assign n3737 = n3506 & n3736;
  assign n3738 = n2048 & ~n3737;
  assign n3739 = n453 ^ n84;
  assign n3740 = ~n3738 & ~n3739;
  assign n3741 = n3735 & n3740;
  assign n3717 = n3470 ^ n2477;
  assign n3718 = n3237 & ~n3717;
  assign n3719 = n3718 ^ n3470;
  assign n3712 = n3235 ^ n2935;
  assign n3713 = n3222 & ~n3712;
  assign n3714 = n3713 ^ n3221;
  assign n3707 = n3258 ^ n2346;
  assign n3708 = n2993 & n3707;
  assign n3703 = n2447 ^ n1337;
  assign n3704 = ~n2962 & n3258;
  assign n3705 = n3704 ^ n2942;
  assign n3706 = ~n3703 & ~n3705;
  assign n3709 = n3708 ^ n3706;
  assign n3700 = n3225 ^ n1283;
  assign n3696 = n1283 & n3258;
  assign n3694 = n2424 ^ n2349;
  assign n3695 = n3694 ^ n3243;
  assign n3697 = n3696 ^ n3695;
  assign n3698 = n3697 ^ n3225;
  assign n3699 = ~n2962 & ~n3698;
  assign n3701 = n3700 ^ n3699;
  assign n3702 = n3701 ^ n2970;
  assign n3710 = n3709 ^ n3702;
  assign n3690 = n2934 ^ n2921;
  assign n3691 = n2922 & ~n3690;
  assign n3692 = n3691 ^ n2934;
  assign n3685 = n2716 ^ n2571;
  assign n3686 = n2572 & ~n3685;
  assign n3687 = n3686 ^ n2506;
  assign n3666 = n555 & ~n2360;
  assign n3665 = n2361 & n2511;
  assign n3667 = n3666 ^ n3665;
  assign n3668 = ~n751 & n3667;
  assign n3669 = n3668 ^ n3666;
  assign n3663 = n584 & ~n2594;
  assign n3664 = n3663 ^ n2359;
  assign n3670 = n3669 ^ n3664;
  assign n3671 = n3670 ^ n3664;
  assign n3672 = n583 & n2361;
  assign n3673 = n3672 ^ n2360;
  assign n3674 = n753 & ~n3673;
  assign n3675 = n3674 ^ n2360;
  assign n3676 = ~n555 & ~n3675;
  assign n3677 = n3676 ^ n3664;
  assign n3678 = n3677 ^ n3664;
  assign n3679 = ~n3671 & ~n3678;
  assign n3680 = n3679 ^ n3664;
  assign n3681 = ~n754 & ~n3680;
  assign n3682 = n3681 ^ n3664;
  assign n3657 = n2570 ^ n2364;
  assign n3658 = ~n2561 & ~n3657;
  assign n3659 = n3658 ^ n2364;
  assign n3660 = ~n583 & ~n3659;
  assign n3661 = n3660 ^ n2362;
  assign n3662 = ~n583 & n3661;
  assign n3683 = n3682 ^ n3662;
  assign n3639 = n2356 ^ n792;
  assign n3640 = n2478 & ~n2495;
  assign n3641 = ~n3639 & n3640;
  assign n3642 = ~n2357 & n2484;
  assign n3643 = n2358 & n2490;
  assign n3644 = ~n3642 & ~n3643;
  assign n3645 = n3644 ^ n753;
  assign n3646 = n2478 & n2745;
  assign n3647 = n3646 ^ n3644;
  assign n3648 = n2604 & ~n2744;
  assign n3649 = n3648 ^ n3646;
  assign n3650 = n3647 & n3649;
  assign n3651 = n3650 ^ n3648;
  assign n3652 = n3651 ^ n3646;
  assign n3653 = n3652 ^ n3648;
  assign n3654 = n3645 & ~n3653;
  assign n3655 = n3654 ^ n3648;
  assign n3656 = ~n3641 & ~n3655;
  assign n3684 = n3683 ^ n3656;
  assign n3688 = n3687 ^ n3684;
  assign n3625 = n2719 & ~n3210;
  assign n3627 = ~n2355 & ~n2739;
  assign n3626 = n2407 & ~n2724;
  assign n3628 = n3627 ^ n3626;
  assign n3629 = ~n3625 & ~n3628;
  assign n3630 = ~n955 & ~n3629;
  assign n3631 = n2719 & ~n3209;
  assign n3632 = n955 & ~n3628;
  assign n3633 = ~n3631 & n3632;
  assign n3634 = n2314 ^ n959;
  assign n3635 = n2719 & n3634;
  assign n3636 = n2938 & n3635;
  assign n3637 = ~n3633 & ~n3636;
  assign n3638 = ~n3630 & n3637;
  assign n3689 = n3688 ^ n3638;
  assign n3693 = n3692 ^ n3689;
  assign n3711 = n3710 ^ n3693;
  assign n3715 = n3714 ^ n3711;
  assign n3619 = x1 & ~n2444;
  assign n3618 = n1387 & n2428;
  assign n3620 = n3619 ^ n3618;
  assign n3600 = n137 ^ n125;
  assign n3601 = n3600 ^ n208;
  assign n3602 = n118 & n3601;
  assign n3603 = n3599 & ~n3602;
  assign n3604 = n1409 & n3603;
  assign n3605 = n593 ^ n372;
  assign n3606 = n3604 & ~n3605;
  assign n3607 = n796 ^ n261;
  assign n3608 = ~n76 & n3607;
  assign n3609 = ~n567 & ~n3608;
  assign n3610 = n2282 ^ n319;
  assign n3611 = n3610 ^ n246;
  assign n3612 = ~n838 & ~n3611;
  assign n3613 = n3609 & n3612;
  assign n3614 = n816 & n3613;
  assign n3615 = n3606 & n3614;
  assign n3616 = n2253 & n3615;
  assign n3595 = ~n2429 & n2444;
  assign n3594 = ~n2405 & ~n2444;
  assign n3596 = n3595 ^ n3594;
  assign n3597 = n25 & ~n3596;
  assign n3617 = n3616 ^ n3597;
  assign n3621 = n3620 ^ n3617;
  assign n3622 = ~x0 & ~n3621;
  assign n3623 = n3622 ^ n3617;
  assign n3624 = n3623 ^ n2476;
  assign n3716 = n3715 ^ n3624;
  assign n3720 = n3719 ^ n3716;
  assign n3742 = n3741 ^ n3720;
  assign n3750 = n3749 ^ n3742;
  assign n3757 = n3756 ^ n3750;
  assign n3886 = ~n76 & n609;
  assign n3887 = n3886 ^ n285;
  assign n3888 = n3887 ^ n227;
  assign n3885 = n498 ^ n304;
  assign n3889 = n3888 ^ n3885;
  assign n3890 = n628 ^ n274;
  assign n3891 = n3890 ^ n342;
  assign n3892 = ~n3889 & ~n3891;
  assign n3893 = n560 ^ n405;
  assign n3894 = n287 ^ n166;
  assign n3895 = n3894 ^ n870;
  assign n3896 = n3895 ^ n657;
  assign n3897 = n3896 ^ n519;
  assign n3898 = ~n3893 & ~n3897;
  assign n3899 = n3892 & n3898;
  assign n3900 = n808 & n3899;
  assign n3901 = n3520 & n3900;
  assign n3881 = n3719 ^ n3624;
  assign n3882 = n3716 & ~n3881;
  assign n3883 = n3882 ^ n3719;
  assign n3876 = n3714 ^ n3710;
  assign n3877 = ~n3711 & ~n3876;
  assign n3878 = n3877 ^ n3714;
  assign n3872 = n3692 ^ n3688;
  assign n3873 = n3689 & ~n3872;
  assign n3874 = n3873 ^ n3638;
  assign n3867 = n3687 ^ n3683;
  assign n3868 = n3684 & n3867;
  assign n3869 = n3868 ^ n3656;
  assign n3858 = n584 & ~n2576;
  assign n3859 = n3858 ^ n2358;
  assign n3860 = n754 & n3859;
  assign n3861 = n2359 & n2536;
  assign n3862 = ~n2360 & n2541;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = ~n3860 & n3863;
  assign n3853 = n3682 ^ n3660;
  assign n3854 = ~n3661 & n3853;
  assign n3855 = n3854 ^ n2362;
  assign n3856 = n3855 ^ n2361;
  assign n3857 = ~n583 & n3856;
  assign n3865 = n3864 ^ n3857;
  assign n3839 = n2355 ^ n792;
  assign n3840 = n2478 & ~n2746;
  assign n3841 = n3839 & n3840;
  assign n3842 = n2356 & n2484;
  assign n3843 = ~n2357 & n2490;
  assign n3844 = ~n3842 & ~n3843;
  assign n3845 = n3844 ^ n753;
  assign n3847 = n2478 & n2747;
  assign n3848 = ~n753 & n3847;
  assign n3846 = n2604 & ~n2741;
  assign n3849 = n3848 ^ n3846;
  assign n3850 = n3845 & ~n3849;
  assign n3851 = n3850 ^ n3846;
  assign n3852 = ~n3841 & ~n3851;
  assign n3866 = n3865 ^ n3852;
  assign n3870 = n3869 ^ n3866;
  assign n3821 = ~n960 & n2940;
  assign n3822 = n3821 ^ n955;
  assign n3823 = n3822 ^ n2346;
  assign n3824 = n2719 & n3823;
  assign n3834 = ~n2407 & ~n2739;
  assign n3835 = n3834 ^ n959;
  assign n3831 = n955 & n2314;
  assign n3832 = n2722 & ~n3831;
  assign n3833 = ~n3127 & ~n3832;
  assign n3836 = n3835 ^ n3833;
  assign n3826 = n2314 & ~n2723;
  assign n3827 = n3826 ^ n2732;
  assign n3828 = n2314 ^ n960;
  assign n3829 = n3827 & ~n3828;
  assign n3825 = ~n2314 & ~n2735;
  assign n3830 = n3829 ^ n3825;
  assign n3837 = n3836 ^ n3830;
  assign n3838 = ~n3824 & n3837;
  assign n3871 = n3870 ^ n3838;
  assign n3875 = n3874 ^ n3871;
  assign n3879 = n3878 ^ n3875;
  assign n3805 = n3616 ^ n1385;
  assign n3806 = x1 & n3805;
  assign n3812 = x22 ^ x1;
  assign n3808 = n3596 & n3616;
  assign n3809 = n3808 ^ n3596;
  assign n3810 = n3809 ^ n3594;
  assign n3811 = n25 & ~n3810;
  assign n3813 = n3812 ^ n3811;
  assign n3807 = n1387 & n2444;
  assign n3814 = n3813 ^ n3807;
  assign n3815 = n3814 ^ n3813;
  assign n3816 = ~n3806 & ~n3815;
  assign n3817 = n3816 ^ n3813;
  assign n3818 = ~x0 & n3817;
  assign n3819 = n3818 ^ n3813;
  assign n3780 = n1337 & n3243;
  assign n3781 = n2428 & ~n3780;
  assign n3782 = n1283 & ~n3225;
  assign n3783 = n3782 ^ n2447;
  assign n3784 = ~n1337 & ~n3783;
  assign n3785 = n3784 ^ n2447;
  assign n3786 = ~n2958 & ~n3785;
  assign n3788 = n2996 & ~n3225;
  assign n3787 = ~n2447 & ~n2960;
  assign n3789 = n3788 ^ n3787;
  assign n3790 = ~n3786 & ~n3789;
  assign n3791 = n3243 & n3790;
  assign n3792 = n3791 ^ n2942;
  assign n3793 = n1283 & ~n3792;
  assign n3794 = n3793 ^ n2942;
  assign n3795 = n3781 & ~n3794;
  assign n3796 = n2430 ^ n2392;
  assign n3797 = n3796 ^ n3244;
  assign n3799 = n3797 ^ n2428;
  assign n3800 = n1283 & ~n3799;
  assign n3801 = ~n2969 & ~n3800;
  assign n3802 = n3801 ^ n3790;
  assign n3798 = ~n2944 & n3797;
  assign n3803 = n3802 ^ n3798;
  assign n3804 = ~n3795 & ~n3803;
  assign n3820 = n3819 ^ n3804;
  assign n3880 = n3879 ^ n3820;
  assign n3884 = n3883 ^ n3880;
  assign n3902 = n3901 ^ n3884;
  assign n3758 = n3591 ^ n3587;
  assign n3768 = n3745 & ~n3758;
  assign n3775 = n3768 ^ n3751;
  assign n3776 = n3775 ^ n3746;
  assign n3777 = n3776 ^ n3741;
  assign n3778 = n3742 & ~n3777;
  assign n3779 = n3778 ^ n3720;
  assign n3903 = n3902 ^ n3779;
  assign n3763 = ~n3483 & ~n3742;
  assign n3759 = ~n3751 & n3758;
  assign n3770 = n3763 ^ n3759;
  assign n3771 = n3743 & ~n3770;
  assign n3769 = n3742 & n3768;
  assign n3772 = n3771 ^ n3769;
  assign n3773 = ~n3747 & ~n3772;
  assign n3764 = n3763 ^ n3752;
  assign n3765 = ~n3744 & ~n3764;
  assign n3760 = ~n3743 & n3759;
  assign n3761 = n3742 & n3760;
  assign n3762 = n3752 & n3761;
  assign n3766 = n3765 ^ n3762;
  assign n3767 = n3747 & n3766;
  assign n3774 = n3773 ^ n3767;
  assign n3904 = n3903 ^ n3774;
  assign n4034 = n3732 ^ n377;
  assign n4035 = n419 ^ n251;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = n533 ^ n400;
  assign n4038 = n4037 ^ n402;
  assign n4039 = ~n1070 & ~n4038;
  assign n4040 = n4036 & n4039;
  assign n4041 = n1988 & n4040;
  assign n4042 = n452 & n3565;
  assign n4043 = n863 & n4042;
  assign n4044 = n4041 & n4043;
  assign n4045 = n1396 & n4044;
  assign n4027 = n3595 & ~n3616;
  assign n4028 = ~n2465 & n4027;
  assign n4029 = n4028 ^ n2465;
  assign n4030 = n4029 ^ n2457;
  assign n4023 = n25 & ~n3616;
  assign n4024 = ~n3595 & n4023;
  assign n4025 = ~n2466 & ~n4024;
  assign n4026 = n4025 ^ n2471;
  assign n4031 = n4030 ^ n4026;
  assign n4018 = n3874 ^ n3838;
  assign n4019 = ~n3871 & n4018;
  assign n4020 = n4019 ^ n3874;
  assign n4012 = n3869 ^ n3865;
  assign n4013 = ~n3866 & n4012;
  assign n4014 = n4013 ^ n3852;
  assign n4006 = n3864 ^ n2361;
  assign n4007 = ~n3856 & n4006;
  assign n4008 = n4007 ^ n2361;
  assign n4009 = n4008 ^ n2360;
  assign n4010 = ~n583 & n4009;
  assign n3999 = n584 & ~n2493;
  assign n4000 = n3999 ^ n2357;
  assign n4001 = n754 & ~n4000;
  assign n4002 = n2358 & n2536;
  assign n4003 = n2359 & n2541;
  assign n4004 = ~n4002 & ~n4003;
  assign n4005 = ~n4001 & n4004;
  assign n4011 = n4010 ^ n4005;
  assign n4015 = n4014 ^ n4011;
  assign n3984 = n2478 & n2937;
  assign n3985 = ~n2355 & n2484;
  assign n3986 = n2356 & n2490;
  assign n3987 = ~n3985 & ~n3986;
  assign n3988 = ~n3984 & n3987;
  assign n3989 = ~n753 & ~n3988;
  assign n3990 = n2938 ^ n2378;
  assign n3991 = n2478 & ~n3990;
  assign n3992 = n753 & n3987;
  assign n3993 = ~n3991 & n3992;
  assign n3994 = ~n2407 & n2478;
  assign n3995 = n3994 ^ n2480;
  assign n3996 = ~n2740 & n3995;
  assign n3997 = ~n3993 & ~n3996;
  assign n3998 = ~n3989 & n3997;
  assign n4016 = n4015 ^ n3998;
  assign n3966 = ~n960 & ~n2972;
  assign n3967 = n3966 ^ n955;
  assign n3968 = n3967 ^ n3225;
  assign n3969 = n2719 & n3968;
  assign n3970 = ~n2346 & n2732;
  assign n3974 = n2346 ^ n955;
  assign n3975 = n3974 ^ n3831;
  assign n3976 = n1163 & n3975;
  assign n3977 = n3976 ^ n3831;
  assign n3978 = ~n2719 & ~n3977;
  assign n3972 = n2314 & n2736;
  assign n3971 = n2346 & ~n2733;
  assign n3973 = n3972 ^ n3971;
  assign n3979 = n3978 ^ n3973;
  assign n3980 = ~n959 & n3979;
  assign n3981 = n3980 ^ n3978;
  assign n3982 = ~n3970 & ~n3981;
  assign n3983 = ~n3969 & n3982;
  assign n4017 = n4016 ^ n3983;
  assign n4021 = n4020 ^ n4017;
  assign n3938 = n1337 & ~n2430;
  assign n3939 = n2444 & ~n3938;
  assign n3941 = n2447 ^ n2428;
  assign n3942 = n1337 & ~n3941;
  assign n3943 = n3942 ^ n2447;
  assign n3944 = n2995 ^ n2958;
  assign n3945 = ~n3943 & ~n3944;
  assign n3947 = ~n2447 & n2996;
  assign n3946 = n2428 & ~n2960;
  assign n3948 = n3947 ^ n3946;
  assign n3949 = ~n3945 & ~n3948;
  assign n3940 = ~n2430 & ~n2942;
  assign n3950 = n3949 ^ n3940;
  assign n3951 = n1283 & n3950;
  assign n3952 = n3951 ^ n3949;
  assign n3953 = n3939 & n3952;
  assign n3954 = ~n2444 & ~n2944;
  assign n3955 = ~n2430 & n3954;
  assign n3956 = n1283 & ~n3949;
  assign n3957 = ~n3955 & ~n3956;
  assign n3958 = ~n3953 & n3957;
  assign n3959 = n2942 ^ n1283;
  assign n3960 = n3596 ^ n2429;
  assign n3961 = n3960 ^ n3949;
  assign n3962 = n2942 & ~n3961;
  assign n3963 = n3962 ^ n3960;
  assign n3964 = n3959 & ~n3963;
  assign n3965 = n3958 & ~n3964;
  assign n4022 = n4021 ^ n3965;
  assign n4032 = n4031 ^ n4022;
  assign n3922 = n3883 ^ n3819;
  assign n3923 = ~n3820 & ~n3922;
  assign n3924 = n3923 ^ n3883;
  assign n3925 = n3875 & ~n3878;
  assign n3926 = n3925 ^ n3879;
  assign n3927 = n3924 & n3926;
  assign n3928 = ~n3804 & ~n3819;
  assign n3929 = n3928 ^ n3820;
  assign n3930 = ~n3926 & ~n3929;
  assign n3931 = ~n3883 & n3930;
  assign n3932 = n3883 & n3928;
  assign n3933 = n3932 ^ n3924;
  assign n3934 = n3925 & ~n3933;
  assign n3935 = n3934 ^ n3932;
  assign n3936 = ~n3931 & ~n3935;
  assign n3937 = ~n3927 & n3936;
  assign n4033 = n4032 ^ n3937;
  assign n4046 = n4045 ^ n4033;
  assign n3905 = n3884 ^ n3779;
  assign n3906 = ~n3902 & n3905;
  assign n3907 = n3906 ^ n3779;
  assign n3908 = n3903 & n3907;
  assign n3909 = n3908 ^ n3907;
  assign n3910 = n3909 ^ n3903;
  assign n3911 = ~n3773 & ~n3910;
  assign n3913 = ~n3747 & n3907;
  assign n3912 = n3907 ^ n3747;
  assign n3914 = n3913 ^ n3912;
  assign n3915 = n3914 ^ n3908;
  assign n3916 = ~n3766 & n3915;
  assign n3917 = n3916 ^ n3908;
  assign n3918 = ~n3911 & ~n3917;
  assign n3919 = n3772 & ~n3908;
  assign n3920 = n3913 & ~n3919;
  assign n3921 = n3918 & ~n3920;
  assign n4047 = n4046 ^ n3921;
  assign n4064 = n520 ^ n365;
  assign n4065 = n1065 ^ n491;
  assign n4066 = ~n4064 & n4065;
  assign n4067 = n291 ^ n277;
  assign n4068 = ~n664 & ~n4067;
  assign n4069 = n4066 & n4068;
  assign n4070 = n997 & n4069;
  assign n4071 = n2193 & n4070;
  assign n4072 = n890 & n4071;
  assign n4159 = n4031 ^ n3965;
  assign n4160 = n4022 & ~n4159;
  assign n4161 = n4160 ^ n4031;
  assign n4156 = ~n2971 & ~n3596;
  assign n4149 = n2942 ^ n2444;
  assign n4150 = n4149 ^ n3596;
  assign n4151 = ~n2942 & ~n4150;
  assign n4152 = n4151 ^ n4149;
  assign n4153 = ~n1337 & n4152;
  assign n4154 = n4153 ^ n4149;
  assign n4148 = ~n2942 & n3616;
  assign n4155 = n4154 ^ n4148;
  assign n4157 = n4156 ^ n4155;
  assign n4143 = n1283 & n2428;
  assign n4144 = n4143 ^ n2444;
  assign n4145 = n2959 & ~n4144;
  assign n4142 = n2444 ^ n1283;
  assign n4146 = n4145 ^ n4142;
  assign n4140 = n2428 & n2996;
  assign n4139 = ~n2444 & ~n2961;
  assign n4141 = n4140 ^ n4139;
  assign n4147 = n4146 ^ n4141;
  assign n4158 = n4157 ^ n4147;
  assign n4166 = n4161 ^ n4158;
  assign n4162 = ~n4158 & ~n4161;
  assign n4167 = n4166 ^ n4162;
  assign n4133 = n2739 & ~n3707;
  assign n4134 = n4133 ^ n2346;
  assign n4125 = n2724 & ~n3258;
  assign n4131 = n959 & n4125;
  assign n4132 = n4131 ^ n3258;
  assign n4135 = n4134 ^ n4132;
  assign n4129 = ~n2447 & n2719;
  assign n4127 = ~n2724 & n3225;
  assign n4126 = n2756 & ~n4125;
  assign n4128 = n4127 ^ n4126;
  assign n4130 = n4129 ^ n4128;
  assign n4136 = n4135 ^ n4130;
  assign n4121 = n4014 ^ n3998;
  assign n4122 = n4015 & ~n4121;
  assign n4123 = n4122 ^ n3998;
  assign n4113 = ~n583 & n4008;
  assign n4114 = n4113 ^ n2360;
  assign n4115 = n4113 ^ n4005;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = n4116 ^ n2360;
  assign n4118 = n4117 ^ n2359;
  assign n4119 = ~n583 & ~n4118;
  assign n4097 = ~n2357 & n2536;
  assign n4098 = n2358 & n2541;
  assign n4099 = ~n4097 & ~n4098;
  assign n4101 = n754 & n2745;
  assign n4100 = n754 & ~n2495;
  assign n4102 = n4101 ^ n4100;
  assign n4103 = n4099 & ~n4102;
  assign n4104 = ~n583 & ~n4103;
  assign n4105 = n583 & n4099;
  assign n4106 = ~n4101 & n4105;
  assign n4107 = n2356 ^ n555;
  assign n4108 = n4100 & n4107;
  assign n4109 = ~n4106 & ~n4108;
  assign n4110 = ~n4104 & n4109;
  assign n4111 = n4110 ^ n2476;
  assign n4082 = n2314 ^ n792;
  assign n4083 = n2478 & n4082;
  assign n4084 = n2938 & n4083;
  assign n4086 = ~n2355 & n2490;
  assign n4085 = n2407 & n2484;
  assign n4087 = n4086 ^ n4085;
  assign n4088 = ~n753 & ~n4087;
  assign n4089 = n4088 ^ n753;
  assign n4090 = n4089 ^ n4087;
  assign n4091 = ~n4084 & n4090;
  assign n4092 = n2604 & ~n3210;
  assign n4093 = n4091 & ~n4092;
  assign n4094 = n2478 & ~n3209;
  assign n4095 = n4088 & ~n4094;
  assign n4096 = n4093 & ~n4095;
  assign n4112 = n4111 ^ n4096;
  assign n4120 = n4119 ^ n4112;
  assign n4124 = n4123 ^ n4120;
  assign n4137 = n4136 ^ n4124;
  assign n4079 = n4020 ^ n4016;
  assign n4080 = n4017 & n4079;
  assign n4081 = n4080 ^ n3983;
  assign n4164 = n4137 ^ n4081;
  assign n4138 = ~n4081 & n4137;
  assign n4165 = n4164 ^ n4138;
  assign n4168 = n4167 ^ n4165;
  assign n4163 = n4162 ^ n4138;
  assign n4169 = n4168 ^ n4163;
  assign n4073 = ~n3932 & ~n4032;
  assign n4074 = ~n3925 & ~n3931;
  assign n4075 = ~n4073 & n4074;
  assign n4076 = ~n3926 & ~n4032;
  assign n4077 = n3924 & ~n4076;
  assign n4078 = ~n4075 & ~n4077;
  assign n4170 = n4169 ^ n4078;
  assign n4172 = n4072 & ~n4170;
  assign n4054 = n4033 & ~n4045;
  assign n4055 = n4054 ^ n4046;
  assign n4056 = ~n3907 & ~n4055;
  assign n4174 = ~n4054 & ~n4056;
  assign n4176 = n4172 & n4174;
  assign n4175 = n4174 ^ n4172;
  assign n4177 = n4176 ^ n4175;
  assign n4171 = n4170 ^ n4072;
  assign n4173 = n4172 ^ n4171;
  assign n4178 = n4177 ^ n4173;
  assign n4179 = n4178 ^ n4176;
  assign n4057 = n3910 & n4056;
  assign n4058 = n3766 & ~n4054;
  assign n4059 = n4057 & n4058;
  assign n4052 = n3766 & n3908;
  assign n4053 = n4046 & n4052;
  assign n4060 = n4059 ^ n4053;
  assign n4061 = n3747 & ~n4060;
  assign n4062 = n4061 ^ n3747;
  assign n4048 = ~n3903 & ~n4046;
  assign n4049 = n4048 ^ n3910;
  assign n4050 = n3772 & ~n4049;
  assign n4051 = ~n3747 & ~n4050;
  assign n4063 = n4062 ^ n4051;
  assign n4180 = n4179 ^ n4063;
  assign n4303 = ~n4173 & n4177;
  assign n4305 = n4303 ^ n4061;
  assign n4306 = n4179 & n4305;
  assign n4304 = n4303 ^ n4178;
  assign n4307 = n4306 ^ n4304;
  assign n4308 = ~n4051 & n4307;
  assign n4309 = n4308 ^ n4305;
  assign n4289 = n641 ^ n196;
  assign n4290 = ~n189 & n4289;
  assign n4291 = n461 ^ n322;
  assign n4292 = n4291 ^ n402;
  assign n4293 = ~n4290 & ~n4292;
  assign n4294 = ~n2090 & n4293;
  assign n4295 = n278 ^ n228;
  assign n4296 = n3501 ^ n471;
  assign n4297 = ~n4295 & ~n4296;
  assign n4298 = n4294 & n4297;
  assign n4299 = n3613 & n4298;
  assign n4300 = n3740 & n4299;
  assign n4301 = n2343 & n4300;
  assign n4284 = n4158 ^ n4078;
  assign n4285 = n4284 ^ n4161;
  assign n4286 = ~n4169 & n4285;
  assign n4287 = n4286 ^ n4163;
  assign n4279 = n4136 ^ n4120;
  assign n4280 = n4124 & n4279;
  assign n4281 = n4280 ^ n4136;
  assign n4273 = n3243 ^ n3225;
  assign n4274 = n2739 & ~n4273;
  assign n4275 = n4274 ^ n3225;
  assign n4272 = ~n2725 & n3243;
  assign n4276 = n4275 ^ n4272;
  assign n4267 = ~n2756 & ~n3243;
  assign n4266 = n2756 ^ n2447;
  assign n4268 = n4267 ^ n4266;
  assign n4269 = n2724 & ~n4268;
  assign n4270 = n4269 ^ n4266;
  assign n4265 = n2428 & n2719;
  assign n4271 = n4270 ^ n4265;
  assign n4277 = n4276 ^ n4271;
  assign n4259 = n792 & n2940;
  assign n4258 = n753 & ~n2941;
  assign n4260 = n4259 ^ n4258;
  assign n4261 = n2478 & n4260;
  assign n4245 = ~n2314 & n2484;
  assign n4244 = n2407 & n2490;
  assign n4246 = n4245 ^ n4244;
  assign n4247 = n4246 ^ n753;
  assign n4248 = n4247 ^ n2346;
  assign n4249 = n2478 ^ n2346;
  assign n4250 = ~n2346 & ~n4249;
  assign n4251 = n4250 ^ n2346;
  assign n4252 = n4248 & ~n4251;
  assign n4253 = n4252 ^ n4250;
  assign n4254 = n4253 ^ n2346;
  assign n4255 = n4254 ^ n2478;
  assign n4256 = ~n4246 & ~n4255;
  assign n4257 = n4256 ^ n4247;
  assign n4262 = n4261 ^ n4257;
  assign n4194 = ~n583 & n2359;
  assign n4236 = ~n2476 & n4110;
  assign n4239 = n4236 ^ n4111;
  assign n4240 = ~n4194 & n4239;
  assign n4237 = n2359 & n4236;
  assign n4238 = n4194 & n4237;
  assign n4241 = n4240 ^ n4238;
  assign n4235 = ~n583 & n2358;
  assign n4242 = n4241 ^ n4235;
  assign n4205 = ~n583 & ~n2357;
  assign n4206 = n4205 ^ n2357;
  assign n4207 = n4206 ^ n2356;
  assign n4208 = ~n555 & ~n4207;
  assign n4209 = n4208 ^ n2356;
  assign n4210 = n1954 & n4209;
  assign n4211 = ~n555 & ~n2356;
  assign n4212 = ~n2357 & ~n2526;
  assign n4213 = ~n2300 & ~n4212;
  assign n4214 = ~n4211 & ~n4213;
  assign n4215 = ~n4210 & ~n4214;
  assign n4216 = n4215 ^ n583;
  assign n4217 = n754 & n2747;
  assign n4218 = n4217 ^ n583;
  assign n4219 = n1955 ^ n583;
  assign n4220 = n4219 ^ n2540;
  assign n4221 = ~n2741 & n4220;
  assign n4222 = n2355 ^ n555;
  assign n4223 = n754 & ~n2746;
  assign n4224 = n4222 & n4223;
  assign n4225 = ~n4221 & ~n4224;
  assign n4226 = n4225 ^ n583;
  assign n4227 = ~n583 & ~n4226;
  assign n4228 = n4227 ^ n583;
  assign n4229 = ~n4218 & ~n4228;
  assign n4230 = n4229 ^ n4227;
  assign n4231 = n4230 ^ n583;
  assign n4232 = n4231 ^ n4225;
  assign n4233 = n4216 & ~n4232;
  assign n4234 = n4233 ^ n4225;
  assign n4243 = n4242 ^ n4234;
  assign n4263 = n4262 ^ n4243;
  assign n4195 = n4096 & n4111;
  assign n4196 = ~n4194 & n4195;
  assign n4197 = n4111 ^ n2359;
  assign n4198 = ~n4117 & n4197;
  assign n4199 = ~n4096 & ~n4198;
  assign n4200 = n2359 & ~n4111;
  assign n4201 = n4117 & ~n4200;
  assign n4202 = ~n583 & ~n4201;
  assign n4203 = ~n4199 & n4202;
  assign n4204 = ~n4196 & ~n4203;
  assign n4264 = n4263 ^ n4204;
  assign n4278 = n4277 ^ n4264;
  assign n4282 = n4281 ^ n4278;
  assign n4182 = ~n2444 & n2996;
  assign n4181 = n2962 & ~n3616;
  assign n4183 = n4182 ^ n4181;
  assign n4184 = ~n1283 & n4183;
  assign n4185 = n1283 & ~n4181;
  assign n4186 = ~n2444 & n3398;
  assign n4187 = n4185 & ~n4186;
  assign n4188 = n2942 & ~n4187;
  assign n4189 = n4185 ^ n2943;
  assign n4190 = ~n3810 & ~n4189;
  assign n4191 = n4190 ^ n2943;
  assign n4192 = ~n4188 & ~n4191;
  assign n4193 = ~n4184 & ~n4192;
  assign n4283 = n4282 ^ n4193;
  assign n4288 = n4287 ^ n4283;
  assign n4302 = n4301 ^ n4288;
  assign n4310 = n4309 ^ n4302;
  assign n4431 = n4303 ^ n4288;
  assign n4432 = n4302 & ~n4431;
  assign n4433 = n4432 ^ n4303;
  assign n4411 = n147 ^ n61;
  assign n4412 = ~n43 & n647;
  assign n4413 = n4412 ^ n258;
  assign n4414 = ~n4411 & n4413;
  assign n4415 = ~n3732 & ~n4414;
  assign n4416 = n3599 & n4415;
  assign n4417 = n1985 ^ n471;
  assign n4418 = n4417 ^ n486;
  assign n4419 = n2250 & ~n4418;
  assign n4420 = n4416 & n4419;
  assign n4421 = n375 ^ n166;
  assign n4422 = n4421 ^ n740;
  assign n4423 = ~n854 & ~n4422;
  assign n4424 = n250 ^ n220;
  assign n4425 = n4424 ^ n320;
  assign n4426 = n4423 & ~n4425;
  assign n4427 = n4420 & n4426;
  assign n4428 = n2185 & n4427;
  assign n4429 = n3499 & n4428;
  assign n4405 = n4277 ^ n4204;
  assign n4406 = ~n4264 & ~n4405;
  assign n4407 = n4406 ^ n4277;
  assign n4399 = n2447 ^ n2430;
  assign n4400 = ~n2739 & n4399;
  assign n4401 = n4400 ^ n2430;
  assign n4398 = ~n2430 & ~n2725;
  assign n4402 = n4401 ^ n4398;
  assign n4396 = ~n2444 & n2719;
  assign n4392 = n2428 ^ n955;
  assign n4391 = n955 & n2430;
  assign n4393 = n4392 ^ n4391;
  assign n4394 = n2724 & n4393;
  assign n4395 = n4394 ^ n4392;
  assign n4397 = n4396 ^ n4395;
  assign n4403 = n4402 ^ n4397;
  assign n4387 = n4262 ^ n4242;
  assign n4388 = n4243 & n4387;
  assign n4389 = n4388 ^ n4262;
  assign n4382 = n4240 ^ n4237;
  assign n4383 = ~n4235 & n4382;
  assign n4381 = n4237 ^ n4205;
  assign n4384 = n4383 ^ n4381;
  assign n4365 = n2355 ^ n583;
  assign n4366 = n2529 ^ n2525;
  assign n4367 = ~n4365 & n4366;
  assign n4371 = ~n583 & ~n2356;
  assign n4372 = ~n2301 & ~n4371;
  assign n4370 = n2539 & n4211;
  assign n4373 = n4372 ^ n4370;
  assign n4368 = ~n583 & ~n2355;
  assign n4369 = n2300 & n4368;
  assign n4374 = n4373 ^ n4369;
  assign n4375 = ~n4367 & ~n4374;
  assign n4376 = n584 & n2740;
  assign n4377 = n4376 ^ n555;
  assign n4378 = n4377 ^ n2407;
  assign n4379 = n754 & n4378;
  assign n4380 = n4375 & ~n4379;
  assign n4385 = n4384 ^ n4380;
  assign n4350 = n2478 & ~n3225;
  assign n4351 = n2972 & n4350;
  assign n4352 = n2346 & n2484;
  assign n4353 = ~n2314 & n2490;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = ~n4351 & n4354;
  assign n4356 = ~n753 & ~n4355;
  assign n4357 = n2478 & ~n2972;
  assign n4360 = n3225 ^ n792;
  assign n4358 = n753 & n4354;
  assign n4359 = ~n4350 & n4358;
  assign n4361 = n4360 ^ n4359;
  assign n4362 = n4357 & ~n4361;
  assign n4363 = n4362 ^ n4359;
  assign n4364 = ~n4356 & ~n4363;
  assign n4386 = n4385 ^ n4364;
  assign n4390 = n4389 ^ n4386;
  assign n4404 = n4403 ^ n4390;
  assign n4408 = n4407 ^ n4404;
  assign n4346 = n4278 ^ n4193;
  assign n4347 = ~n4282 & ~n4346;
  assign n4348 = n4347 ^ n4193;
  assign n4335 = ~n1337 & ~n3616;
  assign n4336 = n4335 ^ n1283;
  assign n4337 = ~n3595 & ~n4336;
  assign n4338 = n4337 ^ n1283;
  assign n4339 = n2957 ^ n1393;
  assign n4340 = ~n4338 & n4339;
  assign n4341 = n2958 ^ n1283;
  assign n4342 = ~n3400 & n4341;
  assign n4343 = ~n3616 & n4342;
  assign n4344 = n4343 ^ n1283;
  assign n4345 = ~n4340 & n4344;
  assign n4349 = n4348 ^ n4345;
  assign n4409 = n4408 ^ n4349;
  assign n4323 = ~n4167 & ~n4168;
  assign n4324 = ~n4283 & ~n4323;
  assign n4325 = n4078 & ~n4324;
  assign n4326 = ~n4162 & n4283;
  assign n4327 = ~n4138 & ~n4326;
  assign n4328 = ~n4325 & n4327;
  assign n4329 = ~n4165 & n4283;
  assign n4330 = n4161 ^ n4078;
  assign n4331 = n4284 & n4330;
  assign n4332 = n4331 ^ n4078;
  assign n4333 = ~n4329 & ~n4332;
  assign n4334 = ~n4328 & ~n4333;
  assign n4410 = n4409 ^ n4334;
  assign n4430 = n4429 ^ n4410;
  assign n4434 = n4433 ^ n4430;
  assign n4311 = ~n4179 & n4302;
  assign n4312 = n4311 ^ n4178;
  assign n4313 = n4060 & ~n4312;
  assign n4314 = n3747 & ~n4313;
  assign n4315 = ~n4177 & ~n4302;
  assign n4316 = n4050 & ~n4176;
  assign n4317 = ~n4315 & n4316;
  assign n4318 = n4302 ^ n4174;
  assign n4319 = ~n4173 & n4318;
  assign n4320 = n4319 ^ n4174;
  assign n4321 = n4317 & ~n4320;
  assign n4322 = ~n4314 & ~n4321;
  assign n4435 = n4434 ^ n4322;
  assign n4531 = n4433 ^ n4410;
  assign n4532 = n4430 & ~n4531;
  assign n4533 = n4532 ^ n4433;
  assign n4522 = ~n4404 & ~n4407;
  assign n4523 = n4522 ^ n4334;
  assign n4524 = n4523 ^ n4408;
  assign n4525 = n4524 ^ n4522;
  assign n4526 = n4409 & n4525;
  assign n4527 = n4526 ^ n4523;
  assign n4520 = n4345 & ~n4348;
  assign n4521 = n4520 ^ n4349;
  assign n4528 = n4527 ^ n4521;
  assign n4514 = n3596 ^ n2428;
  assign n4515 = n2739 & ~n4514;
  assign n4516 = n4515 ^ n2428;
  assign n4511 = n2724 & ~n3596;
  assign n4512 = n959 & n4511;
  assign n4513 = n4512 ^ n3596;
  assign n4517 = n4516 ^ n4513;
  assign n4506 = n2756 & n3596;
  assign n4505 = n2756 ^ n2444;
  assign n4507 = n4506 ^ n4505;
  assign n4508 = n2724 & n4507;
  assign n4509 = n4508 ^ n4505;
  assign n4504 = n2719 & ~n3616;
  assign n4510 = n4509 ^ n4504;
  assign n4518 = n4517 ^ n4510;
  assign n4500 = n4403 ^ n4386;
  assign n4501 = n4390 & n4500;
  assign n4502 = n4501 ^ n4403;
  assign n4496 = n2480 & ~n3258;
  assign n4495 = n2484 & ~n3225;
  assign n4497 = n4496 ^ n4495;
  assign n4486 = n2478 & ~n3258;
  assign n4492 = n4486 ^ n2478;
  assign n4490 = n2346 & n2490;
  assign n4489 = ~n2447 & n2478;
  assign n4491 = n4490 ^ n4489;
  assign n4493 = n4492 ^ n4491;
  assign n4487 = n2478 ^ n753;
  assign n4488 = ~n4486 & ~n4487;
  assign n4494 = n4493 ^ n4488;
  assign n4498 = n4497 ^ n4494;
  assign n4482 = n4384 ^ n4364;
  assign n4483 = ~n4385 & ~n4482;
  assign n4484 = n4483 ^ n4364;
  assign n4449 = n583 & ~n4239;
  assign n4450 = n2358 & n2359;
  assign n4451 = n4110 & n4450;
  assign n4452 = ~n2357 & ~n2476;
  assign n4453 = n4451 & n4452;
  assign n4454 = ~n2356 & n4453;
  assign n4455 = ~n4449 & ~n4454;
  assign n4462 = n2306 ^ n583;
  assign n4460 = n2540 ^ n2529;
  assign n4461 = n4460 ^ n2541;
  assign n4463 = n4462 ^ n4461;
  assign n4464 = n4463 ^ n2541;
  assign n4465 = n2938 & ~n4464;
  assign n4459 = n2407 & n2536;
  assign n4466 = n4465 ^ n4459;
  assign n4457 = n754 & ~n2314;
  assign n4456 = ~n2355 & n2541;
  assign n4458 = n4457 ^ n4456;
  assign n4467 = n4466 ^ n4458;
  assign n4468 = ~n4455 & ~n4467;
  assign n4469 = ~n4194 & ~n4235;
  assign n4470 = ~n4205 & n4469;
  assign n4471 = ~n4110 & n4470;
  assign n4472 = n2476 & ~n4471;
  assign n4473 = n4472 ^ n2476;
  assign n4475 = n2356 & ~n4473;
  assign n4474 = ~n4371 & ~n4473;
  assign n4476 = n4475 ^ n4474;
  assign n4477 = n4467 & ~n4476;
  assign n4478 = n4477 ^ n4475;
  assign n4479 = ~n4453 & n4478;
  assign n4480 = ~n4468 & ~n4479;
  assign n4481 = n4480 ^ n1283;
  assign n4485 = n4484 ^ n4481;
  assign n4499 = n4498 ^ n4485;
  assign n4503 = n4502 ^ n4499;
  assign n4519 = n4518 ^ n4503;
  assign n4529 = n4528 ^ n4519;
  assign n4440 = n226 & ~n3554;
  assign n4441 = ~n288 & ~n4292;
  assign n4442 = ~n317 & n571;
  assign n4443 = n4442 ^ n845;
  assign n4444 = n4443 ^ n415;
  assign n4445 = n4441 & ~n4444;
  assign n4446 = n4420 & n4445;
  assign n4447 = ~n4440 & n4446;
  assign n4448 = n2038 & n4447;
  assign n4530 = n4529 ^ n4448;
  assign n4534 = n4533 ^ n4530;
  assign n4436 = n4321 & n4434;
  assign n4437 = ~n3747 & ~n4436;
  assign n4438 = n4313 & ~n4434;
  assign n4439 = ~n4437 & ~n4438;
  assign n4535 = n4534 ^ n4439;
  assign n4633 = n156 ^ n83;
  assign n4634 = ~n60 & n4633;
  assign n4635 = n629 ^ n175;
  assign n4636 = n4635 ^ n700;
  assign n4637 = ~n4634 & n4636;
  assign n4638 = n1964 & n4637;
  assign n4639 = n3500 & n4638;
  assign n4640 = ~n2233 & ~n2331;
  assign n4641 = n464 ^ n375;
  assign n4642 = n4640 & ~n4641;
  assign n4644 = n565 ^ n418;
  assign n4643 = n988 ^ n870;
  assign n4645 = n4644 ^ n4643;
  assign n4646 = n4642 & ~n4645;
  assign n4647 = n4639 & n4646;
  assign n4648 = n3548 & n4647;
  assign n4627 = n4498 ^ n4481;
  assign n4628 = ~n4485 & n4627;
  assign n4629 = n4628 ^ n4484;
  assign n4620 = ~n2444 & ~n2739;
  assign n4619 = ~n2724 & ~n3616;
  assign n4621 = n4620 ^ n4619;
  assign n4622 = n4621 ^ n955;
  assign n4623 = n4622 ^ n959;
  assign n4624 = n2719 & n3810;
  assign n4625 = ~n4623 & n4624;
  assign n4626 = n4625 ^ n4622;
  assign n4630 = n4629 ^ n4626;
  assign n4615 = n4518 ^ n4499;
  assign n4616 = ~n4503 & ~n4615;
  assign n4617 = n4616 ^ n4502;
  assign n4607 = n1283 ^ n583;
  assign n4608 = n4467 ^ n1283;
  assign n4597 = n4205 & n4451;
  assign n4598 = ~n4472 & ~n4597;
  assign n4609 = n4608 ^ n4598;
  assign n4610 = ~n4607 & n4609;
  assign n4611 = n4610 ^ n4598;
  assign n4596 = n4467 ^ n583;
  assign n4599 = n4598 ^ n4596;
  assign n4600 = n4598 ^ n2476;
  assign n4601 = n4598 ^ n4467;
  assign n4602 = n2356 & n4601;
  assign n4603 = n4602 ^ n4467;
  assign n4604 = n4600 & ~n4603;
  assign n4605 = n4604 ^ n2476;
  assign n4606 = n4599 & n4605;
  assign n4612 = n4611 ^ n4606;
  assign n4589 = n2476 ^ n1283;
  assign n4590 = n4371 ^ n583;
  assign n4591 = n4590 ^ n2476;
  assign n4592 = n4589 & ~n4591;
  assign n4593 = n4592 ^ n1283;
  assign n4594 = n4593 ^ n4368;
  assign n4574 = n754 & n2346;
  assign n4575 = ~n2940 & n4574;
  assign n4577 = ~n2314 & n2536;
  assign n4576 = n2407 & n2541;
  assign n4578 = n4577 ^ n4576;
  assign n4579 = ~n4575 & ~n4578;
  assign n4580 = ~n583 & ~n4579;
  assign n4581 = n2346 ^ n555;
  assign n4582 = n754 & n4581;
  assign n4583 = n2940 & n4582;
  assign n4584 = ~n4580 & ~n4583;
  assign n4585 = n754 & ~n2973;
  assign n4586 = n583 & ~n4578;
  assign n4587 = ~n4585 & n4586;
  assign n4588 = n4584 & ~n4587;
  assign n4595 = n4594 ^ n4588;
  assign n4613 = n4612 ^ n4595;
  assign n4558 = ~n792 & n2428;
  assign n4559 = ~n3796 & ~n4558;
  assign n4560 = n2478 & ~n4559;
  assign n4562 = n2490 & ~n3225;
  assign n4561 = ~n2447 & n2484;
  assign n4563 = n4562 ^ n4561;
  assign n4564 = ~n4560 & ~n4563;
  assign n4565 = ~n753 & ~n4564;
  assign n4566 = n753 & ~n4563;
  assign n4567 = ~n792 & n3243;
  assign n4568 = n4567 ^ n2428;
  assign n4569 = n2478 & n4568;
  assign n4570 = n4566 & ~n4569;
  assign n4571 = n2489 & n3797;
  assign n4572 = ~n4570 & ~n4571;
  assign n4573 = ~n4565 & n4572;
  assign n4614 = n4613 ^ n4573;
  assign n4618 = n4617 ^ n4614;
  assign n4631 = n4630 ^ n4618;
  assign n4545 = n4522 ^ n4408;
  assign n4546 = n4519 & n4545;
  assign n4547 = n4348 ^ n4334;
  assign n4548 = n4349 & n4547;
  assign n4549 = n4548 ^ n4334;
  assign n4550 = ~n4546 & ~n4549;
  assign n4551 = n4521 & n4545;
  assign n4552 = ~n4519 & ~n4551;
  assign n4553 = n4334 & ~n4552;
  assign n4554 = n4519 & ~n4520;
  assign n4555 = ~n4522 & ~n4554;
  assign n4556 = ~n4553 & n4555;
  assign n4557 = ~n4550 & ~n4556;
  assign n4632 = n4631 ^ n4557;
  assign n4649 = n4648 ^ n4632;
  assign n4542 = n4533 ^ n4529;
  assign n4543 = ~n4530 & n4542;
  assign n4544 = n4543 ^ n4533;
  assign n4650 = n4649 ^ n4544;
  assign n4539 = n4438 & n4534;
  assign n4540 = n3747 & ~n4539;
  assign n4536 = n4436 & ~n4534;
  assign n4537 = ~n3747 & ~n4536;
  assign n4538 = n4537 ^ n3747;
  assign n4541 = n4540 ^ n4538;
  assign n4651 = n4650 ^ n4541;
  assign n4742 = n4649 ^ n4540;
  assign n4743 = n4742 ^ n4537;
  assign n4744 = n4650 & ~n4743;
  assign n4745 = n4744 ^ n4537;
  assign n4740 = n4632 & n4648;
  assign n4741 = n4740 ^ n4649;
  assign n4746 = n4745 ^ n4741;
  assign n4719 = n959 & ~n3616;
  assign n4720 = n4719 ^ n955;
  assign n4721 = ~n3595 & ~n4720;
  assign n4722 = n4721 ^ n955;
  assign n4723 = ~n2722 & ~n4722;
  assign n4724 = n2727 ^ n955;
  assign n4725 = ~n3616 & n4724;
  assign n4726 = n4725 ^ n955;
  assign n4727 = n2726 ^ n960;
  assign n4728 = n4727 ^ n4723;
  assign n4729 = n4726 & ~n4728;
  assign n4730 = n4729 ^ n4727;
  assign n4731 = ~n4723 & n4730;
  assign n4732 = n4731 ^ n4723;
  assign n4733 = n4732 ^ n4723;
  assign n4716 = n4612 ^ n4573;
  assign n4717 = n4613 & n4716;
  assign n4718 = n4717 ^ n4573;
  assign n4734 = n4733 ^ n4718;
  assign n4712 = n2407 ^ n2355;
  assign n4713 = ~n583 & n4712;
  assign n4694 = ~n2314 & n2511;
  assign n4695 = ~n1955 & ~n4694;
  assign n4696 = n2346 & n2529;
  assign n4697 = n4696 ^ n1954;
  assign n4698 = ~n4695 & ~n4697;
  assign n4700 = n2355 ^ n2314;
  assign n4701 = ~n583 & n4700;
  assign n4699 = n4368 ^ n2314;
  assign n4702 = n4701 ^ n4699;
  assign n4703 = n4702 ^ n2346;
  assign n4704 = n753 & ~n4703;
  assign n4705 = n4704 ^ n2346;
  assign n4706 = ~n555 & n4705;
  assign n4707 = ~n4698 & ~n4706;
  assign n4708 = n584 & ~n2972;
  assign n4709 = n4708 ^ n3225;
  assign n4710 = n754 & n4709;
  assign n4711 = ~n4707 & ~n4710;
  assign n4714 = n4713 ^ n4711;
  assign n4689 = n4588 ^ n4368;
  assign n4690 = n4593 ^ n4588;
  assign n4691 = ~n4689 & n4690;
  assign n4692 = n4691 ^ n4368;
  assign n4674 = n2478 & ~n3960;
  assign n4676 = n2428 & n2484;
  assign n4675 = ~n2447 & n2490;
  assign n4677 = n4676 ^ n4675;
  assign n4678 = ~n4674 & ~n4677;
  assign n4679 = ~n753 & ~n4678;
  assign n4680 = n3596 ^ n2405;
  assign n4681 = n2478 & n4680;
  assign n4682 = n753 & ~n4677;
  assign n4683 = ~n4681 & n4682;
  assign n4684 = n2444 ^ n792;
  assign n4685 = n2478 & ~n4684;
  assign n4686 = ~n2430 & n4685;
  assign n4687 = ~n4683 & ~n4686;
  assign n4688 = ~n4679 & n4687;
  assign n4693 = n4692 ^ n4688;
  assign n4715 = n4714 ^ n4693;
  assign n4735 = n4734 ^ n4715;
  assign n4664 = ~n4614 & n4617;
  assign n4670 = n4664 ^ n4618;
  assign n4663 = n4626 & ~n4629;
  assign n4672 = n4663 ^ n4630;
  assign n4673 = ~n4670 & n4672;
  assign n4736 = n4735 ^ n4673;
  assign n4671 = ~n4630 & n4670;
  assign n4737 = n4736 ^ n4671;
  assign n4666 = ~n4663 & n4664;
  assign n4665 = n4664 ^ n4663;
  assign n4667 = n4666 ^ n4665;
  assign n4668 = n4618 & n4667;
  assign n4661 = n4630 ^ n4557;
  assign n4662 = n4631 & n4661;
  assign n4669 = n4668 ^ n4662;
  assign n4738 = n4737 ^ n4669;
  assign n4654 = n363 ^ n286;
  assign n4652 = n2074 ^ n175;
  assign n4653 = n4652 ^ n115;
  assign n4655 = n4654 ^ n4653;
  assign n4656 = ~n3728 & n4655;
  assign n4657 = n847 & ~n4425;
  assign n4658 = n4656 & n4657;
  assign n4659 = n3505 & n4658;
  assign n4660 = n2253 & n4659;
  assign n4739 = n4738 ^ n4660;
  assign n4747 = n4746 ^ n4739;
  assign n4835 = n4740 ^ n4544;
  assign n4748 = n4544 & ~n4649;
  assign n4836 = n4835 ^ n4748;
  assign n4837 = n4836 ^ n4660;
  assign n4838 = n4739 & ~n4837;
  assign n4839 = n4838 ^ n4738;
  assign n4826 = ~n103 & ~n2201;
  assign n4827 = n3474 ^ n187;
  assign n4828 = n4827 ^ n267;
  assign n4829 = n4826 & n4828;
  assign n4830 = n3737 & n4829;
  assign n4831 = n686 & n4830;
  assign n4832 = n1151 & n3566;
  assign n4833 = n4831 & n4832;
  assign n4820 = n4714 ^ n4692;
  assign n4821 = n4693 & ~n4820;
  assign n4822 = n4821 ^ n4688;
  assign n4799 = n584 & n3258;
  assign n4800 = n4799 ^ n555;
  assign n4801 = n4800 ^ n2447;
  assign n4802 = n754 & n4801;
  assign n4803 = n2538 & n3225;
  assign n4811 = ~n1955 & n3225;
  assign n4812 = n4811 ^ n2525;
  assign n4809 = ~n2346 & n2539;
  assign n4810 = n4809 ^ n1954;
  assign n4813 = n4812 ^ n4810;
  assign n4805 = ~n583 & n2346;
  assign n4806 = n4805 ^ n583;
  assign n4807 = ~n1955 & ~n4806;
  assign n4804 = n2539 & ~n3225;
  assign n4808 = n4807 ^ n4804;
  assign n4814 = n4813 ^ n4808;
  assign n4815 = n555 & n4814;
  assign n4816 = n4815 ^ n4813;
  assign n4817 = ~n4803 & ~n4816;
  assign n4818 = ~n4802 & n4817;
  assign n4792 = n4711 ^ n583;
  assign n4793 = n4792 ^ n2407;
  assign n4794 = n4711 ^ n2355;
  assign n4795 = ~n4712 & ~n4794;
  assign n4796 = ~n4793 & n4795;
  assign n4797 = n4796 ^ n4792;
  assign n4791 = n4701 ^ n955;
  assign n4798 = n4797 ^ n4791;
  assign n4819 = n4818 ^ n4798;
  assign n4823 = n4822 ^ n4819;
  assign n4787 = n4718 ^ n4715;
  assign n4788 = n4734 & n4787;
  assign n4789 = n4788 ^ n4715;
  assign n4772 = n2478 & ~n3808;
  assign n4774 = n2428 & n2490;
  assign n4773 = ~n2444 & n2484;
  assign n4775 = n4774 ^ n4773;
  assign n4777 = n753 & n4775;
  assign n4776 = n4775 ^ n753;
  assign n4778 = n4777 ^ n4776;
  assign n4779 = ~n4772 & ~n4778;
  assign n4780 = n2604 & n3809;
  assign n4781 = n3616 ^ n792;
  assign n4782 = n2478 & n4781;
  assign n4783 = ~n3596 & n4782;
  assign n4784 = ~n4777 & ~n4783;
  assign n4785 = ~n4780 & n4784;
  assign n4786 = ~n4779 & n4785;
  assign n4790 = n4789 ^ n4786;
  assign n4824 = n4823 ^ n4790;
  assign n4762 = ~n4663 & ~n4735;
  assign n4763 = ~n4666 & ~n4762;
  assign n4764 = ~n4670 & ~n4735;
  assign n4765 = ~n4673 & ~n4764;
  assign n4766 = n4763 & n4765;
  assign n4767 = n4557 & ~n4766;
  assign n4768 = n4672 & ~n4763;
  assign n4769 = ~n4667 & n4764;
  assign n4770 = ~n4768 & ~n4769;
  assign n4771 = ~n4767 & n4770;
  assign n4825 = n4824 ^ n4771;
  assign n4834 = n4833 ^ n4825;
  assign n4840 = n4839 ^ n4834;
  assign n4749 = n4536 & ~n4748;
  assign n4750 = n4740 ^ n4739;
  assign n4751 = n4739 ^ n4544;
  assign n4752 = n4750 & n4751;
  assign n4753 = n4752 ^ n4741;
  assign n4754 = n4739 & n4753;
  assign n4755 = n4754 ^ n4741;
  assign n4756 = n4749 & ~n4755;
  assign n4757 = ~n3747 & ~n4756;
  assign n4758 = n4739 & ~n4741;
  assign n4759 = n4758 ^ n4752;
  assign n4760 = n4539 & n4759;
  assign n4761 = ~n4757 & ~n4760;
  assign n4841 = n4840 ^ n4761;
  assign n4898 = n4839 ^ n4825;
  assign n4899 = ~n4834 & n4898;
  assign n4900 = n4899 ^ n4839;
  assign n4892 = n4790 ^ n4771;
  assign n4893 = ~n4824 & ~n4892;
  assign n4891 = ~n4819 & ~n4822;
  assign n4894 = n4893 ^ n4891;
  assign n4889 = n4786 & ~n4789;
  assign n4890 = n4889 ^ n4790;
  assign n4895 = n4894 ^ n4890;
  assign n4886 = n2479 & n3810;
  assign n4883 = n753 & ~n3810;
  assign n4884 = ~n2603 & ~n4883;
  assign n4881 = ~n2444 & n2490;
  assign n4880 = n2484 & ~n3616;
  assign n4882 = n4881 ^ n4880;
  assign n4885 = n4884 ^ n4882;
  assign n4887 = n4886 ^ n4885;
  assign n4876 = n4818 ^ n4791;
  assign n4877 = n4798 & ~n4876;
  assign n4878 = n4877 ^ n4797;
  assign n4871 = ~n2541 & ~n4273;
  assign n4872 = n4871 ^ n3225;
  assign n4863 = ~n2536 & n3243;
  assign n4869 = ~n555 & n4863;
  assign n4870 = n4869 ^ n3243;
  assign n4873 = n4872 ^ n4870;
  assign n4866 = n2447 & n2536;
  assign n4864 = n2536 ^ n583;
  assign n4865 = ~n4863 & ~n4864;
  assign n4867 = n4866 ^ n4865;
  assign n4862 = n754 & n2428;
  assign n4868 = n4867 ^ n4862;
  assign n4874 = n4873 ^ n4868;
  assign n4854 = n2355 ^ n955;
  assign n4855 = ~n4700 & n4854;
  assign n4856 = n4855 ^ n955;
  assign n4857 = n2346 & ~n4856;
  assign n4858 = n4856 ^ n2346;
  assign n4859 = n4858 ^ n4857;
  assign n4860 = ~n583 & ~n4859;
  assign n4861 = ~n4857 & n4860;
  assign n4875 = n4874 ^ n4861;
  assign n4879 = n4878 ^ n4875;
  assign n4888 = n4887 ^ n4879;
  assign n4896 = n4895 ^ n4888;
  assign n4846 = ~n1044 & n2438;
  assign n4847 = n460 ^ n329;
  assign n4848 = n4847 ^ n359;
  assign n4849 = ~n202 & n4848;
  assign n4850 = ~n991 & ~n1065;
  assign n4851 = n4849 & n4850;
  assign n4852 = n4846 & n4851;
  assign n4853 = n655 & n4852;
  assign n4897 = n4896 ^ n4853;
  assign n4901 = n4900 ^ n4897;
  assign n4842 = n4756 & ~n4840;
  assign n4843 = ~n3747 & ~n4842;
  assign n4844 = n4760 & n4840;
  assign n4845 = ~n4843 & ~n4844;
  assign n4902 = n4901 ^ n4845;
  assign n4969 = n4900 ^ n4896;
  assign n4970 = ~n4897 & n4969;
  assign n4971 = n4970 ^ n4900;
  assign n4957 = ~n792 & ~n3616;
  assign n4958 = n4957 ^ n753;
  assign n4959 = ~n3595 & ~n4958;
  assign n4960 = n4959 ^ n753;
  assign n4961 = ~n2482 & ~n4960;
  assign n4962 = n2488 & ~n3616;
  assign n4963 = n4962 ^ n753;
  assign n4964 = ~n4961 & n4963;
  assign n4942 = n754 & n4680;
  assign n4944 = ~n2447 & n2541;
  assign n4943 = n2428 & n2536;
  assign n4945 = n4944 ^ n4943;
  assign n4947 = n583 & n4945;
  assign n4946 = n4945 ^ n583;
  assign n4948 = n4947 ^ n4946;
  assign n4949 = ~n4942 & ~n4948;
  assign n4950 = ~n3960 & n4220;
  assign n4951 = n2444 ^ n555;
  assign n4952 = n754 & n4951;
  assign n4953 = ~n2430 & n4952;
  assign n4954 = ~n4947 & ~n4953;
  assign n4955 = ~n4950 & n4954;
  assign n4956 = ~n4949 & n4955;
  assign n4965 = n4964 ^ n4956;
  assign n4928 = n4890 & ~n4891;
  assign n4929 = n4888 & ~n4928;
  assign n4930 = ~n4771 & ~n4929;
  assign n4931 = n4891 ^ n4823;
  assign n4932 = ~n4888 & ~n4889;
  assign n4933 = n4931 & ~n4932;
  assign n4934 = ~n4930 & n4933;
  assign n4935 = ~n4888 & ~n4891;
  assign n4936 = n4789 ^ n4771;
  assign n4937 = n4786 ^ n4771;
  assign n4938 = ~n4936 & n4937;
  assign n4939 = n4938 ^ n4771;
  assign n4940 = ~n4935 & n4939;
  assign n4941 = ~n4934 & ~n4940;
  assign n4966 = n4965 ^ n4941;
  assign n4924 = n4887 ^ n4875;
  assign n4925 = ~n4879 & n4924;
  assign n4926 = n4925 ^ n4878;
  assign n4921 = ~n583 & ~n3225;
  assign n4920 = ~n4860 & n4874;
  assign n4922 = n4921 ^ n4920;
  assign n4918 = n4857 & ~n4874;
  assign n4919 = ~n583 & n4918;
  assign n4923 = n4922 ^ n4919;
  assign n4927 = n4926 ^ n4923;
  assign n4967 = n4966 ^ n4927;
  assign n4907 = ~n101 & ~n1042;
  assign n4908 = n419 ^ n174;
  assign n4909 = n4908 ^ n414;
  assign n4910 = ~n4907 & ~n4909;
  assign n4911 = n2121 ^ n335;
  assign n4912 = n4911 ^ n218;
  assign n4913 = ~n1070 & n4912;
  assign n4914 = n3898 & n4913;
  assign n4915 = n2031 & n4914;
  assign n4916 = n477 & n4915;
  assign n4917 = n4910 & n4916;
  assign n4968 = n4967 ^ n4917;
  assign n4972 = n4971 ^ n4968;
  assign n4903 = n4842 & ~n4901;
  assign n4904 = ~n3747 & ~n4903;
  assign n4905 = n4844 & n4901;
  assign n4906 = ~n4904 & ~n4905;
  assign n4973 = n4972 ^ n4906;
  assign n5060 = n4971 ^ n4967;
  assign n5061 = ~n4968 & n5060;
  assign n5062 = n5061 ^ n4971;
  assign n5041 = n4923 & ~n4926;
  assign n5050 = n5041 ^ n4927;
  assign n5051 = ~n4941 & ~n5050;
  assign n5033 = n4956 & ~n4964;
  assign n5040 = n5033 ^ n4965;
  assign n5052 = n5051 ^ n5040;
  assign n5024 = n235 & n3225;
  assign n5025 = ~n583 & ~n5024;
  assign n5026 = n5024 ^ n3225;
  assign n5027 = n5026 ^ n2447;
  assign n5028 = n5025 & n5027;
  assign n5029 = n5028 ^ n753;
  assign n4997 = n3616 ^ n555;
  assign n4998 = ~n3596 & n4997;
  assign n4999 = n4998 ^ n3808;
  assign n5002 = ~n2444 & ~n4461;
  assign n5000 = ~n583 & ~n2428;
  assign n5001 = ~n2302 & ~n5000;
  assign n5003 = n5002 ^ n5001;
  assign n5004 = n4999 & ~n5003;
  assign n5015 = n2539 ^ n555;
  assign n5016 = n2428 & n2539;
  assign n5017 = n5015 & ~n5016;
  assign n5012 = n1954 ^ n555;
  assign n5013 = n1954 & ~n2444;
  assign n5014 = ~n5012 & ~n5013;
  assign n5018 = n5017 ^ n5014;
  assign n5008 = ~n2428 & ~n2526;
  assign n5009 = n555 & n5008;
  assign n5007 = ~n555 & n2525;
  assign n5010 = n5009 ^ n5007;
  assign n5005 = ~n555 & n2444;
  assign n5006 = ~n1955 & n5005;
  assign n5011 = n5010 ^ n5006;
  assign n5019 = n5018 ^ n5011;
  assign n5020 = ~n5004 & n5019;
  assign n5021 = n4998 ^ n3809;
  assign n5022 = n4220 & n5021;
  assign n5023 = n5020 & ~n5022;
  assign n5030 = n5029 ^ n5023;
  assign n4995 = ~n4918 & n4921;
  assign n4996 = ~n4920 & ~n4995;
  assign n5031 = n5030 ^ n4996;
  assign n5042 = ~n5031 & ~n5041;
  assign n5053 = n5042 ^ n5041;
  assign n5054 = ~n5040 & ~n5053;
  assign n5055 = n5054 ^ n5041;
  assign n5056 = ~n5052 & ~n5055;
  assign n5057 = n5056 ^ n5042;
  assign n5045 = n5041 ^ n5031;
  assign n5046 = n5045 ^ n5042;
  assign n5032 = ~n4927 & n5031;
  assign n5047 = n5046 ^ n5032;
  assign n5043 = n5040 & n5042;
  assign n5044 = n5043 ^ n5042;
  assign n5048 = n5047 ^ n5044;
  assign n4994 = n4941 ^ n4927;
  assign n5034 = n5033 ^ n5032;
  assign n5035 = n5034 ^ n4965;
  assign n5036 = ~n5032 & n5035;
  assign n5037 = n5036 ^ n5034;
  assign n5038 = ~n4994 & ~n5037;
  assign n5039 = n5038 ^ n5034;
  assign n5049 = n5048 ^ n5039;
  assign n5058 = n5057 ^ n5049;
  assign n4978 = n495 & ~n3553;
  assign n4980 = n693 ^ n365;
  assign n4979 = n2157 ^ n428;
  assign n4981 = n4980 ^ n4979;
  assign n4982 = n4978 & ~n4981;
  assign n4984 = ~n340 & n502;
  assign n4983 = n498 ^ n374;
  assign n4985 = n4984 ^ n4983;
  assign n4986 = n4985 ^ n976;
  assign n4987 = n486 ^ n281;
  assign n4988 = n4987 ^ n222;
  assign n4989 = ~n4986 & ~n4988;
  assign n4990 = n4982 & n4989;
  assign n4991 = n1021 & n4990;
  assign n4992 = n3519 & n4991;
  assign n4993 = n3740 & n4992;
  assign n5059 = n5058 ^ n4993;
  assign n5063 = n5062 ^ n5059;
  assign n4974 = n4903 & ~n4972;
  assign n4975 = ~n3747 & ~n4974;
  assign n4976 = n4905 & n4972;
  assign n4977 = ~n4975 & ~n4976;
  assign n5064 = n5063 ^ n4977;
  assign n5118 = n5062 ^ n5058;
  assign n5119 = ~n5059 & n5118;
  assign n5120 = n5119 ^ n5062;
  assign n5105 = ~n183 & n4633;
  assign n5106 = n2121 ^ n360;
  assign n5107 = n5106 ^ n301;
  assign n5108 = ~n5105 & ~n5107;
  assign n5109 = n304 ^ n177;
  assign n5110 = n5109 ^ n625;
  assign n5111 = ~n220 & n5110;
  assign n5112 = n5108 & n5111;
  assign n5113 = n963 & n5112;
  assign n5114 = n1401 & n5113;
  assign n5115 = n1974 & n2291;
  assign n5116 = n5114 & n5115;
  assign n5100 = n5023 ^ n4996;
  assign n5101 = ~n5030 & ~n5100;
  assign n5102 = n5101 ^ n4996;
  assign n5095 = ~n753 & ~n5024;
  assign n5096 = n5027 & ~n5095;
  assign n5097 = n5096 ^ n2428;
  assign n5098 = ~n583 & n5097;
  assign n5081 = n584 & n3810;
  assign n5082 = n754 & ~n5081;
  assign n5083 = n555 & ~n3616;
  assign n5084 = ~n2444 & n2514;
  assign n5085 = n1954 & ~n5084;
  assign n5086 = ~n5083 & n5085;
  assign n5087 = ~n583 & n2444;
  assign n5088 = n5087 ^ n583;
  assign n5089 = n5088 ^ n3616;
  assign n5090 = n555 & n5089;
  assign n5091 = n5090 ^ n3616;
  assign n5092 = ~n1955 & n5091;
  assign n5093 = ~n5086 & ~n5092;
  assign n5094 = ~n5082 & n5093;
  assign n5099 = n5098 ^ n5094;
  assign n5103 = n5102 ^ n5099;
  assign n5069 = n5040 & n5051;
  assign n5071 = ~n5033 & ~n5047;
  assign n5070 = n5047 ^ n5033;
  assign n5072 = n5071 ^ n5070;
  assign n5073 = ~n5042 & n5072;
  assign n5074 = ~n4941 & n5073;
  assign n5075 = n5040 ^ n5031;
  assign n5076 = n5045 & ~n5075;
  assign n5077 = n5076 ^ n5041;
  assign n5078 = ~n5071 & ~n5077;
  assign n5079 = ~n5074 & n5078;
  assign n5080 = ~n5069 & n5079;
  assign n5104 = n5103 ^ n5080;
  assign n5117 = n5116 ^ n5104;
  assign n5121 = n5120 ^ n5117;
  assign n5065 = n4974 & ~n5063;
  assign n5066 = ~n3747 & ~n5065;
  assign n5067 = n4976 & n5063;
  assign n5068 = ~n5066 & ~n5067;
  assign n5122 = n5121 ^ n5068;
  assign n5188 = n5120 ^ n5104;
  assign n5189 = n5117 & ~n5188;
  assign n5190 = n5189 ^ n5120;
  assign n5141 = n5102 ^ n5080;
  assign n5142 = n5103 & ~n5141;
  assign n5143 = n5142 ^ n5080;
  assign n5146 = n754 & n3595;
  assign n5147 = ~n3616 & ~n4463;
  assign n5148 = ~n5146 & n5147;
  assign n5171 = ~n2428 & ~n5148;
  assign n5172 = n5094 & n5096;
  assign n5173 = n5087 & ~n5172;
  assign n5174 = n5171 & n5173;
  assign n5154 = n2428 & ~n5088;
  assign n5159 = n5094 ^ n583;
  assign n5144 = n583 & ~n5094;
  assign n5160 = n5159 ^ n5144;
  assign n5155 = n5094 ^ n2428;
  assign n5156 = n5097 & n5155;
  assign n5157 = n5156 ^ n2428;
  assign n5158 = ~n583 & ~n5157;
  assign n5161 = n5160 ^ n5158;
  assign n5162 = n5161 ^ n5094;
  assign n5163 = ~n5154 & n5162;
  assign n5169 = n5163 ^ n5162;
  assign n5175 = n5174 ^ n5169;
  assign n5152 = ~n2428 & n2444;
  assign n5180 = n5148 & ~n5152;
  assign n5181 = n5162 & ~n5180;
  assign n5176 = n5088 ^ n5000;
  assign n5177 = ~n5148 & ~n5176;
  assign n5178 = n5177 ^ n5148;
  assign n5179 = ~n5162 & n5178;
  assign n5182 = n5181 ^ n5179;
  assign n5183 = ~n5175 & n5182;
  assign n5167 = ~n5148 & n5154;
  assign n5149 = n583 & ~n5148;
  assign n5150 = n5149 ^ n583;
  assign n5145 = n5144 ^ n583;
  assign n5151 = n5150 ^ n5145;
  assign n5153 = n5152 ^ n5148;
  assign n5164 = ~n5152 & ~n5163;
  assign n5165 = ~n5153 & ~n5164;
  assign n5166 = ~n5151 & ~n5165;
  assign n5168 = n5167 ^ n5166;
  assign n5170 = n5169 ^ n5168;
  assign n5184 = n5183 ^ n5170;
  assign n5185 = ~n5143 & n5184;
  assign n5186 = n5185 ^ n5170;
  assign n5127 = n966 ^ n320;
  assign n5128 = n1184 & ~n5127;
  assign n5129 = n3491 ^ n336;
  assign n5130 = n5129 ^ n223;
  assign n5131 = n5130 ^ n993;
  assign n5132 = n5131 ^ n115;
  assign n5133 = n5109 ^ n450;
  assign n5134 = n5133 ^ n817;
  assign n5135 = n5132 & ~n5134;
  assign n5136 = n3527 & n5135;
  assign n5137 = n1135 & n5136;
  assign n5138 = n2129 & n5137;
  assign n5139 = n5128 & n5138;
  assign n5140 = n4910 & n5139;
  assign n5187 = n5186 ^ n5140;
  assign n5191 = n5190 ^ n5187;
  assign n5123 = n5067 & ~n5121;
  assign n5124 = n3747 & ~n5123;
  assign n5125 = n5065 & n5121;
  assign n5126 = ~n5124 & ~n5125;
  assign n5192 = n5191 ^ n5126;
  assign n5219 = n5190 ^ n5186;
  assign n5220 = n5187 & ~n5219;
  assign n5221 = n5220 ^ n5190;
  assign n5207 = n61 & n2032;
  assign n5208 = ~n2162 & ~n5207;
  assign n5210 = n352 ^ n348;
  assign n5209 = n3518 ^ n304;
  assign n5211 = n5210 ^ n5209;
  assign n5212 = ~n2331 & ~n5211;
  assign n5213 = n3488 & n5212;
  assign n5214 = ~n4981 & n5213;
  assign n5215 = n3532 & n5214;
  assign n5216 = n1057 & n5215;
  assign n5217 = ~n5208 & n5216;
  assign n5201 = n2428 & ~n5087;
  assign n5202 = n3616 & ~n5201;
  assign n5203 = n2444 & n5009;
  assign n5204 = ~n5202 & ~n5203;
  assign n5205 = ~n5149 & n5204;
  assign n5197 = n5162 & n5177;
  assign n5198 = n5197 ^ n5181;
  assign n5199 = n5143 & ~n5198;
  assign n5200 = ~n5179 & ~n5199;
  assign n5206 = n5205 ^ n5200;
  assign n5218 = n5217 ^ n5206;
  assign n5222 = n5221 ^ n5218;
  assign n5193 = n5125 & n5191;
  assign n5194 = ~n3747 & ~n5193;
  assign n5195 = n5123 & ~n5191;
  assign n5196 = ~n5194 & ~n5195;
  assign n5223 = n5222 ^ n5196;
  assign n5239 = n5221 ^ n5206;
  assign n5240 = ~n5218 & n5239;
  assign n5241 = n5240 ^ n5221;
  assign n5228 = ~n873 & ~n1992;
  assign n5229 = ~n4987 & n5228;
  assign n5230 = n395 ^ n217;
  assign n5231 = ~n537 & ~n5230;
  assign n5232 = ~n137 & ~n485;
  assign n5233 = ~n101 & ~n5232;
  assign n5234 = ~n249 & ~n5233;
  assign n5235 = n5231 & n5234;
  assign n5236 = n5229 & n5235;
  assign n5237 = n747 & n5236;
  assign n5238 = n2343 & n5237;
  assign n5242 = n5241 ^ n5238;
  assign n5224 = n5195 & n5222;
  assign n5225 = n3747 & ~n5224;
  assign n5226 = n5193 & ~n5222;
  assign n5227 = ~n5225 & ~n5226;
  assign n5243 = n5242 ^ n5227;
  assign n5255 = n979 & n1020;
  assign n5257 = n998 ^ n628;
  assign n5256 = n4035 ^ n3485;
  assign n5258 = n5257 ^ n5256;
  assign n5259 = n1189 & ~n5258;
  assign n5260 = n5255 & n5259;
  assign n5261 = n712 & n5260;
  assign n5262 = n1128 & n5261;
  assign n5263 = n3545 & n5262;
  assign n5247 = n5226 & n5242;
  assign n5244 = n5238 & n5241;
  assign n5245 = n5244 ^ n5242;
  assign n5246 = n5245 ^ n5226;
  assign n5248 = n5247 ^ n5246;
  assign n5249 = n5248 ^ n5226;
  assign n5250 = ~n3747 & n5249;
  assign n5252 = n5225 & ~n5245;
  assign n5251 = n5224 & n5244;
  assign n5253 = n5252 ^ n5251;
  assign n5254 = ~n5250 & ~n5253;
  assign n5264 = n5263 ^ n5254;
  assign n5272 = n1013 ^ n498;
  assign n5273 = ~n468 & ~n5272;
  assign n5274 = n298 ^ n72;
  assign n5275 = n5274 ^ n662;
  assign n5276 = n5275 ^ n248;
  assign n5277 = n5273 & n5276;
  assign n5278 = ~n4292 & n5277;
  assign n5279 = n398 & n5278;
  assign n5280 = n1040 & n5279;
  assign n5281 = n5128 & n5280;
  assign n5271 = ~n5249 & ~n5263;
  assign n5282 = n5281 ^ n5271;
  assign n5265 = n5245 & ~n5263;
  assign n5266 = n5224 & ~n5265;
  assign n5267 = ~n5247 & ~n5266;
  assign n5268 = ~n5251 & n5263;
  assign n5269 = ~n5267 & ~n5268;
  assign n5270 = n3747 & ~n5269;
  assign n5283 = n5282 ^ n5270;
  assign n5294 = n5270 ^ n3747;
  assign n5295 = n5294 ^ n5281;
  assign n5296 = n5282 & ~n5295;
  assign n5297 = n5296 ^ n3747;
  assign n5284 = n3600 ^ n72;
  assign n5285 = n184 & n5284;
  assign n5287 = n490 ^ n285;
  assign n5286 = n430 ^ n60;
  assign n5288 = n5287 ^ n5286;
  assign n5289 = ~n5285 & n5288;
  assign n5290 = ~n4296 & n5289;
  assign n5291 = ~n161 & n5290;
  assign n5292 = n981 & n5291;
  assign n5293 = n4639 & n5292;
  assign n5298 = n5297 ^ n5293;
  assign n5306 = n5293 ^ n5281;
  assign n5308 = ~n5271 & ~n5306;
  assign n5305 = n5281 & n5293;
  assign n5307 = n5306 ^ n5305;
  assign n5309 = n5308 ^ n5307;
  assign n5310 = n5271 ^ n3747;
  assign n5311 = n5310 ^ n5270;
  assign n5312 = ~n5309 & n5311;
  assign n5313 = n5312 ^ n3747;
  assign n5299 = ~n106 & ~n169;
  assign n5300 = ~n748 & ~n5299;
  assign n5301 = n574 ^ n373;
  assign n5302 = n551 & ~n5301;
  assign n5303 = n2393 & n5302;
  assign n5304 = ~n5300 & n5303;
  assign n5314 = n5313 ^ n5304;
  assign n5319 = n5304 & n5305;
  assign n5316 = ~n5304 & ~n5307;
  assign n5320 = n5319 ^ n5316;
  assign n5321 = ~n5271 & n5320;
  assign n5322 = n5321 ^ n5316;
  assign n5323 = n5269 & n5322;
  assign n5324 = n3747 & ~n5323;
  assign n5317 = n5271 & n5316;
  assign n5315 = n948 & ~n2400;
  assign n5318 = n5317 ^ n5315;
  assign n5325 = n5324 ^ n5318;
  assign n5326 = ~x21 & ~x22;
  assign n5327 = n948 & n5326;
  assign n5328 = n5315 & ~n5317;
  assign n5329 = n5328 ^ n5318;
  assign n5330 = ~n5294 & n5329;
  assign n5331 = n5330 ^ n3747;
  assign n5332 = ~n5327 & ~n5331;
  assign n5333 = ~n5326 & n5328;
  assign n5334 = n5323 & n5333;
  assign n5335 = ~n5332 & ~n5334;
  assign n5336 = n3747 & ~n5334;
  assign y0 = n3593;
  assign y1 = n3757;
  assign y2 = n3904;
  assign y3 = ~n4047;
  assign y4 = ~n4180;
  assign y5 = n4310;
  assign y6 = ~n4435;
  assign y7 = ~n4535;
  assign y8 = n4651;
  assign y9 = n4747;
  assign y10 = ~n4841;
  assign y11 = ~n4902;
  assign y12 = ~n4973;
  assign y13 = ~n5064;
  assign y14 = n5122;
  assign y15 = ~n5192;
  assign y16 = ~n5223;
  assign y17 = ~n5243;
  assign y18 = ~n5264;
  assign y19 = ~n5283;
  assign y20 = ~n5298;
  assign y21 = ~n5314;
  assign y22 = ~n5325;
  assign y23 = n5335;
  assign y24 = n5336;
endmodule
