module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159;
  wire n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595, n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667, n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497, n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854, n44855, n44856, n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002, n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179, n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286, n45287, n45288, n45289, n45290, n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360, n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433, n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506, n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530, n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538, n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578, n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746, n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754, n45755, n45756, n45757, n45758, n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782, n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790, n45791, n45792, n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864, n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274, n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502, n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562, n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634, n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682, n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706, n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790, n46791, n46792, n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841, n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864, n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898, n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913, n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922, n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080, n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138, n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201, n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258, n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377, n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426, n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594, n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642, n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690, n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826, n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834, n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914, n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954, n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962, n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002, n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066, n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098, n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170, n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194, n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202, n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218, n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266, n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290, n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330, n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346, n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386, n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410, n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474, n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482, n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498, n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506, n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514, n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602, n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618, n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634, n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650, n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666, n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682, n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690, n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746, n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754, n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794, n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866, n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890, n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906, n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922, n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010, n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058, n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074, n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098, n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106, n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114, n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154, n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202, n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210, n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226, n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242, n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250, n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266, n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282, n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290, n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298, n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362, n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370, n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378, n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394, n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402, n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418, n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538, n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570, n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634, n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898, n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970, n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994, n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002, n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058, n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090, n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218, n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274, n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282, n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306, n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346, n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370, n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418, n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450, n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490, n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498, n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690, n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722, n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730, n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738, n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746, n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762, n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770, n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778, n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786, n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794, n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802, n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810, n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818, n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834, n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842, n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850, n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858, n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882, n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890, n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898, n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922, n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930, n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938, n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962, n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978, n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994, n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002, n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010, n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018, n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026, n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066, n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074, n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082, n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090, n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098, n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130, n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138, n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146, n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154, n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210, n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218, n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226, n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234, n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266, n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274, n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282, n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330, n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338, n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346, n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354, n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370, n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426, n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434, n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442, n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450, n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458, n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482, n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490, n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498, n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522, n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530, n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554, n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562, n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570, n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602, n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642, n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706, n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714, n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770, n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778, n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842, n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850, n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914, n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922, n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930, n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976, n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984, n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056, n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092, n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120, n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128, n52129, n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138, n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164, n52165, n52166, n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192, n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202, n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210, n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236, n52237, n52238, n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273, n52274, n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282, n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336, n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346, n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354, n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380, n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408, n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418, n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426, n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452, n52453, n52454, n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498, n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506, n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562, n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570, n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596, n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642, n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668, n52669, n52670, n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682, n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706, n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714, n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722, n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746, n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754, n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786, n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794, n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816, n52817, n52818, n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826, n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866, n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890, n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994, n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002, n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010, n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064, n53065, n53066, n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082, n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122, n53123, n53124, n53125, n53126, n53127, n53128, n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136, n53137, n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154, n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172, n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200, n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209, n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218, n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244, n53245, n53246, n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258, n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282, n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290, n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316, n53317, n53318, n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338, n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346, n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389, n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416, n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434, n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442, n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466, n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474, n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482, n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506, n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514, n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530, n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538, n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546, n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554, n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570, n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578, n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594, n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602, n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610, n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618, n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626, n53627, n53628, n53629, n53630, n53631, n53632, n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640, n53641, n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650, n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690, n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704, n53705, n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722, n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746, n53747, n53748, n53749, n53750, n53751, n53752, n53753, n53754, n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762, n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770, n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778, n53779, n53780, n53781, n53782, n53783, n53784, n53785, n53786, n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794, n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802, n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810, n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818, n53819, n53820, n53821, n53822, n53823, n53824, n53825, n53826, n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834, n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842, n53843, n53844, n53845, n53846, n53847, n53848, n53849, n53850, n53851, n53852, n53853, n53854, n53855, n53856, n53857, n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866, n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874, n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882, n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890, n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898, n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906, n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914, n53915, n53916, n53917, n53918, n53919, n53920, n53921, n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938, n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946, n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954, n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962, n53963, n53964, n53965, n53966, n53967, n53968, n53969, n53970, n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978, n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986, n53987, n53988, n53989, n53990, n53991, n53992, n53993, n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010, n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018, n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026, n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034, n54035, n54036, n54037, n54038, n54039, n54040, n54041, n54042, n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050, n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058, n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066, n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074, n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082, n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090, n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098, n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106, n54107, n54108, n54109, n54110, n54111, n54112, n54113, n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122, n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130, n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138, n54139, n54140, n54141, n54142, n54143, n54144, n54145, n54146, n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154, n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162, n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170, n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185, n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194, n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207, n54208, n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216, n54217, n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234, n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242, n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258, n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266, n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274, n54275, n54276, n54277, n54278, n54279, n54280, n54281, n54282, n54283, n54284, n54285, n54286, n54287, n54288, n54289, n54290, n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298, n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306, n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314, n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322, n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330, n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338, n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346, n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370, n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386, n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394, n54395, n54396, n54397, n54398, n54399, n54400, n54401, n54402, n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410, n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418, n54419, n54420, n54421, n54422, n54423, n54424, n54425, n54426, n54427, n54428, n54429, n54430, n54431, n54432, n54433, n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450, n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458, n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466, n54467, n54468, n54469, n54470, n54471, n54472, n54473, n54474, n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495, n54496, n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504, n54505, n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514, n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522, n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540, n54541, n54542, n54543, n54544, n54545, n54546, n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554, n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568, n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577, n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586, n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594, n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612, n54613, n54614, n54615, n54616, n54617, n54618, n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626, n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640, n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658, n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666, n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682, n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690, n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698, n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714, n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730, n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738, n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746, n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754, n54755, n54756, n54757, n54758, n54759, n54760, n54761, n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778, n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793, n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802, n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810, n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818, n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826, n54827, n54828, n54829, n54830, n54831, n54832, n54833, n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842, n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850, n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865, n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890, n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905, n54906, n54907, n54908, n54909, n54910, n54911, n54912, n54913, n54914, n54915, n54916, n54917, n54918, n54919, n54920, n54921, n54922, n54923, n54924, n54925, n54926, n54927, n54928, n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937, n54938, n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946, n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954, n54955, n54956, n54957, n54958, n54959, n54960, n54961, n54962, n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970, n54971, n54972, n54973, n54974, n54975, n54976, n54977, n54978, n54979, n54980, n54981, n54982, n54983, n54984, n54985, n54986, n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994, n54995, n54996, n54997, n54998, n54999, n55000, n55001, n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009, n55010, n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018, n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026, n55027, n55028, n55029, n55030, n55031, n55032, n55033, n55034, n55035, n55036, n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044, n55045, n55046, n55047, n55048, n55049, n55050, n55051, n55052, n55053, n55054, n55055, n55056, n55057, n55058, n55059, n55060, n55061, n55062, n55063, n55064, n55065, n55066, n55067, n55068, n55069, n55070, n55071, n55072, n55073, n55074, n55075, n55076, n55077, n55078, n55079, n55080, n55081, n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098, n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106, n55107, n55108, n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116, n55117, n55118, n55119, n55120, n55121, n55122, n55123, n55124, n55125, n55126, n55127, n55128, n55129, n55130, n55131, n55132, n55133, n55134, n55135, n55136, n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144, n55145, n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153, n55154, n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162, n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171, n55172, n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180, n55181, n55182, n55183, n55184, n55185, n55186, n55187, n55188, n55189, n55190, n55191, n55192, n55193, n55194, n55195, n55196, n55197, n55198, n55199, n55200, n55201, n55202, n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210, n55211, n55212, n55213, n55214, n55215, n55216, n55217, n55218, n55219, n55220, n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234, n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242, n55243, n55244, n55245, n55246, n55247, n55248, n55249, n55250, n55251, n55252, n55253, n55254, n55255, n55256, n55257, n55258, n55259, n55260, n55261, n55262, n55263, n55264, n55265, n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273, n55274, n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282, n55283, n55284, n55285, n55286, n55287, n55288, n55289, n55290, n55291, n55292, n55293, n55294, n55295, n55296, n55297, n55298, n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306, n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314, n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324, n55325, n55326, n55327, n55328, n55329, n55330, n55331, n55332, n55333, n55334, n55335, n55336, n55337, n55338, n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346, n55347, n55348, n55349, n55350, n55351, n55352, n55353, n55354, n55355, n55356, n55357, n55358, n55359, n55360, n55361, n55362, n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370, n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378, n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386, n55387, n55388, n55389, n55390, n55391, n55392, n55393, n55394, n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404, n55405, n55406, n55407, n55408, n55409, n55410, n55411, n55412, n55413, n55414, n55415, n55416, n55417, n55418, n55419, n55420, n55421, n55422, n55423, n55424, n55425, n55426, n55427, n55428, n55429, n55430, n55431, n55432, n55433, n55434, n55435, n55436, n55437, n55438, n55439, n55440, n55441, n55442, n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450, n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458, n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466, n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474, n55475, n55476, n55477, n55478, n55479, n55480, n55481, n55482, n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55490, n55491, n55492, n55493, n55494, n55495, n55496, n55497, n55498, n55499, n55500, n55501, n55502, n55503, n55504, n55505, n55506, n55507, n55508, n55509, n55510, n55511, n55512, n55513, n55514, n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522, n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530, n55531, n55532, n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540, n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548, n55549, n55550, n55551, n55552, n55553, n55554, n55555, n55556, n55557, n55558, n55559, n55560, n55561, n55562, n55563, n55564, n55565, n55566, n55567, n55568, n55569, n55570, n55571, n55572, n55573, n55574, n55575, n55576, n55577, n55578, n55579, n55580, n55581, n55582, n55583, n55584, n55585, n55586, n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594, n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602, n55603, n55604, n55605, n55606, n55607, n55608, n55609, n55610, n55611, n55612, n55613, n55614, n55615, n55616, n55617, n55618, n55619, n55620, n55621, n55622, n55623, n55624, n55625, n55626, n55627, n55628, n55629, n55630, n55631, n55632, n55633, n55634, n55635, n55636, n55637, n55638, n55639, n55640, n55641, n55642, n55643, n55644, n55645, n55646, n55647, n55648, n55649, n55650, n55651, n55652, n55653, n55654, n55655, n55656, n55657, n55658, n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666, n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674, n55675, n55676, n55677, n55678, n55679, n55680, n55681, n55682, n55683, n55684, n55685, n55686, n55687, n55688, n55689, n55690, n55691, n55692, n55693, n55694, n55695, n55696, n55697, n55698, n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706, n55707, n55708, n55709, n55710, n55711, n55712, n55713, n55714, n55715, n55716, n55717, n55718, n55719, n55720, n55721, n55722, n55723, n55724, n55725, n55726, n55727, n55728, n55729, n55730, n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738, n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746, n55747, n55748, n55749, n55750, n55751, n55752, n55753, n55754, n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762, n55763, n55764, n55765, n55766, n55767, n55768, n55769, n55770, n55771, n55772, n55773, n55774, n55775, n55776, n55777, n55778, n55779, n55780, n55781, n55782, n55783, n55784, n55785, n55786, n55787, n55788, n55789, n55790, n55791, n55792, n55793, n55794, n55795, n55796, n55797, n55798, n55799, n55800, n55801, n55802, n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810, n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818, n55819, n55820, n55821, n55822, n55823, n55824, n55825, n55826, n55827, n55828, n55829, n55830, n55831, n55832, n55833, n55834, n55835, n55836, n55837, n55838, n55839, n55840, n55841, n55842, n55843, n55844, n55845, n55846, n55847, n55848, n55849, n55850, n55851, n55852, n55853, n55854, n55855, n55856, n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864, n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872, n55873, n55874, n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882, n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890, n55891, n55892, n55893, n55894, n55895, n55896, n55897, n55898, n55899, n55900, n55901, n55902, n55903, n55904, n55905, n55906, n55907, n55908, n55909, n55910, n55911, n55912, n55913, n55914, n55915, n55916, n55917, n55918, n55919, n55920, n55921, n55922, n55923, n55924, n55925, n55926, n55927, n55928, n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936, n55937, n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945, n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954, n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962, n55963, n55964, n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972, n55973, n55974, n55975, n55976, n55977, n55978, n55979, n55980, n55981, n55982, n55983, n55984, n55985, n55986, n55987, n55988, n55989, n55990, n55991, n55992, n55993, n55994, n55995, n55996, n55997, n55998, n55999, n56000, n56001, n56002, n56003, n56004, n56005, n56006, n56007, n56008, n56009, n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017, n56018, n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026, n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034, n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042, n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050, n56051, n56052, n56053, n56054, n56055, n56056, n56057, n56058, n56059, n56060, n56061, n56062, n56063, n56064, n56065, n56066, n56067, n56068, n56069, n56070, n56071, n56072, n56073, n56074, n56075, n56076, n56077, n56078, n56079, n56080, n56081, n56082, n56083, n56084, n56085, n56086, n56087, n56088, n56089, n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098, n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106, n56107, n56108, n56109, n56110, n56111, n56112, n56113, n56114, n56115, n56116, n56117, n56118, n56119, n56120, n56121, n56122, n56123, n56124, n56125, n56126, n56127, n56128, n56129, n56130, n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138, n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146, n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162, n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170, n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178, n56179, n56180, n56181, n56182, n56183, n56184, n56185, n56186, n56187, n56188, n56189, n56190, n56191, n56192, n56193, n56194, n56195, n56196, n56197, n56198, n56199, n56200, n56201, n56202, n56203, n56204, n56205, n56206, n56207, n56208, n56209, n56210, n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218, n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226, n56227, n56228, n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242, n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250, n56251, n56252, n56253, n56254, n56255, n56256, n56257, n56258, n56259, n56260, n56261, n56262, n56263, n56264, n56265, n56266, n56267, n56268, n56269, n56270, n56271, n56272, n56273, n56274, n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282, n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290, n56291, n56292, n56293, n56294, n56295, n56296, n56297, n56298, n56299, n56300, n56301, n56302, n56303, n56304, n56305, n56306, n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314, n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322, n56323, n56324, n56325, n56326, n56327, n56328, n56329, n56330, n56331, n56332, n56333, n56334, n56335, n56336, n56337, n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345, n56346, n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354, n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362, n56363, n56364, n56365, n56366, n56367, n56368, n56369, n56370, n56371, n56372, n56373, n56374, n56375, n56376, n56377, n56378, n56379, n56380, n56381, n56382, n56383, n56384, n56385;
  assign n1277 = x499 ^ x147;
  assign n1278 = n1277 ^ x339;
  assign n1279 = n1278 ^ x83;
  assign n1385 = n1279 ^ x242;
  assign n1386 = n1385 ^ x434;
  assign n1387 = n1386 ^ x178;
  assign n2478 = n1387 ^ x337;
  assign n2475 = x434 ^ x82;
  assign n2476 = n2475 ^ x274;
  assign n2477 = n2476 ^ x18;
  assign n2479 = n2478 ^ n2477;
  assign n2480 = n2479 ^ x273;
  assign n1297 = x435 ^ x83;
  assign n1298 = n1297 ^ x275;
  assign n1299 = n1298 ^ x19;
  assign n1405 = n1299 ^ x178;
  assign n1406 = n1405 ^ x370;
  assign n1407 = n1406 ^ x114;
  assign n860 = x471 ^ x119;
  assign n861 = n860 ^ x311;
  assign n862 = n861 ^ x55;
  assign n926 = n862 ^ x214;
  assign n927 = n926 ^ x406;
  assign n928 = n927 ^ x150;
  assign n1010 = n928 ^ x309;
  assign n1011 = n1010 ^ x501;
  assign n1012 = n1011 ^ x245;
  assign n1097 = n1012 ^ x404;
  assign n1092 = x501 ^ x149;
  assign n1093 = n1092 ^ x341;
  assign n1094 = n1093 ^ x85;
  assign n1098 = n1097 ^ n1094;
  assign n1099 = n1098 ^ x340;
  assign n1190 = n1099 ^ x499;
  assign n1185 = n1094 ^ x244;
  assign n1186 = n1185 ^ x436;
  assign n1187 = n1186 ^ x180;
  assign n1191 = n1190 ^ n1187;
  assign n1192 = n1191 ^ x435;
  assign n1295 = n1279 ^ n1192;
  assign n1290 = n1187 ^ x339;
  assign n1285 = x436 ^ x84;
  assign n1286 = n1285 ^ x276;
  assign n1287 = n1286 ^ x20;
  assign n1291 = n1290 ^ n1287;
  assign n1292 = n1291 ^ x275;
  assign n1296 = n1295 ^ n1292;
  assign n1300 = n1299 ^ n1296;
  assign n1403 = n1387 ^ n1300;
  assign n1398 = n1292 ^ x434;
  assign n1393 = n1287 ^ x179;
  assign n1394 = n1393 ^ x371;
  assign n1395 = n1394 ^ x115;
  assign n1399 = n1398 ^ n1395;
  assign n1400 = n1399 ^ x370;
  assign n1404 = n1403 ^ n1400;
  assign n1408 = n1407 ^ n1404;
  assign n26509 = n2480 ^ n1408;
  assign n21350 = n2477 ^ n1400;
  assign n3012 = n1395 ^ x274;
  assign n3013 = n3012 ^ x466;
  assign n3014 = n3013 ^ x210;
  assign n21351 = n21350 ^ n3014;
  assign n21352 = n21351 ^ x465;
  assign n26510 = n26509 ^ n21352;
  assign n3159 = n1407 ^ x273;
  assign n3160 = n3159 ^ x465;
  assign n3161 = n3160 ^ x209;
  assign n26511 = n26510 ^ n3161;
  assign n2511 = n2480 ^ x432;
  assign n2508 = n2477 ^ x177;
  assign n2509 = n2508 ^ x369;
  assign n2510 = n2509 ^ x113;
  assign n2512 = n2511 ^ n2510;
  assign n2513 = n2512 ^ x368;
  assign n28581 = n26511 ^ n2513;
  assign n23484 = n21352 ^ n2510;
  assign n3018 = n3014 ^ x369;
  assign n1432 = x466 ^ x114;
  assign n1433 = n1432 ^ x306;
  assign n1434 = n1433 ^ x50;
  assign n3019 = n3018 ^ n1434;
  assign n3020 = n3019 ^ x305;
  assign n23485 = n23484 ^ n3020;
  assign n2430 = x465 ^ x113;
  assign n2431 = n2430 ^ x305;
  assign n2432 = n2431 ^ x49;
  assign n23486 = n23485 ^ n2432;
  assign n28582 = n28581 ^ n23486;
  assign n3171 = n3161 ^ x368;
  assign n3172 = n3171 ^ n2432;
  assign n3173 = n3172 ^ x304;
  assign n28583 = n28582 ^ n3173;
  assign n2462 = x432 ^ x80;
  assign n2463 = n2462 ^ x272;
  assign n2464 = n2463 ^ x16;
  assign n2553 = n2513 ^ n2464;
  assign n2550 = n2510 ^ x272;
  assign n2551 = n2550 ^ x464;
  assign n2552 = n2551 ^ x208;
  assign n2554 = n2553 ^ n2552;
  assign n2555 = n2554 ^ x463;
  assign n30994 = n28583 ^ n2555;
  assign n25442 = n23486 ^ n2552;
  assign n3027 = n3020 ^ x464;
  assign n3024 = n1434 ^ x209;
  assign n3025 = n3024 ^ x401;
  assign n3026 = n3025 ^ x145;
  assign n3028 = n3027 ^ n3026;
  assign n3029 = n3028 ^ x400;
  assign n25443 = n25442 ^ n3029;
  assign n2486 = n2432 ^ x208;
  assign n2487 = n2486 ^ x400;
  assign n2488 = n2487 ^ x144;
  assign n25444 = n25443 ^ n2488;
  assign n30995 = n30994 ^ n25444;
  assign n3183 = n3173 ^ x463;
  assign n3184 = n3183 ^ n2488;
  assign n3185 = n3184 ^ x399;
  assign n30996 = n30995 ^ n3185;
  assign n2527 = n2464 ^ x175;
  assign n2528 = n2527 ^ x367;
  assign n2529 = n2528 ^ x111;
  assign n2610 = n2555 ^ n2529;
  assign n2607 = n2552 ^ x367;
  assign n2604 = x464 ^ x112;
  assign n2605 = n2604 ^ x304;
  assign n2606 = n2605 ^ x48;
  assign n2608 = n2607 ^ n2606;
  assign n2609 = n2608 ^ x303;
  assign n2611 = n2610 ^ n2609;
  assign n2592 = x463 ^ x111;
  assign n2593 = n2592 ^ x303;
  assign n2594 = n2593 ^ x47;
  assign n2612 = n2611 ^ n2594;
  assign n33176 = n30996 ^ n2612;
  assign n27109 = n25444 ^ n2609;
  assign n3039 = n3029 ^ n2606;
  assign n3036 = n3026 ^ x304;
  assign n3037 = n3036 ^ x496;
  assign n3038 = n3037 ^ x240;
  assign n3040 = n3039 ^ n3038;
  assign n3041 = n3040 ^ x495;
  assign n27110 = n27109 ^ n3041;
  assign n2493 = n2488 ^ x303;
  assign n2494 = n2493 ^ x495;
  assign n2495 = n2494 ^ x239;
  assign n27111 = n27110 ^ n2495;
  assign n33177 = n33176 ^ n27111;
  assign n3195 = n3185 ^ n2594;
  assign n3196 = n3195 ^ n2495;
  assign n3197 = n3196 ^ x494;
  assign n33178 = n33177 ^ n3197;
  assign n2569 = n2529 ^ x270;
  assign n2570 = n2569 ^ x462;
  assign n2571 = n2570 ^ x206;
  assign n2658 = n2612 ^ n2571;
  assign n2655 = n2609 ^ x462;
  assign n2652 = n2606 ^ x207;
  assign n2653 = n2652 ^ x399;
  assign n2654 = n2653 ^ x143;
  assign n2656 = n2655 ^ n2654;
  assign n2657 = n2656 ^ x398;
  assign n2659 = n2658 ^ n2657;
  assign n2649 = n2594 ^ x206;
  assign n2650 = n2649 ^ x398;
  assign n2651 = n2650 ^ x142;
  assign n2660 = n2659 ^ n2651;
  assign n35483 = n33178 ^ n2660;
  assign n29403 = n27111 ^ n2657;
  assign n3056 = n3041 ^ n2654;
  assign n3048 = n3038 ^ x399;
  assign n1548 = x496 ^ x144;
  assign n1549 = n1548 ^ x336;
  assign n1550 = n1549 ^ x80;
  assign n3049 = n3048 ^ n1550;
  assign n3050 = n3049 ^ x335;
  assign n3057 = n3056 ^ n3050;
  assign n2533 = x495 ^ x143;
  assign n2534 = n2533 ^ x335;
  assign n2535 = n2534 ^ x79;
  assign n3058 = n3057 ^ n2535;
  assign n29404 = n29403 ^ n3058;
  assign n2532 = n2495 ^ x398;
  assign n2536 = n2535 ^ n2532;
  assign n2537 = n2536 ^ x334;
  assign n29405 = n29404 ^ n2537;
  assign n35484 = n35483 ^ n29405;
  assign n3207 = n3197 ^ n2651;
  assign n3208 = n3207 ^ n2537;
  assign n2770 = x494 ^ x142;
  assign n2771 = n2770 ^ x334;
  assign n2772 = n2771 ^ x78;
  assign n3209 = n3208 ^ n2772;
  assign n35485 = n35484 ^ n3209;
  assign n2620 = n2571 ^ x365;
  assign n2598 = x462 ^ x110;
  assign n2599 = n2598 ^ x302;
  assign n2600 = n2599 ^ x46;
  assign n2621 = n2620 ^ n2600;
  assign n2622 = n2621 ^ x301;
  assign n2715 = n2660 ^ n2622;
  assign n2709 = n2654 ^ x302;
  assign n2710 = n2709 ^ x494;
  assign n2711 = n2710 ^ x238;
  assign n2712 = n2711 ^ n2657;
  assign n2713 = n2712 ^ n2600;
  assign n2714 = n2713 ^ x493;
  assign n2716 = n2715 ^ n2714;
  assign n2706 = n2651 ^ x301;
  assign n2707 = n2706 ^ x493;
  assign n2708 = n2707 ^ x237;
  assign n2717 = n2716 ^ n2708;
  assign n37764 = n35485 ^ n2717;
  assign n3219 = n3209 ^ n2708;
  assign n2577 = n2537 ^ x493;
  assign n2574 = n2535 ^ x238;
  assign n2575 = n2574 ^ x430;
  assign n2576 = n2575 ^ x174;
  assign n2578 = n2577 ^ n2576;
  assign n2579 = n2578 ^ x429;
  assign n3220 = n3219 ^ n2579;
  assign n2836 = n2772 ^ x237;
  assign n2837 = n2836 ^ x429;
  assign n2838 = n2837 ^ x173;
  assign n3221 = n3220 ^ n2838;
  assign n37765 = n37764 ^ n3221;
  assign n31343 = n29405 ^ n2714;
  assign n3063 = n3058 ^ n2711;
  assign n3060 = n3050 ^ x494;
  assign n1551 = n1550 ^ x239;
  assign n1552 = n1551 ^ x431;
  assign n1553 = n1552 ^ x175;
  assign n3061 = n3060 ^ n1553;
  assign n3062 = n3061 ^ x430;
  assign n3064 = n3063 ^ n3062;
  assign n3065 = n3064 ^ n2576;
  assign n31344 = n31343 ^ n3065;
  assign n31345 = n31344 ^ n2579;
  assign n37766 = n37765 ^ n31345;
  assign n2677 = n2622 ^ x460;
  assign n2669 = n2600 ^ x205;
  assign n2670 = n2669 ^ x397;
  assign n2671 = n2670 ^ x141;
  assign n2678 = n2677 ^ n2671;
  assign n2679 = n2678 ^ x396;
  assign n2778 = n2717 ^ n2679;
  assign n2775 = n2714 ^ n2671;
  assign n2769 = n2711 ^ x397;
  assign n2773 = n2772 ^ n2769;
  assign n2774 = n2773 ^ x333;
  assign n2776 = n2775 ^ n2774;
  assign n2625 = x493 ^ x141;
  assign n2626 = n2625 ^ x333;
  assign n2627 = n2626 ^ x77;
  assign n2777 = n2776 ^ n2627;
  assign n2779 = n2778 ^ n2777;
  assign n2766 = n2708 ^ x396;
  assign n2767 = n2766 ^ n2627;
  assign n2768 = n2767 ^ x332;
  assign n2780 = n2779 ^ n2768;
  assign n39938 = n37766 ^ n2780;
  assign n34000 = n31345 ^ n2777;
  assign n3075 = n3065 ^ n2774;
  assign n3072 = n3062 ^ n2772;
  assign n1554 = n1553 ^ x334;
  assign n1513 = x431 ^ x79;
  assign n1514 = n1513 ^ x271;
  assign n1515 = n1514 ^ x15;
  assign n1555 = n1554 ^ n1515;
  assign n1556 = n1555 ^ x270;
  assign n3073 = n3072 ^ n1556;
  assign n2630 = x430 ^ x78;
  assign n2631 = n2630 ^ x270;
  assign n2632 = n2631 ^ x14;
  assign n3074 = n3073 ^ n2632;
  assign n3076 = n3075 ^ n3074;
  assign n2629 = n2576 ^ x333;
  assign n2633 = n2632 ^ n2629;
  assign n2634 = n2633 ^ x269;
  assign n3077 = n3076 ^ n2634;
  assign n34001 = n34000 ^ n3077;
  assign n2628 = n2627 ^ n2579;
  assign n2635 = n2634 ^ n2628;
  assign n1560 = x429 ^ x77;
  assign n1561 = n1560 ^ x269;
  assign n1562 = n1561 ^ x13;
  assign n2636 = n2635 ^ n1562;
  assign n34002 = n34001 ^ n2636;
  assign n39939 = n39938 ^ n34002;
  assign n3231 = n3221 ^ n2768;
  assign n3232 = n3231 ^ n2636;
  assign n2904 = n2838 ^ x332;
  assign n2905 = n2904 ^ n1562;
  assign n2906 = n2905 ^ x268;
  assign n3233 = n3232 ^ n2906;
  assign n39940 = n39939 ^ n3233;
  assign n1571 = x460 ^ x108;
  assign n1572 = n1571 ^ x300;
  assign n1573 = n1572 ^ x44;
  assign n2734 = n2679 ^ n1573;
  assign n2726 = x492 ^ x300;
  assign n2727 = n2726 ^ n2671;
  assign n2728 = n2727 ^ x236;
  assign n2735 = n2734 ^ n2728;
  assign n2736 = n2735 ^ x491;
  assign n2844 = n2780 ^ n2736;
  assign n2841 = n2777 ^ n2728;
  assign n2835 = n2774 ^ x492;
  assign n2839 = n2838 ^ n2835;
  assign n2840 = n2839 ^ x428;
  assign n2842 = n2841 ^ n2840;
  assign n2682 = n2627 ^ x236;
  assign n2683 = n2682 ^ x428;
  assign n2684 = n2683 ^ x172;
  assign n2843 = n2842 ^ n2684;
  assign n2845 = n2844 ^ n2843;
  assign n2832 = n2768 ^ x491;
  assign n2833 = n2832 ^ n2684;
  assign n2834 = n2833 ^ x427;
  assign n2846 = n2845 ^ n2834;
  assign n42164 = n39940 ^ n2846;
  assign n36310 = n34002 ^ n2843;
  assign n3087 = n3077 ^ n2840;
  assign n3084 = n3074 ^ n2838;
  assign n1557 = n1556 ^ x429;
  assign n1516 = n1515 ^ x174;
  assign n1517 = n1516 ^ x366;
  assign n1518 = n1517 ^ x110;
  assign n1558 = n1557 ^ n1518;
  assign n1559 = n1558 ^ x365;
  assign n3085 = n3084 ^ n1559;
  assign n2687 = n2632 ^ x173;
  assign n2688 = n2687 ^ x365;
  assign n2689 = n2688 ^ x109;
  assign n3086 = n3085 ^ n2689;
  assign n3088 = n3087 ^ n3086;
  assign n2686 = n2634 ^ x428;
  assign n2690 = n2689 ^ n2686;
  assign n2691 = n2690 ^ x364;
  assign n3089 = n3088 ^ n2691;
  assign n36311 = n36310 ^ n3089;
  assign n2685 = n2684 ^ n2636;
  assign n2692 = n2691 ^ n2685;
  assign n1566 = n1562 ^ x172;
  assign n1567 = n1566 ^ x364;
  assign n1568 = n1567 ^ x108;
  assign n2693 = n2692 ^ n1568;
  assign n36312 = n36311 ^ n2693;
  assign n42165 = n42164 ^ n36312;
  assign n30147 = n3233 ^ n2834;
  assign n30148 = n30147 ^ n2693;
  assign n2977 = n2906 ^ x427;
  assign n2978 = n2977 ^ n1568;
  assign n2979 = n2978 ^ x363;
  assign n30149 = n30148 ^ n2979;
  assign n42166 = n42165 ^ n30149;
  assign n2792 = n2728 ^ x395;
  assign n2784 = x492 ^ x140;
  assign n2785 = n2784 ^ x332;
  assign n2786 = n2785 ^ x76;
  assign n2793 = n2792 ^ n2786;
  assign n2794 = n2793 ^ x331;
  assign n2909 = n2843 ^ n2794;
  assign n2903 = n2840 ^ n2786;
  assign n2907 = n2906 ^ n2903;
  assign n2742 = x428 ^ x76;
  assign n2743 = n2742 ^ x268;
  assign n2744 = n2743 ^ x12;
  assign n2908 = n2907 ^ n2744;
  assign n2910 = n2909 ^ n2908;
  assign n2748 = n2684 ^ x331;
  assign n2749 = n2748 ^ n2744;
  assign n2750 = n2749 ^ x267;
  assign n2911 = n2910 ^ n2750;
  assign n2912 = n2911 ^ n2846;
  assign n1498 = x491 ^ x139;
  assign n1499 = n1498 ^ x331;
  assign n1500 = n1499 ^ x75;
  assign n2900 = n2834 ^ n1500;
  assign n2901 = n2900 ^ n2750;
  assign n2897 = x427 ^ x267;
  assign n2898 = n2897 ^ x75;
  assign n2899 = n2898 ^ x11;
  assign n2902 = n2901 ^ n2899;
  assign n2913 = n2912 ^ n2902;
  assign n1580 = n1573 ^ x203;
  assign n1581 = n1580 ^ x395;
  assign n1582 = n1581 ^ x139;
  assign n2800 = n2736 ^ n1582;
  assign n2801 = n2800 ^ n2794;
  assign n2802 = n2801 ^ n1500;
  assign n2914 = n2913 ^ n2802;
  assign n44276 = n42166 ^ n2914;
  assign n38518 = n36312 ^ n2911;
  assign n2751 = n2750 ^ n2693;
  assign n2745 = n2744 ^ n2691;
  assign n2739 = n2689 ^ x268;
  assign n2740 = n2739 ^ x460;
  assign n2741 = n2740 ^ x204;
  assign n2746 = n2745 ^ n2741;
  assign n2747 = n2746 ^ x459;
  assign n2752 = n2751 ^ n2747;
  assign n1575 = n1568 ^ x267;
  assign n1576 = n1575 ^ x459;
  assign n1577 = n1576 ^ x203;
  assign n2753 = n2752 ^ n1577;
  assign n38519 = n38518 ^ n2753;
  assign n3099 = n3089 ^ n2908;
  assign n3096 = n3086 ^ n2906;
  assign n1563 = n1562 ^ n1559;
  assign n1519 = n1518 ^ x269;
  assign n1520 = n1519 ^ x461;
  assign n1521 = n1520 ^ x205;
  assign n1564 = n1563 ^ n1521;
  assign n1565 = n1564 ^ x460;
  assign n3097 = n3096 ^ n1565;
  assign n3098 = n3097 ^ n2741;
  assign n3100 = n3099 ^ n3098;
  assign n3101 = n3100 ^ n2747;
  assign n38520 = n38519 ^ n3101;
  assign n44277 = n44276 ^ n38520;
  assign n32260 = n30149 ^ n2902;
  assign n32261 = n32260 ^ n2753;
  assign n3120 = n2979 ^ n2899;
  assign n3121 = n3120 ^ n1577;
  assign n3122 = n3121 ^ x458;
  assign n32262 = n32261 ^ n3122;
  assign n44278 = n44277 ^ n32262;
  assign n1589 = n1582 ^ x298;
  assign n1590 = n1589 ^ x490;
  assign n1591 = n1590 ^ x234;
  assign n2866 = n2802 ^ n1591;
  assign n2858 = n2794 ^ x490;
  assign n2850 = n2786 ^ x235;
  assign n2851 = n2850 ^ x427;
  assign n2852 = n2851 ^ x171;
  assign n2859 = n2858 ^ n2852;
  assign n2860 = n2859 ^ x426;
  assign n2867 = n2866 ^ n2860;
  assign n1504 = n1500 ^ x234;
  assign n1505 = n1504 ^ x426;
  assign n1506 = n1505 ^ x170;
  assign n2868 = n2867 ^ n1506;
  assign n2985 = n2914 ^ n2868;
  assign n2982 = n2911 ^ n2860;
  assign n2976 = n2908 ^ n2852;
  assign n2980 = n2979 ^ n2976;
  assign n2806 = n2744 ^ x171;
  assign n2807 = n2806 ^ x363;
  assign n2808 = n2807 ^ x107;
  assign n2981 = n2980 ^ n2808;
  assign n2983 = n2982 ^ n2981;
  assign n2805 = n2750 ^ x426;
  assign n2809 = n2808 ^ n2805;
  assign n2810 = n2809 ^ x362;
  assign n2984 = n2983 ^ n2810;
  assign n2986 = n2985 ^ n2984;
  assign n2973 = n2902 ^ n1506;
  assign n2974 = n2973 ^ n2810;
  assign n2970 = n2899 ^ x170;
  assign n2971 = n2970 ^ x362;
  assign n2972 = n2971 ^ x106;
  assign n2975 = n2974 ^ n2972;
  assign n2987 = n2986 ^ n2975;
  assign n46334 = n44278 ^ n2987;
  assign n40735 = n38520 ^ n2984;
  assign n3111 = n3101 ^ n2981;
  assign n3108 = n3098 ^ n2979;
  assign n1569 = n1568 ^ n1565;
  assign n1522 = n1521 ^ x364;
  assign n1488 = x461 ^ x109;
  assign n1489 = n1488 ^ x301;
  assign n1490 = n1489 ^ x45;
  assign n1523 = n1522 ^ n1490;
  assign n1524 = n1523 ^ x300;
  assign n1570 = n1569 ^ n1524;
  assign n1574 = n1573 ^ n1570;
  assign n3109 = n3108 ^ n1574;
  assign n2813 = n2741 ^ x363;
  assign n2814 = n2813 ^ n1573;
  assign n2815 = n2814 ^ x299;
  assign n3110 = n3109 ^ n2815;
  assign n3112 = n3111 ^ n3110;
  assign n2812 = n2808 ^ n2747;
  assign n2816 = n2815 ^ n2812;
  assign n1509 = x459 ^ x107;
  assign n1510 = n1509 ^ x299;
  assign n1511 = n1510 ^ x43;
  assign n2817 = n2816 ^ n1511;
  assign n3113 = n3112 ^ n2817;
  assign n40736 = n40735 ^ n3113;
  assign n2811 = n2810 ^ n2753;
  assign n2818 = n2817 ^ n2811;
  assign n1584 = n1577 ^ x362;
  assign n1585 = n1584 ^ n1511;
  assign n1586 = n1585 ^ x298;
  assign n2819 = n2818 ^ n1586;
  assign n40737 = n40736 ^ n2819;
  assign n46335 = n46334 ^ n40737;
  assign n34724 = n32262 ^ n2975;
  assign n34725 = n34724 ^ n2819;
  assign n23539 = n3122 ^ n2972;
  assign n23540 = n23539 ^ n1586;
  assign n2942 = x458 ^ x106;
  assign n2943 = n2942 ^ x298;
  assign n2944 = n2943 ^ x42;
  assign n23541 = n23540 ^ n2944;
  assign n34726 = n34725 ^ n23541;
  assign n46336 = n46335 ^ n34726;
  assign n1598 = n1591 ^ x393;
  assign n1535 = x490 ^ x138;
  assign n1536 = n1535 ^ x330;
  assign n1537 = n1536 ^ x74;
  assign n1599 = n1598 ^ n1537;
  assign n1600 = n1599 ^ x329;
  assign n2935 = n2868 ^ n1600;
  assign n2925 = n2860 ^ n1537;
  assign n2918 = n2852 ^ x330;
  assign n2919 = n2918 ^ n2899;
  assign n2920 = n2919 ^ x266;
  assign n2926 = n2925 ^ n2920;
  assign n1633 = x426 ^ x74;
  assign n1634 = n1633 ^ x266;
  assign n1635 = n1634 ^ x10;
  assign n2927 = n2926 ^ n1635;
  assign n2936 = n2935 ^ n2927;
  assign n1632 = n1506 ^ x329;
  assign n1636 = n1635 ^ n1632;
  assign n1637 = n1636 ^ x265;
  assign n2937 = n2936 ^ n1637;
  assign n38597 = n2987 ^ n2937;
  assign n26496 = n2975 ^ n1637;
  assign n2874 = n2810 ^ n1635;
  assign n2871 = n2808 ^ x266;
  assign n2872 = n2871 ^ x458;
  assign n2873 = n2872 ^ x202;
  assign n2875 = n2874 ^ n2873;
  assign n2876 = n2875 ^ x457;
  assign n26497 = n26496 ^ n2876;
  assign n16609 = n2972 ^ x265;
  assign n16610 = n16609 ^ x457;
  assign n16611 = n16610 ^ x201;
  assign n26498 = n26497 ^ n16611;
  assign n38598 = n38597 ^ n26498;
  assign n32240 = n2984 ^ n2927;
  assign n3126 = n2981 ^ n2920;
  assign n3127 = n3126 ^ n3122;
  assign n3128 = n3127 ^ n2873;
  assign n32241 = n32240 ^ n3128;
  assign n32242 = n32241 ^ n2876;
  assign n38599 = n38598 ^ n32242;
  assign n48401 = n46336 ^ n38599;
  assign n42883 = n40737 ^ n32242;
  assign n3129 = n3128 ^ n3113;
  assign n2881 = n2873 ^ n2817;
  assign n2878 = n2815 ^ x458;
  assign n2879 = n2878 ^ n1582;
  assign n2880 = n2879 ^ x394;
  assign n2882 = n2881 ^ n2880;
  assign n1530 = n1511 ^ x202;
  assign n1531 = n1530 ^ x394;
  assign n1532 = n1531 ^ x138;
  assign n2883 = n2882 ^ n1532;
  assign n3130 = n3129 ^ n2883;
  assign n3123 = n3122 ^ n3110;
  assign n1578 = n1577 ^ n1574;
  assign n1525 = n1524 ^ x459;
  assign n1491 = n1490 ^ x204;
  assign n1492 = n1491 ^ x396;
  assign n1493 = n1492 ^ x140;
  assign n1526 = n1525 ^ n1493;
  assign n1527 = n1526 ^ x395;
  assign n1579 = n1578 ^ n1527;
  assign n1583 = n1582 ^ n1579;
  assign n3124 = n3123 ^ n1583;
  assign n3125 = n3124 ^ n2880;
  assign n3131 = n3130 ^ n3125;
  assign n42884 = n42883 ^ n3131;
  assign n2877 = n2876 ^ n2819;
  assign n2884 = n2883 ^ n2877;
  assign n1593 = n1586 ^ x457;
  assign n1594 = n1593 ^ n1532;
  assign n1595 = n1594 ^ x393;
  assign n2885 = n2884 ^ n1595;
  assign n42885 = n42884 ^ n2885;
  assign n48402 = n48401 ^ n42885;
  assign n36960 = n34726 ^ n26498;
  assign n25500 = n23541 ^ n16611;
  assign n25501 = n25500 ^ n1595;
  assign n15632 = n2944 ^ x201;
  assign n15633 = n15632 ^ x393;
  assign n15634 = n15633 ^ x137;
  assign n25502 = n25501 ^ n15634;
  assign n36961 = n36960 ^ n25502;
  assign n36962 = n36961 ^ n2885;
  assign n48403 = n48402 ^ n36962;
  assign n1610 = n1600 ^ x488;
  assign n1544 = n1537 ^ x233;
  assign n1545 = n1544 ^ x425;
  assign n1546 = n1545 ^ x169;
  assign n1611 = n1610 ^ n1546;
  assign n1612 = n1611 ^ x424;
  assign n3007 = n2937 ^ n1612;
  assign n2999 = n2927 ^ n1546;
  assign n2991 = n2920 ^ x425;
  assign n2992 = n2991 ^ n2972;
  assign n2993 = n2992 ^ x361;
  assign n3000 = n2999 ^ n2993;
  assign n1675 = n1635 ^ x169;
  assign n1676 = n1675 ^ x361;
  assign n1677 = n1676 ^ x105;
  assign n3001 = n3000 ^ n1677;
  assign n3008 = n3007 ^ n3001;
  assign n1674 = n1637 ^ x424;
  assign n1678 = n1677 ^ n1674;
  assign n1679 = n1678 ^ x360;
  assign n3009 = n3008 ^ n1679;
  assign n40729 = n38599 ^ n3009;
  assign n34719 = n32242 ^ n3001;
  assign n28564 = n3128 ^ n2993;
  assign n28565 = n28564 ^ n23541;
  assign n2941 = n2873 ^ x361;
  assign n2945 = n2944 ^ n2941;
  assign n2946 = n2945 ^ x297;
  assign n28566 = n28565 ^ n2946;
  assign n34720 = n34719 ^ n28566;
  assign n2940 = n2876 ^ n1677;
  assign n2947 = n2946 ^ n2940;
  assign n1602 = x457 ^ x297;
  assign n1603 = n1602 ^ x105;
  assign n1604 = n1603 ^ x41;
  assign n2948 = n2947 ^ n1604;
  assign n34721 = n34720 ^ n2948;
  assign n40730 = n40729 ^ n34721;
  assign n28559 = n26498 ^ n1679;
  assign n28560 = n28559 ^ n2948;
  assign n18663 = n16611 ^ x360;
  assign n18664 = n18663 ^ n1604;
  assign n18665 = n18664 ^ x296;
  assign n28561 = n28560 ^ n18665;
  assign n40731 = n40730 ^ n28561;
  assign n50481 = n48403 ^ n40731;
  assign n44936 = n42885 ^ n34721;
  assign n39318 = n28566 ^ n3131;
  assign n33154 = n23541 ^ n3125;
  assign n1587 = n1586 ^ n1583;
  assign n1494 = n1493 ^ x299;
  assign n1495 = n1494 ^ x491;
  assign n1496 = n1495 ^ x235;
  assign n1512 = n1511 ^ n1496;
  assign n1528 = n1527 ^ n1512;
  assign n1529 = n1528 ^ x490;
  assign n1588 = n1587 ^ n1529;
  assign n1592 = n1591 ^ n1588;
  assign n33155 = n33154 ^ n1592;
  assign n2951 = n2944 ^ n2880;
  assign n2952 = n2951 ^ n1591;
  assign n2953 = n2952 ^ x489;
  assign n33156 = n33155 ^ n2953;
  assign n39319 = n39318 ^ n33156;
  assign n2950 = n2946 ^ n2883;
  assign n2954 = n2953 ^ n2950;
  assign n1539 = n1532 ^ x297;
  assign n1540 = n1539 ^ x489;
  assign n1541 = n1540 ^ x233;
  assign n2955 = n2954 ^ n1541;
  assign n39320 = n39319 ^ n2955;
  assign n44937 = n44936 ^ n39320;
  assign n2949 = n2948 ^ n2885;
  assign n2956 = n2955 ^ n2949;
  assign n1605 = n1604 ^ n1595;
  assign n1606 = n1605 ^ n1541;
  assign n1607 = n1606 ^ x488;
  assign n2957 = n2956 ^ n1607;
  assign n44938 = n44937 ^ n2957;
  assign n50482 = n50481 ^ n44938;
  assign n39215 = n36962 ^ n28561;
  assign n39216 = n39215 ^ n2957;
  assign n27249 = n25502 ^ n18665;
  assign n27250 = n27249 ^ n1607;
  assign n17353 = n15634 ^ x296;
  assign n17354 = n17353 ^ x488;
  assign n17355 = n17354 ^ x232;
  assign n27251 = n27250 ^ n17355;
  assign n39217 = n39216 ^ n27251;
  assign n50483 = n50482 ^ n39217;
  assign n1625 = x328 ^ x136;
  assign n1626 = n1625 ^ x488;
  assign n1627 = n1626 ^ x72;
  assign n1652 = n1627 ^ n1612;
  assign n1644 = n1546 ^ x328;
  assign n1639 = x425 ^ x73;
  assign n1640 = n1639 ^ x265;
  assign n1641 = n1640 ^ x9;
  assign n1645 = n1644 ^ n1641;
  assign n1646 = n1645 ^ x264;
  assign n1653 = n1652 ^ n1646;
  assign n1649 = x424 ^ x72;
  assign n1650 = n1649 ^ x264;
  assign n1651 = n1650 ^ x8;
  assign n1654 = n1653 ^ n1651;
  assign n32231 = n3009 ^ n1654;
  assign n26643 = n3001 ^ n1646;
  assign n21695 = n2993 ^ n1641;
  assign n21696 = n21695 ^ n16611;
  assign n21697 = n21696 ^ x456;
  assign n26644 = n26643 ^ n21697;
  assign n1736 = n1677 ^ x264;
  assign n1737 = n1736 ^ x456;
  assign n1738 = n1737 ^ x200;
  assign n26645 = n26644 ^ n1738;
  assign n32232 = n32231 ^ n26645;
  assign n1735 = n1679 ^ n1651;
  assign n1739 = n1738 ^ n1735;
  assign n1740 = n1739 ^ x455;
  assign n32233 = n32232 ^ n1740;
  assign n42960 = n40731 ^ n32233;
  assign n36955 = n34721 ^ n26645;
  assign n31048 = n28566 ^ n21697;
  assign n31049 = n31048 ^ n25502;
  assign n20375 = n2946 ^ x456;
  assign n20376 = n20375 ^ n15634;
  assign n20377 = n20376 ^ x392;
  assign n31050 = n31049 ^ n20377;
  assign n36956 = n36955 ^ n31050;
  assign n25430 = n2948 ^ n1738;
  assign n25431 = n25430 ^ n20377;
  assign n1614 = n1604 ^ x200;
  assign n1615 = n1614 ^ x392;
  assign n1616 = n1615 ^ x136;
  assign n25432 = n25431 ^ n1616;
  assign n36957 = n36956 ^ n25432;
  assign n42961 = n42960 ^ n36957;
  assign n31063 = n28561 ^ n1740;
  assign n31064 = n31063 ^ n25432;
  assign n20526 = n18665 ^ x455;
  assign n20527 = n20526 ^ n1616;
  assign n20528 = n20527 ^ x391;
  assign n31065 = n31064 ^ n20528;
  assign n42962 = n42961 ^ n31065;
  assign n52561 = n50483 ^ n42962;
  assign n47075 = n44938 ^ n36957;
  assign n41442 = n39320 ^ n31050;
  assign n35470 = n33156 ^ n25502;
  assign n1596 = n1595 ^ n1592;
  assign n1533 = n1532 ^ n1529;
  assign n1497 = n1496 ^ x394;
  assign n1501 = n1500 ^ n1497;
  assign n1502 = n1501 ^ x330;
  assign n1534 = n1533 ^ n1502;
  assign n1538 = n1537 ^ n1534;
  assign n1597 = n1596 ^ n1538;
  assign n1601 = n1600 ^ n1597;
  assign n35471 = n35470 ^ n1601;
  assign n24024 = n15634 ^ n2953;
  assign n24025 = n24024 ^ n1600;
  assign n1619 = x489 ^ x137;
  assign n1620 = n1619 ^ x329;
  assign n1621 = n1620 ^ x73;
  assign n24026 = n24025 ^ n1621;
  assign n35472 = n35471 ^ n24026;
  assign n41443 = n41442 ^ n35472;
  assign n29389 = n20377 ^ n2955;
  assign n29390 = n29389 ^ n24026;
  assign n1618 = n1541 ^ x392;
  assign n1622 = n1621 ^ n1618;
  assign n1623 = n1622 ^ x328;
  assign n29391 = n29390 ^ n1623;
  assign n41444 = n41443 ^ n29391;
  assign n47076 = n47075 ^ n41444;
  assign n35465 = n25432 ^ n2957;
  assign n35466 = n35465 ^ n29391;
  assign n1617 = n1616 ^ n1607;
  assign n1624 = n1623 ^ n1617;
  assign n1628 = n1627 ^ n1624;
  assign n35467 = n35466 ^ n1628;
  assign n47077 = n47076 ^ n35467;
  assign n52562 = n52561 ^ n47077;
  assign n41437 = n39217 ^ n31065;
  assign n41438 = n41437 ^ n35467;
  assign n29384 = n27251 ^ n20528;
  assign n29385 = n29384 ^ n1628;
  assign n19278 = n17355 ^ x391;
  assign n19279 = n19278 ^ n1627;
  assign n19280 = n19279 ^ x327;
  assign n29386 = n29385 ^ n19280;
  assign n41439 = n41438 ^ n29386;
  assign n52563 = n52562 ^ n41439;
  assign n1667 = x423 ^ x231;
  assign n1668 = n1667 ^ n1627;
  assign n1669 = n1668 ^ x167;
  assign n1694 = n1669 ^ n1654;
  assign n1686 = n1646 ^ x423;
  assign n1681 = n1641 ^ x168;
  assign n1682 = n1681 ^ x360;
  assign n1683 = n1682 ^ x104;
  assign n1687 = n1686 ^ n1683;
  assign n1688 = n1687 ^ x359;
  assign n1695 = n1694 ^ n1688;
  assign n1691 = n1651 ^ x167;
  assign n1692 = n1691 ^ x359;
  assign n1693 = n1692 ^ x103;
  assign n1696 = n1695 ^ n1693;
  assign n34837 = n32233 ^ n1696;
  assign n28554 = n26645 ^ n1688;
  assign n23466 = n21697 ^ n1683;
  assign n23467 = n23466 ^ n18665;
  assign n1778 = x456 ^ x104;
  assign n1779 = n1778 ^ x296;
  assign n1780 = n1779 ^ x40;
  assign n23468 = n23467 ^ n1780;
  assign n28555 = n28554 ^ n23468;
  assign n1777 = n1738 ^ x359;
  assign n1781 = n1780 ^ n1777;
  assign n1782 = n1781 ^ x295;
  assign n28556 = n28555 ^ n1782;
  assign n34838 = n34837 ^ n28556;
  assign n1776 = n1740 ^ n1693;
  assign n1783 = n1782 ^ n1776;
  assign n1770 = x455 ^ x39;
  assign n1771 = n1770 ^ x295;
  assign n1772 = n1771 ^ x103;
  assign n1784 = n1783 ^ n1772;
  assign n34839 = n34838 ^ n1784;
  assign n44930 = n42962 ^ n34839;
  assign n39210 = n36957 ^ n28556;
  assign n33147 = n31050 ^ n23468;
  assign n33148 = n33147 ^ n27251;
  assign n22089 = n20377 ^ n1780;
  assign n22090 = n22089 ^ n17355;
  assign n22091 = n22090 ^ x487;
  assign n33149 = n33148 ^ n22091;
  assign n39211 = n39210 ^ n33149;
  assign n27419 = n25432 ^ n1782;
  assign n27420 = n27419 ^ n22091;
  assign n1656 = n1616 ^ x295;
  assign n1657 = n1656 ^ x487;
  assign n1658 = n1657 ^ x231;
  assign n27421 = n27420 ^ n1658;
  assign n39212 = n39211 ^ n27421;
  assign n44931 = n44930 ^ n39212;
  assign n33142 = n31065 ^ n1784;
  assign n33143 = n33142 ^ n27421;
  assign n22230 = n20528 ^ n1772;
  assign n22231 = n22230 ^ n1658;
  assign n22232 = n22231 ^ x486;
  assign n33144 = n33143 ^ n22232;
  assign n44932 = n44931 ^ n33144;
  assign n54614 = n52563 ^ n44932;
  assign n49155 = n47077 ^ n39212;
  assign n43649 = n41444 ^ n33149;
  assign n37752 = n35472 ^ n27251;
  assign n1608 = n1607 ^ n1601;
  assign n1542 = n1541 ^ n1538;
  assign n1503 = n1502 ^ x489;
  assign n1507 = n1506 ^ n1503;
  assign n1508 = n1507 ^ x425;
  assign n1543 = n1542 ^ n1508;
  assign n1547 = n1546 ^ n1543;
  assign n1609 = n1608 ^ n1547;
  assign n1613 = n1612 ^ n1609;
  assign n37753 = n37752 ^ n1613;
  assign n26121 = n24026 ^ n17355;
  assign n26122 = n26121 ^ n1612;
  assign n1661 = n1621 ^ x232;
  assign n1662 = n1661 ^ x424;
  assign n1663 = n1662 ^ x168;
  assign n26123 = n26122 ^ n1663;
  assign n37754 = n37753 ^ n26123;
  assign n43650 = n43649 ^ n37754;
  assign n31786 = n29391 ^ n22091;
  assign n31787 = n31786 ^ n26123;
  assign n1660 = n1623 ^ x487;
  assign n1664 = n1663 ^ n1660;
  assign n1665 = n1664 ^ x423;
  assign n31788 = n31787 ^ n1665;
  assign n43651 = n43650 ^ n31788;
  assign n49156 = n49155 ^ n43651;
  assign n37747 = n35467 ^ n27421;
  assign n37748 = n37747 ^ n31788;
  assign n1659 = n1658 ^ n1628;
  assign n1666 = n1665 ^ n1659;
  assign n1670 = n1669 ^ n1666;
  assign n37749 = n37748 ^ n1670;
  assign n49157 = n49156 ^ n37749;
  assign n54615 = n54614 ^ n49157;
  assign n43635 = n41439 ^ n33144;
  assign n43636 = n43635 ^ n37749;
  assign n31781 = n29386 ^ n22232;
  assign n31782 = n31781 ^ n1670;
  assign n21117 = n19280 ^ x486;
  assign n21118 = n21117 ^ n1669;
  assign n21119 = n21118 ^ x422;
  assign n31783 = n31782 ^ n21119;
  assign n43637 = n43636 ^ n31783;
  assign n54616 = n54615 ^ n43637;
  assign n2211 = x450 ^ x98;
  assign n2212 = n2211 ^ x290;
  assign n2213 = n2212 ^ x34;
  assign n2313 = n2213 ^ x193;
  assign n2314 = n2313 ^ x385;
  assign n2315 = n2314 ^ x129;
  assign n16887 = n2315 ^ x288;
  assign n16888 = n16887 ^ x480;
  assign n16889 = n16888 ^ x224;
  assign n1806 = x422 ^ x70;
  assign n1807 = n1806 ^ x262;
  assign n1808 = n1807 ^ x6;
  assign n1872 = n1808 ^ x165;
  assign n1873 = n1872 ^ x357;
  assign n1874 = n1873 ^ x101;
  assign n1944 = n1874 ^ x260;
  assign n1945 = n1944 ^ x452;
  assign n1946 = n1945 ^ x196;
  assign n2031 = n1946 ^ x355;
  assign n1900 = x452 ^ x36;
  assign n1901 = n1900 ^ x100;
  assign n1902 = n1901 ^ x292;
  assign n2032 = n2031 ^ n1902;
  assign n2033 = n2032 ^ x291;
  assign n2122 = n2033 ^ x450;
  assign n1968 = n1902 ^ x195;
  assign n1969 = n1968 ^ x387;
  assign n1970 = n1969 ^ x131;
  assign n2123 = n2122 ^ n1970;
  assign n2124 = n2123 ^ x386;
  assign n2218 = n2213 ^ n2124;
  assign n2062 = n1970 ^ x290;
  assign n2063 = n2062 ^ x482;
  assign n2064 = n2063 ^ x226;
  assign n2219 = n2218 ^ n2064;
  assign n2220 = n2219 ^ x481;
  assign n2316 = n2315 ^ n2220;
  assign n2155 = n2064 ^ x385;
  assign n2147 = x482 ^ x130;
  assign n2148 = n2147 ^ x322;
  assign n2149 = n2148 ^ x66;
  assign n2156 = n2155 ^ n2149;
  assign n2157 = n2156 ^ x321;
  assign n2317 = n2316 ^ n2157;
  assign n2306 = x481 ^ x129;
  assign n2307 = n2306 ^ x321;
  assign n2308 = n2307 ^ x65;
  assign n2318 = n2317 ^ n2308;
  assign n25771 = n16889 ^ n2318;
  assign n2249 = n2157 ^ x480;
  assign n2239 = x417 ^ x225;
  assign n2240 = n2239 ^ n2149;
  assign n2241 = n2240 ^ x161;
  assign n2250 = n2249 ^ n2241;
  assign n2251 = n2250 ^ x416;
  assign n25772 = n25771 ^ n2251;
  assign n15937 = n2308 ^ x224;
  assign n15938 = n15937 ^ x416;
  assign n15939 = n15938 ^ x160;
  assign n25773 = n25772 ^ n15939;
  assign n18927 = n16889 ^ x415;
  assign n2301 = x480 ^ x128;
  assign n2302 = n2301 ^ x64;
  assign n2303 = n2302 ^ x320;
  assign n18928 = n18927 ^ n2303;
  assign n18929 = n18928 ^ x351;
  assign n27761 = n25773 ^ n18929;
  assign n2356 = x416 ^ x64;
  assign n2357 = n2356 ^ x256;
  assign n2358 = n2357 ^ x0;
  assign n2354 = n2303 ^ n2251;
  assign n2348 = n2241 ^ x320;
  assign n2340 = x417 ^ x65;
  assign n2341 = n2340 ^ x257;
  assign n2342 = n2341 ^ x1;
  assign n2349 = n2348 ^ n2342;
  assign n2350 = n2349 ^ x256;
  assign n2355 = n2354 ^ n2350;
  assign n2359 = n2358 ^ n2355;
  assign n27762 = n27761 ^ n2359;
  assign n17658 = n15939 ^ x351;
  assign n17659 = n17658 ^ n2358;
  assign n17660 = n17659 ^ x287;
  assign n27763 = n27762 ^ n17660;
  assign n20849 = n18929 ^ x510;
  assign n3273 = n2303 ^ x255;
  assign n3274 = n3273 ^ x447;
  assign n3275 = n3274 ^ x191;
  assign n20850 = n20849 ^ n3275;
  assign n20851 = n20850 ^ x446;
  assign n29647 = n27763 ^ n20851;
  assign n24200 = n3275 ^ n2359;
  assign n19666 = n2350 ^ x447;
  assign n14472 = n2342 ^ x160;
  assign n14473 = n14472 ^ x352;
  assign n14474 = n14473 ^ x96;
  assign n19667 = n19666 ^ n14474;
  assign n19668 = n19667 ^ x383;
  assign n24201 = n24200 ^ n19668;
  assign n14476 = n2358 ^ x191;
  assign n14477 = n14476 ^ x383;
  assign n14478 = n14477 ^ x127;
  assign n24202 = n24201 ^ n14478;
  assign n29648 = n29647 ^ n24202;
  assign n19661 = n17660 ^ x446;
  assign n19662 = n19661 ^ n14478;
  assign n19663 = n19662 ^ x382;
  assign n29649 = n29648 ^ n19663;
  assign n633 = x510 ^ x158;
  assign n634 = n633 ^ x350;
  assign n635 = n634 ^ x94;
  assign n22840 = n20851 ^ n635;
  assign n3276 = n3275 ^ x350;
  assign n3240 = x447 ^ x95;
  assign n3241 = n3240 ^ x287;
  assign n3242 = n3241 ^ x31;
  assign n3277 = n3276 ^ n3242;
  assign n3278 = n3277 ^ x286;
  assign n22841 = n22840 ^ n3278;
  assign n539 = x446 ^ x94;
  assign n540 = n539 ^ x286;
  assign n541 = n540 ^ x30;
  assign n22842 = n22841 ^ n541;
  assign n32317 = n29649 ^ n22842;
  assign n26560 = n24202 ^ n3278;
  assign n21378 = n19668 ^ n3242;
  assign n16652 = n14474 ^ x287;
  assign n16653 = n16652 ^ x479;
  assign n16654 = n16653 ^ x223;
  assign n21379 = n21378 ^ n16654;
  assign n21380 = n21379 ^ x478;
  assign n26561 = n26560 ^ n21380;
  assign n16647 = n14478 ^ x286;
  assign n16648 = n16647 ^ x478;
  assign n16649 = n16648 ^ x222;
  assign n26562 = n26561 ^ n16649;
  assign n32318 = n32317 ^ n26562;
  assign n21373 = n19663 ^ n541;
  assign n21374 = n21373 ^ n16649;
  assign n21375 = n21374 ^ x477;
  assign n32319 = n32318 ^ n21375;
  assign n636 = n635 ^ x253;
  assign n637 = n636 ^ x445;
  assign n638 = n637 ^ x189;
  assign n24746 = n22842 ^ n638;
  assign n3279 = n3278 ^ x445;
  assign n3243 = n3242 ^ x190;
  assign n3244 = n3243 ^ x382;
  assign n3245 = n3244 ^ x126;
  assign n3280 = n3279 ^ n3245;
  assign n3281 = n3280 ^ x381;
  assign n24747 = n24746 ^ n3281;
  assign n554 = n541 ^ x189;
  assign n555 = n554 ^ x381;
  assign n556 = n555 ^ x125;
  assign n24748 = n24747 ^ n556;
  assign n34239 = n32319 ^ n24748;
  assign n28646 = n26562 ^ n3281;
  assign n23080 = n21380 ^ n3245;
  assign n18392 = n16654 ^ x382;
  assign n670 = x479 ^ x127;
  assign n671 = n670 ^ x319;
  assign n672 = n671 ^ x63;
  assign n18393 = n18392 ^ n672;
  assign n18394 = n18393 ^ x318;
  assign n23081 = n23080 ^ n18394;
  assign n13560 = x478 ^ x126;
  assign n13561 = n13560 ^ x318;
  assign n13562 = n13561 ^ x62;
  assign n23082 = n23081 ^ n13562;
  assign n28647 = n28646 ^ n23082;
  assign n18387 = n16649 ^ x381;
  assign n18388 = n18387 ^ n13562;
  assign n18389 = n18388 ^ x317;
  assign n28648 = n28647 ^ n18389;
  assign n34240 = n34239 ^ n28648;
  assign n23104 = n21375 ^ n556;
  assign n23105 = n23104 ^ n18389;
  assign n3250 = x477 ^ x125;
  assign n3251 = n3250 ^ x317;
  assign n3252 = n3251 ^ x61;
  assign n23106 = n23105 ^ n3252;
  assign n34241 = n34240 ^ n23106;
  assign n545 = x445 ^ x93;
  assign n546 = n545 ^ x285;
  assign n547 = n546 ^ x29;
  assign n3282 = n3281 ^ n547;
  assign n3246 = n3245 ^ x285;
  assign n3247 = n3246 ^ x477;
  assign n3248 = n3247 ^ x221;
  assign n3283 = n3282 ^ n3248;
  assign n3284 = n3283 ^ x476;
  assign n30504 = n28648 ^ n3284;
  assign n25033 = n23082 ^ n3248;
  assign n20272 = n18394 ^ x477;
  assign n673 = n672 ^ x222;
  assign n674 = n673 ^ x414;
  assign n675 = n674 ^ x158;
  assign n20273 = n20272 ^ n675;
  assign n20274 = n20273 ^ x413;
  assign n25034 = n25033 ^ n20274;
  assign n15239 = n13562 ^ x221;
  assign n15240 = n15239 ^ x413;
  assign n15241 = n15240 ^ x157;
  assign n25035 = n25034 ^ n15241;
  assign n30505 = n30504 ^ n25035;
  assign n20267 = n18389 ^ x476;
  assign n20268 = n20267 ^ n15241;
  assign n20269 = n20268 ^ x412;
  assign n30506 = n30505 ^ n20269;
  assign n36550 = n34241 ^ n30506;
  assign n639 = n638 ^ x348;
  assign n640 = n639 ^ n547;
  assign n641 = n640 ^ x284;
  assign n26537 = n24748 ^ n641;
  assign n26538 = n26537 ^ n3284;
  assign n572 = n556 ^ x284;
  assign n573 = n572 ^ x476;
  assign n574 = n573 ^ x220;
  assign n26539 = n26538 ^ n574;
  assign n36551 = n36550 ^ n26539;
  assign n25002 = n23106 ^ n574;
  assign n25003 = n25002 ^ n20269;
  assign n3256 = n3252 ^ x220;
  assign n3257 = n3256 ^ x412;
  assign n3258 = n3257 ^ x156;
  assign n25004 = n25003 ^ n3258;
  assign n36552 = n36551 ^ n25004;
  assign n642 = n641 ^ x443;
  assign n560 = n547 ^ x188;
  assign n561 = n560 ^ x380;
  assign n562 = n561 ^ x124;
  assign n643 = n642 ^ n562;
  assign n644 = n643 ^ x379;
  assign n28609 = n26539 ^ n644;
  assign n3285 = n3284 ^ n562;
  assign n3249 = n3248 ^ x380;
  assign n3253 = n3252 ^ n3249;
  assign n3254 = n3253 ^ x316;
  assign n3286 = n3285 ^ n3254;
  assign n591 = x476 ^ x124;
  assign n592 = n591 ^ x316;
  assign n593 = n592 ^ x60;
  assign n3287 = n3286 ^ n593;
  assign n28610 = n28609 ^ n3287;
  assign n590 = n574 ^ x379;
  assign n594 = n593 ^ n590;
  assign n595 = n594 ^ x315;
  assign n28611 = n28610 ^ n595;
  assign n38759 = n36552 ^ n28611;
  assign n33235 = n30506 ^ n3287;
  assign n27172 = n25035 ^ n3254;
  assign n22126 = n20274 ^ n3252;
  assign n697 = n675 ^ x317;
  assign n698 = n697 ^ x509;
  assign n699 = n698 ^ x253;
  assign n22127 = n22126 ^ n699;
  assign n22128 = n22127 ^ x508;
  assign n27173 = n27172 ^ n22128;
  assign n16881 = n15241 ^ x316;
  assign n16882 = n16881 ^ x508;
  assign n16883 = n16882 ^ x252;
  assign n27174 = n27173 ^ n16883;
  assign n33236 = n33235 ^ n27174;
  assign n22156 = n20269 ^ n593;
  assign n22157 = n22156 ^ n16883;
  assign n22158 = n22157 ^ x507;
  assign n33237 = n33236 ^ n22158;
  assign n38760 = n38759 ^ n33237;
  assign n27179 = n25004 ^ n595;
  assign n27180 = n27179 ^ n22158;
  assign n3262 = n3258 ^ x315;
  assign n3263 = n3262 ^ x507;
  assign n3264 = n3263 ^ x251;
  assign n27181 = n27180 ^ n3264;
  assign n38761 = n38760 ^ n27181;
  assign n645 = x443 ^ x91;
  assign n646 = n645 ^ x283;
  assign n647 = n646 ^ x27;
  assign n648 = n647 ^ n644;
  assign n578 = n562 ^ x283;
  assign n579 = n578 ^ x475;
  assign n580 = n579 ^ x219;
  assign n649 = n648 ^ n580;
  assign n650 = n649 ^ x474;
  assign n30494 = n28611 ^ n650;
  assign n3288 = n3287 ^ n580;
  assign n3255 = n3254 ^ x475;
  assign n3259 = n3258 ^ n3255;
  assign n3260 = n3259 ^ x411;
  assign n3289 = n3288 ^ n3260;
  assign n618 = n593 ^ x155;
  assign n619 = n618 ^ x411;
  assign n620 = n619 ^ x219;
  assign n3290 = n3289 ^ n620;
  assign n30495 = n30494 ^ n3290;
  assign n617 = n595 ^ x474;
  assign n621 = n620 ^ n617;
  assign n622 = n621 ^ x410;
  assign n30496 = n30495 ^ n622;
  assign n41071 = n38761 ^ n30496;
  assign n35542 = n33237 ^ n3290;
  assign n29024 = n27174 ^ n3260;
  assign n23681 = n22128 ^ n3258;
  assign n703 = n699 ^ x412;
  assign n513 = x509 ^ x157;
  assign n514 = n513 ^ x349;
  assign n515 = n514 ^ x93;
  assign n704 = n703 ^ n515;
  assign n705 = n704 ^ x348;
  assign n23682 = n23681 ^ n705;
  assign n14274 = x508 ^ x156;
  assign n14275 = n14274 ^ x348;
  assign n14276 = n14275 ^ x92;
  assign n23683 = n23682 ^ n14276;
  assign n29025 = n29024 ^ n23683;
  assign n18916 = n16883 ^ x411;
  assign n18917 = n18916 ^ n14276;
  assign n18918 = n18917 ^ x347;
  assign n29026 = n29025 ^ n18918;
  assign n35543 = n35542 ^ n29026;
  assign n23676 = n22158 ^ n620;
  assign n23677 = n23676 ^ n18918;
  assign n715 = x507 ^ x155;
  assign n716 = n715 ^ x347;
  assign n717 = n716 ^ x91;
  assign n23678 = n23677 ^ n717;
  assign n35544 = n35543 ^ n23678;
  assign n41072 = n41071 ^ n35544;
  assign n29019 = n27181 ^ n622;
  assign n29020 = n29019 ^ n23678;
  assign n3268 = n3264 ^ x410;
  assign n3269 = n3268 ^ n717;
  assign n3270 = n3269 ^ x346;
  assign n29021 = n29020 ^ n3270;
  assign n41073 = n41072 ^ n29021;
  assign n656 = x474 ^ x122;
  assign n657 = n656 ^ x314;
  assign n658 = n657 ^ x58;
  assign n651 = n647 ^ x186;
  assign n652 = n651 ^ x378;
  assign n653 = n652 ^ x122;
  assign n654 = n653 ^ n650;
  assign n602 = n580 ^ x378;
  assign n597 = x475 ^ x123;
  assign n598 = n597 ^ x315;
  assign n599 = n598 ^ x59;
  assign n603 = n602 ^ n599;
  assign n604 = n603 ^ x314;
  assign n655 = n654 ^ n604;
  assign n659 = n658 ^ n655;
  assign n33225 = n30496 ^ n659;
  assign n3291 = n3290 ^ n604;
  assign n3261 = n3260 ^ n599;
  assign n3265 = n3264 ^ n3261;
  assign n3266 = n3265 ^ x506;
  assign n3292 = n3291 ^ n3266;
  assign n765 = n620 ^ x314;
  assign n766 = n765 ^ x506;
  assign n767 = n766 ^ x250;
  assign n3293 = n3292 ^ n767;
  assign n33226 = n33225 ^ n3293;
  assign n764 = n658 ^ n622;
  assign n768 = n767 ^ n764;
  assign n769 = n768 ^ x505;
  assign n33227 = n33226 ^ n769;
  assign n43399 = n41073 ^ n33227;
  assign n37831 = n35544 ^ n3293;
  assign n31387 = n29026 ^ n3266;
  assign n25796 = n23683 ^ n3264;
  assign n709 = n705 ^ x507;
  assign n549 = n515 ^ x252;
  assign n550 = n549 ^ x444;
  assign n551 = n550 ^ x188;
  assign n710 = n709 ^ n551;
  assign n711 = n710 ^ x443;
  assign n25797 = n25796 ^ n711;
  assign n15956 = n14276 ^ x251;
  assign n15957 = n15956 ^ x443;
  assign n15958 = n15957 ^ x187;
  assign n25798 = n25797 ^ n15958;
  assign n31388 = n31387 ^ n25798;
  assign n20837 = n18918 ^ x506;
  assign n20838 = n20837 ^ n15958;
  assign n20839 = n20838 ^ x442;
  assign n31389 = n31388 ^ n20839;
  assign n37832 = n37831 ^ n31389;
  assign n25752 = n23678 ^ n767;
  assign n25753 = n25752 ^ n20839;
  assign n724 = n717 ^ x250;
  assign n725 = n724 ^ x442;
  assign n726 = n725 ^ x186;
  assign n25754 = n25753 ^ n726;
  assign n37833 = n37832 ^ n25754;
  assign n43400 = n43399 ^ n37833;
  assign n31382 = n29021 ^ n769;
  assign n31383 = n31382 ^ n25754;
  assign n3299 = n3270 ^ x505;
  assign n3300 = n3299 ^ n726;
  assign n3301 = n3300 ^ x441;
  assign n31384 = n31383 ^ n3301;
  assign n43401 = n43400 ^ n31384;
  assign n665 = n658 ^ x217;
  assign n666 = n665 ^ x409;
  assign n667 = n666 ^ x153;
  assign n660 = n653 ^ x281;
  assign n661 = n660 ^ x473;
  assign n662 = n661 ^ x217;
  assign n663 = n662 ^ n659;
  assign n629 = n604 ^ x473;
  assign n624 = n599 ^ x218;
  assign n625 = n624 ^ x410;
  assign n626 = n625 ^ x154;
  assign n630 = n629 ^ n626;
  assign n631 = n630 ^ x409;
  assign n664 = n663 ^ n631;
  assign n668 = n667 ^ n664;
  assign n35532 = n33227 ^ n668;
  assign n3294 = n3293 ^ n631;
  assign n3267 = n3266 ^ n626;
  assign n3271 = n3270 ^ n3267;
  assign n818 = x506 ^ x154;
  assign n819 = n818 ^ x346;
  assign n820 = n819 ^ x90;
  assign n3272 = n3271 ^ n820;
  assign n3295 = n3294 ^ n3272;
  assign n817 = n767 ^ x409;
  assign n821 = n820 ^ n817;
  assign n822 = n821 ^ x345;
  assign n3296 = n3295 ^ n822;
  assign n35533 = n35532 ^ n3296;
  assign n824 = x505 ^ x153;
  assign n825 = n824 ^ x345;
  assign n826 = n825 ^ x89;
  assign n816 = n769 ^ n667;
  assign n823 = n822 ^ n816;
  assign n827 = n826 ^ n823;
  assign n35534 = n35533 ^ n827;
  assign n45419 = n43401 ^ n35534;
  assign n39988 = n37833 ^ n3296;
  assign n33462 = n31389 ^ n3272;
  assign n27740 = n25798 ^ n3270;
  assign n718 = n717 ^ n711;
  assign n565 = x444 ^ x92;
  assign n566 = n565 ^ x284;
  assign n567 = n566 ^ x28;
  assign n564 = n551 ^ x347;
  assign n568 = n567 ^ n564;
  assign n569 = n568 ^ x283;
  assign n719 = n718 ^ n569;
  assign n720 = n719 ^ n647;
  assign n27741 = n27740 ^ n720;
  assign n17647 = n15958 ^ x346;
  assign n17648 = n17647 ^ n647;
  assign n17649 = n17648 ^ x282;
  assign n27742 = n27741 ^ n17649;
  assign n33463 = n33462 ^ n27742;
  assign n22831 = n20839 ^ n17649;
  assign n22832 = n22831 ^ n820;
  assign n606 = x442 ^ x90;
  assign n607 = n606 ^ x282;
  assign n608 = n607 ^ x26;
  assign n22833 = n22832 ^ n608;
  assign n33464 = n33463 ^ n22833;
  assign n39989 = n39988 ^ n33464;
  assign n27735 = n25754 ^ n822;
  assign n27736 = n27735 ^ n22833;
  assign n733 = n726 ^ x345;
  assign n734 = n733 ^ n608;
  assign n735 = n734 ^ x281;
  assign n27737 = n27736 ^ n735;
  assign n39990 = n39989 ^ n27737;
  assign n45420 = n45419 ^ n39990;
  assign n33537 = n31384 ^ n827;
  assign n33538 = n33537 ^ n27737;
  assign n3308 = n3301 ^ n826;
  assign n3309 = n3308 ^ n735;
  assign n956 = x441 ^ x89;
  assign n957 = n956 ^ x281;
  assign n958 = n957 ^ x25;
  assign n3310 = n3309 ^ n958;
  assign n33539 = n33538 ^ n3310;
  assign n45421 = n45420 ^ n33539;
  assign n784 = n667 ^ x312;
  assign n785 = n784 ^ x504;
  assign n786 = n785 ^ x248;
  assign n758 = n662 ^ x376;
  assign n753 = x473 ^ x121;
  assign n754 = n753 ^ x313;
  assign n755 = n754 ^ x57;
  assign n759 = n758 ^ n755;
  assign n760 = n759 ^ x312;
  assign n782 = n760 ^ n668;
  assign n777 = n755 ^ n631;
  assign n771 = n626 ^ x313;
  assign n772 = n771 ^ x505;
  assign n773 = n772 ^ x249;
  assign n778 = n777 ^ n773;
  assign n779 = n778 ^ x504;
  assign n783 = n782 ^ n779;
  assign n787 = n786 ^ n783;
  assign n37841 = n35534 ^ n787;
  assign n3298 = n3272 ^ n773;
  assign n3302 = n3301 ^ n3298;
  assign n884 = n820 ^ x249;
  assign n885 = n884 ^ x441;
  assign n886 = n885 ^ x185;
  assign n3303 = n3302 ^ n886;
  assign n3297 = n3296 ^ n779;
  assign n3304 = n3303 ^ n3297;
  assign n883 = n822 ^ x504;
  assign n887 = n886 ^ n883;
  assign n888 = n887 ^ x440;
  assign n3305 = n3304 ^ n888;
  assign n37842 = n37841 ^ n3305;
  assign n890 = n826 ^ x248;
  assign n891 = n890 ^ x440;
  assign n892 = n891 ^ x184;
  assign n882 = n827 ^ n786;
  assign n889 = n888 ^ n882;
  assign n893 = n892 ^ n889;
  assign n37843 = n37842 ^ n893;
  assign n47519 = n45421 ^ n37843;
  assign n42207 = n39990 ^ n3305;
  assign n35833 = n33464 ^ n3303;
  assign n30173 = n27742 ^ n3301;
  assign n727 = n726 ^ n720;
  assign n583 = n567 ^ x187;
  assign n584 = n583 ^ x379;
  assign n585 = n584 ^ x123;
  assign n582 = n569 ^ x442;
  assign n586 = n585 ^ n582;
  assign n587 = n586 ^ x378;
  assign n728 = n727 ^ n587;
  assign n729 = n728 ^ n653;
  assign n30174 = n30173 ^ n729;
  assign n19690 = n17649 ^ x441;
  assign n19691 = n19690 ^ n653;
  assign n19692 = n19691 ^ x377;
  assign n30175 = n30174 ^ n19692;
  assign n35834 = n35833 ^ n30175;
  assign n24767 = n22833 ^ n886;
  assign n24768 = n24767 ^ n19692;
  assign n742 = n608 ^ x185;
  assign n743 = n742 ^ x377;
  assign n744 = n743 ^ x121;
  assign n24769 = n24768 ^ n744;
  assign n35835 = n35834 ^ n24769;
  assign n42208 = n42207 ^ n35835;
  assign n30192 = n27737 ^ n888;
  assign n30193 = n30192 ^ n24769;
  assign n741 = n735 ^ x440;
  assign n745 = n744 ^ n741;
  assign n746 = n745 ^ x376;
  assign n30194 = n30193 ^ n746;
  assign n42209 = n42208 ^ n30194;
  assign n47520 = n47519 ^ n42209;
  assign n35828 = n33539 ^ n893;
  assign n35829 = n35828 ^ n30194;
  assign n3317 = n3310 ^ n892;
  assign n3318 = n3317 ^ n746;
  assign n1041 = n958 ^ x184;
  assign n1042 = n1041 ^ x376;
  assign n1043 = n1042 ^ x120;
  assign n3319 = n3318 ^ n1043;
  assign n35830 = n35829 ^ n3319;
  assign n47521 = n47520 ^ n35830;
  assign n844 = n786 ^ x407;
  assign n836 = x504 ^ x152;
  assign n837 = n836 ^ x344;
  assign n838 = n837 ^ x88;
  assign n845 = n844 ^ n838;
  assign n846 = n845 ^ x343;
  assign n809 = n760 ^ x471;
  assign n804 = n755 ^ x216;
  assign n805 = n804 ^ x408;
  assign n806 = n805 ^ x152;
  assign n810 = n809 ^ n806;
  assign n811 = n810 ^ x407;
  assign n842 = n811 ^ n787;
  assign n834 = n806 ^ n779;
  assign n829 = n773 ^ x408;
  assign n830 = n829 ^ n826;
  assign n831 = n830 ^ x344;
  assign n835 = n834 ^ n831;
  assign n839 = n838 ^ n835;
  assign n843 = n842 ^ n839;
  assign n847 = n846 ^ n843;
  assign n39978 = n37843 ^ n847;
  assign n3307 = n3303 ^ n831;
  assign n3311 = n3310 ^ n3307;
  assign n955 = n886 ^ x344;
  assign n959 = n958 ^ n955;
  assign n960 = n959 ^ x280;
  assign n3312 = n3311 ^ n960;
  assign n3306 = n3305 ^ n839;
  assign n3313 = n3312 ^ n3306;
  assign n954 = n888 ^ n838;
  assign n961 = n960 ^ n954;
  assign n789 = x440 ^ x88;
  assign n790 = n789 ^ x280;
  assign n791 = n790 ^ x24;
  assign n962 = n961 ^ n791;
  assign n3314 = n3313 ^ n962;
  assign n39979 = n39978 ^ n3314;
  assign n964 = n892 ^ x343;
  assign n965 = n964 ^ n791;
  assign n966 = n965 ^ x279;
  assign n953 = n893 ^ n846;
  assign n963 = n962 ^ n953;
  assign n967 = n966 ^ n963;
  assign n39980 = n39979 ^ n967;
  assign n49557 = n47521 ^ n39980;
  assign n43971 = n42209 ^ n3314;
  assign n38082 = n35835 ^ n3312;
  assign n32295 = n30175 ^ n3310;
  assign n736 = n735 ^ n729;
  assign n610 = n585 ^ x282;
  assign n611 = n610 ^ x474;
  assign n612 = n611 ^ x218;
  assign n609 = n608 ^ n587;
  assign n613 = n612 ^ n609;
  assign n614 = n613 ^ x473;
  assign n737 = n736 ^ n614;
  assign n738 = n737 ^ n662;
  assign n32296 = n32295 ^ n738;
  assign n21408 = n19692 ^ n958;
  assign n21409 = n21408 ^ n662;
  assign n21410 = n21409 ^ x472;
  assign n32297 = n32296 ^ n21410;
  assign n38083 = n38082 ^ n32297;
  assign n26524 = n24769 ^ n960;
  assign n26525 = n26524 ^ n21410;
  assign n793 = n744 ^ x280;
  assign n794 = n793 ^ x472;
  assign n795 = n794 ^ x216;
  assign n26526 = n26525 ^ n795;
  assign n38084 = n38083 ^ n26526;
  assign n43972 = n43971 ^ n38084;
  assign n32290 = n30194 ^ n962;
  assign n32291 = n32290 ^ n26526;
  assign n792 = n791 ^ n746;
  assign n796 = n795 ^ n792;
  assign n797 = n796 ^ x471;
  assign n32292 = n32291 ^ n797;
  assign n43973 = n43972 ^ n32292;
  assign n49558 = n49557 ^ n43973;
  assign n38077 = n35830 ^ n967;
  assign n38078 = n38077 ^ n32292;
  assign n3326 = n3319 ^ n966;
  assign n3327 = n3326 ^ n797;
  assign n1141 = n1043 ^ x279;
  assign n1142 = n1141 ^ x471;
  assign n1143 = n1142 ^ x215;
  assign n3328 = n3327 ^ n1143;
  assign n38079 = n38078 ^ n3328;
  assign n49559 = n49558 ^ n38079;
  assign n910 = n846 ^ x502;
  assign n902 = n838 ^ x247;
  assign n903 = n902 ^ x439;
  assign n904 = n903 ^ x183;
  assign n911 = n910 ^ n904;
  assign n912 = n911 ^ x438;
  assign n875 = n862 ^ n811;
  assign n870 = n806 ^ x311;
  assign n871 = n870 ^ x503;
  assign n872 = n871 ^ x247;
  assign n876 = n875 ^ n872;
  assign n877 = n876 ^ x502;
  assign n908 = n877 ^ n847;
  assign n900 = n872 ^ n839;
  assign n895 = n831 ^ x503;
  assign n896 = n895 ^ n892;
  assign n897 = n896 ^ x439;
  assign n901 = n900 ^ n897;
  assign n905 = n904 ^ n901;
  assign n909 = n908 ^ n905;
  assign n913 = n912 ^ n909;
  assign n42229 = n39980 ^ n913;
  assign n3316 = n3312 ^ n897;
  assign n3320 = n3319 ^ n3316;
  assign n1040 = n960 ^ x439;
  assign n1044 = n1043 ^ n1040;
  assign n1045 = n1044 ^ x375;
  assign n3321 = n3320 ^ n1045;
  assign n3315 = n3314 ^ n905;
  assign n3322 = n3321 ^ n3315;
  assign n1039 = n962 ^ n904;
  assign n1046 = n1045 ^ n1039;
  assign n849 = n791 ^ x183;
  assign n850 = n849 ^ x375;
  assign n851 = n850 ^ x119;
  assign n1047 = n1046 ^ n851;
  assign n3323 = n3322 ^ n1047;
  assign n42230 = n42229 ^ n3323;
  assign n1049 = n966 ^ x438;
  assign n1050 = n1049 ^ n851;
  assign n1051 = n1050 ^ x374;
  assign n1038 = n967 ^ n912;
  assign n1048 = n1047 ^ n1038;
  assign n1052 = n1051 ^ n1048;
  assign n42231 = n42230 ^ n1052;
  assign n51567 = n49559 ^ n42231;
  assign n45948 = n43973 ^ n3323;
  assign n40300 = n38084 ^ n3321;
  assign n34763 = n32297 ^ n3319;
  assign n749 = n612 ^ x377;
  assign n750 = n749 ^ n658;
  assign n751 = n750 ^ x313;
  assign n748 = n744 ^ n614;
  assign n752 = n751 ^ n748;
  assign n756 = n755 ^ n752;
  assign n747 = n746 ^ n738;
  assign n757 = n756 ^ n747;
  assign n761 = n760 ^ n757;
  assign n34764 = n34763 ^ n761;
  assign n23068 = n21410 ^ n1043;
  assign n23069 = n23068 ^ n760;
  assign n854 = x472 ^ x120;
  assign n855 = n854 ^ x312;
  assign n856 = n855 ^ x56;
  assign n23070 = n23069 ^ n856;
  assign n34765 = n34764 ^ n23070;
  assign n40301 = n40300 ^ n34765;
  assign n28671 = n26526 ^ n1045;
  assign n28672 = n28671 ^ n23070;
  assign n853 = n795 ^ x375;
  assign n857 = n856 ^ n853;
  assign n858 = n857 ^ x311;
  assign n28673 = n28672 ^ n858;
  assign n40302 = n40301 ^ n28673;
  assign n45949 = n45948 ^ n40302;
  assign n34758 = n32292 ^ n1047;
  assign n34759 = n34758 ^ n28673;
  assign n852 = n851 ^ n797;
  assign n859 = n858 ^ n852;
  assign n863 = n862 ^ n859;
  assign n34760 = n34759 ^ n863;
  assign n45950 = n45949 ^ n34760;
  assign n51568 = n51567 ^ n45950;
  assign n40392 = n38079 ^ n1052;
  assign n40393 = n40392 ^ n34760;
  assign n3335 = n3328 ^ n1051;
  assign n3336 = n3335 ^ n863;
  assign n1224 = n1143 ^ x374;
  assign n1225 = n1224 ^ n862;
  assign n1226 = n1225 ^ x310;
  assign n3337 = n3336 ^ n1226;
  assign n40394 = n40393 ^ n3337;
  assign n51569 = n51568 ^ n40394;
  assign n990 = x438 ^ x86;
  assign n991 = n990 ^ x278;
  assign n992 = n991 ^ x22;
  assign n946 = x502 ^ x150;
  assign n947 = n946 ^ x342;
  assign n948 = n947 ^ x86;
  assign n988 = n948 ^ n912;
  assign n980 = n904 ^ x342;
  assign n971 = x439 ^ x87;
  assign n972 = n971 ^ x279;
  assign n973 = n972 ^ x23;
  assign n981 = n980 ^ n973;
  assign n982 = n981 ^ x278;
  assign n989 = n988 ^ n982;
  assign n993 = n992 ^ n989;
  assign n944 = n928 ^ n877;
  assign n932 = x503 ^ x151;
  assign n933 = n932 ^ x343;
  assign n934 = n933 ^ x87;
  assign n931 = n872 ^ x406;
  assign n935 = n934 ^ n931;
  assign n936 = n935 ^ x342;
  assign n945 = n944 ^ n936;
  assign n949 = n948 ^ n945;
  assign n986 = n949 ^ n913;
  assign n978 = n936 ^ n905;
  assign n969 = n934 ^ n897;
  assign n970 = n969 ^ n966;
  assign n974 = n973 ^ n970;
  assign n979 = n978 ^ n974;
  assign n983 = n982 ^ n979;
  assign n987 = n986 ^ n983;
  assign n994 = n993 ^ n987;
  assign n43961 = n42231 ^ n994;
  assign n3325 = n3321 ^ n974;
  assign n3329 = n3328 ^ n3325;
  assign n1140 = n1045 ^ n973;
  assign n1144 = n1143 ^ n1140;
  assign n1145 = n1144 ^ x470;
  assign n3330 = n3329 ^ n1145;
  assign n3324 = n3323 ^ n983;
  assign n3331 = n3330 ^ n3324;
  assign n1139 = n1047 ^ n982;
  assign n1146 = n1145 ^ n1139;
  assign n915 = n851 ^ x278;
  assign n916 = n915 ^ x470;
  assign n917 = n916 ^ x214;
  assign n1147 = n1146 ^ n917;
  assign n3332 = n3331 ^ n1147;
  assign n43962 = n43961 ^ n3332;
  assign n1138 = n1052 ^ n993;
  assign n1148 = n1147 ^ n1138;
  assign n1129 = n1051 ^ n992;
  assign n1130 = n1129 ^ n917;
  assign n1131 = n1130 ^ x469;
  assign n1149 = n1148 ^ n1131;
  assign n43963 = n43962 ^ n1149;
  assign n53699 = n51569 ^ n43963;
  assign n48089 = n45950 ^ n3332;
  assign n42484 = n40302 ^ n3330;
  assign n36997 = n34765 ^ n3328;
  assign n800 = n751 ^ x472;
  assign n801 = n800 ^ n667;
  assign n802 = n801 ^ x408;
  assign n799 = n795 ^ n756;
  assign n803 = n802 ^ n799;
  assign n807 = n806 ^ n803;
  assign n798 = n797 ^ n761;
  assign n808 = n807 ^ n798;
  assign n812 = n811 ^ n808;
  assign n36998 = n36997 ^ n812;
  assign n25056 = n23070 ^ n1143;
  assign n25057 = n25056 ^ n811;
  assign n920 = n856 ^ x215;
  assign n921 = n920 ^ x407;
  assign n922 = n921 ^ x151;
  assign n25058 = n25057 ^ n922;
  assign n36999 = n36998 ^ n25058;
  assign n42485 = n42484 ^ n36999;
  assign n30482 = n28673 ^ n1145;
  assign n30483 = n30482 ^ n25058;
  assign n919 = n858 ^ x470;
  assign n923 = n922 ^ n919;
  assign n924 = n923 ^ x406;
  assign n30484 = n30483 ^ n924;
  assign n42486 = n42485 ^ n30484;
  assign n48090 = n48089 ^ n42486;
  assign n37008 = n34760 ^ n1147;
  assign n918 = n917 ^ n863;
  assign n925 = n924 ^ n918;
  assign n929 = n928 ^ n925;
  assign n37009 = n37008 ^ n929;
  assign n37010 = n37009 ^ n30484;
  assign n48091 = n48090 ^ n37010;
  assign n53700 = n53699 ^ n48091;
  assign n42479 = n40394 ^ n1149;
  assign n42480 = n42479 ^ n37010;
  assign n3345 = n3337 ^ n1131;
  assign n3346 = n3345 ^ n929;
  assign n1332 = n1226 ^ x469;
  assign n1333 = n1332 ^ n928;
  assign n1334 = n1333 ^ x405;
  assign n3347 = n3346 ^ n1334;
  assign n42481 = n42480 ^ n3347;
  assign n53701 = n53700 ^ n42481;
  assign n1843 = n1780 ^ x199;
  assign n1844 = n1843 ^ x391;
  assign n1845 = n1844 ^ x135;
  assign n1842 = n1782 ^ x454;
  assign n1846 = n1845 ^ n1842;
  assign n1847 = n1846 ^ x390;
  assign n1712 = n1693 ^ x262;
  assign n1713 = n1712 ^ x454;
  assign n1714 = n1713 ^ x198;
  assign n1841 = n1784 ^ n1714;
  assign n1848 = n1847 ^ n1841;
  assign n1836 = n1772 ^ x198;
  assign n1837 = n1836 ^ x390;
  assign n1838 = n1837 ^ x134;
  assign n1849 = n1848 ^ n1838;
  assign n35455 = n33144 ^ n1849;
  assign n29379 = n27421 ^ n1847;
  assign n24017 = n22091 ^ n1845;
  assign n24018 = n24017 ^ n19280;
  assign n1717 = x487 ^ x135;
  assign n1718 = n1717 ^ x327;
  assign n1719 = n1718 ^ x71;
  assign n24019 = n24018 ^ n1719;
  assign n29380 = n29379 ^ n24019;
  assign n1720 = n1658 ^ x390;
  assign n1721 = n1720 ^ n1719;
  assign n1722 = n1721 ^ x326;
  assign n29381 = n29380 ^ n1722;
  assign n35456 = n35455 ^ n29381;
  assign n24119 = n22232 ^ n1838;
  assign n24120 = n24119 ^ n1722;
  assign n1994 = x486 ^ x134;
  assign n1995 = n1994 ^ x326;
  assign n1996 = n1995 ^ x70;
  assign n24121 = n24120 ^ n1996;
  assign n35457 = n35456 ^ n24121;
  assign n1915 = n1845 ^ x294;
  assign n1916 = n1915 ^ x486;
  assign n1917 = n1916 ^ x230;
  assign n1790 = x454 ^ x102;
  assign n1791 = n1790 ^ x38;
  assign n1792 = n1791 ^ x294;
  assign n1914 = n1847 ^ n1792;
  assign n1918 = n1917 ^ n1914;
  assign n1919 = n1918 ^ x485;
  assign n1798 = n1714 ^ x357;
  assign n1799 = n1798 ^ n1792;
  assign n1800 = n1799 ^ x293;
  assign n1913 = n1849 ^ n1800;
  assign n1920 = n1919 ^ n1913;
  assign n1908 = n1838 ^ x293;
  assign n1909 = n1908 ^ x485;
  assign n1910 = n1909 ^ x229;
  assign n1921 = n1920 ^ n1910;
  assign n37737 = n35457 ^ n1921;
  assign n31776 = n29381 ^ n1919;
  assign n26114 = n24019 ^ n1917;
  assign n26115 = n26114 ^ n21119;
  assign n1746 = n1719 ^ x230;
  assign n1747 = n1746 ^ x422;
  assign n1748 = n1747 ^ x166;
  assign n26116 = n26115 ^ n1748;
  assign n31777 = n31776 ^ n26116;
  assign n1749 = n1722 ^ x485;
  assign n1750 = n1749 ^ n1748;
  assign n1751 = n1750 ^ x421;
  assign n31778 = n31777 ^ n1751;
  assign n37738 = n37737 ^ n31778;
  assign n26109 = n24121 ^ n1910;
  assign n26110 = n26109 ^ n1751;
  assign n2072 = n1996 ^ x229;
  assign n2073 = n2072 ^ x421;
  assign n2074 = n2073 ^ x165;
  assign n26111 = n26110 ^ n2074;
  assign n37739 = n37738 ^ n26111;
  assign n1993 = n1917 ^ x389;
  assign n1997 = n1996 ^ n1993;
  assign n1998 = n1997 ^ x325;
  assign n1856 = n1792 ^ x197;
  assign n1857 = n1856 ^ x389;
  assign n1858 = n1857 ^ x133;
  assign n1992 = n1919 ^ n1858;
  assign n1999 = n1998 ^ n1992;
  assign n1812 = x485 ^ x133;
  assign n1813 = n1812 ^ x325;
  assign n1814 = n1813 ^ x69;
  assign n2000 = n1999 ^ n1814;
  assign n1864 = n1800 ^ x452;
  assign n1865 = n1864 ^ n1858;
  assign n1866 = n1865 ^ x388;
  assign n1991 = n1921 ^ n1866;
  assign n2001 = n2000 ^ n1991;
  assign n1983 = n1910 ^ x388;
  assign n1984 = n1983 ^ n1814;
  assign n1985 = n1984 ^ x324;
  assign n2002 = n2001 ^ n1985;
  assign n39913 = n37739 ^ n2002;
  assign n33933 = n31778 ^ n2000;
  assign n28153 = n26116 ^ n1998;
  assign n22799 = n21119 ^ n1996;
  assign n1699 = x263 ^ x71;
  assign n1700 = n1699 ^ x423;
  assign n1701 = n1700 ^ x7;
  assign n1698 = n1669 ^ x326;
  assign n1702 = n1701 ^ n1698;
  assign n1703 = n1702 ^ x262;
  assign n22800 = n22799 ^ n1703;
  assign n22801 = n22800 ^ n1808;
  assign n28154 = n28153 ^ n22801;
  assign n1809 = n1748 ^ x325;
  assign n1810 = n1809 ^ n1808;
  assign n1811 = n1810 ^ x261;
  assign n28155 = n28154 ^ n1811;
  assign n33934 = n33933 ^ n28155;
  assign n1815 = n1814 ^ n1751;
  assign n1816 = n1815 ^ n1811;
  assign n1803 = x421 ^ x69;
  assign n1804 = n1803 ^ x261;
  assign n1805 = n1804 ^ x5;
  assign n1817 = n1816 ^ n1805;
  assign n33935 = n33934 ^ n1817;
  assign n39914 = n39913 ^ n33935;
  assign n28148 = n26111 ^ n1985;
  assign n28149 = n28148 ^ n1817;
  assign n2174 = n2074 ^ x324;
  assign n2175 = n2174 ^ n1805;
  assign n2176 = n2175 ^ x260;
  assign n28150 = n28149 ^ n2176;
  assign n39915 = n39914 ^ n28150;
  assign n2080 = n1985 ^ x483;
  assign n1878 = n1814 ^ x228;
  assign n1879 = n1878 ^ x420;
  assign n1880 = n1879 ^ x164;
  assign n2081 = n2080 ^ n1880;
  assign n2082 = n2081 ^ x419;
  assign n2071 = n1998 ^ x484;
  assign n2075 = n2074 ^ n2071;
  assign n2076 = n2075 ^ x420;
  assign n1928 = n1858 ^ x292;
  assign n1929 = n1928 ^ x484;
  assign n1930 = n1929 ^ x228;
  assign n2070 = n2000 ^ n1930;
  assign n2077 = n2076 ^ n2070;
  assign n2078 = n2077 ^ n1880;
  assign n1936 = n1902 ^ n1866;
  assign n1937 = n1936 ^ n1930;
  assign n1938 = n1937 ^ x483;
  assign n2069 = n2002 ^ n1938;
  assign n2079 = n2078 ^ n2069;
  assign n2083 = n2082 ^ n2079;
  assign n42310 = n39915 ^ n2083;
  assign n36279 = n33935 ^ n2078;
  assign n30128 = n28155 ^ n2076;
  assign n24697 = n22801 ^ n2074;
  assign n1763 = n1703 ^ x421;
  assign n1758 = n1701 ^ x166;
  assign n1759 = n1758 ^ x358;
  assign n1760 = n1759 ^ x102;
  assign n1764 = n1763 ^ n1760;
  assign n1765 = n1764 ^ x357;
  assign n24698 = n24697 ^ n1765;
  assign n24699 = n24698 ^ n1874;
  assign n30129 = n30128 ^ n24699;
  assign n1875 = n1811 ^ x420;
  assign n1876 = n1875 ^ n1874;
  assign n1877 = n1876 ^ x356;
  assign n30130 = n30129 ^ n1877;
  assign n36280 = n36279 ^ n30130;
  assign n1881 = n1880 ^ n1817;
  assign n1882 = n1881 ^ n1877;
  assign n1869 = n1805 ^ x164;
  assign n1870 = n1869 ^ x356;
  assign n1871 = n1870 ^ x100;
  assign n1883 = n1882 ^ n1871;
  assign n36281 = n36280 ^ n1883;
  assign n42311 = n42310 ^ n36281;
  assign n30123 = n28150 ^ n2082;
  assign n30124 = n30123 ^ n1883;
  assign n2262 = n2176 ^ x419;
  assign n2263 = n2262 ^ n1871;
  assign n2264 = n2263 ^ x355;
  assign n30125 = n30124 ^ n2264;
  assign n42312 = n42311 ^ n30125;
  assign n1987 = x484 ^ x132;
  assign n1988 = n1987 ^ x324;
  assign n1989 = n1988 ^ x68;
  assign n2173 = n2076 ^ n1989;
  assign n2177 = n2176 ^ n2173;
  assign n1947 = x420 ^ x68;
  assign n1948 = n1947 ^ x260;
  assign n1949 = n1948 ^ x4;
  assign n2178 = n2177 ^ n1949;
  assign n2009 = n1930 ^ x387;
  assign n2010 = n2009 ^ n1989;
  assign n2011 = n2010 ^ x323;
  assign n2172 = n2078 ^ n2011;
  assign n2179 = n2178 ^ n2172;
  assign n1953 = n1880 ^ x323;
  assign n1954 = n1953 ^ n1949;
  assign n1955 = n1954 ^ x259;
  assign n2180 = n2179 ^ n1955;
  assign n2019 = x483 ^ x131;
  assign n2020 = n2019 ^ x323;
  assign n2021 = n2020 ^ x67;
  assign n2017 = n1970 ^ n1938;
  assign n2018 = n2017 ^ n2011;
  assign n2022 = n2021 ^ n2018;
  assign n2171 = n2083 ^ n2022;
  assign n2181 = n2180 ^ n2171;
  assign n2163 = n2082 ^ n2021;
  assign n2164 = n2163 ^ n1955;
  assign n676 = x419 ^ x67;
  assign n677 = n676 ^ x259;
  assign n678 = n677 ^ x3;
  assign n2165 = n2164 ^ n678;
  assign n2182 = n2181 ^ n2165;
  assign n44001 = n42312 ^ n2182;
  assign n38619 = n36281 ^ n2180;
  assign n32746 = n30130 ^ n2178;
  assign n26796 = n24699 ^ n2176;
  assign n1829 = n1805 ^ n1765;
  assign n1824 = n1760 ^ x261;
  assign n1825 = n1824 ^ x453;
  assign n1826 = n1825 ^ x197;
  assign n1830 = n1829 ^ n1826;
  assign n1831 = n1830 ^ x452;
  assign n26797 = n26796 ^ n1831;
  assign n26798 = n26797 ^ n1946;
  assign n32747 = n32746 ^ n26798;
  assign n1950 = n1949 ^ n1877;
  assign n1951 = n1950 ^ n1946;
  assign n1952 = n1951 ^ x451;
  assign n32748 = n32747 ^ n1952;
  assign n38620 = n38619 ^ n32748;
  assign n1956 = n1955 ^ n1883;
  assign n1957 = n1956 ^ n1952;
  assign n1941 = n1871 ^ x259;
  assign n1942 = n1941 ^ x451;
  assign n1943 = n1942 ^ x195;
  assign n1958 = n1957 ^ n1943;
  assign n38621 = n38620 ^ n1958;
  assign n44002 = n44001 ^ n38621;
  assign n32741 = n30125 ^ n2165;
  assign n32742 = n32741 ^ n1958;
  assign n2373 = n2264 ^ n678;
  assign n2374 = n2373 ^ n1943;
  assign n2375 = n2374 ^ x450;
  assign n32743 = n32742 ^ n2375;
  assign n44003 = n44002 ^ n32743;
  assign n1706 = n1683 ^ x263;
  assign n1707 = n1706 ^ x455;
  assign n1708 = n1707 ^ x199;
  assign n1705 = n1701 ^ n1688;
  assign n1709 = n1708 ^ n1705;
  assign n1710 = n1709 ^ x454;
  assign n31059 = n28556 ^ n1710;
  assign n25425 = n23468 ^ n1708;
  assign n25426 = n25425 ^ n20528;
  assign n25427 = n25426 ^ n1845;
  assign n31060 = n31059 ^ n25427;
  assign n31061 = n31060 ^ n1847;
  assign n1788 = n1760 ^ n1710;
  assign n1769 = n1708 ^ x358;
  assign n1773 = n1772 ^ n1769;
  assign n1774 = n1773 ^ x294;
  assign n1789 = n1788 ^ n1774;
  assign n1793 = n1792 ^ n1789;
  assign n33137 = n31061 ^ n1793;
  assign n27431 = n25427 ^ n1774;
  assign n27432 = n27431 ^ n22232;
  assign n27433 = n27432 ^ n1917;
  assign n33138 = n33137 ^ n27433;
  assign n33139 = n33138 ^ n1919;
  assign n1854 = n1826 ^ n1793;
  assign n1835 = n1774 ^ x453;
  assign n1839 = n1838 ^ n1835;
  assign n1840 = n1839 ^ x389;
  assign n1855 = n1854 ^ n1840;
  assign n1859 = n1858 ^ n1855;
  assign n35450 = n33139 ^ n1859;
  assign n29374 = n27433 ^ n1840;
  assign n29375 = n29374 ^ n24121;
  assign n29376 = n29375 ^ n1998;
  assign n35451 = n35450 ^ n29376;
  assign n35452 = n35451 ^ n2000;
  assign n1893 = n1826 ^ x356;
  assign n1888 = x293 ^ x101;
  assign n1889 = n1888 ^ x453;
  assign n1890 = n1889 ^ x37;
  assign n1894 = n1893 ^ n1890;
  assign n1895 = n1894 ^ x292;
  assign n1926 = n1895 ^ n1859;
  assign n1907 = n1890 ^ n1840;
  assign n1911 = n1910 ^ n1907;
  assign n1912 = n1911 ^ x484;
  assign n1927 = n1926 ^ n1912;
  assign n1931 = n1930 ^ n1927;
  assign n37732 = n35452 ^ n1931;
  assign n37733 = n37732 ^ n2078;
  assign n31771 = n29376 ^ n1912;
  assign n31772 = n31771 ^ n26111;
  assign n31773 = n31772 ^ n2076;
  assign n37734 = n37733 ^ n31773;
  assign n1962 = n1890 ^ x196;
  assign n1963 = n1962 ^ x388;
  assign n1964 = n1963 ^ x132;
  assign n1961 = n1895 ^ x451;
  assign n1965 = n1964 ^ n1961;
  assign n1966 = n1965 ^ x387;
  assign n2007 = n1966 ^ n1931;
  assign n1982 = n1964 ^ n1912;
  assign n1986 = n1985 ^ n1982;
  assign n1990 = n1989 ^ n1986;
  assign n2008 = n2007 ^ n1990;
  assign n2012 = n2011 ^ n2008;
  assign n40100 = n37734 ^ n2012;
  assign n34104 = n31773 ^ n1990;
  assign n34105 = n34104 ^ n28150;
  assign n34106 = n34105 ^ n2178;
  assign n40101 = n40100 ^ n34106;
  assign n40102 = n40101 ^ n2180;
  assign n2096 = n2011 ^ x482;
  assign n2086 = n1989 ^ x227;
  assign n2087 = n2086 ^ x419;
  assign n2088 = n2087 ^ x163;
  assign n2097 = n2096 ^ n2088;
  assign n2098 = n2097 ^ x418;
  assign n2026 = x451 ^ x99;
  assign n2027 = n2026 ^ x291;
  assign n2028 = n2027 ^ x35;
  assign n2055 = n2028 ^ n1966;
  assign n2050 = n1964 ^ x291;
  assign n2051 = n2050 ^ x483;
  assign n2052 = n2051 ^ x227;
  assign n2056 = n2055 ^ n2052;
  assign n2057 = n2056 ^ x482;
  assign n2094 = n2057 ^ n2012;
  assign n2084 = n2052 ^ n1990;
  assign n2085 = n2084 ^ n2082;
  assign n2089 = n2088 ^ n2085;
  assign n2095 = n2094 ^ n2089;
  assign n2099 = n2098 ^ n2095;
  assign n41696 = n40102 ^ n2099;
  assign n2261 = n2178 ^ n2088;
  assign n2265 = n2264 ^ n2261;
  assign n2034 = n1949 ^ x163;
  assign n2035 = n2034 ^ x355;
  assign n2036 = n2035 ^ x99;
  assign n2266 = n2265 ^ n2036;
  assign n36401 = n34106 ^ n2266;
  assign n36402 = n36401 ^ n30125;
  assign n36403 = n36402 ^ n2089;
  assign n41697 = n41696 ^ n36403;
  assign n2260 = n2180 ^ n2098;
  assign n2267 = n2266 ^ n2260;
  assign n2040 = n1955 ^ x418;
  assign n2041 = n2040 ^ n2036;
  assign n2042 = n2041 ^ x354;
  assign n2268 = n2267 ^ n2042;
  assign n41698 = n41697 ^ n2268;
  assign n2167 = n2088 ^ x322;
  assign n2168 = n2167 ^ n678;
  assign n2169 = n2168 ^ x258;
  assign n2372 = n2266 ^ n2169;
  assign n2376 = n2375 ^ n2372;
  assign n2118 = n2036 ^ x258;
  assign n2119 = n2118 ^ x450;
  assign n2120 = n2119 ^ x194;
  assign n2377 = n2376 ^ n2120;
  assign n2277 = n2169 ^ x417;
  assign n679 = n678 ^ x162;
  assign n680 = n679 ^ x354;
  assign n681 = n680 ^ x98;
  assign n2278 = n2277 ^ n681;
  assign n2279 = n2278 ^ x353;
  assign n28626 = n2377 ^ n2279;
  assign n23150 = n2375 ^ n681;
  assign n2025 = n1943 ^ x354;
  assign n2029 = n2028 ^ n2025;
  assign n2030 = n2029 ^ x290;
  assign n23151 = n23150 ^ n2030;
  assign n23152 = n23151 ^ n2213;
  assign n28627 = n28626 ^ n23152;
  assign n2214 = n2120 ^ x353;
  assign n2215 = n2214 ^ n2213;
  assign n2216 = n2215 ^ x289;
  assign n28628 = n28627 ^ n2216;
  assign n2385 = n2342 ^ n2279;
  assign n682 = n681 ^ x257;
  assign n683 = n682 ^ x449;
  assign n684 = n683 ^ x193;
  assign n2386 = n2385 ^ n684;
  assign n2387 = n2386 ^ x448;
  assign n30516 = n28628 ^ n2387;
  assign n25017 = n23152 ^ n684;
  assign n2113 = n2028 ^ x194;
  assign n2114 = n2113 ^ x386;
  assign n2115 = n2114 ^ x130;
  assign n2112 = n2030 ^ x449;
  assign n2116 = n2115 ^ n2112;
  assign n2117 = n2116 ^ x385;
  assign n25018 = n25017 ^ n2117;
  assign n25019 = n25018 ^ n2315;
  assign n30517 = n30516 ^ n25019;
  assign n2319 = n2216 ^ x448;
  assign n2320 = n2319 ^ n2315;
  assign n2321 = n2320 ^ x384;
  assign n30518 = n30517 ^ n2321;
  assign n23086 = n14474 ^ n2387;
  assign n685 = n684 ^ x352;
  assign n516 = x449 ^ x97;
  assign n517 = n516 ^ x289;
  assign n518 = n517 ^ x33;
  assign n686 = n685 ^ n518;
  assign n687 = n686 ^ x288;
  assign n23087 = n23086 ^ n687;
  assign n13564 = x448 ^ x96;
  assign n13565 = n13564 ^ x288;
  assign n13566 = n13565 ^ x32;
  assign n23088 = n23087 ^ n13566;
  assign n33254 = n30518 ^ n23088;
  assign n27145 = n25019 ^ n687;
  assign n2206 = n2115 ^ x289;
  assign n2207 = n2206 ^ x481;
  assign n2208 = n2207 ^ x225;
  assign n2205 = n2117 ^ n518;
  assign n2209 = n2208 ^ n2205;
  assign n2210 = n2209 ^ x480;
  assign n27146 = n27145 ^ n2210;
  assign n27147 = n27146 ^ n16889;
  assign n33255 = n33254 ^ n27147;
  assign n22138 = n2321 ^ x511;
  assign n22139 = n22138 ^ n16889;
  assign n22140 = n22139 ^ n13566;
  assign n33256 = n33255 ^ n22140;
  assign n25013 = n23088 ^ n16654;
  assign n688 = n687 ^ x479;
  assign n519 = n518 ^ x192;
  assign n520 = n519 ^ x384;
  assign n521 = n520 ^ x128;
  assign n689 = n688 ^ n521;
  assign n690 = n689 ^ x415;
  assign n25014 = n25013 ^ n690;
  assign n15246 = n13566 ^ x223;
  assign n15247 = n15246 ^ x415;
  assign n15248 = n15247 ^ x159;
  assign n25015 = n25014 ^ n15248;
  assign n35562 = n33256 ^ n25015;
  assign n28807 = n27147 ^ n690;
  assign n2305 = n2208 ^ x384;
  assign n2309 = n2308 ^ n2305;
  assign n2310 = n2309 ^ x320;
  assign n2304 = n2210 ^ n521;
  assign n2311 = n2310 ^ n2304;
  assign n2312 = n2311 ^ n2303;
  assign n28808 = n28807 ^ n2312;
  assign n28809 = n28808 ^ n18929;
  assign n35563 = n35562 ^ n28809;
  assign n23698 = n22140 ^ n15248;
  assign n23699 = n23698 ^ n18929;
  assign n526 = x511 ^ x159;
  assign n527 = n526 ^ x351;
  assign n528 = n527 ^ x95;
  assign n23700 = n23699 ^ n528;
  assign n35564 = n35563 ^ n23700;
  assign n2145 = n2115 ^ n2057;
  assign n2140 = n2052 ^ x386;
  assign n2141 = n2140 ^ n2021;
  assign n2142 = n2141 ^ x322;
  assign n2146 = n2145 ^ n2142;
  assign n2150 = n2149 ^ n2146;
  assign n2237 = n2208 ^ n2150;
  assign n2234 = n2142 ^ x481;
  assign n2105 = n2021 ^ x226;
  assign n2106 = n2105 ^ x418;
  assign n2107 = n2106 ^ x162;
  assign n2235 = n2234 ^ n2107;
  assign n2236 = n2235 ^ x417;
  assign n2238 = n2237 ^ n2236;
  assign n2242 = n2241 ^ n2238;
  assign n3351 = ~x30 & ~x31;
  assign n3352 = x29 & ~n3351;
  assign n3353 = x28 & n3352;
  assign n3354 = ~x27 & ~n3353;
  assign n3355 = ~x26 & n3354;
  assign n3356 = x25 & ~n3355;
  assign n3357 = ~x24 & ~n3356;
  assign n3358 = x23 & ~n3357;
  assign n3359 = x22 & n3358;
  assign n3515 = n3359 ^ x21;
  assign n3508 = n3357 ^ x23;
  assign n3424 = n3354 ^ x26;
  assign n3416 = n3352 ^ x28;
  assign n3360 = x21 & n3359;
  assign n3361 = ~x20 & ~n3360;
  assign n3362 = ~x19 & n3361;
  assign n3363 = x18 & ~n3362;
  assign n3364 = x17 & n3363;
  assign n3365 = ~x16 & ~n3364;
  assign n3366 = x15 & ~n3365;
  assign n3367 = x14 & n3366;
  assign n3368 = ~x13 & ~n3367;
  assign n3369 = x12 & ~n3368;
  assign n3370 = ~x11 & ~n3369;
  assign n3371 = ~x10 & n3370;
  assign n3372 = x9 & ~n3371;
  assign n3373 = ~x8 & ~n3372;
  assign n3374 = ~x7 & n3373;
  assign n3375 = ~x6 & n3374;
  assign n3376 = ~x5 & n3375;
  assign n3380 = ~x4 & n3376;
  assign n3388 = ~x3 & n3380;
  assign n3392 = x2 & ~n3388;
  assign n3393 = x1 & n3392;
  assign n3394 = n3393 ^ x0;
  assign n3389 = n3388 ^ x2;
  assign n3397 = n3392 ^ x1;
  assign n3402 = ~n3389 & n3397;
  assign n3381 = n3380 ^ x3;
  assign n3395 = n3381 & n3389;
  assign n3396 = n3395 ^ n3389;
  assign n3398 = n3397 ^ n3396;
  assign n3399 = n3398 ^ n3395;
  assign n3400 = ~n3398 & n3399;
  assign n3401 = n3400 ^ n3399;
  assign n3403 = n3402 ^ n3401;
  assign n3404 = n3394 & n3403;
  assign n3405 = x31 & n3404;
  assign n3406 = x31 ^ x30;
  assign n3412 = n3405 & n3406;
  assign n3413 = n3351 ^ x29;
  assign n3417 = n3412 & n3413;
  assign n3420 = n3416 & ~n3417;
  assign n3421 = n3353 ^ x27;
  assign n3425 = ~n3420 & n3421;
  assign n3443 = ~n3424 & n3425;
  assign n3444 = n3355 ^ x25;
  assign n3509 = n3443 & n3444;
  assign n3510 = n3356 ^ x24;
  assign n3511 = n3509 & n3510;
  assign n3512 = n3508 & n3511;
  assign n3513 = n3358 ^ x22;
  assign n3514 = n3512 & ~n3513;
  assign n3543 = n3515 ^ n3514;
  assign n3536 = n3513 ^ n3512;
  assign n3537 = n3511 ^ n3508;
  assign n3445 = n3444 ^ n3443;
  assign n3407 = n3406 ^ n3405;
  assign n3408 = n3404 ^ x31;
  assign n3409 = n3394 & ~n3401;
  assign n3410 = n3408 & n3409;
  assign n3411 = n3407 & n3410;
  assign n3414 = n3413 ^ n3412;
  assign n3415 = ~n3411 & ~n3414;
  assign n3418 = n3417 ^ n3416;
  assign n3419 = n3415 & ~n3418;
  assign n3422 = n3421 ^ n3420;
  assign n3423 = n3419 & n3422;
  assign n3426 = n3425 ^ n3424;
  assign n3446 = ~n3423 & ~n3426;
  assign n3538 = ~n3445 & ~n3446;
  assign n3539 = n3510 ^ n3509;
  assign n3540 = ~n3538 & n3539;
  assign n3541 = ~n3537 & ~n3540;
  assign n3542 = ~n3536 & ~n3541;
  assign n3568 = n3543 ^ n3542;
  assign n3569 = n3541 ^ n3536;
  assign n3570 = n3540 ^ n3537;
  assign n3427 = n3426 ^ n3423;
  assign n3428 = n3422 ^ n3419;
  assign n3429 = n3418 ^ n3415;
  assign n3430 = n3414 ^ n3411;
  assign n3377 = n3376 ^ x4;
  assign n3431 = n3377 & n3400;
  assign n3432 = n3431 ^ n3399;
  assign n3433 = n3402 ^ n3394;
  assign n3434 = n3432 & ~n3433;
  assign n3435 = n3409 ^ n3408;
  assign n3436 = ~n3434 & ~n3435;
  assign n3437 = n3410 ^ n3407;
  assign n3438 = n3436 & ~n3437;
  assign n3439 = ~n3430 & ~n3438;
  assign n3440 = n3429 & n3439;
  assign n3441 = n3428 & ~n3440;
  assign n3442 = ~n3427 & n3441;
  assign n3447 = n3446 ^ n3445;
  assign n3571 = ~n3442 & ~n3447;
  assign n3572 = n3539 ^ n3538;
  assign n3573 = n3571 & ~n3572;
  assign n3574 = ~n3570 & n3573;
  assign n3575 = n3569 & n3574;
  assign n3576 = ~n3568 & ~n3575;
  assign n3544 = ~n3542 & n3543;
  assign n3516 = n3514 & ~n3515;
  assign n3507 = n3360 ^ x20;
  assign n3535 = n3516 ^ n3507;
  assign n3567 = n3544 ^ n3535;
  assign n3628 = n3576 ^ n3567;
  assign n3629 = n3628 ^ x47;
  assign n3450 = n3440 ^ n3428;
  assign n3451 = n3450 ^ x54;
  assign n3454 = n3437 ^ n3436;
  assign n3455 = n3454 ^ x57;
  assign n3456 = n3435 ^ n3434;
  assign n3457 = n3456 ^ x58;
  assign n3459 = ~n3377 & n3395;
  assign n3460 = n3459 ^ n3398;
  assign n3461 = n3460 ^ x60;
  assign n3387 = n3377 & n3381;
  assign n3390 = n3389 ^ n3387;
  assign n3462 = n3390 ^ x61;
  assign n3378 = x63 & ~n3377;
  assign n3379 = n3378 ^ x62;
  assign n3382 = n3381 ^ n3377;
  assign n3383 = n3382 ^ n3378;
  assign n3384 = n3379 & ~n3383;
  assign n3385 = n3384 ^ x62;
  assign n3463 = n3390 ^ n3385;
  assign n3464 = n3462 & ~n3463;
  assign n3465 = n3464 ^ x61;
  assign n3466 = n3465 ^ n3460;
  assign n3467 = n3461 & ~n3466;
  assign n3468 = n3467 ^ x60;
  assign n3458 = n3433 ^ n3432;
  assign n3469 = n3468 ^ n3458;
  assign n3470 = n3458 ^ x59;
  assign n3471 = ~n3469 & n3470;
  assign n3472 = n3471 ^ x59;
  assign n3473 = n3472 ^ n3456;
  assign n3474 = n3457 & ~n3473;
  assign n3475 = n3474 ^ x58;
  assign n3476 = n3475 ^ n3454;
  assign n3477 = ~n3455 & n3476;
  assign n3478 = n3477 ^ x57;
  assign n3453 = n3438 ^ n3430;
  assign n3479 = n3478 ^ n3453;
  assign n3480 = n3453 ^ x56;
  assign n3481 = n3479 & ~n3480;
  assign n3482 = n3481 ^ x56;
  assign n3452 = n3439 ^ n3429;
  assign n3483 = n3482 ^ n3452;
  assign n3484 = n3452 ^ x55;
  assign n3485 = n3483 & ~n3484;
  assign n3486 = n3485 ^ x55;
  assign n3487 = n3486 ^ n3450;
  assign n3488 = ~n3451 & n3487;
  assign n3489 = n3488 ^ x54;
  assign n3449 = n3441 ^ n3427;
  assign n3490 = n3489 ^ n3449;
  assign n3491 = n3449 ^ x53;
  assign n3492 = n3490 & ~n3491;
  assign n3493 = n3492 ^ x53;
  assign n3448 = n3447 ^ n3442;
  assign n3494 = n3493 ^ n3448;
  assign n3634 = n3448 ^ x52;
  assign n3635 = n3494 & ~n3634;
  assign n3636 = n3635 ^ x52;
  assign n3633 = n3572 ^ n3571;
  assign n3637 = n3636 ^ n3633;
  assign n3638 = n3633 ^ x51;
  assign n3639 = ~n3637 & n3638;
  assign n3640 = n3639 ^ x51;
  assign n3632 = n3573 ^ n3570;
  assign n3641 = n3640 ^ n3632;
  assign n3642 = n3632 ^ x50;
  assign n3643 = ~n3641 & n3642;
  assign n3644 = n3643 ^ x50;
  assign n3631 = n3574 ^ n3569;
  assign n3645 = n3644 ^ n3631;
  assign n3646 = n3631 ^ x49;
  assign n3647 = n3645 & ~n3646;
  assign n3648 = n3647 ^ x49;
  assign n3630 = n3575 ^ n3568;
  assign n3649 = n3648 ^ n3630;
  assign n3650 = n3630 ^ x48;
  assign n3651 = ~n3649 & n3650;
  assign n3652 = n3651 ^ x48;
  assign n3653 = n3652 ^ n3628;
  assign n3654 = ~n3629 & n3653;
  assign n3655 = n3654 ^ x47;
  assign n3577 = ~n3567 & n3576;
  assign n3545 = ~n3535 & n3544;
  assign n3518 = n3361 ^ x19;
  assign n3517 = n3507 & n3516;
  assign n3534 = n3518 ^ n3517;
  assign n3566 = n3545 ^ n3534;
  assign n3627 = n3577 ^ n3566;
  assign n3656 = n3655 ^ n3627;
  assign n3657 = n3627 ^ x46;
  assign n3658 = ~n3656 & n3657;
  assign n3659 = n3658 ^ x46;
  assign n3519 = n3517 & ~n3518;
  assign n3496 = n3362 ^ x18;
  assign n3547 = n3519 ^ n3496;
  assign n3546 = ~n3534 & ~n3545;
  assign n3579 = n3547 ^ n3546;
  assign n3578 = n3566 & ~n3577;
  assign n3626 = n3579 ^ n3578;
  assign n3660 = n3659 ^ n3626;
  assign n3661 = n3626 ^ x45;
  assign n3662 = ~n3660 & n3661;
  assign n3663 = n3662 ^ x45;
  assign n3521 = n3363 ^ x17;
  assign n3520 = ~n3496 & ~n3519;
  assign n3549 = n3521 ^ n3520;
  assign n3548 = ~n3546 & n3547;
  assign n3581 = n3549 ^ n3548;
  assign n3580 = ~n3578 & ~n3579;
  assign n3625 = n3581 ^ n3580;
  assign n3664 = n3663 ^ n3625;
  assign n3853 = n3664 ^ x44;
  assign n3815 = n3652 ^ n3629;
  assign n3529 = n3370 ^ x10;
  assign n3816 = n3815 ^ n3529;
  assign n3817 = n3649 ^ x48;
  assign n3818 = n3645 ^ x49;
  assign n3819 = n3641 ^ x50;
  assign n3820 = n3637 ^ x51;
  assign n3504 = n3366 ^ x14;
  assign n3821 = n3820 ^ n3504;
  assign n3495 = n3494 ^ x52;
  assign n3778 = n3490 ^ x53;
  assign n3783 = n3486 ^ x54;
  assign n3784 = n3783 ^ n3450;
  assign n3788 = n3483 ^ x55;
  assign n3822 = n3788 ^ n3496;
  assign n3792 = n3479 ^ x56;
  assign n3796 = n3475 ^ x57;
  assign n3797 = n3796 ^ n3454;
  assign n3801 = n3472 ^ x58;
  assign n3802 = n3801 ^ n3456;
  assign n3806 = n3469 ^ x59;
  assign n3823 = n3806 ^ n3513;
  assign n3386 = n3385 ^ x61;
  assign n3391 = n3390 ^ n3386;
  assign n3498 = n3382 ^ n3379;
  assign n3499 = n3377 ^ x63;
  assign n3500 = n3499 ^ n3424;
  assign n3506 = n3364 ^ x16;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = n3506 & n3522;
  assign n3505 = n3365 ^ x15;
  assign n3552 = n3523 ^ n3505;
  assign n3533 = n3522 ^ n3506;
  assign n3550 = n3548 & ~n3549;
  assign n3551 = n3533 & ~n3550;
  assign n3584 = n3552 ^ n3551;
  assign n3565 = n3550 ^ n3533;
  assign n3582 = n3580 & ~n3581;
  assign n3583 = n3565 & n3582;
  assign n3622 = n3584 ^ n3583;
  assign n3623 = n3622 ^ x42;
  assign n3665 = n3625 ^ x44;
  assign n3666 = n3664 & ~n3665;
  assign n3667 = n3666 ^ x44;
  assign n3624 = n3582 ^ n3565;
  assign n3668 = n3667 ^ n3624;
  assign n3669 = n3624 ^ x43;
  assign n3670 = ~n3668 & n3669;
  assign n3671 = n3670 ^ x43;
  assign n3672 = n3671 ^ n3622;
  assign n3673 = ~n3623 & n3672;
  assign n3674 = n3673 ^ x42;
  assign n3585 = n3583 & ~n3584;
  assign n3553 = n3551 & n3552;
  assign n3524 = n3505 & n3523;
  assign n3532 = n3524 ^ n3504;
  assign n3564 = n3553 ^ n3532;
  assign n3621 = n3585 ^ n3564;
  assign n3675 = n3674 ^ n3621;
  assign n3676 = n3621 ^ x41;
  assign n3677 = n3675 & ~n3676;
  assign n3678 = n3677 ^ x41;
  assign n3586 = ~n3564 & n3585;
  assign n3554 = n3532 & ~n3553;
  assign n3525 = ~n3504 & n3524;
  assign n3503 = n3367 ^ x13;
  assign n3531 = n3525 ^ n3503;
  assign n3563 = n3554 ^ n3531;
  assign n3620 = n3586 ^ n3563;
  assign n3679 = n3678 ^ n3620;
  assign n3680 = n3620 ^ x40;
  assign n3681 = ~n3679 & n3680;
  assign n3682 = n3681 ^ x40;
  assign n3587 = n3563 & ~n3586;
  assign n3526 = n3503 & n3525;
  assign n3502 = n3368 ^ x12;
  assign n3556 = n3526 ^ n3502;
  assign n3555 = ~n3531 & n3554;
  assign n3562 = n3556 ^ n3555;
  assign n3619 = n3587 ^ n3562;
  assign n3683 = n3682 ^ n3619;
  assign n3684 = n3619 ^ x39;
  assign n3685 = ~n3683 & n3684;
  assign n3686 = n3685 ^ x39;
  assign n3588 = ~n3562 & ~n3587;
  assign n3527 = n3502 & n3526;
  assign n3501 = n3369 ^ x11;
  assign n3558 = n3527 ^ n3501;
  assign n3557 = n3555 & ~n3556;
  assign n3561 = n3558 ^ n3557;
  assign n3618 = n3588 ^ n3561;
  assign n3687 = n3686 ^ n3618;
  assign n3688 = n3618 ^ x38;
  assign n3689 = ~n3687 & n3688;
  assign n3690 = n3689 ^ x38;
  assign n3589 = n3561 & ~n3588;
  assign n3559 = n3557 & ~n3558;
  assign n3528 = n3501 & n3527;
  assign n3530 = n3529 ^ n3528;
  assign n3560 = n3559 ^ n3530;
  assign n3617 = n3589 ^ n3560;
  assign n3691 = n3690 ^ n3617;
  assign n3692 = n3617 ^ x37;
  assign n3693 = ~n3691 & n3692;
  assign n3694 = n3693 ^ x37;
  assign n3593 = n3371 ^ x9;
  assign n3592 = ~n3528 & n3529;
  assign n3594 = n3593 ^ n3592;
  assign n3591 = ~n3530 & n3559;
  assign n3595 = n3594 ^ n3591;
  assign n3590 = ~n3560 & ~n3589;
  assign n3616 = n3595 ^ n3590;
  assign n3695 = n3694 ^ n3616;
  assign n3696 = n3616 ^ x36;
  assign n3697 = n3695 & ~n3696;
  assign n3698 = n3697 ^ x36;
  assign n3600 = n3591 & n3594;
  assign n3598 = n3372 ^ x8;
  assign n3597 = ~n3592 & n3593;
  assign n3599 = n3598 ^ n3597;
  assign n3601 = n3600 ^ n3599;
  assign n3596 = ~n3590 & ~n3595;
  assign n3615 = n3601 ^ n3596;
  assign n3699 = n3698 ^ n3615;
  assign n3700 = n3615 ^ x35;
  assign n3701 = ~n3699 & n3700;
  assign n3702 = n3701 ^ x35;
  assign n3606 = n3599 & ~n3600;
  assign n3604 = n3373 ^ x7;
  assign n3603 = n3597 & n3598;
  assign n3605 = n3604 ^ n3603;
  assign n3607 = n3606 ^ n3605;
  assign n3602 = n3596 & ~n3601;
  assign n3614 = n3607 ^ n3602;
  assign n3703 = n3702 ^ n3614;
  assign n3704 = n3614 ^ x34;
  assign n3705 = ~n3703 & n3704;
  assign n3706 = n3705 ^ x34;
  assign n3611 = n3374 ^ x6;
  assign n3609 = n3606 ^ n3604;
  assign n3610 = n3605 & n3609;
  assign n3612 = n3611 ^ n3610;
  assign n3608 = ~n3602 & ~n3607;
  assign n3613 = n3612 ^ n3608;
  assign n3707 = n3706 ^ n3613;
  assign n3708 = n3707 ^ x33;
  assign n3709 = n3699 ^ x35;
  assign n3710 = n3406 & n3709;
  assign n3711 = n3703 ^ x34;
  assign n3712 = n3710 & n3711;
  assign n3713 = ~n3708 & n3712;
  assign n3718 = n3613 ^ x33;
  assign n3719 = n3707 & ~n3718;
  assign n3720 = n3719 ^ x33;
  assign n3716 = n3375 ^ x5;
  assign n3714 = ~n3611 & n3613;
  assign n3715 = n3714 ^ n3611;
  assign n3717 = n3716 ^ n3715;
  assign n3721 = n3720 ^ n3717;
  assign n3722 = n3721 ^ x32;
  assign n3723 = n3713 & n3722;
  assign n3724 = n3723 ^ n3499;
  assign n3725 = n3500 & n3724;
  assign n3726 = n3725 ^ n3424;
  assign n3824 = ~n3498 & n3726;
  assign n3825 = ~n3391 & n3824;
  assign n3826 = n3465 ^ n3461;
  assign n3827 = ~n3825 & n3826;
  assign n3828 = n3827 ^ n3806;
  assign n3829 = ~n3823 & ~n3828;
  assign n3830 = n3829 ^ n3513;
  assign n3831 = n3802 & ~n3830;
  assign n3832 = n3797 & ~n3831;
  assign n3833 = ~n3792 & ~n3832;
  assign n3834 = n3833 ^ n3788;
  assign n3835 = ~n3822 & n3834;
  assign n3836 = n3835 ^ n3496;
  assign n3837 = n3784 & ~n3836;
  assign n3838 = ~n3778 & ~n3837;
  assign n3839 = n3495 & ~n3838;
  assign n3840 = n3839 ^ n3820;
  assign n3841 = ~n3821 & n3840;
  assign n3842 = n3841 ^ n3504;
  assign n3843 = n3819 & ~n3842;
  assign n3844 = ~n3818 & n3843;
  assign n3845 = ~n3817 & ~n3844;
  assign n3846 = n3845 ^ n3815;
  assign n3847 = n3816 & ~n3846;
  assign n3848 = n3847 ^ n3529;
  assign n3849 = n3656 ^ x46;
  assign n3850 = n3848 & ~n3849;
  assign n3851 = n3660 ^ x45;
  assign n3852 = n3850 & ~n3851;
  assign n3868 = n3853 ^ n3852;
  assign n3869 = n3851 ^ n3850;
  assign n3870 = n3849 ^ n3848;
  assign n3871 = n3838 ^ n3495;
  assign n3872 = n3837 ^ n3778;
  assign n3873 = n3836 ^ n3784;
  assign n3874 = n3833 ^ n3822;
  assign n3875 = n3832 ^ n3792;
  assign n3876 = n3830 ^ n3802;
  assign n3877 = n3826 ^ n3825;
  assign n3878 = n3824 ^ n3391;
  assign n3727 = n3726 ^ n3498;
  assign n3728 = n3712 ^ n3708;
  assign n3729 = n3709 ^ n3406;
  assign n3730 = n3711 ^ n3710;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = n3728 & n3731;
  assign n3733 = n3722 ^ n3713;
  assign n3734 = n3732 & ~n3733;
  assign n3735 = n3723 ^ n3500;
  assign n3736 = n3734 & ~n3735;
  assign n3879 = ~n3727 & n3736;
  assign n3880 = ~n3878 & n3879;
  assign n3881 = ~n3877 & ~n3880;
  assign n3882 = n3827 ^ n3823;
  assign n3883 = n3881 & ~n3882;
  assign n3884 = n3876 & ~n3883;
  assign n3885 = n3831 ^ n3797;
  assign n3886 = n3884 & ~n3885;
  assign n3887 = ~n3875 & n3886;
  assign n3888 = ~n3874 & ~n3887;
  assign n3889 = ~n3873 & ~n3888;
  assign n3890 = ~n3872 & n3889;
  assign n3891 = n3871 & ~n3890;
  assign n3892 = n3839 ^ n3821;
  assign n3893 = ~n3891 & ~n3892;
  assign n3894 = n3842 ^ n3819;
  assign n3895 = ~n3893 & ~n3894;
  assign n3896 = n3843 ^ n3818;
  assign n3897 = ~n3895 & n3896;
  assign n3898 = n3844 ^ n3817;
  assign n3899 = n3897 & n3898;
  assign n3900 = n3845 ^ n3816;
  assign n3901 = n3899 & n3900;
  assign n3902 = n3870 & ~n3901;
  assign n3903 = ~n3869 & ~n3902;
  assign n3904 = ~n3868 & ~n3903;
  assign n3854 = n3852 & n3853;
  assign n3866 = n3854 ^ n3611;
  assign n3813 = n3668 ^ x43;
  assign n3867 = n3866 ^ n3813;
  assign n3957 = n3904 ^ n3867;
  assign n3920 = n3901 ^ n3870;
  assign n3921 = n3896 ^ n3895;
  assign n3922 = n3894 ^ n3893;
  assign n3923 = n3892 ^ n3891;
  assign n3924 = n3890 ^ n3871;
  assign n3925 = n3889 ^ n3872;
  assign n3926 = n3888 ^ n3873;
  assign n3927 = n3887 ^ n3874;
  assign n3928 = n3885 ^ n3884;
  assign n3929 = n3880 ^ n3877;
  assign n3737 = n3736 ^ n3727;
  assign n3738 = n3695 ^ x36;
  assign n3739 = ~n3729 & ~n3738;
  assign n3740 = n3730 ^ n3729;
  assign n3741 = n3739 & ~n3740;
  assign n3742 = n3731 ^ n3728;
  assign n3743 = ~n3741 & n3742;
  assign n3744 = n3733 ^ n3732;
  assign n3745 = n3743 & ~n3744;
  assign n3746 = n3735 ^ n3734;
  assign n3747 = ~n3745 & n3746;
  assign n3930 = n3737 & n3747;
  assign n3931 = n3879 ^ n3878;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = ~n3929 & n3932;
  assign n3934 = n3882 ^ n3881;
  assign n3935 = ~n3933 & ~n3934;
  assign n3936 = n3883 ^ n3876;
  assign n3937 = n3935 & n3936;
  assign n3938 = ~n3928 & ~n3937;
  assign n3939 = n3886 ^ n3875;
  assign n3940 = n3938 & ~n3939;
  assign n3941 = ~n3927 & n3940;
  assign n3942 = n3926 & n3941;
  assign n3943 = n3925 & ~n3942;
  assign n3944 = ~n3924 & n3943;
  assign n3945 = n3923 & ~n3944;
  assign n3946 = n3922 & ~n3945;
  assign n3947 = n3921 & n3946;
  assign n3948 = n3898 ^ n3897;
  assign n3949 = n3947 & ~n3948;
  assign n3950 = n3900 ^ n3899;
  assign n3951 = n3949 & ~n3950;
  assign n3952 = ~n3920 & n3951;
  assign n3953 = n3902 ^ n3869;
  assign n3954 = ~n3952 & n3953;
  assign n3955 = n3903 ^ n3868;
  assign n3956 = ~n3954 & n3955;
  assign n3976 = n3957 ^ n3956;
  assign n3977 = n3976 ^ x70;
  assign n3981 = n3950 ^ n3949;
  assign n3982 = n3981 ^ x74;
  assign n3983 = n3948 ^ n3947;
  assign n3984 = n3983 ^ x75;
  assign n3988 = n3943 ^ n3924;
  assign n3989 = n3988 ^ x79;
  assign n3749 = n3746 ^ n3745;
  assign n3750 = n3749 ^ x90;
  assign n3754 = x95 & n3738;
  assign n3755 = n3754 ^ x94;
  assign n3756 = n3738 ^ n3729;
  assign n3757 = n3756 ^ n3754;
  assign n3758 = n3755 & ~n3757;
  assign n3759 = n3758 ^ x94;
  assign n3753 = n3740 ^ n3739;
  assign n3760 = n3759 ^ n3753;
  assign n3761 = n3753 ^ x93;
  assign n3762 = n3760 & ~n3761;
  assign n3763 = n3762 ^ x93;
  assign n3752 = n3742 ^ n3741;
  assign n3764 = n3763 ^ n3752;
  assign n3765 = n3752 ^ x92;
  assign n3766 = ~n3764 & n3765;
  assign n3767 = n3766 ^ x92;
  assign n3751 = n3744 ^ n3743;
  assign n3768 = n3767 ^ n3751;
  assign n3769 = n3751 ^ x91;
  assign n3770 = ~n3768 & n3769;
  assign n3771 = n3770 ^ x91;
  assign n3772 = n3771 ^ n3749;
  assign n3773 = ~n3750 & n3772;
  assign n3774 = n3773 ^ x90;
  assign n3748 = n3747 ^ n3737;
  assign n3775 = n3774 ^ n3748;
  assign n3999 = n3748 ^ x89;
  assign n4000 = ~n3775 & n3999;
  assign n4001 = n4000 ^ x89;
  assign n3998 = n3931 ^ n3930;
  assign n4002 = n4001 ^ n3998;
  assign n4003 = n3998 ^ x88;
  assign n4004 = n4002 & ~n4003;
  assign n4005 = n4004 ^ x88;
  assign n3997 = n3932 ^ n3929;
  assign n4006 = n4005 ^ n3997;
  assign n4007 = n3997 ^ x87;
  assign n4008 = ~n4006 & n4007;
  assign n4009 = n4008 ^ x87;
  assign n3996 = n3934 ^ n3933;
  assign n4010 = n4009 ^ n3996;
  assign n4011 = n3996 ^ x86;
  assign n4012 = ~n4010 & n4011;
  assign n4013 = n4012 ^ x86;
  assign n3995 = n3936 ^ n3935;
  assign n4014 = n4013 ^ n3995;
  assign n4015 = n3995 ^ x85;
  assign n4016 = ~n4014 & n4015;
  assign n4017 = n4016 ^ x85;
  assign n3994 = n3937 ^ n3928;
  assign n4018 = n4017 ^ n3994;
  assign n4019 = n3994 ^ x84;
  assign n4020 = n4018 & ~n4019;
  assign n4021 = n4020 ^ x84;
  assign n3993 = n3939 ^ n3938;
  assign n4022 = n4021 ^ n3993;
  assign n4023 = n3993 ^ x83;
  assign n4024 = ~n4022 & n4023;
  assign n4025 = n4024 ^ x83;
  assign n3992 = n3940 ^ n3927;
  assign n4026 = n4025 ^ n3992;
  assign n4027 = n3992 ^ x82;
  assign n4028 = ~n4026 & n4027;
  assign n4029 = n4028 ^ x82;
  assign n3991 = n3941 ^ n3926;
  assign n4030 = n4029 ^ n3991;
  assign n4031 = n3991 ^ x81;
  assign n4032 = n4030 & ~n4031;
  assign n4033 = n4032 ^ x81;
  assign n3990 = n3942 ^ n3925;
  assign n4034 = n4033 ^ n3990;
  assign n4035 = n3990 ^ x80;
  assign n4036 = n4034 & ~n4035;
  assign n4037 = n4036 ^ x80;
  assign n4038 = n4037 ^ n3988;
  assign n4039 = ~n3989 & n4038;
  assign n4040 = n4039 ^ x79;
  assign n3987 = n3944 ^ n3923;
  assign n4041 = n4040 ^ n3987;
  assign n4042 = n3987 ^ x78;
  assign n4043 = ~n4041 & n4042;
  assign n4044 = n4043 ^ x78;
  assign n3986 = n3945 ^ n3922;
  assign n4045 = n4044 ^ n3986;
  assign n4046 = n3986 ^ x77;
  assign n4047 = n4045 & ~n4046;
  assign n4048 = n4047 ^ x77;
  assign n3985 = n3946 ^ n3921;
  assign n4049 = n4048 ^ n3985;
  assign n4050 = n3985 ^ x76;
  assign n4051 = ~n4049 & n4050;
  assign n4052 = n4051 ^ x76;
  assign n4053 = n4052 ^ n3983;
  assign n4054 = ~n3984 & n4053;
  assign n4055 = n4054 ^ x75;
  assign n4056 = n4055 ^ n3981;
  assign n4057 = ~n3982 & n4056;
  assign n4058 = n4057 ^ x74;
  assign n3980 = n3951 ^ n3920;
  assign n4059 = n4058 ^ n3980;
  assign n4060 = n3980 ^ x73;
  assign n4061 = n4059 & ~n4060;
  assign n4062 = n4061 ^ x73;
  assign n3979 = n3953 ^ n3952;
  assign n4063 = n4062 ^ n3979;
  assign n4064 = n3979 ^ x72;
  assign n4065 = ~n4063 & n4064;
  assign n4066 = n4065 ^ x72;
  assign n3978 = n3955 ^ n3954;
  assign n4067 = n4066 ^ n3978;
  assign n4068 = n3978 ^ x71;
  assign n4069 = n4067 & ~n4068;
  assign n4070 = n4069 ^ x71;
  assign n4071 = n4070 ^ n3976;
  assign n4072 = ~n3977 & n4071;
  assign n4073 = n4072 ^ x70;
  assign n3905 = n3867 & n3904;
  assign n3814 = n3813 ^ n3611;
  assign n3855 = n3854 ^ n3813;
  assign n3856 = ~n3814 & n3855;
  assign n3857 = n3856 ^ n3611;
  assign n3811 = n3671 ^ x42;
  assign n3812 = n3811 ^ n3622;
  assign n3865 = n3857 ^ n3812;
  assign n3959 = n3905 ^ n3865;
  assign n3958 = ~n3956 & ~n3957;
  assign n3975 = n3959 ^ n3958;
  assign n4074 = n4073 ^ n3975;
  assign n4075 = n3975 ^ x69;
  assign n4076 = n4074 & ~n4075;
  assign n4077 = n4076 ^ x69;
  assign n3906 = n3865 & n3905;
  assign n3858 = ~n3812 & ~n3857;
  assign n3810 = n3675 ^ x41;
  assign n3864 = n3858 ^ n3810;
  assign n3961 = n3906 ^ n3864;
  assign n3960 = ~n3958 & n3959;
  assign n3974 = n3961 ^ n3960;
  assign n4078 = n4077 ^ n3974;
  assign n4102 = n4078 ^ x68;
  assign n4101 = ~n3413 & ~n3499;
  assign n4174 = n4102 ^ n4101;
  assign n4518 = n4174 ^ x127;
  assign n3794 = n3760 ^ x93;
  assign n5224 = n3794 ^ n3391;
  assign n5225 = ~n4518 & ~n5224;
  assign n5226 = n5225 ^ n3391;
  assign n4523 = n4070 ^ n3977;
  assign n5031 = n3738 ^ n3377;
  assign n5032 = ~n4523 & ~n5031;
  assign n5033 = n5032 ^ n3377;
  assign n4214 = n3504 & n3817;
  assign n4213 = n4014 ^ x85;
  assign n4215 = n4214 ^ n4213;
  assign n4205 = n3505 & ~n3818;
  assign n4204 = n4010 ^ x86;
  assign n4206 = n4205 ^ n4204;
  assign n4195 = ~n3506 & n3819;
  assign n4194 = n4006 ^ x87;
  assign n4196 = n4195 ^ n4194;
  assign n4142 = n4002 ^ x88;
  assign n4141 = n3521 & n3820;
  assign n4143 = n4142 ^ n4141;
  assign n3776 = n3775 ^ x89;
  assign n3497 = ~n3495 & n3496;
  assign n3777 = n3776 ^ n3497;
  assign n3780 = n3771 ^ x90;
  assign n3781 = n3780 ^ n3749;
  assign n3779 = n3518 & ~n3778;
  assign n3782 = n3781 ^ n3779;
  assign n3786 = n3768 ^ x91;
  assign n3785 = ~n3507 & ~n3784;
  assign n3787 = n3786 ^ n3785;
  assign n3790 = n3764 ^ x92;
  assign n3789 = n3515 & ~n3788;
  assign n3791 = n3790 ^ n3789;
  assign n3793 = ~n3513 & ~n3792;
  assign n3795 = n3794 ^ n3793;
  assign n3799 = n3756 ^ n3755;
  assign n3798 = n3508 & ~n3797;
  assign n3800 = n3799 ^ n3798;
  assign n3804 = n3738 ^ x95;
  assign n3803 = ~n3510 & n3802;
  assign n3805 = n3804 ^ n3803;
  assign n3962 = ~n3960 & n3961;
  assign n3907 = ~n3864 & ~n3906;
  assign n3860 = n3679 ^ x40;
  assign n3859 = n3810 & ~n3858;
  assign n3863 = n3860 ^ n3859;
  assign n3919 = n3907 ^ n3863;
  assign n3972 = n3962 ^ n3919;
  assign n3973 = n3972 ^ x67;
  assign n4079 = n3974 ^ x68;
  assign n4080 = ~n4078 & n4079;
  assign n4081 = n4080 ^ x68;
  assign n4082 = n4081 ^ n3972;
  assign n4083 = n3973 & ~n4082;
  assign n4084 = n4083 ^ x67;
  assign n3908 = ~n3863 & n3907;
  assign n3861 = n3859 & ~n3860;
  assign n3808 = n3683 ^ x39;
  assign n3809 = n3808 ^ n3389;
  assign n3862 = n3861 ^ n3809;
  assign n3964 = n3908 ^ n3862;
  assign n3963 = ~n3919 & n3962;
  assign n3971 = n3964 ^ n3963;
  assign n4085 = n4084 ^ n3971;
  assign n4086 = n3971 ^ x66;
  assign n4087 = n4085 & ~n4086;
  assign n4088 = n4087 ^ x66;
  assign n3965 = ~n3963 & n3964;
  assign n3913 = n3687 ^ x38;
  assign n3910 = n3861 ^ n3808;
  assign n3911 = n3809 & n3910;
  assign n3912 = n3911 ^ n3389;
  assign n3914 = n3913 ^ n3912;
  assign n3909 = ~n3862 & ~n3908;
  assign n3918 = n3914 ^ n3909;
  assign n3966 = n3965 ^ n3918;
  assign n4089 = n4088 ^ n3966;
  assign n4090 = n3966 ^ x65;
  assign n4091 = ~n4089 & n4090;
  assign n4092 = n4091 ^ x65;
  assign n3967 = n3918 ^ n3912;
  assign n3968 = n3966 & ~n3967;
  assign n3969 = n3968 ^ x64;
  assign n3916 = n3691 ^ x37;
  assign n3915 = n3909 & ~n3914;
  assign n3917 = n3916 ^ n3915;
  assign n3970 = n3969 ^ n3917;
  assign n4093 = n4092 ^ n3970;
  assign n3807 = ~n3444 & n3806;
  assign n4094 = n4093 ^ n3807;
  assign n4096 = n4089 ^ x65;
  assign n4095 = n3424 & n3826;
  assign n4097 = n4096 ^ n4095;
  assign n4099 = n3391 & ~n3421;
  assign n4098 = n4085 ^ x66;
  assign n4100 = n4099 ^ n4098;
  assign n4104 = n3416 & n3498;
  assign n4103 = n4101 & n4102;
  assign n4105 = n4104 ^ n4103;
  assign n4106 = n4081 ^ x67;
  assign n4107 = n4106 ^ n3972;
  assign n4108 = n4107 ^ n4104;
  assign n4109 = n4105 & ~n4108;
  assign n4110 = n4109 ^ n4103;
  assign n4111 = n4110 ^ n4098;
  assign n4112 = ~n4100 & n4111;
  assign n4113 = n4112 ^ n4099;
  assign n4114 = n4113 ^ n4096;
  assign n4115 = n4097 & ~n4114;
  assign n4116 = n4115 ^ n4095;
  assign n4117 = n4116 ^ n4093;
  assign n4118 = ~n4094 & n4117;
  assign n4119 = n4118 ^ n3807;
  assign n4120 = n4119 ^ n3804;
  assign n4121 = n3805 & ~n4120;
  assign n4122 = n4121 ^ n3803;
  assign n4123 = n4122 ^ n3799;
  assign n4124 = ~n3800 & ~n4123;
  assign n4125 = n4124 ^ n3798;
  assign n4126 = n4125 ^ n3794;
  assign n4127 = n3795 & ~n4126;
  assign n4128 = n4127 ^ n3793;
  assign n4129 = n4128 ^ n3790;
  assign n4130 = n3791 & n4129;
  assign n4131 = n4130 ^ n3789;
  assign n4132 = n4131 ^ n3786;
  assign n4133 = n3787 & ~n4132;
  assign n4134 = n4133 ^ n3785;
  assign n4135 = n4134 ^ n3781;
  assign n4136 = ~n3782 & n4135;
  assign n4137 = n4136 ^ n3779;
  assign n4138 = n4137 ^ n3776;
  assign n4139 = ~n3777 & ~n4138;
  assign n4140 = n4139 ^ n3497;
  assign n4191 = n4142 ^ n4140;
  assign n4192 = ~n4143 & ~n4191;
  assign n4193 = n4192 ^ n4141;
  assign n4201 = n4194 ^ n4193;
  assign n4202 = n4196 & ~n4201;
  assign n4203 = n4202 ^ n4195;
  assign n4210 = n4205 ^ n4203;
  assign n4211 = ~n4206 & n4210;
  assign n4212 = n4211 ^ n4204;
  assign n4311 = n4213 ^ n4212;
  assign n4312 = n4215 & ~n4311;
  assign n4313 = n4312 ^ n4214;
  assign n4309 = n4018 ^ x84;
  assign n4308 = n3503 & ~n3815;
  assign n4310 = n4309 ^ n4308;
  assign n4328 = n4313 ^ n4310;
  assign n4216 = n4215 ^ n4212;
  assign n4144 = n4143 ^ n4140;
  assign n4145 = n4134 ^ n3782;
  assign n4146 = n4128 ^ n3791;
  assign n4147 = n4125 ^ n3795;
  assign n4148 = n4119 ^ n3805;
  assign n4149 = n4107 ^ n4105;
  assign n4150 = n4110 ^ n4100;
  assign n4151 = n4149 & ~n4150;
  assign n4152 = n4113 ^ n4097;
  assign n4153 = n4151 & n4152;
  assign n4154 = n4116 ^ n4094;
  assign n4155 = n4153 & ~n4154;
  assign n4156 = ~n4148 & ~n4155;
  assign n4157 = n4122 ^ n3800;
  assign n4158 = n4156 & n4157;
  assign n4159 = n4147 & n4158;
  assign n4160 = ~n4146 & ~n4159;
  assign n4161 = n4131 ^ n3787;
  assign n4162 = ~n4160 & ~n4161;
  assign n4163 = ~n4145 & ~n4162;
  assign n4164 = n4137 ^ n3777;
  assign n4165 = ~n4163 & n4164;
  assign n4190 = n4144 & ~n4165;
  assign n4197 = n4196 ^ n4193;
  assign n4200 = ~n4190 & ~n4197;
  assign n4207 = n4206 ^ n4203;
  assign n4217 = n4200 & n4207;
  assign n4329 = n4216 & ~n4217;
  assign n4330 = ~n4328 & ~n4329;
  assign n4314 = n4313 ^ n4309;
  assign n4315 = n4310 & n4314;
  assign n4316 = n4315 ^ n4308;
  assign n4306 = ~n3502 & n3849;
  assign n4305 = n4022 ^ x83;
  assign n4307 = n4306 ^ n4305;
  assign n4327 = n4316 ^ n4307;
  assign n4344 = n4330 ^ n4327;
  assign n4345 = n4329 ^ n4328;
  assign n4166 = n4165 ^ n4144;
  assign n4167 = n4164 ^ n4163;
  assign n4168 = n4162 ^ n4145;
  assign n4169 = n4159 ^ n4146;
  assign n4170 = n4158 ^ n4147;
  assign n4171 = n4155 ^ n4148;
  assign n4172 = n4154 ^ n4153;
  assign n4173 = n4150 ^ n4149;
  assign n4175 = ~n4149 & n4174;
  assign n4176 = ~n4173 & n4175;
  assign n4177 = n4152 ^ n4151;
  assign n4178 = ~n4176 & ~n4177;
  assign n4179 = n4172 & n4178;
  assign n4180 = ~n4171 & ~n4179;
  assign n4181 = n4157 ^ n4156;
  assign n4182 = n4180 & ~n4181;
  assign n4183 = n4170 & ~n4182;
  assign n4184 = ~n4169 & n4183;
  assign n4185 = n4161 ^ n4160;
  assign n4186 = ~n4184 & ~n4185;
  assign n4187 = n4168 & n4186;
  assign n4188 = ~n4167 & ~n4187;
  assign n4189 = n4166 & n4188;
  assign n4198 = n4197 ^ n4190;
  assign n4199 = n4189 & n4198;
  assign n4208 = n4207 ^ n4200;
  assign n4209 = n4199 & n4208;
  assign n4218 = n4217 ^ n4216;
  assign n4346 = ~n4209 & ~n4218;
  assign n4347 = ~n4345 & n4346;
  assign n4348 = n4344 & ~n4347;
  assign n4317 = n4316 ^ n4305;
  assign n4318 = n4307 & n4317;
  assign n4319 = n4318 ^ n4306;
  assign n4303 = ~n3501 & n3851;
  assign n4302 = n4026 ^ x82;
  assign n4304 = n4303 ^ n4302;
  assign n4332 = n4319 ^ n4304;
  assign n4331 = n4327 & n4330;
  assign n4343 = n4332 ^ n4331;
  assign n4368 = n4348 ^ n4343;
  assign n4419 = n4368 ^ x109;
  assign n4370 = n4347 ^ n4344;
  assign n4414 = n4370 ^ x110;
  assign n4372 = n4346 ^ n4345;
  assign n4415 = n4372 ^ x111;
  assign n4373 = ~x111 & n4372;
  assign n4416 = n4415 ^ n4373;
  assign n4417 = n4414 & ~n4416;
  assign n4371 = ~x110 & ~n4370;
  assign n4418 = n4417 ^ n4371;
  assign n4219 = n4218 ^ n4209;
  assign n4220 = n4219 ^ x112;
  assign n4221 = n4208 ^ n4199;
  assign n4222 = n4221 ^ x113;
  assign n4223 = n4198 ^ n4189;
  assign n4224 = n4223 ^ x114;
  assign n4225 = n4188 ^ n4166;
  assign n4226 = n4225 ^ x115;
  assign n4227 = n4182 ^ n4170;
  assign n4228 = n4227 ^ x120;
  assign n4229 = n4181 ^ n4180;
  assign n4230 = n4229 ^ x121;
  assign n4231 = n4179 ^ n4171;
  assign n4232 = n4231 ^ x122;
  assign n4233 = n4178 ^ n4172;
  assign n4234 = n4233 ^ x123;
  assign n4235 = n4176 ^ n4151;
  assign n4236 = n4235 ^ n4152;
  assign n4237 = n4236 ^ x124;
  assign n4238 = n4175 ^ n4173;
  assign n4239 = n4238 ^ x125;
  assign n4240 = x127 & ~n4174;
  assign n4241 = n4240 ^ x126;
  assign n4242 = n4174 ^ n4149;
  assign n4243 = n4242 ^ n4240;
  assign n4244 = n4241 & n4243;
  assign n4245 = n4244 ^ x126;
  assign n4246 = n4245 ^ n4238;
  assign n4247 = ~n4239 & n4246;
  assign n4248 = n4247 ^ x125;
  assign n4249 = n4248 ^ n4236;
  assign n4250 = ~n4237 & n4249;
  assign n4251 = n4250 ^ x124;
  assign n4252 = n4251 ^ n4233;
  assign n4253 = ~n4234 & n4252;
  assign n4254 = n4253 ^ x123;
  assign n4255 = n4254 ^ n4231;
  assign n4256 = n4232 & ~n4255;
  assign n4257 = n4256 ^ x122;
  assign n4258 = n4257 ^ n4229;
  assign n4259 = ~n4230 & n4258;
  assign n4260 = n4259 ^ x121;
  assign n4261 = n4260 ^ n4227;
  assign n4262 = n4228 & ~n4261;
  assign n4263 = n4262 ^ x120;
  assign n4264 = n4186 ^ n4168;
  assign n4265 = ~x117 & ~n4264;
  assign n4266 = n4185 ^ n4184;
  assign n4267 = ~x118 & ~n4266;
  assign n4268 = n4183 ^ n4169;
  assign n4270 = x119 & n4268;
  assign n4269 = n4268 ^ x119;
  assign n4271 = n4270 ^ n4269;
  assign n4272 = ~n4267 & n4271;
  assign n4273 = n4187 ^ n4167;
  assign n4274 = ~x116 & n4273;
  assign n4275 = n4272 & ~n4274;
  assign n4276 = ~n4265 & n4275;
  assign n4277 = n4263 & n4276;
  assign n4278 = n4273 ^ x116;
  assign n4279 = n4264 ^ x117;
  assign n4280 = n4266 ^ x118;
  assign n4281 = ~n4270 & n4280;
  assign n4282 = n4281 ^ n4267;
  assign n4283 = n4282 ^ n4264;
  assign n4284 = n4279 & n4283;
  assign n4285 = n4284 ^ x117;
  assign n4286 = ~n4278 & n4285;
  assign n4287 = n4286 ^ n4278;
  assign n4288 = n4287 ^ n4274;
  assign n4289 = ~n4277 & ~n4288;
  assign n4290 = n4289 ^ n4225;
  assign n4291 = ~n4226 & ~n4290;
  assign n4292 = n4291 ^ x115;
  assign n4293 = n4292 ^ n4223;
  assign n4294 = ~n4224 & n4293;
  assign n4295 = n4294 ^ x114;
  assign n4296 = n4295 ^ n4221;
  assign n4297 = ~n4222 & n4296;
  assign n4298 = n4297 ^ x113;
  assign n4299 = n4298 ^ n4219;
  assign n4300 = n4220 & ~n4299;
  assign n4301 = n4300 ^ x112;
  assign n4374 = ~n4371 & ~n4373;
  assign n4982 = n4301 & n4374;
  assign n4983 = n4418 & ~n4982;
  assign n4984 = n4983 ^ n4368;
  assign n4985 = n4419 & n4984;
  assign n4986 = n4985 ^ x109;
  assign n4333 = ~n4331 & n4332;
  assign n4324 = n3529 & ~n3853;
  assign n4323 = n4030 ^ x81;
  assign n4325 = n4324 ^ n4323;
  assign n4320 = n4319 ^ n4302;
  assign n4321 = n4304 & ~n4320;
  assign n4322 = n4321 ^ n4303;
  assign n4326 = n4325 ^ n4322;
  assign n4350 = n4333 ^ n4326;
  assign n4349 = ~n4343 & ~n4348;
  assign n4375 = n4350 ^ n4349;
  assign n4413 = n4375 ^ x108;
  assign n4987 = n4986 ^ n4413;
  assign n4526 = n4067 ^ x71;
  assign n4979 = n3916 ^ n3716;
  assign n4980 = ~n4526 & n4979;
  assign n4981 = n4980 ^ n3716;
  assign n4988 = n4987 ^ n4981;
  assign n4528 = n4063 ^ x72;
  assign n4990 = n3913 ^ n3611;
  assign n4991 = n4528 & n4990;
  assign n4992 = n4991 ^ n3611;
  assign n4989 = n4983 ^ n4419;
  assign n4993 = n4992 ^ n4989;
  assign n4535 = n4055 ^ n3982;
  assign n5000 = n3860 ^ n3598;
  assign n5001 = ~n4535 & ~n5000;
  assign n5002 = n5001 ^ n3598;
  assign n4999 = n4415 ^ n4301;
  assign n5003 = n5002 ^ n4999;
  assign n4538 = n4052 ^ n3984;
  assign n5004 = n3810 ^ n3593;
  assign n5005 = ~n4538 & n5004;
  assign n5006 = n5005 ^ n3593;
  assign n4901 = n4298 ^ n4220;
  assign n5007 = n5006 ^ n4901;
  assign n4444 = n4049 ^ x76;
  assign n4892 = n3812 ^ n3529;
  assign n4893 = n4444 & ~n4892;
  assign n4894 = n4893 ^ n3529;
  assign n4891 = n4295 ^ n4222;
  assign n4895 = n4894 ^ n4891;
  assign n4397 = n4045 ^ x77;
  assign n4714 = n3813 ^ n3501;
  assign n4715 = ~n4397 & ~n4714;
  assign n4716 = n4715 ^ n3501;
  assign n4713 = n4292 ^ n4224;
  assign n4717 = n4716 ^ n4713;
  assign n4383 = n4041 ^ x78;
  assign n4457 = n3853 ^ n3502;
  assign n4458 = n4383 & n4457;
  assign n4459 = n4458 ^ n3502;
  assign n4455 = n4289 ^ x115;
  assign n4456 = n4455 ^ n4225;
  assign n4460 = n4459 ^ n4456;
  assign n4464 = n4263 & n4272;
  assign n4465 = n4282 & ~n4464;
  assign n4466 = n4465 ^ n4264;
  assign n4467 = n4279 & n4466;
  assign n4468 = n4467 ^ x117;
  assign n4469 = n4468 ^ n4278;
  assign n4357 = n4037 ^ n3989;
  assign n4461 = n3851 ^ n3503;
  assign n4462 = ~n4357 & ~n4461;
  assign n4463 = n4462 ^ n3503;
  assign n4470 = n4469 ^ n4463;
  assign n4340 = n4034 ^ x80;
  assign n4472 = n3849 ^ n3504;
  assign n4473 = ~n4340 & n4472;
  assign n4474 = n4473 ^ n3504;
  assign n4471 = n4465 ^ n4279;
  assign n4475 = n4474 ^ n4471;
  assign n4479 = n3815 ^ n3505;
  assign n4480 = ~n4323 & n4479;
  assign n4481 = n4480 ^ n3505;
  assign n4476 = n4263 & n4269;
  assign n4477 = n4476 ^ n4270;
  assign n4478 = n4477 ^ n4280;
  assign n4482 = n4481 ^ n4478;
  assign n4484 = n3817 ^ n3506;
  assign n4485 = n4302 & ~n4484;
  assign n4486 = n4485 ^ n3506;
  assign n4483 = n4269 ^ n4263;
  assign n4487 = n4486 ^ n4483;
  assign n4489 = n3818 ^ n3521;
  assign n4490 = n4305 & ~n4489;
  assign n4491 = n4490 ^ n3521;
  assign n4488 = n4260 ^ n4228;
  assign n4492 = n4491 ^ n4488;
  assign n4687 = n4257 ^ n4230;
  assign n4496 = n4254 ^ n4232;
  assign n4493 = n3820 ^ n3518;
  assign n4494 = n4213 & n4493;
  assign n4495 = n4494 ^ n3518;
  assign n4497 = n4496 ^ n4495;
  assign n4676 = n4251 ^ n4234;
  assign n4500 = n3778 ^ n3515;
  assign n4501 = n4194 & ~n4500;
  assign n4502 = n4501 ^ n3515;
  assign n4498 = n4248 ^ x124;
  assign n4499 = n4498 ^ n4236;
  assign n4503 = n4502 ^ n4499;
  assign n4507 = n4245 ^ x125;
  assign n4508 = n4507 ^ n4238;
  assign n4504 = n3784 ^ n3513;
  assign n4505 = ~n4142 & ~n4504;
  assign n4506 = n4505 ^ n3513;
  assign n4509 = n4508 ^ n4506;
  assign n4513 = n4242 ^ n4241;
  assign n4510 = n3788 ^ n3508;
  assign n4511 = n3776 & n4510;
  assign n4512 = n4511 ^ n3508;
  assign n4514 = n4513 ^ n4512;
  assign n4515 = n3792 ^ n3510;
  assign n4516 = ~n3781 & n4515;
  assign n4517 = n4516 ^ n3510;
  assign n4519 = n4518 ^ n4517;
  assign n4627 = n3797 ^ n3444;
  assign n4628 = n3786 & n4627;
  assign n4629 = n4628 ^ n3444;
  assign n4529 = ~n3397 & n3709;
  assign n4530 = n4529 ^ n4528;
  assign n4532 = n3389 & ~n3738;
  assign n4531 = n4059 ^ x73;
  assign n4533 = n4532 ^ n4531;
  assign n4534 = n3381 & n3916;
  assign n4536 = n4535 ^ n4534;
  assign n4537 = n3377 & n3913;
  assign n4539 = n4538 ^ n4537;
  assign n4443 = ~n3716 & n3808;
  assign n4445 = n4444 ^ n4443;
  assign n4395 = ~n3611 & n3860;
  assign n4439 = n4397 ^ n4395;
  assign n4382 = ~n3604 & ~n3810;
  assign n4384 = n4383 ^ n4382;
  assign n4358 = ~n3598 & ~n3812;
  assign n4359 = n4358 ^ n4357;
  assign n4338 = n3593 & n3813;
  assign n4353 = n4340 ^ n4338;
  assign n4335 = n4323 ^ n4322;
  assign n4336 = ~n4325 & n4335;
  assign n4337 = n4336 ^ n4324;
  assign n4354 = n4340 ^ n4337;
  assign n4355 = n4353 & n4354;
  assign n4356 = n4355 ^ n4338;
  assign n4379 = n4357 ^ n4356;
  assign n4380 = ~n4359 & ~n4379;
  assign n4381 = n4380 ^ n4358;
  assign n4392 = n4383 ^ n4381;
  assign n4393 = ~n4384 & ~n4392;
  assign n4394 = n4393 ^ n4382;
  assign n4440 = n4397 ^ n4394;
  assign n4441 = n4439 & ~n4440;
  assign n4442 = n4441 ^ n4395;
  assign n4540 = n4444 ^ n4442;
  assign n4541 = ~n4445 & n4540;
  assign n4542 = n4541 ^ n4443;
  assign n4543 = n4542 ^ n4538;
  assign n4544 = ~n4539 & ~n4543;
  assign n4545 = n4544 ^ n4537;
  assign n4546 = n4545 ^ n4535;
  assign n4547 = ~n4536 & n4546;
  assign n4548 = n4547 ^ n4534;
  assign n4549 = n4548 ^ n4531;
  assign n4550 = n4533 & n4549;
  assign n4551 = n4550 ^ n4532;
  assign n4552 = n4551 ^ n4528;
  assign n4553 = ~n4530 & n4552;
  assign n4554 = n4553 ^ n4529;
  assign n4525 = ~n3394 & n3711;
  assign n4527 = n4526 ^ n4525;
  assign n4562 = n4554 ^ n4527;
  assign n4563 = n4551 ^ n4530;
  assign n4564 = n4548 ^ n4533;
  assign n4565 = n4545 ^ n4536;
  assign n4566 = n4542 ^ n4539;
  assign n4446 = n4445 ^ n4442;
  assign n4385 = n4384 ^ n4381;
  assign n4360 = n4359 ^ n4356;
  assign n4334 = ~n4326 & n4333;
  assign n4339 = n4338 ^ n4337;
  assign n4341 = n4340 ^ n4339;
  assign n4361 = ~n4334 & ~n4341;
  assign n4386 = ~n4360 & n4361;
  assign n4391 = n4385 & n4386;
  assign n4396 = n4395 ^ n4394;
  assign n4398 = n4397 ^ n4396;
  assign n4447 = n4391 & n4398;
  assign n4567 = ~n4446 & n4447;
  assign n4568 = ~n4566 & n4567;
  assign n4569 = ~n4565 & ~n4568;
  assign n4570 = ~n4564 & ~n4569;
  assign n4571 = ~n4563 & n4570;
  assign n4585 = ~n4562 & n4571;
  assign n4555 = n4554 ^ n4525;
  assign n4556 = n4527 & ~n4555;
  assign n4557 = n4556 ^ n4554;
  assign n4522 = x31 & ~n3708;
  assign n4524 = n4523 ^ n4522;
  assign n4583 = n4557 ^ n4524;
  assign n4591 = n4585 ^ n4583;
  assign n4572 = n4571 ^ n4562;
  assign n4573 = n4569 ^ n4564;
  assign n4399 = n4398 ^ n4391;
  assign n4387 = n4386 ^ n4385;
  assign n4342 = n4341 ^ n4334;
  assign n4351 = n4349 & ~n4350;
  assign n4352 = ~n4342 & n4351;
  assign n4362 = n4361 ^ n4360;
  assign n4388 = n4352 & n4362;
  assign n4400 = ~n4387 & n4388;
  assign n4438 = n4399 & ~n4400;
  assign n4448 = n4447 ^ n4446;
  assign n4574 = ~n4438 & n4448;
  assign n4575 = n4567 ^ n4566;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = n4568 ^ n4565;
  assign n4578 = ~n4576 & n4577;
  assign n4579 = n4573 & ~n4578;
  assign n4580 = n4570 ^ n4563;
  assign n4581 = n4579 & ~n4580;
  assign n4582 = n4572 & ~n4581;
  assign n4592 = n4591 ^ n4582;
  assign n4593 = n4592 ^ x97;
  assign n4594 = n4581 ^ n4572;
  assign n4595 = n4594 ^ x98;
  assign n4596 = n4580 ^ n4579;
  assign n4597 = n4596 ^ x99;
  assign n4599 = n4577 ^ n4576;
  assign n4600 = n4599 ^ x101;
  assign n4601 = n4575 ^ n4574;
  assign n4602 = n4601 ^ x102;
  assign n4449 = n4448 ^ n4438;
  assign n4603 = n4449 ^ x103;
  assign n4363 = n4362 ^ n4352;
  assign n4364 = ~x106 & ~n4363;
  assign n4365 = n4351 ^ n4342;
  assign n4366 = ~x107 & n4365;
  assign n4367 = ~n4364 & ~n4366;
  assign n4369 = ~x109 & ~n4368;
  assign n4376 = ~x108 & n4375;
  assign n4377 = n4374 & ~n4376;
  assign n4378 = ~n4369 & n4377;
  assign n4389 = n4388 ^ n4387;
  assign n4390 = ~x105 & n4389;
  assign n4401 = n4400 ^ n4399;
  assign n4402 = ~x104 & ~n4401;
  assign n4403 = ~n4390 & ~n4402;
  assign n4404 = n4378 & n4403;
  assign n4405 = n4367 & n4404;
  assign n4406 = n4301 & n4405;
  assign n4407 = n4401 ^ x104;
  assign n4408 = n4363 ^ x106;
  assign n4409 = n4365 ^ x107;
  assign n4410 = n4409 ^ n4366;
  assign n4411 = n4408 & ~n4410;
  assign n4412 = n4411 ^ n4364;
  assign n4420 = n4418 & n4419;
  assign n4421 = n4420 ^ n4369;
  assign n4422 = n4421 ^ n4375;
  assign n4423 = ~n4413 & ~n4422;
  assign n4424 = n4423 ^ x108;
  assign n4425 = n4367 & n4424;
  assign n4426 = n4389 ^ x105;
  assign n4427 = n4426 ^ n4390;
  assign n4428 = ~n4425 & ~n4427;
  assign n4429 = n4412 & n4428;
  assign n4430 = n4429 ^ n4401;
  assign n4431 = n4430 ^ n4401;
  assign n4432 = ~n4390 & ~n4431;
  assign n4433 = n4432 ^ n4401;
  assign n4434 = n4407 & ~n4433;
  assign n4435 = n4434 ^ x104;
  assign n4436 = ~n4406 & ~n4435;
  assign n4604 = n4449 ^ n4436;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = n4605 ^ x103;
  assign n4607 = n4606 ^ n4601;
  assign n4608 = ~n4602 & n4607;
  assign n4609 = n4608 ^ x102;
  assign n4610 = n4609 ^ n4599;
  assign n4611 = ~n4600 & n4610;
  assign n4612 = n4611 ^ x101;
  assign n4598 = n4578 ^ n4573;
  assign n4613 = n4612 ^ n4598;
  assign n4614 = n4598 ^ x100;
  assign n4615 = ~n4613 & n4614;
  assign n4616 = n4615 ^ x100;
  assign n4617 = n4616 ^ n4596;
  assign n4618 = n4597 & ~n4617;
  assign n4619 = n4618 ^ x99;
  assign n4620 = n4619 ^ n4594;
  assign n4621 = ~n4595 & n4620;
  assign n4622 = n4621 ^ x98;
  assign n4623 = n4622 ^ n4592;
  assign n4624 = n4593 & ~n4623;
  assign n4625 = n4624 ^ x97;
  assign n4584 = n4583 ^ n4582;
  assign n4586 = n4585 ^ n4582;
  assign n4587 = ~n4584 & n4586;
  assign n4588 = n4587 ^ n4583;
  assign n4589 = n4588 ^ x96;
  assign n4558 = n4557 ^ n4523;
  assign n4559 = n4524 & ~n4558;
  assign n4560 = n4559 ^ n4522;
  assign n4520 = ~n3406 & n3722;
  assign n4451 = n4074 ^ x69;
  assign n4521 = n4520 ^ n4451;
  assign n4561 = n4560 ^ n4521;
  assign n4590 = n4589 ^ n4561;
  assign n4626 = n4625 ^ n4590;
  assign n4630 = n4629 ^ n4626;
  assign n4632 = n3802 ^ n3424;
  assign n4633 = n3790 & n4632;
  assign n4634 = n4633 ^ n3424;
  assign n4631 = n4622 ^ n4593;
  assign n4635 = n4634 ^ n4631;
  assign n4641 = n3826 ^ n3416;
  assign n4642 = n3799 & n4641;
  assign n4643 = n4642 ^ n3416;
  assign n4639 = n4616 ^ x99;
  assign n4640 = n4639 ^ n4596;
  assign n4644 = n4643 ^ n4640;
  assign n4645 = n4613 ^ x100;
  assign n4646 = n3413 ^ n3391;
  assign n4647 = n3804 & ~n4646;
  assign n4648 = n4647 ^ n3413;
  assign n4649 = n4645 & ~n4648;
  assign n4650 = n4649 ^ n4640;
  assign n4651 = ~n4644 & n4650;
  assign n4652 = n4651 ^ n4649;
  assign n4636 = n3806 ^ n3421;
  assign n4637 = ~n3794 & ~n4636;
  assign n4638 = n4637 ^ n3421;
  assign n4653 = n4652 ^ n4638;
  assign n4654 = n4619 ^ n4595;
  assign n4655 = n4654 ^ n4652;
  assign n4656 = ~n4653 & n4655;
  assign n4657 = n4656 ^ n4638;
  assign n4658 = n4657 ^ n4634;
  assign n4659 = n4635 & n4658;
  assign n4660 = n4659 ^ n4631;
  assign n4661 = n4660 ^ n4629;
  assign n4662 = n4630 & ~n4661;
  assign n4663 = n4662 ^ n4660;
  assign n4664 = n4663 ^ n4517;
  assign n4665 = n4519 & n4664;
  assign n4666 = n4665 ^ n4518;
  assign n4667 = n4666 ^ n4512;
  assign n4668 = n4514 & ~n4667;
  assign n4669 = n4668 ^ n4513;
  assign n4670 = n4669 ^ n4508;
  assign n4671 = ~n4509 & ~n4670;
  assign n4672 = n4671 ^ n4506;
  assign n4673 = n4672 ^ n4499;
  assign n4674 = ~n4503 & n4673;
  assign n4675 = n4674 ^ n4502;
  assign n4677 = n4676 ^ n4675;
  assign n4678 = n3507 ^ n3495;
  assign n4679 = n4204 & n4678;
  assign n4680 = n4679 ^ n3507;
  assign n4681 = n4680 ^ n4676;
  assign n4682 = n4677 & n4681;
  assign n4683 = n4682 ^ n4680;
  assign n4684 = n4683 ^ n4496;
  assign n4685 = n4497 & n4684;
  assign n4686 = n4685 ^ n4495;
  assign n4688 = n4687 ^ n4686;
  assign n4689 = n3819 ^ n3496;
  assign n4690 = ~n4309 & ~n4689;
  assign n4691 = n4690 ^ n3496;
  assign n4692 = n4691 ^ n4687;
  assign n4693 = n4688 & n4692;
  assign n4694 = n4693 ^ n4691;
  assign n4695 = n4694 ^ n4488;
  assign n4696 = n4492 & n4695;
  assign n4697 = n4696 ^ n4491;
  assign n4698 = n4697 ^ n4483;
  assign n4699 = ~n4487 & ~n4698;
  assign n4700 = n4699 ^ n4486;
  assign n4701 = n4700 ^ n4478;
  assign n4702 = ~n4482 & n4701;
  assign n4703 = n4702 ^ n4481;
  assign n4704 = n4703 ^ n4471;
  assign n4705 = ~n4475 & ~n4704;
  assign n4706 = n4705 ^ n4474;
  assign n4707 = n4706 ^ n4469;
  assign n4708 = n4470 & n4707;
  assign n4709 = n4708 ^ n4463;
  assign n4710 = n4709 ^ n4456;
  assign n4711 = ~n4460 & n4710;
  assign n4712 = n4711 ^ n4459;
  assign n4888 = n4713 ^ n4712;
  assign n4889 = n4717 & ~n4888;
  assign n4890 = n4889 ^ n4716;
  assign n5008 = n4891 ^ n4890;
  assign n5009 = ~n4895 & ~n5008;
  assign n5010 = n5009 ^ n4894;
  assign n5011 = n5010 ^ n4901;
  assign n5012 = ~n5007 & ~n5011;
  assign n5013 = n5012 ^ n5006;
  assign n5014 = n5013 ^ n5002;
  assign n5015 = n5003 & ~n5014;
  assign n5016 = n5015 ^ n4999;
  assign n4994 = n4372 ^ n4301;
  assign n4995 = ~n4415 & n4994;
  assign n4996 = n4995 ^ x111;
  assign n4997 = n4996 ^ x110;
  assign n4998 = n4997 ^ n4370;
  assign n5017 = n5016 ^ n4998;
  assign n5018 = n3808 ^ n3604;
  assign n5019 = ~n4531 & n5018;
  assign n5020 = n5019 ^ n3604;
  assign n5021 = n5020 ^ n4998;
  assign n5022 = n5017 & n5021;
  assign n5023 = n5022 ^ n5020;
  assign n5024 = n5023 ^ n4992;
  assign n5025 = ~n4993 & ~n5024;
  assign n5026 = n5025 ^ n4989;
  assign n5027 = n5026 ^ n4987;
  assign n5028 = ~n4988 & ~n5027;
  assign n5029 = n5028 ^ n4981;
  assign n4965 = n4301 & n4378;
  assign n4966 = ~n4424 & ~n4965;
  assign n4978 = n4966 ^ n4409;
  assign n5030 = n5029 ^ n4978;
  assign n5054 = n5033 ^ n5030;
  assign n5044 = n5026 ^ n4981;
  assign n5045 = n5044 ^ n4987;
  assign n5046 = n5020 ^ n5017;
  assign n5047 = n5010 ^ n5007;
  assign n5048 = n5013 ^ n5003;
  assign n5049 = ~n5047 & ~n5048;
  assign n5050 = n5046 & ~n5049;
  assign n5051 = n5023 ^ n4993;
  assign n5052 = n5050 & n5051;
  assign n5053 = ~n5045 & n5052;
  assign n5071 = n5054 ^ n5053;
  assign n5072 = n5052 ^ n5045;
  assign n5073 = n5049 ^ n5046;
  assign n4718 = n4717 ^ n4712;
  assign n4719 = n4706 ^ n4463;
  assign n4720 = n4719 ^ n4469;
  assign n4740 = n4703 ^ n4475;
  assign n4721 = n4691 ^ n4688;
  assign n4722 = n4680 ^ n4677;
  assign n4723 = n4669 ^ n4509;
  assign n4724 = n4666 ^ n4514;
  assign n4725 = n4724 ^ n4723;
  assign n4726 = n4723 & ~n4725;
  assign n4727 = n4726 ^ n4724;
  assign n4728 = n4672 ^ n4503;
  assign n4729 = ~n4727 & ~n4728;
  assign n4730 = n4722 & n4729;
  assign n4731 = n4683 ^ n4497;
  assign n4732 = n4730 & ~n4731;
  assign n4733 = ~n4721 & ~n4732;
  assign n4734 = n4694 ^ n4492;
  assign n4735 = ~n4733 & ~n4734;
  assign n4736 = n4697 ^ n4487;
  assign n4737 = n4735 & ~n4736;
  assign n4738 = n4700 ^ n4482;
  assign n4739 = ~n4737 & ~n4738;
  assign n4741 = n4740 ^ n4739;
  assign n4742 = n4738 ^ n4737;
  assign n4743 = n4736 ^ n4735;
  assign n4744 = n4732 ^ n4721;
  assign n4745 = n4731 ^ n4730;
  assign n4746 = n4728 ^ n4727;
  assign n4747 = n4663 ^ n4519;
  assign n4748 = n4660 ^ n4630;
  assign n4749 = n4648 ^ n4645;
  assign n4750 = n4649 ^ n4643;
  assign n4751 = n4750 ^ n4640;
  assign n4752 = ~n4749 & n4751;
  assign n4753 = n4654 ^ n4653;
  assign n4754 = n4752 & n4753;
  assign n4755 = n4657 ^ n4635;
  assign n4756 = ~n4754 & n4755;
  assign n4757 = n4748 & n4756;
  assign n4758 = n4747 & ~n4757;
  assign n4759 = n4726 & n4758;
  assign n4760 = n4759 ^ n4725;
  assign n4761 = ~n4746 & ~n4760;
  assign n4762 = n4729 ^ n4722;
  assign n4763 = ~n4761 & n4762;
  assign n4764 = ~n4745 & n4763;
  assign n4765 = n4744 & ~n4764;
  assign n4766 = n4734 ^ n4733;
  assign n4767 = n4765 & ~n4766;
  assign n4768 = n4743 & n4767;
  assign n4769 = n4742 & n4768;
  assign n4770 = n4769 ^ n4739;
  assign n4771 = ~n4741 & n4770;
  assign n4772 = n4771 ^ n4739;
  assign n4773 = ~n4720 & n4772;
  assign n4774 = n4709 ^ n4460;
  assign n4775 = n4773 & ~n4774;
  assign n4887 = ~n4718 & ~n4775;
  assign n4896 = n4895 ^ n4890;
  assign n5074 = n4887 & n4896;
  assign n5075 = n5047 & n5074;
  assign n5076 = n5048 ^ n5047;
  assign n5077 = n5075 & n5076;
  assign n5078 = n5073 & n5077;
  assign n5079 = n5051 ^ n5050;
  assign n5080 = ~n5078 & n5079;
  assign n5081 = n5072 & ~n5080;
  assign n5082 = n5071 & ~n5081;
  assign n5055 = ~n5053 & n5054;
  assign n5034 = n5033 ^ n4978;
  assign n5035 = ~n5030 & n5034;
  assign n5036 = n5035 ^ n5033;
  assign n4974 = n3709 ^ n3381;
  assign n4975 = ~n4451 & n4974;
  assign n4976 = n4975 ^ n3381;
  assign n5042 = n5036 ^ n4976;
  assign n4970 = n4966 ^ n4365;
  assign n4971 = ~n4409 & ~n4970;
  assign n4972 = n4971 ^ x107;
  assign n4973 = n4972 ^ n4408;
  assign n5043 = n5042 ^ n4973;
  assign n5070 = n5055 ^ n5043;
  assign n5117 = n5082 ^ n5070;
  assign n5118 = n5117 ^ x133;
  assign n5119 = n5079 ^ n5078;
  assign n5120 = n5119 ^ x136;
  assign n4897 = n4896 ^ n4887;
  assign n5128 = ~x140 & ~n4897;
  assign n4898 = n4897 ^ x140;
  assign n4776 = n4775 ^ n4718;
  assign n4777 = n4776 ^ x141;
  assign n4778 = n4774 ^ n4773;
  assign n4779 = n4778 ^ x142;
  assign n4780 = n4739 ^ n4720;
  assign n4781 = n4780 ^ n4771;
  assign n4783 = n4781 ^ x143;
  assign n4782 = ~x143 & ~n4781;
  assign n4784 = n4783 ^ n4782;
  assign n4785 = n4784 ^ n4778;
  assign n4786 = n4779 & n4785;
  assign n4787 = n4786 ^ x142;
  assign n5123 = n4787 ^ n4776;
  assign n5124 = n4777 & ~n5123;
  assign n5125 = n5124 ^ x141;
  assign n5126 = n4898 & n5125;
  assign n5127 = n5126 ^ n4898;
  assign n5129 = n5128 ^ n5127;
  assign n5130 = n5074 ^ n5047;
  assign n5131 = ~x139 & ~n5130;
  assign n5132 = n5076 ^ n5075;
  assign n5133 = ~x138 & ~n5132;
  assign n5134 = ~n5131 & ~n5133;
  assign n5135 = ~n5129 & n5134;
  assign n5121 = n5077 ^ n5073;
  assign n5136 = n5121 ^ x137;
  assign n5137 = n5132 ^ x138;
  assign n5138 = n5130 ^ x139;
  assign n5139 = n5138 ^ n5131;
  assign n5140 = n5137 & n5139;
  assign n5141 = n5140 ^ n5133;
  assign n5142 = n5136 & n5141;
  assign n5143 = ~n5135 & n5142;
  assign n5122 = ~x137 & ~n5121;
  assign n5144 = n5143 ^ n5122;
  assign n5145 = n5144 ^ n5119;
  assign n5146 = n5120 & n5145;
  assign n5147 = n5146 ^ x136;
  assign n5148 = n5081 ^ n5071;
  assign n5149 = ~x134 & ~n5148;
  assign n5150 = n5080 ^ n5072;
  assign n5152 = x135 & ~n5150;
  assign n5151 = n5150 ^ x135;
  assign n5153 = n5152 ^ n5151;
  assign n5154 = ~n5149 & ~n5153;
  assign n5155 = n5147 & n5154;
  assign n5156 = n5155 ^ n5117;
  assign n5157 = n5156 ^ n5117;
  assign n5158 = n5148 ^ x134;
  assign n5159 = ~n5152 & n5158;
  assign n5160 = n5159 ^ n5149;
  assign n5161 = ~n5157 & n5160;
  assign n5162 = n5161 ^ n5117;
  assign n5163 = ~n5118 & ~n5162;
  assign n5164 = n5163 ^ x133;
  assign n4788 = n4724 & n4758;
  assign n4789 = n4788 ^ n4725;
  assign n4790 = n4789 ^ x152;
  assign n4791 = n4758 ^ n4724;
  assign n4792 = n4791 ^ x153;
  assign n4793 = n4757 ^ n4747;
  assign n4794 = n4793 ^ x154;
  assign n4795 = n4756 ^ n4748;
  assign n4796 = n4795 ^ x155;
  assign n4797 = n4755 ^ n4754;
  assign n4798 = n4797 ^ x156;
  assign n4799 = n4753 ^ n4752;
  assign n4800 = n4799 ^ x157;
  assign n4801 = x159 & n4749;
  assign n4802 = n4801 ^ x158;
  assign n4803 = n4751 ^ n4749;
  assign n4804 = n4803 ^ n4801;
  assign n4805 = n4802 & n4804;
  assign n4806 = n4805 ^ x158;
  assign n4807 = n4806 ^ n4799;
  assign n4808 = n4800 & ~n4807;
  assign n4809 = n4808 ^ x157;
  assign n4810 = n4809 ^ n4797;
  assign n4811 = n4798 & ~n4810;
  assign n4812 = n4811 ^ x156;
  assign n4813 = n4812 ^ n4795;
  assign n4814 = ~n4796 & n4813;
  assign n4815 = n4814 ^ x155;
  assign n4816 = n4815 ^ n4793;
  assign n4817 = ~n4794 & n4816;
  assign n4818 = n4817 ^ x154;
  assign n4819 = n4818 ^ n4791;
  assign n4820 = n4792 & ~n4819;
  assign n4821 = n4820 ^ x153;
  assign n4822 = n4821 ^ n4789;
  assign n4823 = ~n4790 & n4822;
  assign n4824 = n4823 ^ x152;
  assign n4825 = n4767 ^ n4743;
  assign n4826 = ~x146 & n4825;
  assign n4827 = n4766 ^ n4765;
  assign n4829 = n4827 ^ x147;
  assign n4828 = x147 & n4827;
  assign n4830 = n4829 ^ n4828;
  assign n4831 = ~n4826 & n4830;
  assign n4832 = n4763 ^ n4745;
  assign n4833 = ~x149 & n4832;
  assign n4834 = n4764 ^ n4744;
  assign n4835 = ~x148 & ~n4834;
  assign n4836 = n4762 ^ n4761;
  assign n4837 = ~x150 & n4836;
  assign n4838 = n4760 ^ n4746;
  assign n4840 = n4838 ^ x151;
  assign n4839 = x151 & ~n4838;
  assign n4841 = n4840 ^ n4839;
  assign n4842 = ~n4837 & ~n4841;
  assign n4843 = ~n4835 & n4842;
  assign n4844 = ~n4833 & n4843;
  assign n4845 = n4769 ^ n4741;
  assign n4846 = ~x144 & ~n4845;
  assign n4847 = n4768 ^ n4742;
  assign n4849 = x145 & ~n4847;
  assign n4848 = n4847 ^ x145;
  assign n4850 = n4849 ^ n4848;
  assign n4851 = ~n4846 & ~n4850;
  assign n4852 = n4844 & n4851;
  assign n4853 = n4831 & n4852;
  assign n4854 = n4824 & n4853;
  assign n4855 = n4845 ^ x144;
  assign n4856 = n4825 ^ x146;
  assign n4857 = ~n4828 & ~n4856;
  assign n4858 = n4857 ^ n4826;
  assign n4859 = n4834 ^ x148;
  assign n4860 = n4832 ^ x149;
  assign n4861 = n4836 ^ x150;
  assign n4862 = ~n4839 & ~n4861;
  assign n4863 = n4862 ^ n4837;
  assign n4864 = n4863 ^ n4832;
  assign n4865 = ~n4860 & ~n4864;
  assign n4866 = n4865 ^ x149;
  assign n4867 = n4859 & n4866;
  assign n4868 = n4867 ^ n4859;
  assign n4869 = n4868 ^ n4835;
  assign n4870 = n4831 & ~n4869;
  assign n4871 = ~n4849 & ~n4870;
  assign n4872 = n4858 & n4871;
  assign n4873 = n4872 ^ n4845;
  assign n4874 = n4873 ^ n4845;
  assign n4875 = ~n4850 & ~n4874;
  assign n4876 = n4875 ^ n4845;
  assign n4877 = n4855 & ~n4876;
  assign n4878 = n4877 ^ x144;
  assign n4879 = ~n4854 & ~n4878;
  assign n5165 = ~x141 & ~n4776;
  assign n4880 = ~x142 & ~n4778;
  assign n4881 = ~n4782 & ~n4880;
  assign n5166 = n4881 & ~n5128;
  assign n5167 = ~n5165 & n5166;
  assign n5168 = ~x136 & ~n5119;
  assign n5169 = ~n5122 & ~n5168;
  assign n5170 = n5167 & n5169;
  assign n5171 = n5134 & n5170;
  assign n5172 = ~x133 & n5117;
  assign n5173 = n5171 & ~n5172;
  assign n5174 = n5154 & n5173;
  assign n5175 = ~n4879 & n5174;
  assign n5176 = ~n5164 & ~n5175;
  assign n5056 = n5043 & n5055;
  assign n4977 = n4976 ^ n4973;
  assign n5037 = n5036 ^ n4973;
  assign n5038 = n4977 & ~n5037;
  assign n5039 = n5038 ^ n4976;
  assign n4967 = n4367 & ~n4966;
  assign n4968 = n4412 & ~n4967;
  assign n4969 = n4968 ^ n4426;
  assign n5040 = n5039 ^ n4969;
  assign n4962 = n3711 ^ n3389;
  assign n4963 = n4102 & ~n4962;
  assign n4964 = n4963 ^ n3389;
  assign n5041 = n5040 ^ n4964;
  assign n5084 = n5056 ^ n5041;
  assign n5083 = n5070 & ~n5082;
  assign n5115 = n5084 ^ n5083;
  assign n5116 = n5115 ^ x132;
  assign n5223 = n5176 ^ n5116;
  assign n5412 = n5226 ^ n5223;
  assign n5587 = n5412 ^ n3413;
  assign n6053 = n5587 ^ x191;
  assign n4950 = n4806 ^ n4800;
  assign n6688 = n4950 ^ n4508;
  assign n6689 = n6053 & ~n6688;
  assign n6690 = n6689 ^ n4508;
  assign n5871 = ~n4879 & n5171;
  assign n5872 = ~n5147 & ~n5871;
  assign n5913 = n5872 ^ n5150;
  assign n5914 = ~n5151 & ~n5913;
  assign n5915 = n5914 ^ x135;
  assign n5916 = n5915 ^ n5158;
  assign n6375 = n4645 ^ n4102;
  assign n6376 = n5916 & n6375;
  assign n6377 = n6376 ^ n4102;
  assign n4905 = n4824 & n4842;
  assign n4906 = n4863 & ~n4905;
  assign n5288 = n4906 ^ n4832;
  assign n5289 = ~n4860 & ~n5288;
  assign n5290 = n5289 ^ x149;
  assign n5291 = n5290 ^ n4859;
  assign n5292 = n4397 ^ n3851;
  assign n5293 = ~n4999 & ~n5292;
  assign n5294 = n5293 ^ n3851;
  assign n5295 = n5291 & n5294;
  assign n4907 = n4906 ^ n4860;
  assign n4902 = n4383 ^ n3849;
  assign n4903 = n4901 & n4902;
  assign n4904 = n4903 ^ n3849;
  assign n4908 = n4907 ^ n4904;
  assign n4912 = n4838 ^ n4824;
  assign n4913 = ~n4840 & n4912;
  assign n4914 = n4913 ^ x151;
  assign n4915 = n4914 ^ n4861;
  assign n4909 = n4357 ^ n3815;
  assign n4910 = ~n4891 & n4909;
  assign n4911 = n4910 ^ n3815;
  assign n4916 = n4915 ^ n4911;
  assign n4920 = n4840 ^ n4824;
  assign n4917 = n4340 ^ n3817;
  assign n4918 = ~n4713 & ~n4917;
  assign n4919 = n4918 ^ n3817;
  assign n4921 = n4920 ^ n4919;
  assign n4925 = n4821 ^ n4790;
  assign n4922 = n4323 ^ n3818;
  assign n4923 = n4456 & n4922;
  assign n4924 = n4923 ^ n3818;
  assign n4926 = n4925 ^ n4924;
  assign n4930 = n4818 ^ n4792;
  assign n4927 = n4302 ^ n3819;
  assign n4928 = ~n4469 & n4927;
  assign n4929 = n4928 ^ n3819;
  assign n4931 = n4930 ^ n4929;
  assign n4935 = n4815 ^ n4794;
  assign n4932 = n4305 ^ n3820;
  assign n4933 = ~n4471 & n4932;
  assign n4934 = n4933 ^ n3820;
  assign n4936 = n4935 ^ n4934;
  assign n4940 = n4812 ^ n4796;
  assign n4937 = n4309 ^ n3495;
  assign n4938 = n4478 & n4937;
  assign n4939 = n4938 ^ n3495;
  assign n4941 = n4940 ^ n4939;
  assign n4943 = n4213 ^ n3778;
  assign n4944 = n4483 & ~n4943;
  assign n4945 = n4944 ^ n3778;
  assign n4942 = n4809 ^ n4798;
  assign n4946 = n4945 ^ n4942;
  assign n4947 = n4204 ^ n3784;
  assign n4948 = n4488 & ~n4947;
  assign n4949 = n4948 ^ n3784;
  assign n4951 = n4950 ^ n4949;
  assign n4955 = n4803 ^ n4802;
  assign n4952 = n4194 ^ n3788;
  assign n4953 = ~n4687 & ~n4952;
  assign n4954 = n4953 ^ n3788;
  assign n4956 = n4955 ^ n4954;
  assign n4960 = n4749 ^ x159;
  assign n4957 = n4142 ^ n3792;
  assign n4958 = n4496 & n4957;
  assign n4959 = n4958 ^ n3792;
  assign n4961 = n4960 ^ n4959;
  assign n5204 = n3797 ^ n3776;
  assign n5205 = ~n4676 & ~n5204;
  assign n5206 = n5205 ^ n3797;
  assign n5104 = n3499 ^ x31;
  assign n5105 = n4096 & n5104;
  assign n5106 = n5105 ^ x31;
  assign n5090 = n3722 ^ n3394;
  assign n5091 = ~n4098 & ~n5090;
  assign n5092 = n5091 ^ n3394;
  assign n4437 = n4436 ^ x103;
  assign n4450 = n4449 ^ n4437;
  assign n5093 = n5092 ^ n4450;
  assign n5061 = ~n4426 & ~n4968;
  assign n5062 = n5061 ^ n4427;
  assign n5063 = n5062 ^ n4407;
  assign n5058 = n4969 ^ n4964;
  assign n5059 = ~n5040 & ~n5058;
  assign n5060 = n5059 ^ n4964;
  assign n5064 = n5063 ^ n5060;
  assign n5065 = n3708 ^ n3397;
  assign n5066 = n4107 & ~n5065;
  assign n5067 = n5066 ^ n3397;
  assign n5087 = n5067 ^ n5063;
  assign n5088 = n5064 & n5087;
  assign n5089 = n5088 ^ n5067;
  assign n5100 = n5089 ^ n4450;
  assign n5101 = ~n5093 & ~n5100;
  assign n5102 = n5101 ^ n5092;
  assign n5099 = n4606 ^ n4602;
  assign n5103 = n5102 ^ n5099;
  assign n5107 = n5106 ^ n5103;
  assign n5094 = n5093 ^ n5089;
  assign n5057 = n5041 & ~n5056;
  assign n5068 = n5067 ^ n5064;
  assign n5095 = n5057 & n5068;
  assign n5098 = ~n5094 & ~n5095;
  assign n5108 = n5107 ^ n5098;
  assign n5069 = n5068 ^ n5057;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = n5069 & n5085;
  assign n5096 = n5095 ^ n5094;
  assign n5097 = ~n5086 & n5096;
  assign n5198 = n5098 ^ n5097;
  assign n5199 = n5108 & n5198;
  assign n5200 = n5199 ^ n5097;
  assign n5193 = n3498 ^ n3406;
  assign n5194 = ~n4093 & ~n5193;
  assign n5195 = n5194 ^ n3406;
  assign n5192 = n4609 ^ n4600;
  assign n5196 = n5195 ^ n5192;
  assign n5189 = n5106 ^ n5099;
  assign n5190 = ~n5103 & n5189;
  assign n5191 = n5190 ^ n5106;
  assign n5197 = n5196 ^ n5191;
  assign n5201 = n5200 ^ n5197;
  assign n5202 = n5201 ^ x128;
  assign n5109 = n5108 ^ n5097;
  assign n5110 = n5109 ^ x129;
  assign n5111 = n5096 ^ n5086;
  assign n5112 = n5111 ^ x130;
  assign n5113 = n5085 ^ n5069;
  assign n5114 = n5113 ^ x131;
  assign n5177 = n5176 ^ n5115;
  assign n5178 = ~n5116 & ~n5177;
  assign n5179 = n5178 ^ x132;
  assign n5180 = n5179 ^ n5113;
  assign n5181 = ~n5114 & n5180;
  assign n5182 = n5181 ^ x131;
  assign n5183 = n5182 ^ n5111;
  assign n5184 = ~n5112 & n5183;
  assign n5185 = n5184 ^ x130;
  assign n5186 = n5185 ^ n5109;
  assign n5187 = ~n5110 & n5186;
  assign n5188 = n5187 ^ x129;
  assign n5203 = n5202 ^ n5188;
  assign n5207 = n5206 ^ n5203;
  assign n5211 = n5185 ^ n5110;
  assign n5208 = n3802 ^ n3781;
  assign n5209 = ~n4499 & ~n5208;
  assign n5210 = n5209 ^ n3802;
  assign n5212 = n5211 ^ n5210;
  assign n5216 = n5182 ^ n5112;
  assign n5213 = n3806 ^ n3786;
  assign n5214 = ~n4508 & n5213;
  assign n5215 = n5214 ^ n3806;
  assign n5217 = n5216 ^ n5215;
  assign n5219 = n3826 ^ n3790;
  assign n5220 = ~n4513 & n5219;
  assign n5221 = n5220 ^ n3826;
  assign n5218 = n5179 ^ n5114;
  assign n5222 = n5221 ^ n5218;
  assign n5227 = n5223 & n5226;
  assign n5228 = n5227 ^ n5218;
  assign n5229 = n5222 & ~n5228;
  assign n5230 = n5229 ^ n5227;
  assign n5231 = n5230 ^ n5215;
  assign n5232 = n5217 & n5231;
  assign n5233 = n5232 ^ n5230;
  assign n5234 = n5233 ^ n5211;
  assign n5235 = ~n5212 & n5234;
  assign n5236 = n5235 ^ n5210;
  assign n5237 = n5236 ^ n5206;
  assign n5238 = ~n5207 & n5237;
  assign n5239 = n5238 ^ n5203;
  assign n5240 = n5239 ^ n4960;
  assign n5241 = ~n4961 & ~n5240;
  assign n5242 = n5241 ^ n4959;
  assign n5243 = n5242 ^ n4955;
  assign n5244 = n4956 & ~n5243;
  assign n5245 = n5244 ^ n4954;
  assign n5246 = n5245 ^ n4950;
  assign n5247 = ~n4951 & n5246;
  assign n5248 = n5247 ^ n4949;
  assign n5249 = n5248 ^ n4942;
  assign n5250 = ~n4946 & n5249;
  assign n5251 = n5250 ^ n4945;
  assign n5252 = n5251 ^ n4939;
  assign n5253 = n4941 & ~n5252;
  assign n5254 = n5253 ^ n4940;
  assign n5255 = n5254 ^ n4935;
  assign n5256 = ~n4936 & ~n5255;
  assign n5257 = n5256 ^ n4934;
  assign n5258 = n5257 ^ n4930;
  assign n5259 = n4931 & ~n5258;
  assign n5260 = n5259 ^ n4929;
  assign n5261 = n5260 ^ n4925;
  assign n5262 = n4926 & n5261;
  assign n5263 = n5262 ^ n4924;
  assign n5264 = n5263 ^ n4920;
  assign n5265 = ~n4921 & ~n5264;
  assign n5266 = n5265 ^ n4919;
  assign n5267 = n5266 ^ n4915;
  assign n5268 = n4916 & n5267;
  assign n5269 = n5268 ^ n4911;
  assign n5270 = n5269 ^ n4907;
  assign n5271 = n4908 & n5270;
  assign n5272 = n5271 ^ n4904;
  assign n5296 = n5294 ^ n5291;
  assign n5297 = n5296 ^ n5295;
  assign n5464 = n5272 & n5297;
  assign n5469 = ~n5295 & ~n5464;
  assign n5284 = n4444 ^ n3853;
  assign n5285 = n4998 & ~n5284;
  assign n5286 = n5285 ^ n3853;
  assign n5273 = n4824 & n4844;
  assign n5274 = n4869 & ~n5273;
  assign n5283 = n5274 ^ n4829;
  assign n5342 = n5286 ^ n5283;
  assign n5470 = n5469 ^ n5342;
  assign n5510 = n5470 ^ n3502;
  assign n5472 = n5296 ^ n5272;
  assign n5473 = ~n3503 & n5472;
  assign n5511 = n5473 ^ n5470;
  assign n5512 = n5510 & n5511;
  assign n5513 = n5512 ^ n3502;
  assign n5471 = n3502 & n5470;
  assign n5386 = n5269 ^ n4908;
  assign n5387 = n5386 ^ n3504;
  assign n5388 = n5266 ^ n4916;
  assign n5389 = n5388 ^ n3505;
  assign n5390 = n5263 ^ n4921;
  assign n5391 = n5390 ^ n3506;
  assign n5392 = n5260 ^ n4926;
  assign n5393 = n5392 ^ n3521;
  assign n5394 = n5257 ^ n4931;
  assign n5395 = n5394 ^ n3496;
  assign n5396 = n5254 ^ n4936;
  assign n5397 = n5396 ^ n3518;
  assign n5398 = n5251 ^ n4941;
  assign n5399 = n5398 ^ n3507;
  assign n5400 = n5245 ^ n4951;
  assign n5401 = n5400 ^ n3513;
  assign n5402 = n5242 ^ n4956;
  assign n5403 = n5402 ^ n3508;
  assign n5404 = n5239 ^ n4961;
  assign n5405 = n5404 ^ n3510;
  assign n5406 = n5236 ^ n5207;
  assign n5407 = n5406 ^ n3444;
  assign n5408 = n5233 ^ n5212;
  assign n5409 = n5408 ^ n3424;
  assign n5410 = n5230 ^ n5217;
  assign n5411 = n5410 ^ n3421;
  assign n5413 = ~n3413 & n5412;
  assign n5414 = n5413 ^ n3416;
  assign n5415 = n5227 ^ n5221;
  assign n5416 = n5415 ^ n5218;
  assign n5417 = n5416 ^ n5413;
  assign n5418 = n5414 & n5417;
  assign n5419 = n5418 ^ n3416;
  assign n5420 = n5419 ^ n5410;
  assign n5421 = n5411 & n5420;
  assign n5422 = n5421 ^ n3421;
  assign n5423 = n5422 ^ n5408;
  assign n5424 = ~n5409 & ~n5423;
  assign n5425 = n5424 ^ n3424;
  assign n5426 = n5425 ^ n5406;
  assign n5427 = n5407 & n5426;
  assign n5428 = n5427 ^ n3444;
  assign n5429 = n5428 ^ n5404;
  assign n5430 = n5405 & ~n5429;
  assign n5431 = n5430 ^ n3510;
  assign n5432 = n5431 ^ n5402;
  assign n5433 = n5403 & ~n5432;
  assign n5434 = n5433 ^ n3508;
  assign n5435 = n5434 ^ n5400;
  assign n5436 = n5401 & n5435;
  assign n5437 = n5436 ^ n3513;
  assign n5438 = n5437 ^ n3515;
  assign n5439 = n5248 ^ n4946;
  assign n5440 = n5439 ^ n5437;
  assign n5441 = n5438 & ~n5440;
  assign n5442 = n5441 ^ n3515;
  assign n5443 = n5442 ^ n5398;
  assign n5444 = n5399 & n5443;
  assign n5445 = n5444 ^ n3507;
  assign n5446 = n5445 ^ n5396;
  assign n5447 = n5397 & n5446;
  assign n5448 = n5447 ^ n3518;
  assign n5449 = n5448 ^ n5394;
  assign n5450 = ~n5395 & ~n5449;
  assign n5451 = n5450 ^ n3496;
  assign n5452 = n5451 ^ n5392;
  assign n5453 = n5393 & n5452;
  assign n5454 = n5453 ^ n3521;
  assign n5455 = n5454 ^ n5390;
  assign n5456 = ~n5391 & ~n5455;
  assign n5457 = n5456 ^ n3506;
  assign n5458 = n5457 ^ n5388;
  assign n5459 = ~n5389 & n5458;
  assign n5460 = n5459 ^ n3505;
  assign n5461 = n5460 ^ n5386;
  assign n5462 = ~n5387 & ~n5461;
  assign n5463 = n5462 ^ n3504;
  assign n5474 = n5472 ^ n3503;
  assign n5475 = n5474 ^ n5473;
  assign n5566 = n5463 & ~n5475;
  assign n5567 = ~n5471 & n5566;
  assign n5568 = n5513 & ~n5567;
  assign n5343 = ~n5295 & n5342;
  assign n5287 = n5283 & n5286;
  assign n5344 = n5343 ^ n5287;
  assign n5465 = ~n5287 & n5464;
  assign n5466 = n5344 & ~n5465;
  assign n5279 = n4538 ^ n3813;
  assign n5280 = ~n4989 & ~n5279;
  assign n5281 = n5280 ^ n3813;
  assign n5275 = n5274 ^ n4827;
  assign n5276 = n4829 & n5275;
  assign n5277 = n5276 ^ x147;
  assign n5278 = n5277 ^ n4856;
  assign n5341 = n5281 ^ n5278;
  assign n5467 = n5466 ^ n5341;
  assign n5509 = n5467 ^ n3501;
  assign n5575 = n5568 ^ n5509;
  assign n5573 = ~n5473 & ~n5566;
  assign n5574 = n5573 ^ n5510;
  assign n5578 = n5460 ^ n5387;
  assign n5579 = n5457 ^ n5389;
  assign n5580 = n5451 ^ n5393;
  assign n5581 = n5448 ^ n5395;
  assign n5582 = n5445 ^ n5397;
  assign n5583 = n5442 ^ n5399;
  assign n5584 = n5434 ^ n5401;
  assign n5585 = n5428 ^ n5405;
  assign n5586 = n5425 ^ n5407;
  assign n5588 = n5416 ^ n5414;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = n5419 ^ n5411;
  assign n5591 = n5589 & n5590;
  assign n5592 = n5422 ^ n5409;
  assign n5593 = ~n5591 & ~n5592;
  assign n5594 = ~n5586 & n5593;
  assign n5595 = ~n5585 & n5594;
  assign n5596 = n5595 ^ n5585;
  assign n5597 = n5431 ^ n5403;
  assign n5598 = n5597 ^ n5596;
  assign n5599 = ~n5596 & ~n5598;
  assign n5600 = n5599 ^ n5584;
  assign n5601 = n5584 & n5600;
  assign n5602 = n5439 ^ n3515;
  assign n5603 = n5602 ^ n5437;
  assign n5604 = n5601 & ~n5603;
  assign n5605 = n5583 & n5604;
  assign n5606 = n5605 ^ n5583;
  assign n5607 = ~n5582 & n5606;
  assign n5608 = n5607 ^ n5581;
  assign n5609 = n5581 & n5608;
  assign n5610 = n5580 & n5609;
  assign n5611 = n5454 ^ n5391;
  assign n5612 = n5610 & n5611;
  assign n5613 = ~n5579 & n5612;
  assign n5614 = n5613 ^ n5578;
  assign n5615 = n5578 & n5614;
  assign n5616 = n5474 ^ n5463;
  assign n5650 = n5615 & ~n5616;
  assign n5651 = n5574 & ~n5650;
  assign n5652 = n5575 & ~n5651;
  assign n5569 = n5568 ^ n5467;
  assign n5570 = ~n5509 & n5569;
  assign n5571 = n5570 ^ n3501;
  assign n5476 = n5466 ^ n5278;
  assign n5477 = ~n5341 & ~n5476;
  assign n5478 = n5477 ^ n5281;
  assign n5301 = n4831 & ~n5274;
  assign n5302 = n4858 & ~n5301;
  assign n5303 = n5302 ^ n4848;
  assign n5298 = n4535 ^ n3812;
  assign n5299 = ~n4987 & n5298;
  assign n5300 = n5299 ^ n3812;
  assign n5340 = n5303 ^ n5300;
  assign n5479 = n5478 ^ n5340;
  assign n5508 = n5479 ^ n3529;
  assign n5572 = n5571 ^ n5508;
  assign n5653 = n5652 ^ n5572;
  assign n5654 = n5653 ^ x172;
  assign n5655 = n5651 ^ n5575;
  assign n5656 = n5655 ^ x173;
  assign n5657 = n5650 ^ n5574;
  assign n5658 = n5657 ^ x174;
  assign n5659 = n5616 ^ n5615;
  assign n5660 = n5659 ^ x175;
  assign n5661 = n5614 ^ x176;
  assign n5662 = n5612 ^ n5579;
  assign n5663 = n5662 ^ x177;
  assign n5664 = n5611 ^ n5610;
  assign n5665 = n5664 ^ x178;
  assign n5666 = n5609 ^ n5580;
  assign n5667 = n5666 ^ x179;
  assign n5668 = n5600 ^ x184;
  assign n5669 = n5592 ^ n5591;
  assign n5670 = n5669 ^ x188;
  assign n5671 = x191 & n5587;
  assign n5672 = n5671 ^ x190;
  assign n5673 = n5588 ^ n5587;
  assign n5674 = n5673 ^ n5671;
  assign n5675 = n5672 & ~n5674;
  assign n5676 = n5675 ^ x190;
  assign n5677 = n5676 ^ x189;
  assign n5678 = n5590 ^ n5589;
  assign n5679 = n5678 ^ n5676;
  assign n5680 = n5677 & ~n5679;
  assign n5681 = n5680 ^ x189;
  assign n5682 = n5681 ^ n5669;
  assign n5683 = ~n5670 & n5682;
  assign n5684 = n5683 ^ x188;
  assign n5685 = n5594 ^ n5585;
  assign n5686 = ~x186 & ~n5685;
  assign n5687 = n5593 ^ n5586;
  assign n5689 = n5687 ^ x187;
  assign n5688 = x187 & n5687;
  assign n5690 = n5689 ^ n5688;
  assign n5691 = ~n5686 & n5690;
  assign n5692 = n5684 & n5691;
  assign n5693 = n5685 ^ x186;
  assign n5694 = n5688 ^ n5685;
  assign n5695 = n5693 & ~n5694;
  assign n5696 = n5695 ^ x186;
  assign n5697 = ~n5692 & ~n5696;
  assign n5698 = n5697 ^ x185;
  assign n5699 = n5697 ^ n5598;
  assign n5700 = ~n5698 & n5699;
  assign n5701 = n5700 ^ x185;
  assign n5702 = n5701 ^ n5600;
  assign n5703 = n5668 & ~n5702;
  assign n5704 = n5703 ^ x184;
  assign n5705 = n5604 ^ n5583;
  assign n5706 = ~x182 & n5705;
  assign n5707 = n5603 ^ n5601;
  assign n5709 = x183 & n5707;
  assign n5708 = n5707 ^ x183;
  assign n5710 = n5709 ^ n5708;
  assign n5711 = ~n5706 & n5710;
  assign n5712 = n5606 ^ n5582;
  assign n5713 = ~x181 & n5712;
  assign n5714 = n5711 & ~n5713;
  assign n5715 = ~x180 & ~n5608;
  assign n5716 = n5714 & ~n5715;
  assign n5717 = n5704 & n5716;
  assign n5718 = n5608 ^ x180;
  assign n5719 = n5712 ^ x181;
  assign n5720 = n5709 ^ x182;
  assign n5721 = n5709 ^ n5705;
  assign n5722 = n5720 & n5721;
  assign n5723 = n5722 ^ x182;
  assign n5724 = n5723 ^ n5712;
  assign n5725 = ~n5719 & n5724;
  assign n5726 = n5725 ^ x181;
  assign n5727 = n5726 ^ n5608;
  assign n5728 = n5718 & ~n5727;
  assign n5729 = n5728 ^ x180;
  assign n5730 = ~n5717 & ~n5729;
  assign n5731 = n5730 ^ n5666;
  assign n5732 = ~n5667 & ~n5731;
  assign n5733 = n5732 ^ x179;
  assign n5734 = n5733 ^ n5664;
  assign n5735 = ~n5665 & n5734;
  assign n5736 = n5735 ^ x178;
  assign n5737 = n5736 ^ n5662;
  assign n5738 = n5663 & ~n5737;
  assign n5739 = n5738 ^ x177;
  assign n5740 = n5739 ^ n5614;
  assign n5741 = ~n5661 & n5740;
  assign n5742 = n5741 ^ x176;
  assign n5743 = n5742 ^ n5659;
  assign n5744 = ~n5660 & n5743;
  assign n5745 = n5744 ^ x175;
  assign n5746 = n5745 ^ n5657;
  assign n5747 = n5658 & ~n5746;
  assign n5748 = n5747 ^ x174;
  assign n5749 = n5748 ^ n5655;
  assign n5750 = ~n5656 & n5749;
  assign n5751 = n5750 ^ x173;
  assign n5752 = n5751 ^ n5653;
  assign n5753 = n5654 & ~n5752;
  assign n5754 = n5753 ^ x172;
  assign n6263 = n5754 ^ x171;
  assign n5576 = ~n5574 & n5575;
  assign n5577 = n5572 & n5576;
  assign n5514 = n5513 ^ n5467;
  assign n5515 = ~n5509 & n5514;
  assign n5516 = n5515 ^ n3501;
  assign n5517 = n5516 ^ n5479;
  assign n5518 = ~n5508 & ~n5517;
  assign n5519 = n5518 ^ n3529;
  assign n5468 = n3501 & ~n5467;
  assign n5480 = ~n3529 & n5479;
  assign n5481 = ~n5475 & ~n5480;
  assign n5482 = ~n5471 & n5481;
  assign n5483 = ~n5468 & n5482;
  assign n5554 = n5463 & n5483;
  assign n5555 = ~n5519 & ~n5554;
  assign n5345 = n5344 ^ n5278;
  assign n5346 = ~n5341 & ~n5345;
  assign n5347 = n5346 ^ n5281;
  assign n5348 = n5347 ^ n5300;
  assign n5349 = ~n5340 & n5348;
  assign n5350 = n5349 ^ n5303;
  assign n5282 = n5278 & ~n5281;
  assign n5304 = n5300 & ~n5303;
  assign n5305 = n5297 & ~n5304;
  assign n5306 = ~n5287 & n5305;
  assign n5307 = ~n5282 & n5306;
  assign n5484 = n5272 & n5307;
  assign n5485 = ~n5350 & ~n5484;
  assign n5312 = n4531 ^ n3810;
  assign n5313 = n4978 & n5312;
  assign n5314 = n5313 ^ n3810;
  assign n5308 = n5302 ^ n4847;
  assign n5309 = ~n4848 & ~n5308;
  assign n5310 = n5309 ^ x145;
  assign n5311 = n5310 ^ n4855;
  assign n5316 = n5314 ^ n5311;
  assign n5486 = n5485 ^ n5316;
  assign n5488 = n5486 ^ n3593;
  assign n5565 = n5555 ^ n5488;
  assign n5647 = n5577 ^ n5565;
  assign n5617 = n5575 & ~n5616;
  assign n5618 = n5572 & n5617;
  assign n5619 = n5615 & n5618;
  assign n5620 = ~n5577 & n5619;
  assign n5648 = n5647 ^ n5620;
  assign n6264 = n6263 ^ n5648;
  assign n6378 = n6377 ^ n6264;
  assign n5323 = n4783 & ~n4879;
  assign n5324 = n5323 ^ n4784;
  assign n5325 = n5324 ^ n4779;
  assign n6379 = n4987 ^ n4444;
  assign n6380 = ~n5325 & ~n6379;
  assign n6381 = n6380 ^ n4444;
  assign n6316 = n5730 ^ x179;
  assign n6317 = n6316 ^ n5666;
  assign n6382 = n6381 ^ n6317;
  assign n6096 = n5704 & n5711;
  assign n6097 = ~n5723 & ~n6096;
  assign n6165 = n6097 ^ n5712;
  assign n6166 = ~n5719 & ~n6165;
  assign n6167 = n6166 ^ x181;
  assign n6168 = n6167 ^ n5718;
  assign n6098 = n6097 ^ n5719;
  assign n6087 = n5705 ^ x182;
  assign n6085 = n5704 & n5708;
  assign n6086 = n6085 ^ n5709;
  assign n6088 = n6087 ^ n6086;
  assign n6014 = n5708 ^ n5704;
  assign n6011 = n4901 ^ n4340;
  assign n6012 = ~n5278 & ~n6011;
  assign n6013 = n6012 ^ n4340;
  assign n6015 = n6014 ^ n6013;
  assign n6019 = n5701 ^ n5668;
  assign n6016 = n4891 ^ n4323;
  assign n6017 = ~n5283 & n6016;
  assign n6018 = n6017 ^ n4323;
  assign n6020 = n6019 ^ n6018;
  assign n6021 = n4713 ^ n4302;
  assign n6022 = n5291 & ~n6021;
  assign n6023 = n6022 ^ n4302;
  assign n5991 = n5598 ^ x185;
  assign n5992 = n5991 ^ n5697;
  assign n6024 = n6023 ^ n5992;
  assign n6025 = n4456 ^ n4305;
  assign n6026 = n4907 & n6025;
  assign n6027 = n6026 ^ n4305;
  assign n5998 = n5684 & n5689;
  assign n5999 = n5998 ^ n5688;
  assign n6000 = n5999 ^ n5693;
  assign n6028 = n6027 ^ n6000;
  assign n6032 = n5689 ^ n5684;
  assign n6029 = n4469 ^ n4309;
  assign n6030 = ~n4915 & n6029;
  assign n6031 = n6030 ^ n4309;
  assign n6033 = n6032 ^ n6031;
  assign n6037 = n5681 ^ n5670;
  assign n6034 = n4471 ^ n4213;
  assign n6035 = ~n4920 & ~n6034;
  assign n6036 = n6035 ^ n4213;
  assign n6038 = n6037 ^ n6036;
  assign n6042 = n5678 ^ x189;
  assign n6043 = n6042 ^ n5676;
  assign n6039 = n4478 ^ n4204;
  assign n6040 = ~n4925 & n6039;
  assign n6041 = n6040 ^ n4204;
  assign n6044 = n6043 ^ n6041;
  assign n6048 = n5673 ^ n5672;
  assign n6045 = n4483 ^ n4194;
  assign n6046 = n4930 & n6045;
  assign n6047 = n6046 ^ n4194;
  assign n6049 = n6048 ^ n6047;
  assign n6050 = n4488 ^ n4142;
  assign n6051 = ~n4935 & ~n6050;
  assign n6052 = n6051 ^ n4142;
  assign n6054 = n6053 ^ n6052;
  assign n5981 = n4687 ^ n3776;
  assign n5982 = ~n4940 & ~n5981;
  assign n5983 = n5982 ^ n3776;
  assign n5843 = n4096 ^ n3708;
  assign n5844 = n4640 & ~n5843;
  assign n5845 = n5844 ^ n3708;
  assign n5377 = ~n4879 & n5167;
  assign n5378 = n5129 & ~n5377;
  assign n5787 = n5134 & ~n5378;
  assign n5788 = n5141 & ~n5787;
  assign n5839 = n5788 ^ n5121;
  assign n5840 = n5136 & n5839;
  assign n5841 = n5840 ^ x137;
  assign n5842 = n5841 ^ n5120;
  assign n5846 = n5845 ^ n5842;
  assign n5315 = n5311 & ~n5314;
  assign n5317 = n5316 ^ n5315;
  assign n5318 = n4528 ^ n3860;
  assign n5319 = n4973 & n5318;
  assign n5320 = n5319 ^ n3860;
  assign n5321 = n4879 ^ n4783;
  assign n5322 = ~n5320 & n5321;
  assign n5326 = n4526 ^ n3808;
  assign n5327 = n4969 & ~n5326;
  assign n5328 = n5327 ^ n3808;
  assign n5329 = n5325 & ~n5328;
  assign n4882 = ~n4879 & n4881;
  assign n4883 = ~n4787 & ~n4882;
  assign n5330 = n4883 ^ n4777;
  assign n5331 = n4523 ^ n3913;
  assign n5332 = n5063 & ~n5331;
  assign n5333 = n5332 ^ n3913;
  assign n5334 = n5330 & ~n5333;
  assign n5335 = ~n5329 & ~n5334;
  assign n5336 = ~n5322 & n5335;
  assign n5337 = ~n5317 & n5336;
  assign n5338 = n5307 & n5337;
  assign n5339 = n5272 & n5338;
  assign n5351 = n5337 & n5350;
  assign n5352 = n5333 ^ n5330;
  assign n5353 = n5328 ^ n5325;
  assign n5354 = n5321 ^ n5320;
  assign n5355 = ~n5315 & ~n5354;
  assign n5356 = n5355 ^ n5322;
  assign n5357 = n5356 ^ n5325;
  assign n5358 = ~n5353 & ~n5357;
  assign n5359 = n5358 ^ n5328;
  assign n5360 = n5359 ^ n5330;
  assign n5361 = ~n5352 & ~n5360;
  assign n5362 = n5361 ^ n5330;
  assign n5363 = ~n5351 & n5362;
  assign n5364 = ~n5339 & n5363;
  assign n5543 = n5378 ^ n5130;
  assign n5544 = n5138 & n5543;
  assign n5545 = n5544 ^ x139;
  assign n5546 = n5545 ^ n5137;
  assign n5547 = n4107 ^ n3709;
  assign n5548 = ~n5192 & n5547;
  assign n5549 = n5548 ^ n3709;
  assign n5826 = ~n5546 & ~n5549;
  assign n4452 = n4451 ^ n3916;
  assign n4453 = n4450 & ~n4452;
  assign n4454 = n4453 ^ n3916;
  assign n4884 = n4883 ^ n4776;
  assign n4885 = n4777 & n4884;
  assign n4886 = n4885 ^ x141;
  assign n4899 = n4898 ^ n4886;
  assign n5370 = ~n4454 & ~n4899;
  assign n5374 = n4102 ^ n3738;
  assign n5375 = ~n5099 & ~n5374;
  assign n5376 = n5375 ^ n3738;
  assign n5379 = n5378 ^ n5138;
  assign n5539 = n5376 & n5379;
  assign n5784 = n4098 ^ n3711;
  assign n5785 = n4645 & ~n5784;
  assign n5786 = n5785 ^ n3711;
  assign n5789 = n5788 ^ n5136;
  assign n5827 = ~n5786 & n5789;
  assign n5828 = ~n5539 & ~n5827;
  assign n5829 = ~n5370 & n5828;
  assign n5830 = ~n5826 & n5829;
  assign n5831 = ~n5364 & n5830;
  assign n5790 = n5789 ^ n5786;
  assign n5550 = n5549 ^ n5546;
  assign n4900 = n4899 ^ n4454;
  assign n5371 = n5370 ^ n4900;
  assign n5380 = n5379 ^ n5376;
  assign n5538 = n5371 & n5380;
  assign n5540 = n5539 ^ n5538;
  assign n5832 = n5546 ^ n5540;
  assign n5833 = n5550 & n5832;
  assign n5834 = n5833 ^ n5549;
  assign n5835 = n5834 ^ n5789;
  assign n5836 = ~n5790 & n5835;
  assign n5837 = n5836 ^ n5786;
  assign n5838 = ~n5831 & ~n5837;
  assign n5878 = n5842 ^ n5838;
  assign n5879 = ~n5846 & n5878;
  assign n5880 = n5879 ^ n5845;
  assign n5874 = n4093 ^ n3722;
  assign n5875 = ~n4654 & ~n5874;
  assign n5876 = n5875 ^ n3722;
  assign n5873 = n5872 ^ n5151;
  assign n5877 = n5876 ^ n5873;
  assign n5881 = n5880 ^ n5877;
  assign n5882 = n5881 ^ n3394;
  assign n5847 = n5846 ^ n5838;
  assign n5848 = n5847 ^ n3397;
  assign n5487 = ~n3593 & n5486;
  assign n5489 = n5488 ^ n5487;
  assign n5490 = ~n5317 & ~n5485;
  assign n5491 = ~n5315 & ~n5490;
  assign n5492 = n5491 ^ n5354;
  assign n5493 = n3598 & ~n5492;
  assign n5494 = ~n5322 & n5490;
  assign n5495 = n5356 & ~n5494;
  assign n5496 = n5495 ^ n5353;
  assign n5497 = ~n3604 & ~n5496;
  assign n5498 = n5495 ^ n5328;
  assign n5499 = ~n5353 & n5498;
  assign n5500 = n5499 ^ n5325;
  assign n5501 = n5500 ^ n5352;
  assign n5502 = ~n3611 & ~n5501;
  assign n5503 = ~n5497 & ~n5502;
  assign n5504 = ~n5493 & n5503;
  assign n5505 = ~n5489 & n5504;
  assign n5506 = n5483 & n5505;
  assign n5507 = n5463 & n5506;
  assign n5520 = n5505 & n5519;
  assign n5521 = n5501 ^ n3611;
  assign n5522 = n5496 ^ n3604;
  assign n5523 = n5492 ^ n3598;
  assign n5524 = n5492 ^ n5487;
  assign n5525 = ~n5523 & ~n5524;
  assign n5526 = n5525 ^ n3598;
  assign n5527 = n5526 ^ n5496;
  assign n5528 = n5522 & n5527;
  assign n5529 = n5528 ^ n3604;
  assign n5530 = n5529 ^ n5501;
  assign n5531 = n5521 & n5530;
  assign n5532 = n5531 ^ n5501;
  assign n5533 = ~n5520 & ~n5532;
  assign n5534 = ~n5507 & n5533;
  assign n5372 = ~n5364 & ~n5370;
  assign n5541 = n5372 & ~n5539;
  assign n5542 = n5540 & ~n5541;
  assign n5551 = n5550 ^ n5542;
  assign n5813 = ~n3381 & n5551;
  assign n5373 = n5371 & ~n5372;
  assign n5381 = n5380 ^ n5373;
  assign n5385 = ~n3377 & n5381;
  assign n5365 = n5364 ^ n4900;
  assign n5367 = ~n3716 & n5365;
  assign n5781 = n5546 ^ n5542;
  assign n5782 = n5550 & n5781;
  assign n5783 = n5782 ^ n5549;
  assign n5791 = n5790 ^ n5783;
  assign n5814 = n3389 & n5791;
  assign n5815 = ~n5367 & ~n5814;
  assign n5816 = ~n5385 & n5815;
  assign n5817 = ~n5813 & n5816;
  assign n5818 = ~n5534 & n5817;
  assign n5792 = n5791 ^ n3389;
  assign n5552 = n5551 ^ n3381;
  assign n5366 = n5365 ^ n3716;
  assign n5368 = n5367 ^ n5366;
  assign n5369 = n5368 ^ n3377;
  assign n5382 = n5381 ^ n5368;
  assign n5383 = n5369 & n5382;
  assign n5384 = n5383 ^ n3377;
  assign n5819 = n5551 ^ n5384;
  assign n5820 = ~n5552 & n5819;
  assign n5821 = n5820 ^ n3381;
  assign n5822 = n5821 ^ n5791;
  assign n5823 = n5792 & n5822;
  assign n5824 = n5823 ^ n3389;
  assign n5825 = ~n5818 & n5824;
  assign n5868 = n5847 ^ n5825;
  assign n5869 = n5848 & n5868;
  assign n5870 = n5869 ^ n3397;
  assign n5923 = n5881 ^ n5870;
  assign n5924 = n5882 & n5923;
  assign n5925 = n5924 ^ n3394;
  assign n5918 = n5880 ^ n5876;
  assign n5919 = n5877 & n5918;
  assign n5920 = n5919 ^ n5873;
  assign n5910 = n3804 ^ n3499;
  assign n5911 = n4631 & ~n5910;
  assign n5912 = n5911 ^ n3499;
  assign n5917 = n5916 ^ n5912;
  assign n5921 = n5920 ^ n5917;
  assign n5922 = n5921 ^ x31;
  assign n5926 = n5925 ^ n5922;
  assign n5883 = n5882 ^ n5870;
  assign n5535 = ~n5367 & ~n5534;
  assign n5536 = ~n5385 & n5535;
  assign n5537 = ~n5384 & ~n5536;
  assign n5777 = n5537 ^ n3381;
  assign n5778 = n5551 ^ n5537;
  assign n5779 = ~n5777 & ~n5778;
  assign n5780 = n5779 ^ n3381;
  assign n5793 = n5792 ^ n5780;
  assign n5553 = n5552 ^ n5537;
  assign n5556 = ~n5489 & ~n5555;
  assign n5557 = ~n5493 & n5556;
  assign n5558 = n5526 & ~n5557;
  assign n5559 = n5558 ^ n5496;
  assign n5560 = n5522 & n5559;
  assign n5561 = n5560 ^ n3604;
  assign n5562 = n5561 ^ n5521;
  assign n5563 = ~n5487 & ~n5556;
  assign n5564 = n5563 ^ n5523;
  assign n5621 = n5620 ^ n5577;
  assign n5622 = n5565 & ~n5621;
  assign n5623 = n5622 ^ n5565;
  assign n5624 = n5564 & n5623;
  assign n5625 = n5558 ^ n5522;
  assign n5626 = n5625 ^ n5624;
  assign n5627 = n5624 & n5626;
  assign n5628 = ~n5562 & ~n5627;
  assign n5629 = n5534 ^ n5366;
  assign n5630 = n5628 & n5629;
  assign n5631 = n5630 ^ n5629;
  assign n5633 = n5381 ^ n3377;
  assign n5632 = ~n5368 & ~n5535;
  assign n5634 = n5633 ^ n5632;
  assign n5635 = ~n5631 & ~n5634;
  assign n5794 = n5553 & ~n5635;
  assign n5812 = ~n5793 & ~n5794;
  assign n5849 = n5848 ^ n5825;
  assign n5867 = n5812 & n5849;
  assign n5884 = n5883 ^ n5867;
  assign n5909 = n5883 & n5884;
  assign n5927 = n5926 ^ n5909;
  assign n5975 = n5927 ^ x161;
  assign n5885 = n5884 ^ x162;
  assign n5850 = n5849 ^ n5812;
  assign n5851 = n5850 ^ x163;
  assign n5795 = n5794 ^ n5793;
  assign n5808 = n5795 ^ x164;
  assign n5636 = n5635 ^ n5553;
  assign n5637 = n5636 ^ x165;
  assign n5638 = n5634 ^ n5631;
  assign n5639 = n5638 ^ x166;
  assign n5640 = n5629 ^ n5628;
  assign n5641 = n5640 ^ x167;
  assign n5642 = n5627 ^ n5562;
  assign n5643 = n5642 ^ x168;
  assign n5644 = n5626 ^ x169;
  assign n5645 = n5623 ^ n5564;
  assign n5646 = n5645 ^ x170;
  assign n5649 = n5648 ^ x171;
  assign n5755 = n5754 ^ n5648;
  assign n5756 = n5649 & ~n5755;
  assign n5757 = n5756 ^ x171;
  assign n5758 = n5757 ^ n5645;
  assign n5759 = n5646 & ~n5758;
  assign n5760 = n5759 ^ x170;
  assign n5761 = n5760 ^ n5626;
  assign n5762 = ~n5644 & n5761;
  assign n5763 = n5762 ^ x169;
  assign n5764 = n5763 ^ n5642;
  assign n5765 = ~n5643 & n5764;
  assign n5766 = n5765 ^ x168;
  assign n5767 = n5766 ^ n5640;
  assign n5768 = ~n5641 & n5767;
  assign n5769 = n5768 ^ x167;
  assign n5770 = n5769 ^ n5638;
  assign n5771 = ~n5639 & n5770;
  assign n5772 = n5771 ^ x166;
  assign n5773 = n5772 ^ n5636;
  assign n5774 = ~n5637 & n5773;
  assign n5775 = n5774 ^ x165;
  assign n5809 = n5795 ^ n5775;
  assign n5810 = ~n5808 & n5809;
  assign n5811 = n5810 ^ x164;
  assign n5864 = n5850 ^ n5811;
  assign n5865 = ~n5851 & n5864;
  assign n5866 = n5865 ^ x163;
  assign n5905 = n5884 ^ n5866;
  assign n5906 = ~n5885 & n5905;
  assign n5907 = n5906 ^ x162;
  assign n5976 = n5927 ^ n5907;
  assign n5977 = n5975 & ~n5976;
  assign n5978 = n5977 ^ x161;
  assign n5979 = n5978 ^ x160;
  assign n5969 = n5925 ^ x31;
  assign n5970 = n5925 ^ n5921;
  assign n5971 = n5969 & ~n5970;
  assign n5972 = n5971 ^ x31;
  assign n5964 = n5920 ^ n5916;
  assign n5965 = ~n5917 & ~n5964;
  assign n5966 = n5965 ^ n5912;
  assign n5960 = n5154 & ~n5872;
  assign n5961 = n5160 & ~n5960;
  assign n5962 = n5961 ^ n5118;
  assign n5957 = n3799 ^ n3498;
  assign n5958 = n4626 & n5957;
  assign n5959 = n5958 ^ n3498;
  assign n5963 = n5962 ^ n5959;
  assign n5967 = n5966 ^ n5963;
  assign n5968 = n5967 ^ n3406;
  assign n5973 = n5972 ^ n5968;
  assign n5956 = ~n5909 & n5926;
  assign n5974 = n5973 ^ n5956;
  assign n5980 = n5979 ^ n5974;
  assign n5984 = n5983 ^ n5980;
  assign n5908 = n5907 ^ x161;
  assign n5928 = n5927 ^ n5908;
  assign n5902 = n4496 ^ n3781;
  assign n5903 = n4942 & ~n5902;
  assign n5904 = n5903 ^ n3781;
  assign n5929 = n5928 ^ n5904;
  assign n5886 = n5885 ^ n5866;
  assign n5861 = n4676 ^ n3786;
  assign n5862 = n4950 & ~n5861;
  assign n5863 = n5862 ^ n3786;
  assign n5887 = n5886 ^ n5863;
  assign n5852 = n5851 ^ n5811;
  assign n5804 = n4499 ^ n3790;
  assign n5805 = ~n4955 & ~n5804;
  assign n5806 = n5805 ^ n3790;
  assign n5857 = n5852 ^ n5806;
  assign n5776 = n5775 ^ x164;
  assign n5796 = n5795 ^ n5776;
  assign n5797 = n4508 ^ n3794;
  assign n5798 = n4960 & n5797;
  assign n5799 = n5798 ^ n3794;
  assign n5803 = ~n5796 & ~n5799;
  assign n5858 = n5852 ^ n5803;
  assign n5859 = n5857 & ~n5858;
  assign n5860 = n5859 ^ n5803;
  assign n5899 = n5886 ^ n5860;
  assign n5900 = ~n5887 & n5899;
  assign n5901 = n5900 ^ n5863;
  assign n5953 = n5928 ^ n5901;
  assign n5954 = ~n5929 & ~n5953;
  assign n5955 = n5954 ^ n5904;
  assign n6055 = n5980 ^ n5955;
  assign n6056 = n5984 & n6055;
  assign n6057 = n6056 ^ n5983;
  assign n6058 = n6057 ^ n6053;
  assign n6059 = ~n6054 & ~n6058;
  assign n6060 = n6059 ^ n6052;
  assign n6061 = n6060 ^ n6048;
  assign n6062 = n6049 & n6061;
  assign n6063 = n6062 ^ n6047;
  assign n6064 = n6063 ^ n6043;
  assign n6065 = n6044 & ~n6064;
  assign n6066 = n6065 ^ n6041;
  assign n6067 = n6066 ^ n6037;
  assign n6068 = ~n6038 & n6067;
  assign n6069 = n6068 ^ n6036;
  assign n6070 = n6069 ^ n6032;
  assign n6071 = ~n6033 & ~n6070;
  assign n6072 = n6071 ^ n6031;
  assign n6073 = n6072 ^ n6000;
  assign n6074 = n6028 & n6073;
  assign n6075 = n6074 ^ n6027;
  assign n6076 = n6075 ^ n5992;
  assign n6077 = ~n6024 & n6076;
  assign n6078 = n6077 ^ n6023;
  assign n6079 = n6078 ^ n6019;
  assign n6080 = ~n6020 & ~n6079;
  assign n6081 = n6080 ^ n6018;
  assign n6082 = n6081 ^ n6014;
  assign n6083 = ~n6015 & n6082;
  assign n6084 = n6083 ^ n6013;
  assign n6089 = n6088 ^ n6084;
  assign n6090 = n4999 ^ n4357;
  assign n6091 = n5303 & n6090;
  assign n6092 = n6091 ^ n4357;
  assign n6093 = n6092 ^ n6088;
  assign n6094 = ~n6089 & n6093;
  assign n6095 = n6094 ^ n6092;
  assign n6099 = n6098 ^ n6095;
  assign n6008 = n4998 ^ n4383;
  assign n6009 = n5311 & n6008;
  assign n6010 = n6009 ^ n4383;
  assign n6162 = n6098 ^ n6010;
  assign n6163 = n6099 & n6162;
  assign n6164 = n6163 ^ n6010;
  assign n6169 = n6168 ^ n6164;
  assign n6159 = n4989 ^ n4397;
  assign n6160 = ~n5321 & n6159;
  assign n6161 = n6160 ^ n4397;
  assign n6383 = n6168 ^ n6161;
  assign n6384 = ~n6169 & ~n6383;
  assign n6385 = n6384 ^ n6161;
  assign n6386 = n6385 ^ n6317;
  assign n6387 = n6382 & n6386;
  assign n6388 = n6387 ^ n6381;
  assign n6309 = n5733 ^ n5665;
  assign n6389 = n6388 ^ n6309;
  assign n6390 = n4978 ^ n4538;
  assign n6391 = ~n5330 & ~n6390;
  assign n6392 = n6391 ^ n4538;
  assign n6393 = n6392 ^ n6309;
  assign n6394 = n6389 & n6393;
  assign n6395 = n6394 ^ n6392;
  assign n6303 = n5736 ^ n5663;
  assign n6396 = n6395 ^ n6303;
  assign n6397 = n4973 ^ n4535;
  assign n6398 = n4899 & ~n6397;
  assign n6399 = n6398 ^ n4535;
  assign n6400 = n6399 ^ n6303;
  assign n6401 = n6396 & ~n6400;
  assign n6402 = n6401 ^ n6399;
  assign n6297 = n5739 ^ n5661;
  assign n6403 = n6402 ^ n6297;
  assign n6404 = n4969 ^ n4531;
  assign n6405 = ~n5379 & ~n6404;
  assign n6406 = n6405 ^ n4531;
  assign n6407 = n6406 ^ n6297;
  assign n6408 = ~n6403 & n6407;
  assign n6409 = n6408 ^ n6406;
  assign n6290 = n5742 ^ n5660;
  assign n6410 = n6409 ^ n6290;
  assign n6411 = n5063 ^ n4528;
  assign n6412 = n5546 & n6411;
  assign n6413 = n6412 ^ n4528;
  assign n6414 = n6413 ^ n6290;
  assign n6415 = ~n6410 & ~n6414;
  assign n6416 = n6415 ^ n6413;
  assign n6284 = n5745 ^ n5658;
  assign n6417 = n6416 ^ n6284;
  assign n6418 = n4526 ^ n4450;
  assign n6419 = ~n5789 & ~n6418;
  assign n6420 = n6419 ^ n4526;
  assign n6421 = n6420 ^ n6284;
  assign n6422 = ~n6417 & ~n6421;
  assign n6423 = n6422 ^ n6420;
  assign n6277 = n5748 ^ n5656;
  assign n6424 = n6423 ^ n6277;
  assign n6425 = n5099 ^ n4523;
  assign n6426 = n5842 & n6425;
  assign n6427 = n6426 ^ n4523;
  assign n6428 = n6427 ^ n6277;
  assign n6429 = ~n6424 & n6428;
  assign n6430 = n6429 ^ n6427;
  assign n6271 = n5751 ^ n5654;
  assign n6431 = n6430 ^ n6271;
  assign n6432 = n5192 ^ n4451;
  assign n6433 = n5873 & n6432;
  assign n6434 = n6433 ^ n4451;
  assign n6435 = n6434 ^ n6271;
  assign n6436 = n6431 & ~n6435;
  assign n6437 = n6436 ^ n6434;
  assign n6438 = n6437 ^ n6264;
  assign n6439 = n6378 & n6438;
  assign n6440 = n6439 ^ n6377;
  assign n6371 = n4640 ^ n4107;
  assign n6372 = n5962 & n6371;
  assign n6373 = n6372 ^ n4107;
  assign n6460 = n6440 ^ n6373;
  assign n6004 = n5757 ^ n5646;
  assign n6461 = n6460 ^ n6004;
  assign n6462 = n6461 ^ n3709;
  assign n6463 = n6437 ^ n6377;
  assign n6464 = n6463 ^ n6264;
  assign n6465 = n6464 ^ n3738;
  assign n6466 = n6434 ^ n6431;
  assign n6467 = n6466 ^ n3916;
  assign n6468 = n6427 ^ n6424;
  assign n6469 = n6468 ^ n3913;
  assign n6470 = n6420 ^ n6417;
  assign n6471 = n6470 ^ n3808;
  assign n6472 = n6413 ^ n6410;
  assign n6473 = n6472 ^ n3860;
  assign n6474 = n6406 ^ n6403;
  assign n6475 = n6474 ^ n3810;
  assign n6476 = n6399 ^ n6396;
  assign n6477 = n6476 ^ n3812;
  assign n6478 = n6392 ^ n6389;
  assign n6479 = n6478 ^ n3813;
  assign n6480 = n6385 ^ n6382;
  assign n6481 = n6480 ^ n3853;
  assign n6170 = n6169 ^ n6161;
  assign n6482 = n6170 ^ n3851;
  assign n6100 = n6099 ^ n6010;
  assign n6101 = n6100 ^ n3849;
  assign n6102 = n6092 ^ n6089;
  assign n6103 = n6102 ^ n3815;
  assign n6104 = n6081 ^ n6015;
  assign n6105 = n6104 ^ n3817;
  assign n6106 = n6078 ^ n6020;
  assign n6107 = n6106 ^ n3818;
  assign n6108 = n6075 ^ n6024;
  assign n6109 = n6108 ^ n3819;
  assign n6110 = n6072 ^ n6028;
  assign n6111 = n6110 ^ n3820;
  assign n6112 = n6069 ^ n6033;
  assign n6113 = n6112 ^ n3495;
  assign n6114 = n6066 ^ n6038;
  assign n6115 = n6114 ^ n3778;
  assign n6116 = n6063 ^ n6044;
  assign n6117 = n6116 ^ n3784;
  assign n6118 = n6060 ^ n6049;
  assign n6119 = n6118 ^ n3788;
  assign n6120 = n6057 ^ n6054;
  assign n6121 = n6120 ^ n3792;
  assign n5985 = n5984 ^ n5955;
  assign n5986 = n5985 ^ n3797;
  assign n5930 = n5929 ^ n5901;
  assign n5949 = n5930 ^ n3802;
  assign n5888 = n5887 ^ n5860;
  assign n5889 = n5888 ^ n3806;
  assign n5800 = n5799 ^ n5796;
  assign n5801 = n3391 & n5800;
  assign n5802 = n5801 ^ n3826;
  assign n5807 = n5806 ^ n5803;
  assign n5853 = n5852 ^ n5807;
  assign n5854 = n5853 ^ n5801;
  assign n5855 = n5802 & n5854;
  assign n5856 = n5855 ^ n3826;
  assign n5895 = n5888 ^ n5856;
  assign n5896 = ~n5889 & n5895;
  assign n5897 = n5896 ^ n3806;
  assign n5950 = n5930 ^ n5897;
  assign n5951 = ~n5949 & n5950;
  assign n5952 = n5951 ^ n3802;
  assign n6122 = n5985 ^ n5952;
  assign n6123 = n5986 & n6122;
  assign n6124 = n6123 ^ n3797;
  assign n6125 = n6124 ^ n6120;
  assign n6126 = n6121 & ~n6125;
  assign n6127 = n6126 ^ n3792;
  assign n6128 = n6127 ^ n6118;
  assign n6129 = n6119 & ~n6128;
  assign n6130 = n6129 ^ n3788;
  assign n6131 = n6130 ^ n6116;
  assign n6132 = ~n6117 & n6131;
  assign n6133 = n6132 ^ n3784;
  assign n6134 = n6133 ^ n6114;
  assign n6135 = n6115 & ~n6134;
  assign n6136 = n6135 ^ n3778;
  assign n6137 = n6136 ^ n6112;
  assign n6138 = n6113 & ~n6137;
  assign n6139 = n6138 ^ n3495;
  assign n6140 = n6139 ^ n6110;
  assign n6141 = ~n6111 & ~n6140;
  assign n6142 = n6141 ^ n3820;
  assign n6143 = n6142 ^ n6108;
  assign n6144 = ~n6109 & n6143;
  assign n6145 = n6144 ^ n3819;
  assign n6146 = n6145 ^ n6106;
  assign n6147 = n6107 & n6146;
  assign n6148 = n6147 ^ n3818;
  assign n6149 = n6148 ^ n6104;
  assign n6150 = n6105 & n6149;
  assign n6151 = n6150 ^ n3817;
  assign n6152 = n6151 ^ n6102;
  assign n6153 = n6103 & n6152;
  assign n6154 = n6153 ^ n3815;
  assign n6155 = n6154 ^ n6100;
  assign n6156 = ~n6101 & ~n6155;
  assign n6157 = n6156 ^ n3849;
  assign n6483 = n6170 ^ n6157;
  assign n6484 = ~n6482 & n6483;
  assign n6485 = n6484 ^ n3851;
  assign n6486 = n6485 ^ n6480;
  assign n6487 = n6481 & n6486;
  assign n6488 = n6487 ^ n3853;
  assign n6489 = n6488 ^ n6478;
  assign n6490 = n6479 & n6489;
  assign n6491 = n6490 ^ n3813;
  assign n6492 = n6491 ^ n6476;
  assign n6493 = ~n6477 & ~n6492;
  assign n6494 = n6493 ^ n3812;
  assign n6495 = n6494 ^ n6474;
  assign n6496 = n6475 & ~n6495;
  assign n6497 = n6496 ^ n3810;
  assign n6498 = n6497 ^ n6472;
  assign n6499 = n6473 & n6498;
  assign n6500 = n6499 ^ n3860;
  assign n6501 = n6500 ^ n6470;
  assign n6502 = ~n6471 & n6501;
  assign n6503 = n6502 ^ n3808;
  assign n6504 = n6503 ^ n6468;
  assign n6505 = ~n6469 & n6504;
  assign n6506 = n6505 ^ n3913;
  assign n6507 = n6506 ^ n6466;
  assign n6508 = n6467 & ~n6507;
  assign n6509 = n6508 ^ n3916;
  assign n6510 = n6509 ^ n6464;
  assign n6511 = n6465 & n6510;
  assign n6512 = n6511 ^ n3738;
  assign n6513 = n6512 ^ n6461;
  assign n6514 = n6462 & n6513;
  assign n6515 = n6514 ^ n3709;
  assign n6555 = n6515 ^ n3711;
  assign n6374 = n6373 ^ n6004;
  assign n6441 = n6440 ^ n6004;
  assign n6442 = n6374 & ~n6441;
  assign n6443 = n6442 ^ n6373;
  assign n6367 = n4654 ^ n4098;
  assign n6368 = n5223 & n6367;
  assign n6369 = n6368 ^ n4098;
  assign n6365 = n5760 ^ x169;
  assign n6366 = n6365 ^ n5626;
  assign n6370 = n6369 ^ n6366;
  assign n6458 = n6443 ^ n6370;
  assign n6556 = n6555 ^ n6458;
  assign n6524 = n6512 ^ n3709;
  assign n6525 = n6524 ^ n6461;
  assign n6526 = n6497 ^ n3860;
  assign n6527 = n6526 ^ n6472;
  assign n6528 = n6491 ^ n3812;
  assign n6529 = n6528 ^ n6476;
  assign n6530 = n6488 ^ n3813;
  assign n6531 = n6530 ^ n6478;
  assign n6532 = n6485 ^ n3853;
  assign n6533 = n6532 ^ n6480;
  assign n6158 = n6157 ^ n3851;
  assign n6171 = n6170 ^ n6158;
  assign n6172 = n6151 ^ n6103;
  assign n6173 = n6142 ^ n3819;
  assign n6174 = n6173 ^ n6108;
  assign n6175 = n6136 ^ n3495;
  assign n6176 = n6175 ^ n6112;
  assign n6177 = n6127 ^ n6119;
  assign n6178 = n6124 ^ n3792;
  assign n6179 = n6178 ^ n6120;
  assign n5890 = n5889 ^ n5856;
  assign n5891 = n5853 ^ n5802;
  assign n5892 = n5800 ^ n3391;
  assign n5893 = ~n5891 & n5892;
  assign n5894 = ~n5890 & n5893;
  assign n5898 = n5897 ^ n3802;
  assign n5931 = n5930 ^ n5898;
  assign n5948 = ~n5894 & n5931;
  assign n5987 = n5986 ^ n5952;
  assign n6180 = n5948 & ~n5987;
  assign n6181 = ~n6179 & ~n6180;
  assign n6182 = ~n6177 & n6181;
  assign n6183 = n6130 ^ n3784;
  assign n6184 = n6183 ^ n6116;
  assign n6185 = ~n6182 & ~n6184;
  assign n6186 = n6133 ^ n6115;
  assign n6187 = n6185 & n6186;
  assign n6188 = ~n6176 & ~n6187;
  assign n6189 = n6139 ^ n6111;
  assign n6190 = n6188 & n6189;
  assign n6191 = n6174 & ~n6190;
  assign n6192 = n6145 ^ n6107;
  assign n6193 = n6191 & ~n6192;
  assign n6194 = n6148 ^ n3817;
  assign n6195 = n6194 ^ n6104;
  assign n6196 = n6193 & n6195;
  assign n6197 = ~n6172 & n6196;
  assign n6198 = n6154 ^ n3849;
  assign n6199 = n6198 ^ n6100;
  assign n6200 = ~n6197 & n6199;
  assign n6534 = ~n6171 & n6200;
  assign n6535 = ~n6533 & ~n6534;
  assign n6536 = ~n6531 & ~n6535;
  assign n6537 = ~n6529 & n6536;
  assign n6538 = n6494 ^ n3810;
  assign n6539 = n6538 ^ n6474;
  assign n6540 = n6537 & ~n6539;
  assign n6541 = ~n6527 & n6540;
  assign n6542 = n6500 ^ n3808;
  assign n6543 = n6542 ^ n6470;
  assign n6544 = n6541 & ~n6543;
  assign n6545 = n6503 ^ n3913;
  assign n6546 = n6545 ^ n6468;
  assign n6547 = ~n6544 & n6546;
  assign n6548 = n6506 ^ n3916;
  assign n6549 = n6548 ^ n6466;
  assign n6550 = ~n6547 & n6549;
  assign n6551 = n6509 ^ n3738;
  assign n6552 = n6551 ^ n6464;
  assign n6553 = ~n6550 & ~n6552;
  assign n6554 = ~n6525 & ~n6553;
  assign n6649 = n6556 ^ n6554;
  assign n6595 = n6553 ^ n6525;
  assign n6596 = n6595 ^ x197;
  assign n6597 = n6552 ^ n6550;
  assign n6598 = n6597 ^ x198;
  assign n6599 = n6549 ^ n6547;
  assign n6600 = n6599 ^ x199;
  assign n6601 = n6546 ^ n6544;
  assign n6602 = n6601 ^ x200;
  assign n6603 = n6543 ^ n6541;
  assign n6604 = n6603 ^ x201;
  assign n6605 = n6540 ^ n6527;
  assign n6606 = n6605 ^ x202;
  assign n6607 = n6539 ^ n6537;
  assign n6608 = n6607 ^ x203;
  assign n6609 = n6536 ^ n6529;
  assign n6610 = n6609 ^ x204;
  assign n6611 = n6535 ^ n6531;
  assign n6612 = n6611 ^ x205;
  assign n6613 = n6534 ^ n6533;
  assign n6614 = n6613 ^ x206;
  assign n6202 = n6199 ^ n6197;
  assign n6203 = n6202 ^ x208;
  assign n6204 = n6196 ^ n6172;
  assign n6205 = n6204 ^ x209;
  assign n6206 = n6195 ^ n6193;
  assign n6207 = n6206 ^ x210;
  assign n6208 = n6192 ^ n6191;
  assign n6209 = n6208 ^ x211;
  assign n6210 = n6190 ^ n6174;
  assign n6211 = n6210 ^ x212;
  assign n6212 = n6189 ^ n6188;
  assign n6213 = n6212 ^ x213;
  assign n6214 = n6187 ^ n6176;
  assign n6215 = n6214 ^ x214;
  assign n6216 = n6186 ^ n6185;
  assign n6217 = n6216 ^ x215;
  assign n6218 = n6184 ^ n6182;
  assign n6219 = n6218 ^ x216;
  assign n6220 = n6181 ^ n6177;
  assign n6221 = n6220 ^ x217;
  assign n6222 = n6180 ^ n6179;
  assign n6223 = n6222 ^ x218;
  assign n5988 = n5987 ^ n5948;
  assign n5989 = n5988 ^ x219;
  assign n5932 = n5931 ^ n5894;
  assign n5933 = n5932 ^ x220;
  assign n5934 = n5893 ^ n5890;
  assign n5935 = n5934 ^ x221;
  assign n5936 = x223 & ~n5892;
  assign n5937 = n5936 ^ x222;
  assign n5938 = n5892 ^ n5891;
  assign n5939 = n5938 ^ n5936;
  assign n5940 = n5937 & n5939;
  assign n5941 = n5940 ^ x222;
  assign n5942 = n5941 ^ n5934;
  assign n5943 = ~n5935 & n5942;
  assign n5944 = n5943 ^ x221;
  assign n5945 = n5944 ^ n5932;
  assign n5946 = n5933 & ~n5945;
  assign n5947 = n5946 ^ x220;
  assign n6224 = n5988 ^ n5947;
  assign n6225 = n5989 & ~n6224;
  assign n6226 = n6225 ^ x219;
  assign n6227 = n6226 ^ n6222;
  assign n6228 = n6223 & ~n6227;
  assign n6229 = n6228 ^ x218;
  assign n6230 = n6229 ^ n6220;
  assign n6231 = ~n6221 & n6230;
  assign n6232 = n6231 ^ x217;
  assign n6233 = n6232 ^ n6218;
  assign n6234 = ~n6219 & n6233;
  assign n6235 = n6234 ^ x216;
  assign n6236 = n6235 ^ n6216;
  assign n6237 = ~n6217 & n6236;
  assign n6238 = n6237 ^ x215;
  assign n6239 = n6238 ^ n6214;
  assign n6240 = n6215 & ~n6239;
  assign n6241 = n6240 ^ x214;
  assign n6242 = n6241 ^ n6212;
  assign n6243 = n6213 & ~n6242;
  assign n6244 = n6243 ^ x213;
  assign n6245 = n6244 ^ n6210;
  assign n6246 = n6211 & ~n6245;
  assign n6247 = n6246 ^ x212;
  assign n6248 = n6247 ^ n6208;
  assign n6249 = n6209 & ~n6248;
  assign n6250 = n6249 ^ x211;
  assign n6251 = n6250 ^ n6206;
  assign n6252 = ~n6207 & n6251;
  assign n6253 = n6252 ^ x210;
  assign n6254 = n6253 ^ n6204;
  assign n6255 = n6205 & ~n6254;
  assign n6256 = n6255 ^ x209;
  assign n6257 = n6256 ^ n6202;
  assign n6258 = ~n6203 & n6257;
  assign n6259 = n6258 ^ x208;
  assign n6201 = n6200 ^ n6171;
  assign n6260 = n6259 ^ n6201;
  assign n6615 = n6201 ^ x207;
  assign n6616 = n6260 & ~n6615;
  assign n6617 = n6616 ^ x207;
  assign n6618 = n6617 ^ n6613;
  assign n6619 = ~n6614 & n6618;
  assign n6620 = n6619 ^ x206;
  assign n6621 = n6620 ^ n6611;
  assign n6622 = n6612 & ~n6621;
  assign n6623 = n6622 ^ x205;
  assign n6624 = n6623 ^ n6609;
  assign n6625 = ~n6610 & n6624;
  assign n6626 = n6625 ^ x204;
  assign n6627 = n6626 ^ n6607;
  assign n6628 = ~n6608 & n6627;
  assign n6629 = n6628 ^ x203;
  assign n6630 = n6629 ^ n6605;
  assign n6631 = ~n6606 & n6630;
  assign n6632 = n6631 ^ x202;
  assign n6633 = n6632 ^ n6603;
  assign n6634 = ~n6604 & n6633;
  assign n6635 = n6634 ^ x201;
  assign n6636 = n6635 ^ n6601;
  assign n6637 = n6602 & ~n6636;
  assign n6638 = n6637 ^ x200;
  assign n6639 = n6638 ^ n6599;
  assign n6640 = ~n6600 & n6639;
  assign n6641 = n6640 ^ x199;
  assign n6642 = n6641 ^ n6597;
  assign n6643 = ~n6598 & n6642;
  assign n6644 = n6643 ^ x198;
  assign n6645 = n6644 ^ n6595;
  assign n6646 = n6596 & ~n6645;
  assign n6647 = n6646 ^ x197;
  assign n6648 = n6647 ^ x196;
  assign n6687 = n6649 ^ n6648;
  assign n6808 = n6690 ^ n6687;
  assign n6904 = n6808 ^ n3794;
  assign n7120 = x255 & n6904;
  assign n7121 = n7120 ^ x254;
  assign n6691 = ~n6687 & ~n6690;
  assign n6683 = n4942 ^ n4499;
  assign n6684 = n6048 & ~n6683;
  assign n6685 = n6684 ^ n4499;
  assign n6811 = n6691 ^ n6685;
  assign n6650 = n6649 ^ n6647;
  assign n6651 = n6648 & n6650;
  assign n6652 = n6651 ^ x196;
  assign n6459 = n6458 ^ n3711;
  assign n6516 = n6515 ^ n6458;
  assign n6517 = n6459 & ~n6516;
  assign n6518 = n6517 ^ n3711;
  assign n6444 = n6443 ^ n6366;
  assign n6445 = n6370 & n6444;
  assign n6446 = n6445 ^ n6369;
  assign n6361 = n4631 ^ n4096;
  assign n6362 = ~n5218 & n6361;
  assign n6363 = n6362 ^ n4096;
  assign n6455 = n6446 ^ n6363;
  assign n6359 = n5763 ^ x168;
  assign n6360 = n6359 ^ n5642;
  assign n6456 = n6455 ^ n6360;
  assign n6457 = n6456 ^ n3708;
  assign n6558 = n6518 ^ n6457;
  assign n6557 = ~n6554 & ~n6556;
  assign n6593 = n6558 ^ n6557;
  assign n6594 = n6593 ^ x195;
  assign n6682 = n6652 ^ n6594;
  assign n6812 = n6811 ^ n6682;
  assign n6809 = ~n3794 & n6808;
  assign n6810 = n6809 ^ n3790;
  assign n6905 = n6812 ^ n6810;
  assign n7122 = n6905 ^ n6904;
  assign n7123 = n7122 ^ n7120;
  assign n7124 = n7121 & n7123;
  assign n7125 = n7124 ^ x254;
  assign n6813 = n6812 ^ n6809;
  assign n6814 = n6810 & ~n6813;
  assign n6815 = n6814 ^ n3790;
  assign n6907 = n6815 ^ n3786;
  assign n6686 = n6685 ^ n6682;
  assign n6692 = n6691 ^ n6682;
  assign n6693 = ~n6686 & ~n6692;
  assign n6694 = n6693 ^ n6691;
  assign n6678 = n4940 ^ n4676;
  assign n6679 = n6043 & n6678;
  assign n6680 = n6679 ^ n4676;
  assign n6559 = n6557 & n6558;
  assign n6519 = n6518 ^ n6456;
  assign n6520 = ~n6457 & ~n6519;
  assign n6521 = n6520 ^ n3708;
  assign n6522 = n6521 ^ n3722;
  assign n6451 = n4626 ^ n4093;
  assign n6452 = ~n5216 & ~n6451;
  assign n6453 = n6452 ^ n4093;
  assign n6364 = n6363 ^ n6360;
  assign n6447 = n6446 ^ n6360;
  assign n6448 = ~n6364 & ~n6447;
  assign n6449 = n6448 ^ n6363;
  assign n6358 = n5766 ^ n5641;
  assign n6450 = n6449 ^ n6358;
  assign n6454 = n6453 ^ n6450;
  assign n6523 = n6522 ^ n6454;
  assign n6657 = n6559 ^ n6523;
  assign n6653 = n6652 ^ n6593;
  assign n6654 = ~n6594 & n6653;
  assign n6655 = n6654 ^ x195;
  assign n6656 = n6655 ^ x194;
  assign n6677 = n6657 ^ n6656;
  assign n6681 = n6680 ^ n6677;
  assign n6806 = n6694 ^ n6681;
  assign n6908 = n6907 ^ n6806;
  assign n6906 = ~n6904 & n6905;
  assign n7118 = n6908 ^ n6906;
  assign n7119 = n7118 ^ x253;
  assign n7370 = n7125 ^ n7119;
  assign n6321 = n6232 ^ x216;
  assign n6322 = n6321 ^ n6218;
  assign n7366 = n6088 ^ n4915;
  assign n7367 = ~n6322 & n7366;
  assign n7368 = n7367 ^ n4915;
  assign n7445 = n7370 ^ n7368;
  assign n6324 = n6229 ^ n6221;
  assign n7307 = n6014 ^ n4920;
  assign n7308 = ~n6324 & ~n7307;
  assign n7309 = n7308 ^ n4920;
  assign n7306 = n7122 ^ n7121;
  assign n7310 = n7309 ^ n7306;
  assign n6329 = n6226 ^ x218;
  assign n6330 = n6329 ^ n6222;
  assign n7268 = n6019 ^ n4925;
  assign n7269 = n6330 & ~n7268;
  assign n7270 = n7269 ^ n4925;
  assign n7267 = n6904 ^ x255;
  assign n7271 = n7270 ^ n7267;
  assign n7020 = n6635 ^ x200;
  assign n7021 = n7020 ^ n6601;
  assign n7008 = n6632 ^ n6604;
  assign n7004 = n5216 ^ n4654;
  assign n7005 = ~n5796 & n7004;
  assign n7006 = n7005 ^ n4654;
  assign n7015 = n7008 ^ n7006;
  assign n6990 = n6629 ^ x202;
  assign n6991 = n6990 ^ n6605;
  assign n6578 = n5772 ^ n5637;
  assign n6986 = n5218 ^ n4640;
  assign n6987 = ~n6578 & ~n6986;
  assign n6988 = n6987 ^ n4640;
  assign n7000 = n6991 ^ n6988;
  assign n6973 = n6626 ^ n6608;
  assign n6561 = n5769 ^ x166;
  assign n6562 = n6561 ^ n5638;
  assign n6970 = n5223 ^ n4645;
  assign n6971 = ~n6562 & n6970;
  assign n6972 = n6971 ^ n4645;
  assign n6974 = n6973 ^ n6972;
  assign n6957 = n6623 ^ x204;
  assign n6958 = n6957 ^ n6609;
  assign n6954 = n5962 ^ n5192;
  assign n6955 = ~n6358 & ~n6954;
  assign n6956 = n6955 ^ n5192;
  assign n6959 = n6958 ^ n6956;
  assign n6885 = n6620 ^ n6612;
  assign n6882 = n5916 ^ n5099;
  assign n6883 = ~n6360 & ~n6882;
  assign n6884 = n6883 ^ n5099;
  assign n6886 = n6885 ^ n6884;
  assign n6757 = n5873 ^ n4450;
  assign n6758 = ~n6366 & n6757;
  assign n6759 = n6758 ^ n4450;
  assign n6755 = n6617 ^ x206;
  assign n6756 = n6755 ^ n6613;
  assign n6760 = n6759 ^ n6756;
  assign n6261 = n6260 ^ x207;
  assign n6005 = n5842 ^ n5063;
  assign n6006 = n6004 & n6005;
  assign n6007 = n6006 ^ n5063;
  assign n6262 = n6261 ^ n6007;
  assign n6268 = n6256 ^ x208;
  assign n6269 = n6268 ^ n6202;
  assign n6265 = n5789 ^ n4969;
  assign n6266 = n6264 & ~n6265;
  assign n6267 = n6266 ^ n4969;
  assign n6270 = n6269 ^ n6267;
  assign n6275 = n6253 ^ n6205;
  assign n6272 = n5546 ^ n4973;
  assign n6273 = n6271 & n6272;
  assign n6274 = n6273 ^ n4973;
  assign n6276 = n6275 ^ n6274;
  assign n6281 = n6250 ^ x210;
  assign n6282 = n6281 ^ n6206;
  assign n6278 = n5379 ^ n4978;
  assign n6279 = ~n6277 & ~n6278;
  assign n6280 = n6279 ^ n4978;
  assign n6283 = n6282 ^ n6280;
  assign n6288 = n6247 ^ n6209;
  assign n6285 = n4987 ^ n4899;
  assign n6286 = n6284 & ~n6285;
  assign n6287 = n6286 ^ n4987;
  assign n6289 = n6288 ^ n6287;
  assign n6294 = n6244 ^ x212;
  assign n6295 = n6294 ^ n6210;
  assign n6291 = n5330 ^ n4989;
  assign n6292 = ~n6290 & n6291;
  assign n6293 = n6292 ^ n4989;
  assign n6296 = n6295 ^ n6293;
  assign n6301 = n6241 ^ n6213;
  assign n6298 = n5325 ^ n4998;
  assign n6299 = ~n6297 & ~n6298;
  assign n6300 = n6299 ^ n4998;
  assign n6302 = n6301 ^ n6300;
  assign n6307 = n6238 ^ n6215;
  assign n6304 = n5321 ^ n4999;
  assign n6305 = n6303 & n6304;
  assign n6306 = n6305 ^ n4999;
  assign n6308 = n6307 ^ n6306;
  assign n6313 = n6235 ^ x215;
  assign n6314 = n6313 ^ n6216;
  assign n6310 = n5311 ^ n4901;
  assign n6311 = ~n6309 & n6310;
  assign n6312 = n6311 ^ n4901;
  assign n6315 = n6314 ^ n6312;
  assign n6318 = n5303 ^ n4891;
  assign n6319 = n6317 & ~n6318;
  assign n6320 = n6319 ^ n4891;
  assign n6323 = n6322 ^ n6320;
  assign n6325 = n5278 ^ n4713;
  assign n6326 = n6168 & n6325;
  assign n6327 = n6326 ^ n4713;
  assign n6328 = n6327 ^ n6324;
  assign n6331 = n5283 ^ n4456;
  assign n6332 = n6098 & ~n6331;
  assign n6333 = n6332 ^ n4456;
  assign n6334 = n6333 ^ n6330;
  assign n6335 = n5291 ^ n4469;
  assign n6336 = ~n6088 & ~n6335;
  assign n6337 = n6336 ^ n4469;
  assign n5990 = n5989 ^ n5947;
  assign n6338 = n6337 ^ n5990;
  assign n6339 = n4907 ^ n4471;
  assign n6340 = n6014 & ~n6339;
  assign n6341 = n6340 ^ n4471;
  assign n5996 = n5944 ^ x220;
  assign n5997 = n5996 ^ n5932;
  assign n6342 = n6341 ^ n5997;
  assign n6344 = n4915 ^ n4478;
  assign n6345 = n6019 & ~n6344;
  assign n6346 = n6345 ^ n4478;
  assign n6343 = n5941 ^ n5935;
  assign n6347 = n6346 ^ n6343;
  assign n6351 = n5938 ^ n5937;
  assign n6348 = n4920 ^ n4483;
  assign n6349 = ~n5992 & ~n6348;
  assign n6350 = n6349 ^ n4483;
  assign n6352 = n6351 ^ n6350;
  assign n6356 = n5892 ^ x223;
  assign n6353 = n4925 ^ n4488;
  assign n6354 = n6000 & ~n6353;
  assign n6355 = n6354 ^ n4488;
  assign n6357 = n6356 ^ n6355;
  assign n6668 = n4930 ^ n4687;
  assign n6669 = n6032 & ~n6668;
  assign n6670 = n6669 ^ n4687;
  assign n6658 = n6657 ^ n6655;
  assign n6659 = n6656 & ~n6658;
  assign n6660 = n6659 ^ x194;
  assign n6661 = n6660 ^ x193;
  assign n6571 = n6454 ^ n3722;
  assign n6572 = n6521 ^ n6454;
  assign n6573 = n6571 & n6572;
  assign n6574 = n6573 ^ n3722;
  assign n6567 = n4518 ^ n3804;
  assign n6568 = ~n5211 & ~n6567;
  assign n6569 = n6568 ^ n3804;
  assign n6563 = n6453 ^ n6358;
  assign n6564 = n6450 & n6563;
  assign n6565 = n6564 ^ n6453;
  assign n6566 = n6565 ^ n6562;
  assign n6570 = n6569 ^ n6566;
  assign n6575 = n6574 ^ n6570;
  assign n6576 = n6575 ^ n3499;
  assign n6560 = ~n6523 & ~n6559;
  assign n6662 = n6576 ^ n6560;
  assign n6663 = n6662 ^ n6660;
  assign n6664 = n6661 & ~n6663;
  assign n6665 = n6664 ^ x193;
  assign n6666 = n6665 ^ x192;
  assign n6589 = n6570 ^ n3499;
  assign n6590 = ~n6575 & ~n6589;
  assign n6591 = n6590 ^ n3499;
  assign n6583 = n6569 ^ n6562;
  assign n6584 = ~n6566 & ~n6583;
  assign n6585 = n6584 ^ n6569;
  assign n6579 = n4513 ^ n3799;
  assign n6580 = n5203 & ~n6579;
  assign n6581 = n6580 ^ n3799;
  assign n6582 = n6581 ^ n6578;
  assign n6586 = n6585 ^ n6582;
  assign n6587 = n6586 ^ n3498;
  assign n6577 = ~n6560 & n6576;
  assign n6588 = n6587 ^ n6577;
  assign n6592 = n6591 ^ n6588;
  assign n6667 = n6666 ^ n6592;
  assign n6671 = n6670 ^ n6667;
  assign n6673 = n4935 ^ n4496;
  assign n6674 = ~n6037 & ~n6673;
  assign n6675 = n6674 ^ n4496;
  assign n6672 = n6662 ^ n6661;
  assign n6676 = n6675 ^ n6672;
  assign n6695 = n6694 ^ n6677;
  assign n6696 = ~n6681 & ~n6695;
  assign n6697 = n6696 ^ n6680;
  assign n6698 = n6697 ^ n6672;
  assign n6699 = n6676 & n6698;
  assign n6700 = n6699 ^ n6675;
  assign n6701 = n6700 ^ n6667;
  assign n6702 = n6671 & n6701;
  assign n6703 = n6702 ^ n6670;
  assign n6704 = n6703 ^ n6356;
  assign n6705 = ~n6357 & ~n6704;
  assign n6706 = n6705 ^ n6355;
  assign n6707 = n6706 ^ n6351;
  assign n6708 = ~n6352 & n6707;
  assign n6709 = n6708 ^ n6350;
  assign n6710 = n6709 ^ n6343;
  assign n6711 = ~n6347 & n6710;
  assign n6712 = n6711 ^ n6346;
  assign n6713 = n6712 ^ n5997;
  assign n6714 = ~n6342 & ~n6713;
  assign n6715 = n6714 ^ n6341;
  assign n6716 = n6715 ^ n5990;
  assign n6717 = ~n6338 & n6716;
  assign n6718 = n6717 ^ n6337;
  assign n6719 = n6718 ^ n6330;
  assign n6720 = n6334 & n6719;
  assign n6721 = n6720 ^ n6333;
  assign n6722 = n6721 ^ n6324;
  assign n6723 = n6328 & n6722;
  assign n6724 = n6723 ^ n6327;
  assign n6725 = n6724 ^ n6322;
  assign n6726 = n6323 & ~n6725;
  assign n6727 = n6726 ^ n6320;
  assign n6728 = n6727 ^ n6314;
  assign n6729 = ~n6315 & ~n6728;
  assign n6730 = n6729 ^ n6312;
  assign n6731 = n6730 ^ n6307;
  assign n6732 = ~n6308 & ~n6731;
  assign n6733 = n6732 ^ n6306;
  assign n6734 = n6733 ^ n6301;
  assign n6735 = n6302 & n6734;
  assign n6736 = n6735 ^ n6300;
  assign n6737 = n6736 ^ n6295;
  assign n6738 = ~n6296 & ~n6737;
  assign n6739 = n6738 ^ n6293;
  assign n6740 = n6739 ^ n6288;
  assign n6741 = ~n6289 & n6740;
  assign n6742 = n6741 ^ n6287;
  assign n6743 = n6742 ^ n6282;
  assign n6744 = ~n6283 & ~n6743;
  assign n6745 = n6744 ^ n6280;
  assign n6746 = n6745 ^ n6275;
  assign n6747 = n6276 & ~n6746;
  assign n6748 = n6747 ^ n6274;
  assign n6749 = n6748 ^ n6269;
  assign n6750 = ~n6270 & n6749;
  assign n6751 = n6750 ^ n6267;
  assign n6752 = n6751 ^ n6261;
  assign n6753 = ~n6262 & n6752;
  assign n6754 = n6753 ^ n6007;
  assign n6879 = n6756 ^ n6754;
  assign n6880 = ~n6760 & n6879;
  assign n6881 = n6880 ^ n6759;
  assign n6951 = n6885 ^ n6881;
  assign n6952 = ~n6886 & ~n6951;
  assign n6953 = n6952 ^ n6884;
  assign n6967 = n6958 ^ n6953;
  assign n6968 = n6959 & ~n6967;
  assign n6969 = n6968 ^ n6956;
  assign n6983 = n6973 ^ n6969;
  assign n6984 = ~n6974 & ~n6983;
  assign n6985 = n6984 ^ n6972;
  assign n7001 = n6991 ^ n6985;
  assign n7002 = ~n7000 & n7001;
  assign n7003 = n7002 ^ n6988;
  assign n7016 = n7008 ^ n7003;
  assign n7017 = n7015 & n7016;
  assign n7018 = n7017 ^ n7006;
  assign n7012 = n5211 ^ n4631;
  assign n7013 = ~n5852 & ~n7012;
  assign n7014 = n7013 ^ n4631;
  assign n7019 = n7018 ^ n7014;
  assign n7022 = n7021 ^ n7019;
  assign n7041 = n7022 ^ n4096;
  assign n7007 = n7006 ^ n7003;
  assign n7009 = n7008 ^ n7007;
  assign n7023 = n7009 ^ n4098;
  assign n6989 = n6988 ^ n6985;
  assign n6992 = n6991 ^ n6989;
  assign n6995 = n6992 ^ n4107;
  assign n6975 = n6974 ^ n6969;
  assign n6976 = n6975 ^ n4102;
  assign n6960 = n6959 ^ n6953;
  assign n6961 = n6960 ^ n4451;
  assign n6887 = n6886 ^ n6881;
  assign n6888 = n6887 ^ n4523;
  assign n6761 = n6760 ^ n6754;
  assign n6762 = n6761 ^ n4526;
  assign n6763 = n6751 ^ n6262;
  assign n6764 = n6763 ^ n4528;
  assign n6765 = n6748 ^ n6270;
  assign n6766 = n6765 ^ n4531;
  assign n6767 = n6745 ^ n6276;
  assign n6768 = n6767 ^ n4535;
  assign n6769 = n6742 ^ n6283;
  assign n6770 = n6769 ^ n4538;
  assign n6771 = n6739 ^ n6289;
  assign n6772 = n6771 ^ n4444;
  assign n6773 = n6736 ^ n6296;
  assign n6774 = n6773 ^ n4397;
  assign n6775 = n6733 ^ n6300;
  assign n6776 = n6775 ^ n6301;
  assign n6777 = n6776 ^ n4383;
  assign n6778 = n6730 ^ n6306;
  assign n6779 = n6778 ^ n6307;
  assign n6780 = n6779 ^ n4357;
  assign n6781 = n6727 ^ n6312;
  assign n6782 = n6781 ^ n6314;
  assign n6783 = n6782 ^ n4340;
  assign n6784 = n6724 ^ n6320;
  assign n6785 = n6784 ^ n6322;
  assign n6786 = n6785 ^ n4323;
  assign n6787 = n6721 ^ n6327;
  assign n6788 = n6787 ^ n6324;
  assign n6789 = n6788 ^ n4302;
  assign n6790 = n6718 ^ n6334;
  assign n6791 = n6790 ^ n4305;
  assign n6792 = n6715 ^ n6338;
  assign n6793 = n6792 ^ n4309;
  assign n6794 = n6712 ^ n6342;
  assign n6795 = n6794 ^ n4213;
  assign n6796 = n6709 ^ n6347;
  assign n6797 = n6796 ^ n4204;
  assign n6798 = n6706 ^ n6352;
  assign n6799 = n6798 ^ n4194;
  assign n6800 = n6703 ^ n6357;
  assign n6801 = n6800 ^ n4142;
  assign n6802 = n6700 ^ n6671;
  assign n6803 = n6802 ^ n3776;
  assign n6804 = n6697 ^ n6676;
  assign n6805 = n6804 ^ n3781;
  assign n6807 = n6806 ^ n3786;
  assign n6816 = n6815 ^ n6806;
  assign n6817 = ~n6807 & n6816;
  assign n6818 = n6817 ^ n3786;
  assign n6819 = n6818 ^ n6804;
  assign n6820 = n6805 & n6819;
  assign n6821 = n6820 ^ n3781;
  assign n6822 = n6821 ^ n6802;
  assign n6823 = n6803 & n6822;
  assign n6824 = n6823 ^ n3776;
  assign n6825 = n6824 ^ n6800;
  assign n6826 = ~n6801 & ~n6825;
  assign n6827 = n6826 ^ n4142;
  assign n6828 = n6827 ^ n6798;
  assign n6829 = ~n6799 & ~n6828;
  assign n6830 = n6829 ^ n4194;
  assign n6831 = n6830 ^ n6796;
  assign n6832 = ~n6797 & n6831;
  assign n6833 = n6832 ^ n4204;
  assign n6834 = n6833 ^ n6794;
  assign n6835 = ~n6795 & n6834;
  assign n6836 = n6835 ^ n4213;
  assign n6837 = n6836 ^ n6792;
  assign n6838 = ~n6793 & ~n6837;
  assign n6839 = n6838 ^ n4309;
  assign n6840 = n6839 ^ n6790;
  assign n6841 = ~n6791 & ~n6840;
  assign n6842 = n6841 ^ n4305;
  assign n6843 = n6842 ^ n6788;
  assign n6844 = n6789 & ~n6843;
  assign n6845 = n6844 ^ n4302;
  assign n6846 = n6845 ^ n6785;
  assign n6847 = n6786 & n6846;
  assign n6848 = n6847 ^ n4323;
  assign n6849 = n6848 ^ n6782;
  assign n6850 = ~n6783 & n6849;
  assign n6851 = n6850 ^ n4340;
  assign n6852 = n6851 ^ n6779;
  assign n6853 = n6780 & ~n6852;
  assign n6854 = n6853 ^ n4357;
  assign n6855 = n6854 ^ n6776;
  assign n6856 = ~n6777 & ~n6855;
  assign n6857 = n6856 ^ n4383;
  assign n6858 = n6857 ^ n6773;
  assign n6859 = n6774 & n6858;
  assign n6860 = n6859 ^ n4397;
  assign n6861 = n6860 ^ n6771;
  assign n6862 = n6772 & n6861;
  assign n6863 = n6862 ^ n4444;
  assign n6864 = n6863 ^ n6769;
  assign n6865 = ~n6770 & ~n6864;
  assign n6866 = n6865 ^ n4538;
  assign n6867 = n6866 ^ n6767;
  assign n6868 = ~n6768 & n6867;
  assign n6869 = n6868 ^ n4535;
  assign n6870 = n6869 ^ n6765;
  assign n6871 = n6766 & ~n6870;
  assign n6872 = n6871 ^ n4531;
  assign n6873 = n6872 ^ n6763;
  assign n6874 = ~n6764 & ~n6873;
  assign n6875 = n6874 ^ n4528;
  assign n6876 = n6875 ^ n6761;
  assign n6877 = n6762 & n6876;
  assign n6878 = n6877 ^ n4526;
  assign n6948 = n6887 ^ n6878;
  assign n6949 = n6888 & ~n6948;
  assign n6950 = n6949 ^ n4523;
  assign n6964 = n6960 ^ n6950;
  assign n6965 = n6961 & ~n6964;
  assign n6966 = n6965 ^ n4451;
  assign n6979 = n6975 ^ n6966;
  assign n6980 = n6976 & n6979;
  assign n6981 = n6980 ^ n4102;
  assign n6996 = n6992 ^ n6981;
  assign n6997 = ~n6995 & n6996;
  assign n6998 = n6997 ^ n4107;
  assign n7024 = n7009 ^ n6998;
  assign n7025 = ~n7023 & ~n7024;
  assign n7026 = n7025 ^ n4098;
  assign n7042 = n7026 ^ n7022;
  assign n7043 = ~n7041 & ~n7042;
  assign n7044 = n7043 ^ n4096;
  assign n7045 = n7044 ^ n4093;
  assign n7037 = n5203 ^ n4626;
  assign n7038 = ~n5886 & n7037;
  assign n7039 = n7038 ^ n4626;
  assign n7034 = n6638 ^ x199;
  assign n7035 = n7034 ^ n6599;
  assign n7030 = n7021 ^ n7014;
  assign n7031 = n7021 ^ n7018;
  assign n7032 = n7030 & n7031;
  assign n7033 = n7032 ^ n7014;
  assign n7036 = n7035 ^ n7033;
  assign n7040 = n7039 ^ n7036;
  assign n7046 = n7045 ^ n7040;
  assign n6889 = n6888 ^ n6878;
  assign n6890 = n6863 ^ n4538;
  assign n6891 = n6890 ^ n6769;
  assign n6892 = n6857 ^ n6774;
  assign n6893 = n6848 ^ n4340;
  assign n6894 = n6893 ^ n6782;
  assign n6895 = n6842 ^ n6789;
  assign n6896 = n6833 ^ n4213;
  assign n6897 = n6896 ^ n6794;
  assign n6898 = n6830 ^ n6797;
  assign n6899 = n6827 ^ n4194;
  assign n6900 = n6899 ^ n6798;
  assign n6901 = n6821 ^ n3776;
  assign n6902 = n6901 ^ n6802;
  assign n6903 = n6818 ^ n6805;
  assign n6909 = n6906 & ~n6908;
  assign n6910 = ~n6903 & ~n6909;
  assign n6911 = n6902 & n6910;
  assign n6912 = n6824 ^ n6801;
  assign n6913 = ~n6911 & ~n6912;
  assign n6914 = n6900 & n6913;
  assign n6915 = n6898 & ~n6914;
  assign n6916 = n6897 & n6915;
  assign n6917 = n6836 ^ n6793;
  assign n6918 = ~n6916 & ~n6917;
  assign n6919 = n6839 ^ n4305;
  assign n6920 = n6919 ^ n6790;
  assign n6921 = n6918 & n6920;
  assign n6922 = ~n6895 & ~n6921;
  assign n6923 = n6845 ^ n4323;
  assign n6924 = n6923 ^ n6785;
  assign n6925 = n6922 & ~n6924;
  assign n6926 = ~n6894 & n6925;
  assign n6927 = n6851 ^ n4357;
  assign n6928 = n6927 ^ n6779;
  assign n6929 = n6926 & n6928;
  assign n6930 = n6854 ^ n4383;
  assign n6931 = n6930 ^ n6776;
  assign n6932 = ~n6929 & n6931;
  assign n6933 = n6892 & n6932;
  assign n6934 = n6860 ^ n6772;
  assign n6935 = ~n6933 & n6934;
  assign n6936 = ~n6891 & ~n6935;
  assign n6937 = n6866 ^ n6768;
  assign n6938 = n6936 & n6937;
  assign n6939 = n6869 ^ n4531;
  assign n6940 = n6939 ^ n6765;
  assign n6941 = n6938 & ~n6940;
  assign n6942 = n6872 ^ n6764;
  assign n6943 = n6941 & n6942;
  assign n6944 = n6875 ^ n4526;
  assign n6945 = n6944 ^ n6761;
  assign n6946 = n6943 & n6945;
  assign n6947 = n6889 & ~n6946;
  assign n6962 = n6961 ^ n6950;
  assign n6963 = ~n6947 & ~n6962;
  assign n6977 = n6976 ^ n6966;
  assign n6978 = ~n6963 & n6977;
  assign n6982 = n6981 ^ n4107;
  assign n6993 = n6992 ^ n6982;
  assign n6994 = ~n6978 & ~n6993;
  assign n6999 = n6998 ^ n4098;
  assign n7010 = n7009 ^ n6999;
  assign n7011 = ~n6994 & n7010;
  assign n7027 = n7026 ^ n4096;
  assign n7028 = n7027 ^ n7022;
  assign n7029 = n7011 & ~n7028;
  assign n7065 = n7046 ^ n7029;
  assign n7066 = n7065 ^ x226;
  assign n7067 = n7028 ^ n7011;
  assign n7068 = n7067 ^ x227;
  assign n7069 = n7010 ^ n6994;
  assign n7070 = n7069 ^ x228;
  assign n7071 = n6993 ^ n6978;
  assign n7072 = n7071 ^ x229;
  assign n7073 = n6977 ^ n6963;
  assign n7074 = n7073 ^ x230;
  assign n7075 = n6962 ^ n6947;
  assign n7076 = n7075 ^ x231;
  assign n7077 = n6946 ^ n6889;
  assign n7078 = n7077 ^ x232;
  assign n7079 = n6945 ^ n6943;
  assign n7080 = n7079 ^ x233;
  assign n7081 = n6942 ^ n6941;
  assign n7082 = n7081 ^ x234;
  assign n7083 = n6940 ^ n6938;
  assign n7084 = n7083 ^ x235;
  assign n7085 = n6937 ^ n6936;
  assign n7086 = n7085 ^ x236;
  assign n7087 = n6935 ^ n6891;
  assign n7088 = n7087 ^ x237;
  assign n7089 = n6934 ^ n6933;
  assign n7090 = n7089 ^ x238;
  assign n7092 = n6931 ^ n6929;
  assign n7093 = n7092 ^ x240;
  assign n7094 = n6928 ^ n6926;
  assign n7095 = n7094 ^ x241;
  assign n7096 = n6925 ^ n6894;
  assign n7097 = n7096 ^ x242;
  assign n7098 = n6924 ^ n6922;
  assign n7099 = n7098 ^ x243;
  assign n7100 = n6921 ^ n6895;
  assign n7101 = n7100 ^ x244;
  assign n7102 = n6920 ^ n6918;
  assign n7103 = n7102 ^ x245;
  assign n7104 = n6917 ^ n6916;
  assign n7105 = n7104 ^ x246;
  assign n7106 = n6915 ^ n6897;
  assign n7107 = n7106 ^ x247;
  assign n7108 = n6914 ^ n6898;
  assign n7109 = n7108 ^ x248;
  assign n7110 = n6913 ^ n6900;
  assign n7111 = n7110 ^ x249;
  assign n7112 = n6912 ^ n6911;
  assign n7113 = n7112 ^ x250;
  assign n7114 = n6910 ^ n6902;
  assign n7115 = n7114 ^ x251;
  assign n7116 = n6909 ^ n6903;
  assign n7117 = n7116 ^ x252;
  assign n7126 = n7125 ^ n7118;
  assign n7127 = ~n7119 & n7126;
  assign n7128 = n7127 ^ x253;
  assign n7129 = n7128 ^ n7116;
  assign n7130 = ~n7117 & n7129;
  assign n7131 = n7130 ^ x252;
  assign n7132 = n7131 ^ n7114;
  assign n7133 = ~n7115 & n7132;
  assign n7134 = n7133 ^ x251;
  assign n7135 = n7134 ^ n7112;
  assign n7136 = n7113 & ~n7135;
  assign n7137 = n7136 ^ x250;
  assign n7138 = n7137 ^ n7110;
  assign n7139 = n7111 & ~n7138;
  assign n7140 = n7139 ^ x249;
  assign n7141 = n7140 ^ n7108;
  assign n7142 = n7109 & ~n7141;
  assign n7143 = n7142 ^ x248;
  assign n7144 = n7143 ^ n7106;
  assign n7145 = ~n7107 & n7144;
  assign n7146 = n7145 ^ x247;
  assign n7147 = n7146 ^ n7104;
  assign n7148 = n7105 & ~n7147;
  assign n7149 = n7148 ^ x246;
  assign n7150 = n7149 ^ n7102;
  assign n7151 = n7103 & ~n7150;
  assign n7152 = n7151 ^ x245;
  assign n7153 = n7152 ^ n7100;
  assign n7154 = ~n7101 & n7153;
  assign n7155 = n7154 ^ x244;
  assign n7156 = n7155 ^ n7098;
  assign n7157 = n7099 & ~n7156;
  assign n7158 = n7157 ^ x243;
  assign n7159 = n7158 ^ n7096;
  assign n7160 = n7097 & ~n7159;
  assign n7161 = n7160 ^ x242;
  assign n7162 = n7161 ^ n7094;
  assign n7163 = ~n7095 & n7162;
  assign n7164 = n7163 ^ x241;
  assign n7165 = n7164 ^ n7092;
  assign n7166 = ~n7093 & n7165;
  assign n7167 = n7166 ^ x240;
  assign n7091 = n6932 ^ n6892;
  assign n7168 = n7167 ^ n7091;
  assign n7169 = n7091 ^ x239;
  assign n7170 = ~n7168 & n7169;
  assign n7171 = n7170 ^ x239;
  assign n7172 = n7171 ^ n7089;
  assign n7173 = n7090 & ~n7172;
  assign n7174 = n7173 ^ x238;
  assign n7175 = n7174 ^ n7087;
  assign n7176 = n7088 & ~n7175;
  assign n7177 = n7176 ^ x237;
  assign n7178 = n7177 ^ n7085;
  assign n7179 = n7086 & ~n7178;
  assign n7180 = n7179 ^ x236;
  assign n7181 = n7180 ^ n7083;
  assign n7182 = ~n7084 & n7181;
  assign n7183 = n7182 ^ x235;
  assign n7184 = n7183 ^ n7081;
  assign n7185 = n7082 & ~n7184;
  assign n7186 = n7185 ^ x234;
  assign n7187 = n7186 ^ n7079;
  assign n7188 = n7080 & ~n7187;
  assign n7189 = n7188 ^ x233;
  assign n7190 = n7189 ^ n7077;
  assign n7191 = n7078 & ~n7190;
  assign n7192 = n7191 ^ x232;
  assign n7193 = n7192 ^ n7075;
  assign n7194 = n7076 & ~n7193;
  assign n7195 = n7194 ^ x231;
  assign n7196 = n7195 ^ n7073;
  assign n7197 = n7074 & ~n7196;
  assign n7198 = n7197 ^ x230;
  assign n7199 = n7198 ^ n7071;
  assign n7200 = n7072 & ~n7199;
  assign n7201 = n7200 ^ x229;
  assign n7202 = n7201 ^ n7069;
  assign n7203 = n7070 & ~n7202;
  assign n7204 = n7203 ^ x228;
  assign n7205 = n7204 ^ n7067;
  assign n7206 = n7068 & ~n7205;
  assign n7207 = n7206 ^ x227;
  assign n7208 = n7207 ^ n7065;
  assign n7209 = ~n7066 & n7208;
  assign n7210 = n7209 ^ x226;
  assign n7211 = n7210 ^ x225;
  assign n7058 = n7040 ^ n4093;
  assign n7059 = n7044 ^ n7040;
  assign n7060 = n7058 & n7059;
  assign n7061 = n7060 ^ n4093;
  assign n7062 = n7061 ^ n3804;
  assign n7054 = n4960 ^ n4518;
  assign n7055 = n5928 & ~n7054;
  assign n7056 = n7055 ^ n4518;
  assign n7051 = n6641 ^ x198;
  assign n7052 = n7051 ^ n6597;
  assign n7048 = n7039 ^ n7035;
  assign n7049 = n7036 & ~n7048;
  assign n7050 = n7049 ^ n7039;
  assign n7053 = n7052 ^ n7050;
  assign n7057 = n7056 ^ n7053;
  assign n7063 = n7062 ^ n7057;
  assign n7047 = ~n7029 & n7046;
  assign n7064 = n7063 ^ n7047;
  assign n7212 = n7211 ^ n7064;
  assign n6001 = n6000 ^ n4935;
  assign n6002 = n5997 & ~n6001;
  assign n6003 = n6002 ^ n4935;
  assign n7213 = n7212 ^ n6003;
  assign n7216 = n6032 ^ n4940;
  assign n7217 = ~n6343 & ~n7216;
  assign n7218 = n7217 ^ n4940;
  assign n7214 = n7207 ^ x226;
  assign n7215 = n7214 ^ n7065;
  assign n7219 = n7218 ^ n7215;
  assign n7221 = n6037 ^ n4942;
  assign n7222 = ~n6351 & ~n7221;
  assign n7223 = n7222 ^ n4942;
  assign n7220 = n7204 ^ n7068;
  assign n7224 = n7223 ^ n7220;
  assign n7225 = n7201 ^ x228;
  assign n7226 = n7225 ^ n7069;
  assign n7227 = n6043 ^ n4950;
  assign n7228 = ~n6356 & n7227;
  assign n7229 = n7228 ^ n4950;
  assign n7230 = n7226 & n7229;
  assign n7231 = n7230 ^ n7220;
  assign n7232 = ~n7224 & n7231;
  assign n7233 = n7232 ^ n7230;
  assign n7234 = n7233 ^ n7215;
  assign n7235 = n7219 & n7234;
  assign n7236 = n7235 ^ n7218;
  assign n7237 = n7236 ^ n7212;
  assign n7238 = ~n7213 & n7237;
  assign n7239 = n7238 ^ n6003;
  assign n5993 = n5992 ^ n4930;
  assign n5994 = n5990 & ~n5993;
  assign n5995 = n5994 ^ n4930;
  assign n7240 = n7239 ^ n5995;
  assign n7258 = n7064 ^ x225;
  assign n7259 = n7210 ^ n7064;
  assign n7260 = n7258 & ~n7259;
  assign n7261 = n7260 ^ x225;
  assign n7262 = n7261 ^ x224;
  assign n7253 = n7057 ^ n3804;
  assign n7254 = n7061 ^ n7057;
  assign n7255 = n7253 & n7254;
  assign n7256 = n7255 ^ n3804;
  assign n7251 = ~n7047 & n7063;
  assign n7247 = n7056 ^ n7052;
  assign n7248 = n7053 & n7247;
  assign n7249 = n7248 ^ n7056;
  assign n7244 = n6644 ^ n6596;
  assign n7241 = n4955 ^ n4513;
  assign n7242 = n5980 & n7241;
  assign n7243 = n7242 ^ n4513;
  assign n7245 = n7244 ^ n7243;
  assign n7246 = n7245 ^ n3799;
  assign n7250 = n7249 ^ n7246;
  assign n7252 = n7251 ^ n7250;
  assign n7257 = n7256 ^ n7252;
  assign n7263 = n7262 ^ n7257;
  assign n7264 = n7263 ^ n7239;
  assign n7265 = ~n7240 & ~n7264;
  assign n7266 = n7265 ^ n5995;
  assign n7303 = n7267 ^ n7266;
  assign n7304 = ~n7271 & ~n7303;
  assign n7305 = n7304 ^ n7270;
  assign n7363 = n7306 ^ n7305;
  assign n7364 = n7310 & ~n7363;
  assign n7365 = n7364 ^ n7309;
  assign n7446 = n7370 ^ n7365;
  assign n7447 = n7445 & ~n7446;
  assign n7448 = n7447 ^ n7368;
  assign n7442 = n7128 ^ x252;
  assign n7443 = n7442 ^ n7116;
  assign n7439 = n6098 ^ n4907;
  assign n7440 = ~n6314 & n7439;
  assign n7441 = n7440 ^ n4907;
  assign n7444 = n7443 ^ n7441;
  assign n7520 = n7448 ^ n7444;
  assign n7521 = n7520 ^ n4471;
  assign n7369 = n7368 ^ n7365;
  assign n7371 = n7370 ^ n7369;
  assign n7372 = n7371 ^ n4478;
  assign n7311 = n7310 ^ n7305;
  assign n7359 = n7311 ^ n4483;
  assign n7272 = n7271 ^ n7266;
  assign n7273 = n7272 ^ n4488;
  assign n7274 = n7263 ^ n5995;
  assign n7275 = n7274 ^ n7239;
  assign n7276 = n7275 ^ n4687;
  assign n7277 = n7236 ^ n6003;
  assign n7278 = n7277 ^ n7212;
  assign n7279 = n7278 ^ n4496;
  assign n7280 = n7233 ^ n7219;
  assign n7281 = n7280 ^ n4676;
  assign n7282 = n7229 ^ n7226;
  assign n7283 = ~n4508 & n7282;
  assign n7284 = n7283 ^ n4499;
  assign n7285 = n7230 ^ n7223;
  assign n7286 = n7285 ^ n7220;
  assign n7287 = n7286 ^ n7283;
  assign n7288 = ~n7284 & ~n7287;
  assign n7289 = n7288 ^ n4499;
  assign n7290 = n7289 ^ n7280;
  assign n7291 = ~n7281 & n7290;
  assign n7292 = n7291 ^ n4676;
  assign n7293 = n7292 ^ n7278;
  assign n7294 = n7279 & n7293;
  assign n7295 = n7294 ^ n4496;
  assign n7296 = n7295 ^ n7275;
  assign n7297 = ~n7276 & ~n7296;
  assign n7298 = n7297 ^ n4687;
  assign n7299 = n7298 ^ n7272;
  assign n7300 = ~n7273 & ~n7299;
  assign n7301 = n7300 ^ n4488;
  assign n7360 = n7311 ^ n7301;
  assign n7361 = ~n7359 & n7360;
  assign n7362 = n7361 ^ n4483;
  assign n7522 = n7371 ^ n7362;
  assign n7523 = ~n7372 & n7522;
  assign n7524 = n7523 ^ n4478;
  assign n7525 = n7524 ^ n7520;
  assign n7526 = ~n7521 & ~n7525;
  assign n7527 = n7526 ^ n4471;
  assign n7449 = n7448 ^ n7443;
  assign n7450 = ~n7444 & ~n7449;
  assign n7451 = n7450 ^ n7441;
  assign n7435 = n6168 ^ n5291;
  assign n7436 = n6307 & n7435;
  assign n7437 = n7436 ^ n5291;
  assign n7517 = n7451 ^ n7437;
  assign n7434 = n7131 ^ n7115;
  assign n7518 = n7517 ^ n7434;
  assign n7519 = n7518 ^ n4469;
  assign n7586 = n7527 ^ n7519;
  assign n7587 = n7524 ^ n4471;
  assign n7588 = n7587 ^ n7520;
  assign n7302 = n7301 ^ n4483;
  assign n7312 = n7311 ^ n7302;
  assign n7313 = n7298 ^ n7273;
  assign n7314 = n7295 ^ n4687;
  assign n7315 = n7314 ^ n7275;
  assign n7316 = n7292 ^ n7279;
  assign n7317 = n7282 ^ n4508;
  assign n7318 = n7286 ^ n7284;
  assign n7319 = ~n7317 & ~n7318;
  assign n7320 = n7289 ^ n4676;
  assign n7321 = n7320 ^ n7280;
  assign n7322 = n7319 & n7321;
  assign n7323 = n7316 & ~n7322;
  assign n7324 = n7315 & n7323;
  assign n7325 = n7313 & ~n7324;
  assign n7358 = ~n7312 & n7325;
  assign n7373 = n7372 ^ n7362;
  assign n7589 = ~n7358 & n7373;
  assign n7590 = n7588 & n7589;
  assign n7591 = ~n7586 & ~n7590;
  assign n7528 = n7527 ^ n7518;
  assign n7529 = n7519 & ~n7528;
  assign n7530 = n7529 ^ n4469;
  assign n7592 = n7530 ^ n4456;
  assign n7438 = n7437 ^ n7434;
  assign n7452 = n7451 ^ n7434;
  assign n7453 = ~n7438 & n7452;
  assign n7454 = n7453 ^ n7437;
  assign n7431 = n7134 ^ x250;
  assign n7432 = n7431 ^ n7112;
  assign n7428 = n6317 ^ n5283;
  assign n7429 = n6301 & ~n7428;
  assign n7430 = n7429 ^ n5283;
  assign n7433 = n7432 ^ n7430;
  assign n7515 = n7454 ^ n7433;
  assign n7593 = n7592 ^ n7515;
  assign n7594 = n7591 & n7593;
  assign n7516 = n7515 ^ n4456;
  assign n7531 = n7530 ^ n7515;
  assign n7532 = ~n7516 & ~n7531;
  assign n7533 = n7532 ^ n4456;
  assign n7455 = n7454 ^ n7432;
  assign n7456 = ~n7433 & ~n7455;
  assign n7457 = n7456 ^ n7430;
  assign n7424 = n6309 ^ n5278;
  assign n7425 = n6295 & n7424;
  assign n7426 = n7425 ^ n5278;
  assign n7512 = n7457 ^ n7426;
  assign n7423 = n7137 ^ n7111;
  assign n7513 = n7512 ^ n7423;
  assign n7514 = n7513 ^ n4713;
  assign n7585 = n7533 ^ n7514;
  assign n7721 = n7594 ^ n7585;
  assign n7722 = n7721 ^ x276;
  assign n7723 = n7593 ^ n7591;
  assign n7724 = n7723 ^ x277;
  assign n7725 = n7590 ^ n7586;
  assign n7726 = n7725 ^ x278;
  assign n7727 = n7589 ^ n7588;
  assign n7728 = n7727 ^ x279;
  assign n7374 = n7373 ^ n7358;
  assign n7729 = n7374 ^ x280;
  assign n7326 = n7325 ^ n7312;
  assign n7327 = n7326 ^ x281;
  assign n7328 = n7324 ^ n7313;
  assign n7329 = n7328 ^ x282;
  assign n7330 = n7323 ^ n7315;
  assign n7331 = n7330 ^ x283;
  assign n7332 = n7322 ^ n7316;
  assign n7333 = n7332 ^ x284;
  assign n7334 = n7321 ^ n7319;
  assign n7335 = n7334 ^ x285;
  assign n7336 = x287 & n7317;
  assign n7337 = n7336 ^ x286;
  assign n7338 = n7318 ^ n7317;
  assign n7339 = n7338 ^ n7336;
  assign n7340 = n7337 & ~n7339;
  assign n7341 = n7340 ^ x286;
  assign n7342 = n7341 ^ n7334;
  assign n7343 = n7335 & ~n7342;
  assign n7344 = n7343 ^ x285;
  assign n7345 = n7344 ^ n7332;
  assign n7346 = n7333 & ~n7345;
  assign n7347 = n7346 ^ x284;
  assign n7348 = n7347 ^ n7330;
  assign n7349 = ~n7331 & n7348;
  assign n7350 = n7349 ^ x283;
  assign n7351 = n7350 ^ n7328;
  assign n7352 = ~n7329 & n7351;
  assign n7353 = n7352 ^ x282;
  assign n7354 = n7353 ^ n7326;
  assign n7355 = ~n7327 & n7354;
  assign n7356 = n7355 ^ x281;
  assign n7730 = n7374 ^ n7356;
  assign n7731 = n7729 & ~n7730;
  assign n7732 = n7731 ^ x280;
  assign n7733 = n7732 ^ n7727;
  assign n7734 = ~n7728 & n7733;
  assign n7735 = n7734 ^ x279;
  assign n7736 = n7735 ^ n7725;
  assign n7737 = n7726 & ~n7736;
  assign n7738 = n7737 ^ x278;
  assign n7739 = n7738 ^ n7723;
  assign n7740 = n7724 & ~n7739;
  assign n7741 = n7740 ^ x277;
  assign n7742 = n7741 ^ n7721;
  assign n7743 = n7722 & ~n7742;
  assign n7744 = n7743 ^ x276;
  assign n7534 = n7533 ^ n7513;
  assign n7535 = ~n7514 & ~n7534;
  assign n7536 = n7535 ^ n4713;
  assign n7596 = n7536 ^ n4891;
  assign n7427 = n7426 ^ n7423;
  assign n7458 = n7457 ^ n7423;
  assign n7459 = ~n7427 & n7458;
  assign n7460 = n7459 ^ n7426;
  assign n7420 = n7140 ^ x248;
  assign n7421 = n7420 ^ n7108;
  assign n7417 = n6303 ^ n5303;
  assign n7418 = n6288 & n7417;
  assign n7419 = n7418 ^ n5303;
  assign n7422 = n7421 ^ n7419;
  assign n7510 = n7460 ^ n7422;
  assign n7597 = n7596 ^ n7510;
  assign n7595 = n7585 & ~n7594;
  assign n7719 = n7597 ^ n7595;
  assign n7720 = n7719 ^ x275;
  assign n7986 = n7744 ^ n7720;
  assign n7617 = n7171 ^ x238;
  assign n7618 = n7617 ^ n7089;
  assign n7983 = n6958 ^ n6271;
  assign n7984 = n7618 & ~n7983;
  assign n7985 = n7984 ^ n6271;
  assign n7987 = n7986 ^ n7985;
  assign n7570 = n7168 ^ x239;
  assign n7990 = n6885 ^ n6277;
  assign n7991 = n7570 & ~n7990;
  assign n7992 = n7991 ^ n6277;
  assign n7988 = n7741 ^ x276;
  assign n7989 = n7988 ^ n7721;
  assign n7993 = n7992 ^ n7989;
  assign n7488 = n7164 ^ x240;
  assign n7489 = n7488 ^ n7092;
  assign n7995 = n6756 ^ n6284;
  assign n7996 = ~n7489 & ~n7995;
  assign n7997 = n7996 ^ n6284;
  assign n7994 = n7738 ^ n7724;
  assign n7998 = n7997 ^ n7994;
  assign n8002 = n7735 ^ n7726;
  assign n7383 = n7161 ^ n7095;
  assign n7999 = n6290 ^ n6261;
  assign n8000 = ~n7383 & n7999;
  assign n8001 = n8000 ^ n6290;
  assign n8003 = n8002 ^ n8001;
  assign n7388 = n7158 ^ x242;
  assign n7389 = n7388 ^ n7096;
  assign n8006 = n6297 ^ n6269;
  assign n8007 = n7389 & n8006;
  assign n8008 = n8007 ^ n6297;
  assign n8004 = n7732 ^ x279;
  assign n8005 = n8004 ^ n7727;
  assign n8009 = n8008 ^ n8005;
  assign n7391 = n7155 ^ n7099;
  assign n8010 = n6303 ^ n6275;
  assign n8011 = n7391 & n8010;
  assign n8012 = n8011 ^ n6303;
  assign n7357 = n7356 ^ x280;
  assign n7375 = n7374 ^ n7357;
  assign n8013 = n8012 ^ n7375;
  assign n7399 = n7152 ^ x244;
  assign n7400 = n7399 ^ n7100;
  assign n8014 = n6309 ^ n6282;
  assign n8015 = ~n7400 & n8014;
  assign n8016 = n8015 ^ n6309;
  assign n7899 = n7353 ^ n7327;
  assign n8017 = n8016 ^ n7899;
  assign n7405 = n7149 ^ n7103;
  assign n8018 = n6317 ^ n6288;
  assign n8019 = n7405 & n8018;
  assign n8020 = n8019 ^ n6317;
  assign n7905 = n7350 ^ x282;
  assign n7906 = n7905 ^ n7328;
  assign n8021 = n8020 ^ n7906;
  assign n7376 = n7146 ^ n7105;
  assign n8023 = n6295 ^ n6168;
  assign n8024 = n7376 & n8023;
  assign n8025 = n8024 ^ n6168;
  assign n8022 = n7347 ^ n7331;
  assign n8026 = n8025 ^ n8022;
  assign n7414 = n7143 ^ x247;
  assign n7415 = n7414 ^ n7106;
  assign n8029 = n6301 ^ n6098;
  assign n8030 = ~n7415 & n8029;
  assign n8031 = n8030 ^ n6098;
  assign n8027 = n7344 ^ x284;
  assign n8028 = n8027 ^ n7332;
  assign n8032 = n8031 ^ n8028;
  assign n8034 = n6307 ^ n6088;
  assign n8035 = n7421 & ~n8034;
  assign n8036 = n8035 ^ n6088;
  assign n8033 = n7341 ^ n7335;
  assign n8037 = n8036 ^ n8033;
  assign n8040 = n6322 ^ n6019;
  assign n8041 = n7432 & ~n8040;
  assign n8042 = n8041 ^ n6019;
  assign n8039 = n7317 ^ x287;
  assign n8043 = n8042 ^ n8039;
  assign n7806 = n7186 ^ n7080;
  assign n7802 = n5886 ^ n5216;
  assign n7803 = ~n6687 & n7802;
  assign n7804 = n7803 ^ n5216;
  assign n7838 = n7806 ^ n7804;
  assign n7688 = n7183 ^ x234;
  assign n7689 = n7688 ^ n7081;
  assign n7684 = n5852 ^ n5218;
  assign n7685 = n7244 & n7684;
  assign n7686 = n7685 ^ n5218;
  assign n7798 = n7689 ^ n7686;
  assign n7671 = n7180 ^ n7084;
  assign n7667 = n5796 ^ n5223;
  assign n7668 = ~n7052 & ~n7667;
  assign n7669 = n7668 ^ n5223;
  assign n7680 = n7671 ^ n7669;
  assign n7652 = n6578 ^ n5962;
  assign n7653 = ~n7035 & ~n7652;
  assign n7654 = n7653 ^ n5962;
  assign n7650 = n7177 ^ x236;
  assign n7651 = n7650 ^ n7085;
  assign n7655 = n7654 ^ n7651;
  assign n7638 = n7174 ^ n7088;
  assign n7634 = n6562 ^ n5916;
  assign n7635 = n7021 & ~n7634;
  assign n7636 = n7635 ^ n5916;
  assign n7646 = n7638 ^ n7636;
  assign n7485 = n6366 ^ n5789;
  assign n7486 = ~n6973 & n7485;
  assign n7487 = n7486 ^ n5789;
  assign n7490 = n7489 ^ n7487;
  assign n7380 = n6004 ^ n5546;
  assign n7381 = ~n6958 & n7380;
  assign n7382 = n7381 ^ n5546;
  assign n7384 = n7383 ^ n7382;
  assign n7385 = n6264 ^ n5379;
  assign n7386 = n6885 & ~n7385;
  assign n7387 = n7386 ^ n5379;
  assign n7390 = n7389 ^ n7387;
  assign n7392 = n6271 ^ n4899;
  assign n7393 = ~n6756 & n7392;
  assign n7394 = n7393 ^ n4899;
  assign n7395 = n7394 ^ n7391;
  assign n7396 = n6277 ^ n5330;
  assign n7397 = ~n6261 & n7396;
  assign n7398 = n7397 ^ n5330;
  assign n7401 = n7400 ^ n7398;
  assign n7402 = n6284 ^ n5325;
  assign n7403 = ~n6269 & ~n7402;
  assign n7404 = n7403 ^ n5325;
  assign n7406 = n7405 ^ n7404;
  assign n7407 = n6290 ^ n5321;
  assign n7408 = n6275 & n7407;
  assign n7409 = n7408 ^ n5321;
  assign n7410 = n7409 ^ n7376;
  assign n7411 = n6297 ^ n5311;
  assign n7412 = ~n6282 & ~n7411;
  assign n7413 = n7412 ^ n5311;
  assign n7416 = n7415 ^ n7413;
  assign n7461 = n7460 ^ n7421;
  assign n7462 = n7422 & n7461;
  assign n7463 = n7462 ^ n7419;
  assign n7464 = n7463 ^ n7415;
  assign n7465 = ~n7416 & n7464;
  assign n7466 = n7465 ^ n7413;
  assign n7467 = n7466 ^ n7376;
  assign n7468 = ~n7410 & ~n7467;
  assign n7469 = n7468 ^ n7409;
  assign n7470 = n7469 ^ n7405;
  assign n7471 = ~n7406 & n7470;
  assign n7472 = n7471 ^ n7404;
  assign n7473 = n7472 ^ n7400;
  assign n7474 = n7401 & ~n7473;
  assign n7475 = n7474 ^ n7398;
  assign n7476 = n7475 ^ n7391;
  assign n7477 = n7395 & n7476;
  assign n7478 = n7477 ^ n7394;
  assign n7479 = n7478 ^ n7389;
  assign n7480 = ~n7390 & ~n7479;
  assign n7481 = n7480 ^ n7387;
  assign n7482 = n7481 ^ n7383;
  assign n7483 = ~n7384 & ~n7482;
  assign n7484 = n7483 ^ n7382;
  assign n7567 = n7489 ^ n7484;
  assign n7568 = n7490 & n7567;
  assign n7569 = n7568 ^ n7487;
  assign n7571 = n7570 ^ n7569;
  assign n7564 = n6360 ^ n5842;
  assign n7565 = ~n6991 & ~n7564;
  assign n7566 = n7565 ^ n5842;
  assign n7619 = n7570 ^ n7566;
  assign n7620 = n7571 & n7619;
  assign n7621 = n7620 ^ n7566;
  assign n7622 = n7621 ^ n7618;
  assign n7614 = n6358 ^ n5873;
  assign n7615 = ~n7008 & ~n7614;
  assign n7616 = n7615 ^ n5873;
  assign n7631 = n7618 ^ n7616;
  assign n7632 = ~n7622 & n7631;
  assign n7633 = n7632 ^ n7616;
  assign n7647 = n7638 ^ n7633;
  assign n7648 = n7646 & ~n7647;
  assign n7649 = n7648 ^ n7636;
  assign n7664 = n7651 ^ n7649;
  assign n7665 = n7655 & ~n7664;
  assign n7666 = n7665 ^ n7654;
  assign n7681 = n7671 ^ n7666;
  assign n7682 = ~n7680 & n7681;
  assign n7683 = n7682 ^ n7669;
  assign n7799 = n7689 ^ n7683;
  assign n7800 = ~n7798 & ~n7799;
  assign n7801 = n7800 ^ n7686;
  assign n7839 = n7806 ^ n7801;
  assign n7840 = ~n7838 & n7839;
  assign n7841 = n7840 ^ n7804;
  assign n7835 = n5928 ^ n5211;
  assign n7836 = ~n6682 & ~n7835;
  assign n7837 = n7836 ^ n5211;
  assign n7842 = n7841 ^ n7837;
  assign n7833 = n7189 ^ x232;
  assign n7834 = n7833 ^ n7077;
  assign n7843 = n7842 ^ n7834;
  assign n7875 = n7843 ^ n4631;
  assign n7805 = n7804 ^ n7801;
  assign n7807 = n7806 ^ n7805;
  assign n7828 = n7807 ^ n4654;
  assign n7687 = n7686 ^ n7683;
  assign n7690 = n7689 ^ n7687;
  assign n7793 = n7690 ^ n4640;
  assign n7670 = n7669 ^ n7666;
  assign n7672 = n7671 ^ n7670;
  assign n7675 = n7672 ^ n4645;
  assign n7656 = n7655 ^ n7649;
  assign n7657 = n7656 ^ n5192;
  assign n7637 = n7636 ^ n7633;
  assign n7639 = n7638 ^ n7637;
  assign n7642 = n7639 ^ n5099;
  assign n7623 = n7622 ^ n7616;
  assign n7626 = n7623 ^ n4450;
  assign n7572 = n7571 ^ n7566;
  assign n7573 = n7572 ^ n5063;
  assign n7491 = n7490 ^ n7484;
  assign n7492 = n7491 ^ n4969;
  assign n7493 = n7481 ^ n7384;
  assign n7494 = n7493 ^ n4973;
  assign n7495 = n7478 ^ n7390;
  assign n7496 = n7495 ^ n4978;
  assign n7497 = n7475 ^ n7394;
  assign n7498 = n7497 ^ n7391;
  assign n7499 = n7498 ^ n4987;
  assign n7500 = n7472 ^ n7401;
  assign n7501 = n7500 ^ n4989;
  assign n7502 = n7469 ^ n7404;
  assign n7503 = n7502 ^ n7405;
  assign n7504 = n7503 ^ n4998;
  assign n7505 = n7466 ^ n7410;
  assign n7506 = n7505 ^ n4999;
  assign n7507 = n7463 ^ n7413;
  assign n7508 = n7507 ^ n7415;
  assign n7509 = n7508 ^ n4901;
  assign n7511 = n7510 ^ n4891;
  assign n7537 = n7536 ^ n7510;
  assign n7538 = n7511 & ~n7537;
  assign n7539 = n7538 ^ n4891;
  assign n7540 = n7539 ^ n7508;
  assign n7541 = ~n7509 & ~n7540;
  assign n7542 = n7541 ^ n4901;
  assign n7543 = n7542 ^ n7505;
  assign n7544 = n7506 & n7543;
  assign n7545 = n7544 ^ n4999;
  assign n7546 = n7545 ^ n7503;
  assign n7547 = n7504 & n7546;
  assign n7548 = n7547 ^ n4998;
  assign n7549 = n7548 ^ n7500;
  assign n7550 = n7501 & n7549;
  assign n7551 = n7550 ^ n4989;
  assign n7552 = n7551 ^ n7498;
  assign n7553 = n7499 & ~n7552;
  assign n7554 = n7553 ^ n4987;
  assign n7555 = n7554 ^ n7495;
  assign n7556 = ~n7496 & ~n7555;
  assign n7557 = n7556 ^ n4978;
  assign n7558 = n7557 ^ n7493;
  assign n7559 = n7494 & ~n7558;
  assign n7560 = n7559 ^ n4973;
  assign n7561 = n7560 ^ n7491;
  assign n7562 = n7492 & ~n7561;
  assign n7563 = n7562 ^ n4969;
  assign n7610 = n7572 ^ n7563;
  assign n7611 = ~n7573 & n7610;
  assign n7612 = n7611 ^ n5063;
  assign n7627 = n7623 ^ n7612;
  assign n7628 = n7626 & ~n7627;
  assign n7629 = n7628 ^ n4450;
  assign n7643 = n7639 ^ n7629;
  assign n7644 = ~n7642 & ~n7643;
  assign n7645 = n7644 ^ n5099;
  assign n7660 = n7656 ^ n7645;
  assign n7661 = ~n7657 & n7660;
  assign n7662 = n7661 ^ n5192;
  assign n7676 = n7672 ^ n7662;
  assign n7677 = ~n7675 & ~n7676;
  assign n7678 = n7677 ^ n4645;
  assign n7794 = n7690 ^ n7678;
  assign n7795 = ~n7793 & n7794;
  assign n7796 = n7795 ^ n4640;
  assign n7829 = n7807 ^ n7796;
  assign n7830 = ~n7828 & ~n7829;
  assign n7831 = n7830 ^ n4654;
  assign n7876 = n7843 ^ n7831;
  assign n7877 = n7875 & n7876;
  assign n7878 = n7877 ^ n4631;
  assign n7879 = n7878 ^ n4626;
  assign n7871 = n5980 ^ n5203;
  assign n7872 = n6677 & n7871;
  assign n7873 = n7872 ^ n5203;
  assign n7866 = n7837 ^ n7834;
  assign n7867 = n7841 ^ n7834;
  assign n7868 = ~n7866 & n7867;
  assign n7869 = n7868 ^ n7837;
  assign n7865 = n7192 ^ n7076;
  assign n7870 = n7869 ^ n7865;
  assign n7874 = n7873 ^ n7870;
  assign n7880 = n7879 ^ n7874;
  assign n7832 = n7831 ^ n4631;
  assign n7844 = n7843 ^ n7832;
  assign n7574 = n7573 ^ n7563;
  assign n7575 = n7560 ^ n4969;
  assign n7576 = n7575 ^ n7491;
  assign n7577 = n7554 ^ n4978;
  assign n7578 = n7577 ^ n7495;
  assign n7579 = n7551 ^ n4987;
  assign n7580 = n7579 ^ n7498;
  assign n7581 = n7548 ^ n7501;
  assign n7582 = n7545 ^ n7504;
  assign n7583 = n7542 ^ n4999;
  assign n7584 = n7583 ^ n7505;
  assign n7598 = n7595 & n7597;
  assign n7599 = n7539 ^ n7509;
  assign n7600 = n7598 & ~n7599;
  assign n7601 = ~n7584 & n7600;
  assign n7602 = ~n7582 & ~n7601;
  assign n7603 = n7581 & n7602;
  assign n7604 = n7580 & ~n7603;
  assign n7605 = n7578 & ~n7604;
  assign n7606 = n7557 ^ n7494;
  assign n7607 = n7605 & n7606;
  assign n7608 = n7576 & n7607;
  assign n7609 = ~n7574 & n7608;
  assign n7613 = n7612 ^ n4450;
  assign n7624 = n7623 ^ n7613;
  assign n7625 = n7609 & n7624;
  assign n7630 = n7629 ^ n5099;
  assign n7640 = n7639 ^ n7630;
  assign n7641 = ~n7625 & n7640;
  assign n7658 = n7657 ^ n7645;
  assign n7659 = ~n7641 & n7658;
  assign n7663 = n7662 ^ n4645;
  assign n7673 = n7672 ^ n7663;
  assign n7674 = ~n7659 & ~n7673;
  assign n7679 = n7678 ^ n4640;
  assign n7691 = n7690 ^ n7679;
  assign n7792 = ~n7674 & ~n7691;
  assign n7797 = n7796 ^ n4654;
  assign n7808 = n7807 ^ n7797;
  assign n7845 = ~n7792 & n7808;
  assign n7864 = n7844 & n7845;
  assign n7881 = n7880 ^ n7864;
  assign n7882 = n7881 ^ x258;
  assign n7846 = n7845 ^ n7844;
  assign n7860 = n7846 ^ x259;
  assign n7809 = n7808 ^ n7792;
  assign n7823 = n7809 ^ x260;
  assign n7692 = n7691 ^ n7674;
  assign n7693 = n7692 ^ x261;
  assign n7694 = n7673 ^ n7659;
  assign n7695 = n7694 ^ x262;
  assign n7696 = n7658 ^ n7641;
  assign n7697 = n7696 ^ x263;
  assign n7698 = n7640 ^ n7625;
  assign n7699 = n7698 ^ x264;
  assign n7700 = n7624 ^ n7609;
  assign n7701 = n7700 ^ x265;
  assign n7702 = n7608 ^ n7574;
  assign n7703 = n7702 ^ x266;
  assign n7704 = n7607 ^ n7576;
  assign n7705 = n7704 ^ x267;
  assign n7706 = n7606 ^ n7605;
  assign n7707 = n7706 ^ x268;
  assign n7708 = n7604 ^ n7578;
  assign n7709 = n7708 ^ x269;
  assign n7710 = n7603 ^ n7580;
  assign n7711 = n7710 ^ x270;
  assign n7713 = n7601 ^ n7582;
  assign n7714 = n7713 ^ x272;
  assign n7715 = n7600 ^ n7584;
  assign n7716 = n7715 ^ x273;
  assign n7717 = n7599 ^ n7598;
  assign n7718 = n7717 ^ x274;
  assign n7745 = n7744 ^ n7719;
  assign n7746 = ~n7720 & n7745;
  assign n7747 = n7746 ^ x275;
  assign n7748 = n7747 ^ n7717;
  assign n7749 = n7718 & ~n7748;
  assign n7750 = n7749 ^ x274;
  assign n7751 = n7750 ^ n7715;
  assign n7752 = n7716 & ~n7751;
  assign n7753 = n7752 ^ x273;
  assign n7754 = n7753 ^ n7713;
  assign n7755 = n7714 & ~n7754;
  assign n7756 = n7755 ^ x272;
  assign n7712 = n7602 ^ n7581;
  assign n7757 = n7756 ^ n7712;
  assign n7758 = n7712 ^ x271;
  assign n7759 = ~n7757 & n7758;
  assign n7760 = n7759 ^ x271;
  assign n7761 = n7760 ^ n7710;
  assign n7762 = n7711 & ~n7761;
  assign n7763 = n7762 ^ x270;
  assign n7764 = n7763 ^ n7708;
  assign n7765 = ~n7709 & n7764;
  assign n7766 = n7765 ^ x269;
  assign n7767 = n7766 ^ n7706;
  assign n7768 = n7707 & ~n7767;
  assign n7769 = n7768 ^ x268;
  assign n7770 = n7769 ^ n7704;
  assign n7771 = n7705 & ~n7770;
  assign n7772 = n7771 ^ x267;
  assign n7773 = n7772 ^ n7702;
  assign n7774 = ~n7703 & n7773;
  assign n7775 = n7774 ^ x266;
  assign n7776 = n7775 ^ n7700;
  assign n7777 = n7701 & ~n7776;
  assign n7778 = n7777 ^ x265;
  assign n7779 = n7778 ^ n7698;
  assign n7780 = n7699 & ~n7779;
  assign n7781 = n7780 ^ x264;
  assign n7782 = n7781 ^ n7696;
  assign n7783 = ~n7697 & n7782;
  assign n7784 = n7783 ^ x263;
  assign n7785 = n7784 ^ n7694;
  assign n7786 = ~n7695 & n7785;
  assign n7787 = n7786 ^ x262;
  assign n7788 = n7787 ^ n7692;
  assign n7789 = n7693 & ~n7788;
  assign n7790 = n7789 ^ x261;
  assign n7824 = n7809 ^ n7790;
  assign n7825 = n7823 & ~n7824;
  assign n7826 = n7825 ^ x260;
  assign n7861 = n7846 ^ n7826;
  assign n7862 = ~n7860 & n7861;
  assign n7863 = n7862 ^ x259;
  assign n8066 = n7881 ^ n7863;
  assign n8067 = n7882 & ~n8066;
  assign n8068 = n8067 ^ x258;
  assign n8069 = n8068 ^ x257;
  assign n8059 = n7874 ^ n4626;
  assign n8060 = n7878 ^ n7874;
  assign n8061 = ~n8059 & n8060;
  assign n8062 = n8061 ^ n4626;
  assign n8063 = n8062 ^ n4518;
  assign n8055 = n6053 ^ n4960;
  assign n8056 = n6672 & n8055;
  assign n8057 = n8056 ^ n4960;
  assign n8051 = n7873 ^ n7865;
  assign n8052 = n7870 & n8051;
  assign n8053 = n8052 ^ n7873;
  assign n7938 = n7195 ^ x230;
  assign n7939 = n7938 ^ n7073;
  assign n8054 = n8053 ^ n7939;
  assign n8058 = n8057 ^ n8054;
  assign n8064 = n8063 ^ n8058;
  assign n8050 = ~n7864 & ~n7880;
  assign n8065 = n8064 ^ n8050;
  assign n8070 = n8069 ^ n8065;
  assign n8047 = n6330 ^ n6000;
  assign n8048 = ~n7443 & n8047;
  assign n8049 = n8048 ^ n6000;
  assign n8071 = n8070 ^ n8049;
  assign n7827 = n7826 ^ x259;
  assign n7847 = n7846 ^ n7827;
  assign n7819 = n6037 ^ n5997;
  assign n7820 = ~n7306 & ~n7819;
  assign n7821 = n7820 ^ n6037;
  assign n7887 = n7847 ^ n7821;
  assign n7791 = n7790 ^ x260;
  assign n7810 = n7809 ^ n7791;
  assign n7811 = n6343 ^ n6043;
  assign n7812 = n7267 & ~n7811;
  assign n7813 = n7812 ^ n6043;
  assign n7818 = n7810 & n7813;
  assign n7888 = n7847 ^ n7818;
  assign n7889 = ~n7887 & ~n7888;
  assign n7890 = n7889 ^ n7818;
  assign n7884 = n6032 ^ n5990;
  assign n7885 = ~n7370 & n7884;
  assign n7886 = n7885 ^ n6032;
  assign n7891 = n7890 ^ n7886;
  assign n7883 = n7882 ^ n7863;
  assign n8072 = n7890 ^ n7883;
  assign n8073 = n7891 & ~n8072;
  assign n8074 = n8073 ^ n7886;
  assign n8075 = n8074 ^ n8070;
  assign n8076 = n8071 & ~n8075;
  assign n8077 = n8076 ^ n8049;
  assign n8044 = n6324 ^ n5992;
  assign n8045 = ~n7434 & n8044;
  assign n8046 = n8045 ^ n5992;
  assign n8078 = n8077 ^ n8046;
  assign n8095 = n8065 ^ x257;
  assign n8096 = n8068 ^ n8065;
  assign n8097 = n8095 & ~n8096;
  assign n8098 = n8097 ^ x257;
  assign n8099 = n8098 ^ x256;
  assign n8090 = n8058 ^ n4518;
  assign n8091 = n8062 ^ n8058;
  assign n8092 = ~n8090 & ~n8091;
  assign n8093 = n8092 ^ n4518;
  assign n8088 = ~n8050 & n8064;
  assign n8084 = n8057 ^ n7939;
  assign n8085 = ~n8054 & n8084;
  assign n8086 = n8085 ^ n8057;
  assign n8079 = n6048 ^ n4955;
  assign n8080 = ~n6667 & ~n8079;
  assign n8081 = n8080 ^ n4955;
  assign n7932 = n7198 ^ n7072;
  assign n8082 = n8081 ^ n7932;
  assign n8083 = n8082 ^ n4513;
  assign n8087 = n8086 ^ n8083;
  assign n8089 = n8088 ^ n8087;
  assign n8094 = n8093 ^ n8089;
  assign n8100 = n8099 ^ n8094;
  assign n8101 = n8100 ^ n8077;
  assign n8102 = ~n8078 & ~n8101;
  assign n8103 = n8102 ^ n8046;
  assign n8104 = n8103 ^ n8039;
  assign n8105 = n8043 & n8104;
  assign n8106 = n8105 ^ n8042;
  assign n8038 = n7338 ^ n7337;
  assign n8107 = n8106 ^ n8038;
  assign n8108 = n6314 ^ n6014;
  assign n8109 = n7423 & ~n8108;
  assign n8110 = n8109 ^ n6014;
  assign n8111 = n8110 ^ n8038;
  assign n8112 = ~n8107 & n8111;
  assign n8113 = n8112 ^ n8110;
  assign n8114 = n8113 ^ n8033;
  assign n8115 = ~n8037 & ~n8114;
  assign n8116 = n8115 ^ n8036;
  assign n8117 = n8116 ^ n8028;
  assign n8118 = n8032 & n8117;
  assign n8119 = n8118 ^ n8031;
  assign n8120 = n8119 ^ n8022;
  assign n8121 = ~n8026 & n8120;
  assign n8122 = n8121 ^ n8025;
  assign n8123 = n8122 ^ n7906;
  assign n8124 = ~n8021 & n8123;
  assign n8125 = n8124 ^ n8020;
  assign n8126 = n8125 ^ n7899;
  assign n8127 = n8017 & n8126;
  assign n8128 = n8127 ^ n8016;
  assign n8129 = n8128 ^ n7375;
  assign n8130 = n8013 & n8129;
  assign n8131 = n8130 ^ n8012;
  assign n8132 = n8131 ^ n8005;
  assign n8133 = n8009 & n8132;
  assign n8134 = n8133 ^ n8008;
  assign n8135 = n8134 ^ n8002;
  assign n8136 = ~n8003 & n8135;
  assign n8137 = n8136 ^ n8001;
  assign n8138 = n8137 ^ n7994;
  assign n8139 = n7998 & n8138;
  assign n8140 = n8139 ^ n7997;
  assign n8141 = n8140 ^ n7989;
  assign n8142 = ~n7993 & ~n8141;
  assign n8143 = n8142 ^ n7992;
  assign n8144 = n8143 ^ n7986;
  assign n8145 = ~n7987 & ~n8144;
  assign n8146 = n8145 ^ n7985;
  assign n7979 = n6973 ^ n6264;
  assign n7980 = n7638 & ~n7979;
  assign n7981 = n7980 ^ n6264;
  assign n7977 = n7747 ^ x274;
  assign n7978 = n7977 ^ n7717;
  assign n7982 = n7981 ^ n7978;
  assign n8224 = n8146 ^ n7982;
  assign n8225 = n8224 ^ n5379;
  assign n8226 = n8143 ^ n7987;
  assign n8227 = n8226 ^ n4899;
  assign n8228 = n8140 ^ n7992;
  assign n8229 = n8228 ^ n7989;
  assign n8230 = n8229 ^ n5330;
  assign n8231 = n8137 ^ n7998;
  assign n8232 = n8231 ^ n5325;
  assign n8233 = n8134 ^ n8003;
  assign n8234 = n8233 ^ n5321;
  assign n8235 = n8131 ^ n8009;
  assign n8236 = n8235 ^ n5311;
  assign n8237 = n8128 ^ n8013;
  assign n8238 = n8237 ^ n5303;
  assign n8239 = n8125 ^ n8017;
  assign n8240 = n8239 ^ n5278;
  assign n8241 = n8122 ^ n8021;
  assign n8242 = n8241 ^ n5283;
  assign n8243 = n8119 ^ n8025;
  assign n8244 = n8243 ^ n8022;
  assign n8245 = n8244 ^ n5291;
  assign n8246 = n8116 ^ n8031;
  assign n8247 = n8246 ^ n8028;
  assign n8248 = n8247 ^ n4907;
  assign n8249 = n8113 ^ n8036;
  assign n8250 = n8249 ^ n8033;
  assign n8251 = n8250 ^ n4915;
  assign n8252 = n8110 ^ n8107;
  assign n8253 = n8252 ^ n4920;
  assign n8254 = n8103 ^ n8042;
  assign n8255 = n8254 ^ n8039;
  assign n8256 = n8255 ^ n4925;
  assign n8257 = n8100 ^ n8078;
  assign n8258 = n8257 ^ n4930;
  assign n8259 = n8074 ^ n8049;
  assign n8260 = n8259 ^ n8070;
  assign n8261 = n8260 ^ n4935;
  assign n7892 = n7891 ^ n7883;
  assign n8262 = n7892 ^ n4940;
  assign n7814 = n7813 ^ n7810;
  assign n7849 = n4950 & n7814;
  assign n7850 = n7849 ^ n4942;
  assign n7822 = n7821 ^ n7818;
  assign n7848 = n7847 ^ n7822;
  assign n7856 = n7849 ^ n7848;
  assign n7857 = n7850 & ~n7856;
  assign n7858 = n7857 ^ n4942;
  assign n8263 = n7892 ^ n7858;
  assign n8264 = ~n8262 & ~n8263;
  assign n8265 = n8264 ^ n4940;
  assign n8266 = n8265 ^ n8260;
  assign n8267 = ~n8261 & n8266;
  assign n8268 = n8267 ^ n4935;
  assign n8269 = n8268 ^ n8257;
  assign n8270 = ~n8258 & ~n8269;
  assign n8271 = n8270 ^ n4930;
  assign n8272 = n8271 ^ n8255;
  assign n8273 = n8256 & n8272;
  assign n8274 = n8273 ^ n4925;
  assign n8275 = n8274 ^ n8252;
  assign n8276 = ~n8253 & n8275;
  assign n8277 = n8276 ^ n4920;
  assign n8278 = n8277 ^ n8250;
  assign n8279 = n8251 & ~n8278;
  assign n8280 = n8279 ^ n4915;
  assign n8281 = n8280 ^ n8247;
  assign n8282 = ~n8248 & ~n8281;
  assign n8283 = n8282 ^ n4907;
  assign n8284 = n8283 ^ n8244;
  assign n8285 = ~n8245 & n8284;
  assign n8286 = n8285 ^ n5291;
  assign n8287 = n8286 ^ n8241;
  assign n8288 = n8242 & n8287;
  assign n8289 = n8288 ^ n5283;
  assign n8290 = n8289 ^ n8239;
  assign n8291 = ~n8240 & n8290;
  assign n8292 = n8291 ^ n5278;
  assign n8293 = n8292 ^ n8237;
  assign n8294 = ~n8238 & ~n8293;
  assign n8295 = n8294 ^ n5303;
  assign n8296 = n8295 ^ n8235;
  assign n8297 = n8236 & ~n8296;
  assign n8298 = n8297 ^ n5311;
  assign n8299 = n8298 ^ n8233;
  assign n8300 = ~n8234 & ~n8299;
  assign n8301 = n8300 ^ n5321;
  assign n8302 = n8301 ^ n8231;
  assign n8303 = n8232 & ~n8302;
  assign n8304 = n8303 ^ n5325;
  assign n8305 = n8304 ^ n8229;
  assign n8306 = n8230 & ~n8305;
  assign n8307 = n8306 ^ n5330;
  assign n8308 = n8307 ^ n8226;
  assign n8309 = n8227 & n8308;
  assign n8310 = n8309 ^ n4899;
  assign n8311 = n8310 ^ n8224;
  assign n8312 = ~n8225 & ~n8311;
  assign n8313 = n8312 ^ n5379;
  assign n8147 = n8146 ^ n7978;
  assign n8148 = n7982 & ~n8147;
  assign n8149 = n8148 ^ n7981;
  assign n7975 = n7750 ^ n7716;
  assign n7972 = n6991 ^ n6004;
  assign n7973 = n7651 & ~n7972;
  assign n7974 = n7973 ^ n6004;
  assign n7976 = n7975 ^ n7974;
  assign n8222 = n8149 ^ n7976;
  assign n8223 = n8222 ^ n5546;
  assign n8402 = n8313 ^ n8223;
  assign n8358 = n8310 ^ n5379;
  assign n8359 = n8358 ^ n8224;
  assign n8360 = n8307 ^ n8227;
  assign n8361 = n8295 ^ n8236;
  assign n8362 = n8292 ^ n5303;
  assign n8363 = n8362 ^ n8237;
  assign n8364 = n8289 ^ n8240;
  assign n8365 = n8277 ^ n4915;
  assign n8366 = n8365 ^ n8250;
  assign n8367 = n8274 ^ n4920;
  assign n8368 = n8367 ^ n8252;
  assign n7859 = n7858 ^ n4940;
  assign n7893 = n7892 ^ n7859;
  assign n7815 = n7814 ^ n4950;
  assign n7851 = n7850 ^ n7848;
  assign n7894 = n7815 & n7851;
  assign n8369 = ~n7893 & n7894;
  assign n8370 = n8265 ^ n8261;
  assign n8371 = ~n8369 & ~n8370;
  assign n8372 = n8268 ^ n4930;
  assign n8373 = n8372 ^ n8257;
  assign n8374 = n8371 & ~n8373;
  assign n8375 = n8271 ^ n4925;
  assign n8376 = n8375 ^ n8255;
  assign n8377 = ~n8374 & n8376;
  assign n8378 = n8368 & n8377;
  assign n8379 = n8366 & ~n8378;
  assign n8380 = n8280 ^ n4907;
  assign n8381 = n8380 ^ n8247;
  assign n8382 = n8379 & ~n8381;
  assign n8383 = n8283 ^ n5291;
  assign n8384 = n8383 ^ n8244;
  assign n8385 = ~n8382 & ~n8384;
  assign n8386 = n8286 ^ n5283;
  assign n8387 = n8386 ^ n8241;
  assign n8388 = n8385 & n8387;
  assign n8389 = ~n8364 & ~n8388;
  assign n8390 = ~n8363 & n8389;
  assign n8391 = ~n8361 & n8390;
  assign n8392 = n8298 ^ n5321;
  assign n8393 = n8392 ^ n8233;
  assign n8394 = n8391 & n8393;
  assign n8395 = n8301 ^ n5325;
  assign n8396 = n8395 ^ n8231;
  assign n8397 = ~n8394 & ~n8396;
  assign n8398 = n8304 ^ n8230;
  assign n8399 = n8397 & ~n8398;
  assign n8400 = n8360 & ~n8399;
  assign n8401 = ~n8359 & ~n8400;
  assign n8449 = n8402 ^ n8401;
  assign n8450 = n8449 ^ x300;
  assign n8451 = n8400 ^ n8359;
  assign n8452 = n8451 ^ x301;
  assign n8453 = n8399 ^ n8360;
  assign n8454 = n8453 ^ x302;
  assign n8456 = n8396 ^ n8394;
  assign n8457 = n8456 ^ x304;
  assign n8458 = n8393 ^ n8391;
  assign n8459 = n8458 ^ x305;
  assign n8460 = n8390 ^ n8361;
  assign n8461 = n8460 ^ x306;
  assign n8462 = n8389 ^ n8363;
  assign n8463 = n8462 ^ x307;
  assign n8465 = n8387 ^ n8385;
  assign n8466 = n8465 ^ x309;
  assign n8467 = n8384 ^ n8382;
  assign n8468 = n8467 ^ x310;
  assign n8469 = n8381 ^ n8379;
  assign n8470 = n8469 ^ x311;
  assign n8471 = n8378 ^ n8366;
  assign n8472 = n8471 ^ x312;
  assign n8473 = n8377 ^ n8368;
  assign n8474 = n8473 ^ x313;
  assign n8475 = n8376 ^ n8374;
  assign n8476 = n8475 ^ x314;
  assign n8477 = n8373 ^ n8371;
  assign n8478 = n8477 ^ x315;
  assign n8479 = n8370 ^ n8369;
  assign n8480 = n8479 ^ x316;
  assign n7895 = n7894 ^ n7893;
  assign n7896 = n7895 ^ x317;
  assign n7816 = x319 & ~n7815;
  assign n7817 = n7816 ^ x318;
  assign n7852 = n7851 ^ n7815;
  assign n7853 = n7852 ^ n7816;
  assign n7854 = n7817 & ~n7853;
  assign n7855 = n7854 ^ x318;
  assign n8481 = n7895 ^ n7855;
  assign n8482 = ~n7896 & n8481;
  assign n8483 = n8482 ^ x317;
  assign n8484 = n8483 ^ n8479;
  assign n8485 = ~n8480 & n8484;
  assign n8486 = n8485 ^ x316;
  assign n8487 = n8486 ^ n8477;
  assign n8488 = n8478 & ~n8487;
  assign n8489 = n8488 ^ x315;
  assign n8490 = n8489 ^ n8475;
  assign n8491 = ~n8476 & n8490;
  assign n8492 = n8491 ^ x314;
  assign n8493 = n8492 ^ n8473;
  assign n8494 = n8474 & ~n8493;
  assign n8495 = n8494 ^ x313;
  assign n8496 = n8495 ^ n8471;
  assign n8497 = n8472 & ~n8496;
  assign n8498 = n8497 ^ x312;
  assign n8499 = n8498 ^ n8469;
  assign n8500 = n8470 & ~n8499;
  assign n8501 = n8500 ^ x311;
  assign n8502 = n8501 ^ n8467;
  assign n8503 = n8468 & ~n8502;
  assign n8504 = n8503 ^ x310;
  assign n8505 = n8504 ^ n8465;
  assign n8506 = n8466 & ~n8505;
  assign n8507 = n8506 ^ x309;
  assign n8464 = n8388 ^ n8364;
  assign n8508 = n8507 ^ n8464;
  assign n8509 = n8464 ^ x308;
  assign n8510 = n8508 & ~n8509;
  assign n8511 = n8510 ^ x308;
  assign n8512 = n8511 ^ n8462;
  assign n8513 = n8463 & ~n8512;
  assign n8514 = n8513 ^ x307;
  assign n8515 = n8514 ^ n8460;
  assign n8516 = n8461 & ~n8515;
  assign n8517 = n8516 ^ x306;
  assign n8518 = n8517 ^ n8458;
  assign n8519 = ~n8459 & n8518;
  assign n8520 = n8519 ^ x305;
  assign n8521 = n8520 ^ n8456;
  assign n8522 = n8457 & ~n8521;
  assign n8523 = n8522 ^ x304;
  assign n8455 = n8398 ^ n8397;
  assign n8524 = n8523 ^ n8455;
  assign n8525 = n8455 ^ x303;
  assign n8526 = n8524 & ~n8525;
  assign n8527 = n8526 ^ x303;
  assign n8528 = n8527 ^ n8453;
  assign n8529 = n8454 & ~n8528;
  assign n8530 = n8529 ^ x302;
  assign n8531 = n8530 ^ n8451;
  assign n8532 = n8452 & ~n8531;
  assign n8533 = n8532 ^ x301;
  assign n8534 = n8533 ^ n8449;
  assign n8535 = ~n8450 & n8534;
  assign n8536 = n8535 ^ x300;
  assign n8403 = n8401 & ~n8402;
  assign n8314 = n8313 ^ n8222;
  assign n8315 = n8223 & n8314;
  assign n8316 = n8315 ^ n5546;
  assign n8356 = n8316 ^ n5789;
  assign n8150 = n8149 ^ n7975;
  assign n8151 = n7976 & ~n8150;
  assign n8152 = n8151 ^ n7974;
  assign n7969 = n7753 ^ x272;
  assign n7970 = n7969 ^ n7713;
  assign n7966 = n7008 ^ n6366;
  assign n7967 = ~n7671 & n7966;
  assign n7968 = n7967 ^ n6366;
  assign n7971 = n7970 ^ n7968;
  assign n8220 = n8152 ^ n7971;
  assign n8357 = n8356 ^ n8220;
  assign n8447 = n8403 ^ n8357;
  assign n8448 = n8447 ^ x299;
  assign n8904 = n8536 ^ n8448;
  assign n7925 = n7775 ^ n7701;
  assign n9412 = n7925 ^ n7806;
  assign n9413 = n8904 & n9412;
  assign n9414 = n9413 ^ n7806;
  assign n8855 = n8495 ^ x312;
  assign n8856 = n8855 ^ n8471;
  assign n8852 = n7383 ^ n6275;
  assign n8853 = ~n7986 & ~n8852;
  assign n8854 = n8853 ^ n6275;
  assign n8857 = n8856 ^ n8854;
  assign n8776 = n8492 ^ n8474;
  assign n8773 = n7389 ^ n6282;
  assign n8774 = n7989 & ~n8773;
  assign n8775 = n8774 ^ n6282;
  assign n8777 = n8776 ^ n8775;
  assign n8708 = n8489 ^ x314;
  assign n8709 = n8708 ^ n8475;
  assign n8705 = n7391 ^ n6288;
  assign n8706 = n7994 & n8705;
  assign n8707 = n8706 ^ n6288;
  assign n8710 = n8709 ^ n8707;
  assign n8675 = n8486 ^ n8478;
  assign n8672 = n7400 ^ n6295;
  assign n8673 = n8002 & ~n8672;
  assign n8674 = n8673 ^ n6295;
  assign n8676 = n8675 ^ n8674;
  assign n8622 = n7405 ^ n6301;
  assign n8623 = ~n8005 & n8622;
  assign n8624 = n8623 ^ n6301;
  assign n8620 = n8483 ^ x316;
  assign n8621 = n8620 ^ n8479;
  assign n8625 = n8624 ^ n8621;
  assign n7897 = n7896 ^ n7855;
  assign n7377 = n7376 ^ n6307;
  assign n7378 = n7375 & n7377;
  assign n7379 = n7378 ^ n6307;
  assign n7898 = n7897 ^ n7379;
  assign n7903 = n7852 ^ n7817;
  assign n7900 = n7415 ^ n6314;
  assign n7901 = ~n7899 & n7900;
  assign n7902 = n7901 ^ n6314;
  assign n7904 = n7903 ^ n7902;
  assign n7910 = n7815 ^ x319;
  assign n7907 = n7421 ^ n6322;
  assign n7908 = ~n7906 & ~n7907;
  assign n7909 = n7908 ^ n6322;
  assign n7911 = n7910 ^ n7909;
  assign n8573 = n7423 ^ n6324;
  assign n8574 = ~n8022 & ~n8573;
  assign n8575 = n8574 ^ n6324;
  assign n7926 = n6677 ^ n5886;
  assign n7927 = n7226 & ~n7926;
  assign n7928 = n7927 ^ n5886;
  assign n7929 = n7928 ^ n7925;
  assign n7933 = n6682 ^ n5852;
  assign n7934 = n7932 & n7933;
  assign n7935 = n7934 ^ n5852;
  assign n7930 = n7772 ^ x266;
  assign n7931 = n7930 ^ n7702;
  assign n7936 = n7935 ^ n7931;
  assign n7940 = n6687 ^ n5796;
  assign n7941 = n7939 & n7940;
  assign n7942 = n7941 ^ n5796;
  assign n7937 = n7769 ^ n7705;
  assign n7943 = n7942 ^ n7937;
  assign n7947 = n7766 ^ x268;
  assign n7948 = n7947 ^ n7706;
  assign n7944 = n7244 ^ n6578;
  assign n7945 = n7865 & ~n7944;
  assign n7946 = n7945 ^ n6578;
  assign n7949 = n7948 ^ n7946;
  assign n7953 = n7763 ^ n7709;
  assign n7950 = n7052 ^ n6562;
  assign n7951 = n7834 & n7950;
  assign n7952 = n7951 ^ n6562;
  assign n7954 = n7953 ^ n7952;
  assign n7958 = n7760 ^ x270;
  assign n7959 = n7958 ^ n7710;
  assign n7955 = n7035 ^ n6358;
  assign n7956 = n7806 & n7955;
  assign n7957 = n7956 ^ n6358;
  assign n7960 = n7959 ^ n7957;
  assign n7964 = n7757 ^ x271;
  assign n7961 = n7021 ^ n6360;
  assign n7962 = n7689 & ~n7961;
  assign n7963 = n7962 ^ n6360;
  assign n7965 = n7964 ^ n7963;
  assign n8153 = n8152 ^ n7970;
  assign n8154 = ~n7971 & ~n8153;
  assign n8155 = n8154 ^ n7968;
  assign n8156 = n8155 ^ n7964;
  assign n8157 = ~n7965 & n8156;
  assign n8158 = n8157 ^ n7963;
  assign n8159 = n8158 ^ n7959;
  assign n8160 = ~n7960 & n8159;
  assign n8161 = n8160 ^ n7957;
  assign n8162 = n8161 ^ n7953;
  assign n8163 = n7954 & ~n8162;
  assign n8164 = n8163 ^ n7952;
  assign n8165 = n8164 ^ n7948;
  assign n8166 = ~n7949 & n8165;
  assign n8167 = n8166 ^ n7946;
  assign n8168 = n8167 ^ n7937;
  assign n8169 = ~n7943 & n8168;
  assign n8170 = n8169 ^ n7942;
  assign n8171 = n8170 ^ n7931;
  assign n8172 = n7936 & ~n8171;
  assign n8173 = n8172 ^ n7935;
  assign n8174 = n8173 ^ n7925;
  assign n8175 = ~n7929 & n8174;
  assign n8176 = n8175 ^ n7928;
  assign n7921 = n6672 ^ n5928;
  assign n7922 = n7220 & n7921;
  assign n7923 = n7922 ^ n5928;
  assign n8200 = n8176 ^ n7923;
  assign n7919 = n7778 ^ x264;
  assign n7920 = n7919 ^ n7698;
  assign n8201 = n8200 ^ n7920;
  assign n8202 = n8201 ^ n5211;
  assign n8203 = n8173 ^ n7928;
  assign n8204 = n8203 ^ n7925;
  assign n8205 = n8204 ^ n5216;
  assign n8206 = n8170 ^ n7935;
  assign n8207 = n8206 ^ n7931;
  assign n8208 = n8207 ^ n5218;
  assign n8209 = n8167 ^ n7942;
  assign n8210 = n8209 ^ n7937;
  assign n8211 = n8210 ^ n5223;
  assign n8212 = n8164 ^ n7949;
  assign n8213 = n8212 ^ n5962;
  assign n8214 = n8161 ^ n7954;
  assign n8215 = n8214 ^ n5916;
  assign n8216 = n8158 ^ n7960;
  assign n8217 = n8216 ^ n5873;
  assign n8218 = n8155 ^ n7965;
  assign n8219 = n8218 ^ n5842;
  assign n8221 = n8220 ^ n5789;
  assign n8317 = n8316 ^ n8220;
  assign n8318 = n8221 & n8317;
  assign n8319 = n8318 ^ n5789;
  assign n8320 = n8319 ^ n8218;
  assign n8321 = n8219 & n8320;
  assign n8322 = n8321 ^ n5842;
  assign n8323 = n8322 ^ n8216;
  assign n8324 = n8217 & ~n8323;
  assign n8325 = n8324 ^ n5873;
  assign n8326 = n8325 ^ n8214;
  assign n8327 = ~n8215 & n8326;
  assign n8328 = n8327 ^ n5916;
  assign n8329 = n8328 ^ n8212;
  assign n8330 = n8213 & ~n8329;
  assign n8331 = n8330 ^ n5962;
  assign n8332 = n8331 ^ n8210;
  assign n8333 = n8211 & ~n8332;
  assign n8334 = n8333 ^ n5223;
  assign n8335 = n8334 ^ n8207;
  assign n8336 = n8208 & n8335;
  assign n8337 = n8336 ^ n5218;
  assign n8338 = n8337 ^ n8204;
  assign n8339 = ~n8205 & n8338;
  assign n8340 = n8339 ^ n5216;
  assign n8341 = n8340 ^ n8201;
  assign n8342 = n8202 & ~n8341;
  assign n8343 = n8342 ^ n5211;
  assign n8349 = n8343 ^ n5203;
  assign n8181 = n6667 ^ n5980;
  assign n8182 = ~n7215 & ~n8181;
  assign n8183 = n8182 ^ n5980;
  assign n7924 = n7923 ^ n7920;
  assign n8177 = n8176 ^ n7920;
  assign n8178 = n7924 & n8177;
  assign n8179 = n8178 ^ n7923;
  assign n7918 = n7781 ^ n7697;
  assign n8180 = n8179 ^ n7918;
  assign n8198 = n8183 ^ n8180;
  assign n8350 = n8349 ^ n8198;
  assign n8351 = n8340 ^ n5211;
  assign n8352 = n8351 ^ n8201;
  assign n8353 = n8337 ^ n5216;
  assign n8354 = n8353 ^ n8204;
  assign n8355 = n8331 ^ n8211;
  assign n8404 = n8357 & n8403;
  assign n8405 = n8319 ^ n8219;
  assign n8406 = n8404 & ~n8405;
  assign n8407 = n8322 ^ n5873;
  assign n8408 = n8407 ^ n8216;
  assign n8409 = n8406 & n8408;
  assign n8410 = n8325 ^ n8215;
  assign n8411 = ~n8409 & n8410;
  assign n8412 = n8328 ^ n8213;
  assign n8413 = ~n8411 & n8412;
  assign n8414 = ~n8355 & ~n8413;
  assign n8415 = n8334 ^ n5218;
  assign n8416 = n8415 ^ n8207;
  assign n8417 = ~n8414 & n8416;
  assign n8418 = ~n8354 & ~n8417;
  assign n8419 = n8352 & n8418;
  assign n8420 = n8350 & ~n8419;
  assign n8199 = n8198 ^ n5203;
  assign n8344 = n8343 ^ n8198;
  assign n8345 = ~n8199 & ~n8344;
  assign n8346 = n8345 ^ n5203;
  assign n8347 = n8346 ^ n4960;
  assign n8190 = n6356 ^ n6053;
  assign n8191 = n7212 & ~n8190;
  assign n8192 = n8191 ^ n6053;
  assign n8187 = n7784 ^ x262;
  assign n8188 = n8187 ^ n7694;
  assign n8184 = n8183 ^ n7918;
  assign n8185 = n8180 & ~n8184;
  assign n8186 = n8185 ^ n8183;
  assign n8189 = n8188 ^ n8186;
  assign n8197 = n8192 ^ n8189;
  assign n8348 = n8347 ^ n8197;
  assign n8428 = n8420 ^ n8348;
  assign n8429 = n8428 ^ x289;
  assign n8431 = n8418 ^ n8352;
  assign n8432 = n8431 ^ x291;
  assign n8433 = n8417 ^ n8354;
  assign n8434 = n8433 ^ x292;
  assign n8435 = n8416 ^ n8414;
  assign n8436 = n8435 ^ x293;
  assign n8437 = n8413 ^ n8355;
  assign n8438 = n8437 ^ x294;
  assign n8439 = n8412 ^ n8411;
  assign n8440 = n8439 ^ x295;
  assign n8441 = n8410 ^ n8409;
  assign n8442 = n8441 ^ x296;
  assign n8443 = n8408 ^ n8406;
  assign n8444 = n8443 ^ x297;
  assign n8445 = n8405 ^ n8404;
  assign n8446 = n8445 ^ x298;
  assign n8537 = n8536 ^ n8447;
  assign n8538 = n8448 & ~n8537;
  assign n8539 = n8538 ^ x299;
  assign n8540 = n8539 ^ n8445;
  assign n8541 = ~n8446 & n8540;
  assign n8542 = n8541 ^ x298;
  assign n8543 = n8542 ^ n8443;
  assign n8544 = n8444 & ~n8543;
  assign n8545 = n8544 ^ x297;
  assign n8546 = n8545 ^ n8441;
  assign n8547 = n8442 & ~n8546;
  assign n8548 = n8547 ^ x296;
  assign n8549 = n8548 ^ n8439;
  assign n8550 = ~n8440 & n8549;
  assign n8551 = n8550 ^ x295;
  assign n8552 = n8551 ^ n8437;
  assign n8553 = ~n8438 & n8552;
  assign n8554 = n8553 ^ x294;
  assign n8555 = n8554 ^ n8435;
  assign n8556 = ~n8436 & n8555;
  assign n8557 = n8556 ^ x293;
  assign n8558 = n8557 ^ n8433;
  assign n8559 = ~n8434 & n8558;
  assign n8560 = n8559 ^ x292;
  assign n8561 = n8560 ^ n8431;
  assign n8562 = ~n8432 & n8561;
  assign n8563 = n8562 ^ x291;
  assign n8430 = n8419 ^ n8350;
  assign n8564 = n8563 ^ n8430;
  assign n8565 = n8430 ^ x290;
  assign n8566 = n8564 & ~n8565;
  assign n8567 = n8566 ^ x290;
  assign n8568 = n8567 ^ n8428;
  assign n8569 = n8429 & ~n8568;
  assign n8570 = n8569 ^ x289;
  assign n8571 = n8570 ^ x288;
  assign n8423 = n8197 ^ n4960;
  assign n8424 = n8346 ^ n8197;
  assign n8425 = ~n8423 & n8424;
  assign n8426 = n8425 ^ n4960;
  assign n8421 = n8348 & ~n8420;
  assign n8193 = n8192 ^ n8188;
  assign n8194 = n8189 & ~n8193;
  assign n8195 = n8194 ^ n8192;
  assign n7915 = n7787 ^ n7693;
  assign n7912 = n6351 ^ n6048;
  assign n7913 = ~n7263 & ~n7912;
  assign n7914 = n7913 ^ n6048;
  assign n7916 = n7915 ^ n7914;
  assign n7917 = n7916 ^ n4955;
  assign n8196 = n8195 ^ n7917;
  assign n8422 = n8421 ^ n8196;
  assign n8427 = n8426 ^ n8422;
  assign n8572 = n8571 ^ n8427;
  assign n8576 = n8575 ^ n8572;
  assign n8579 = n7432 ^ n6330;
  assign n8580 = n8028 & n8579;
  assign n8581 = n8580 ^ n6330;
  assign n8577 = n8567 ^ x289;
  assign n8578 = n8577 ^ n8428;
  assign n8582 = n8581 ^ n8578;
  assign n8584 = n7434 ^ n5990;
  assign n8585 = n8033 & ~n8584;
  assign n8586 = n8585 ^ n5990;
  assign n8583 = n8564 ^ x290;
  assign n8587 = n8586 ^ n8583;
  assign n8591 = n8560 ^ n8432;
  assign n8588 = n7443 ^ n5997;
  assign n8589 = n8038 & ~n8588;
  assign n8590 = n8589 ^ n5997;
  assign n8592 = n8591 ^ n8590;
  assign n8593 = n8557 ^ x292;
  assign n8594 = n8593 ^ n8433;
  assign n8595 = n7370 ^ n6343;
  assign n8596 = n8039 & n8595;
  assign n8597 = n8596 ^ n6343;
  assign n8598 = ~n8594 & ~n8597;
  assign n8599 = n8598 ^ n8591;
  assign n8600 = n8592 & ~n8599;
  assign n8601 = n8600 ^ n8598;
  assign n8602 = n8601 ^ n8583;
  assign n8603 = ~n8587 & n8602;
  assign n8604 = n8603 ^ n8586;
  assign n8605 = n8604 ^ n8578;
  assign n8606 = n8582 & ~n8605;
  assign n8607 = n8606 ^ n8581;
  assign n8608 = n8607 ^ n8572;
  assign n8609 = ~n8576 & ~n8608;
  assign n8610 = n8609 ^ n8575;
  assign n8611 = n8610 ^ n7910;
  assign n8612 = n7911 & ~n8611;
  assign n8613 = n8612 ^ n7909;
  assign n8614 = n8613 ^ n7903;
  assign n8615 = ~n7904 & n8614;
  assign n8616 = n8615 ^ n7902;
  assign n8617 = n8616 ^ n7897;
  assign n8618 = ~n7898 & ~n8617;
  assign n8619 = n8618 ^ n7379;
  assign n8669 = n8621 ^ n8619;
  assign n8670 = ~n8625 & n8669;
  assign n8671 = n8670 ^ n8624;
  assign n8702 = n8675 ^ n8671;
  assign n8703 = n8676 & ~n8702;
  assign n8704 = n8703 ^ n8674;
  assign n8770 = n8709 ^ n8704;
  assign n8771 = ~n8710 & n8770;
  assign n8772 = n8771 ^ n8707;
  assign n8858 = n8776 ^ n8772;
  assign n8859 = ~n8777 & ~n8858;
  assign n8860 = n8859 ^ n8775;
  assign n8861 = n8860 ^ n8856;
  assign n8862 = n8857 & n8861;
  assign n8863 = n8862 ^ n8854;
  assign n8848 = n7489 ^ n6269;
  assign n8849 = n7978 & n8848;
  assign n8850 = n8849 ^ n6269;
  assign n8846 = n8498 ^ x311;
  assign n8847 = n8846 ^ n8469;
  assign n8851 = n8850 ^ n8847;
  assign n8931 = n8863 ^ n8851;
  assign n8932 = n8931 ^ n6297;
  assign n8933 = n8860 ^ n8857;
  assign n8934 = n8933 ^ n6303;
  assign n8778 = n8777 ^ n8772;
  assign n8779 = n8778 ^ n6309;
  assign n8711 = n8710 ^ n8704;
  assign n8712 = n8711 ^ n6317;
  assign n8677 = n8676 ^ n8671;
  assign n8678 = n8677 ^ n6168;
  assign n8626 = n8625 ^ n8619;
  assign n8627 = n8626 ^ n6098;
  assign n8628 = n8616 ^ n7898;
  assign n8629 = n8628 ^ n6088;
  assign n8630 = n8613 ^ n7904;
  assign n8631 = n8630 ^ n6014;
  assign n8632 = n8610 ^ n7911;
  assign n8633 = n8632 ^ n6019;
  assign n8634 = n8607 ^ n8576;
  assign n8635 = n8634 ^ n5992;
  assign n8636 = n8604 ^ n8582;
  assign n8637 = n8636 ^ n6000;
  assign n8638 = n8601 ^ n8587;
  assign n8639 = n8638 ^ n6032;
  assign n8640 = n8597 ^ n8594;
  assign n8641 = n6043 & n8640;
  assign n8642 = n8641 ^ n6037;
  assign n8643 = n8598 ^ n8590;
  assign n8644 = n8643 ^ n8591;
  assign n8645 = n8644 ^ n8641;
  assign n8646 = ~n8642 & n8645;
  assign n8647 = n8646 ^ n6037;
  assign n8648 = n8647 ^ n8638;
  assign n8649 = ~n8639 & ~n8648;
  assign n8650 = n8649 ^ n6032;
  assign n8651 = n8650 ^ n8636;
  assign n8652 = n8637 & ~n8651;
  assign n8653 = n8652 ^ n6000;
  assign n8654 = n8653 ^ n8634;
  assign n8655 = n8635 & n8654;
  assign n8656 = n8655 ^ n5992;
  assign n8657 = n8656 ^ n8632;
  assign n8658 = ~n8633 & ~n8657;
  assign n8659 = n8658 ^ n6019;
  assign n8660 = n8659 ^ n8630;
  assign n8661 = n8631 & ~n8660;
  assign n8662 = n8661 ^ n6014;
  assign n8663 = n8662 ^ n8628;
  assign n8664 = ~n8629 & ~n8663;
  assign n8665 = n8664 ^ n6088;
  assign n8666 = n8665 ^ n8626;
  assign n8667 = ~n8627 & ~n8666;
  assign n8668 = n8667 ^ n6098;
  assign n8699 = n8677 ^ n8668;
  assign n8700 = n8678 & ~n8699;
  assign n8701 = n8700 ^ n6168;
  assign n8767 = n8711 ^ n8701;
  assign n8768 = ~n8712 & n8767;
  assign n8769 = n8768 ^ n6317;
  assign n8935 = n8778 ^ n8769;
  assign n8936 = n8779 & n8935;
  assign n8937 = n8936 ^ n6309;
  assign n8938 = n8937 ^ n8933;
  assign n8939 = ~n8934 & ~n8938;
  assign n8940 = n8939 ^ n6303;
  assign n8941 = n8940 ^ n8931;
  assign n8942 = n8932 & n8941;
  assign n8943 = n8942 ^ n6297;
  assign n8864 = n8863 ^ n8847;
  assign n8865 = ~n8851 & ~n8864;
  assign n8866 = n8865 ^ n8850;
  assign n8842 = n7570 ^ n6261;
  assign n8843 = n7975 & ~n8842;
  assign n8844 = n8843 ^ n6261;
  assign n8840 = n8501 ^ x310;
  assign n8841 = n8840 ^ n8467;
  assign n8845 = n8844 ^ n8841;
  assign n8929 = n8866 ^ n8845;
  assign n8930 = n8929 ^ n6290;
  assign n9002 = n8943 ^ n8930;
  assign n8679 = n8678 ^ n8668;
  assign n8680 = n8665 ^ n8627;
  assign n8681 = n8662 ^ n8629;
  assign n8682 = n8659 ^ n8631;
  assign n8683 = n8653 ^ n8635;
  assign n8684 = n8640 ^ n6043;
  assign n8685 = n8644 ^ n8642;
  assign n8686 = n8684 & n8685;
  assign n8687 = n8647 ^ n6032;
  assign n8688 = n8687 ^ n8638;
  assign n8689 = n8686 & n8688;
  assign n8690 = n8650 ^ n8637;
  assign n8691 = ~n8689 & ~n8690;
  assign n8692 = ~n8683 & n8691;
  assign n8693 = n8656 ^ n8633;
  assign n8694 = ~n8692 & n8693;
  assign n8695 = n8682 & n8694;
  assign n8696 = n8681 & ~n8695;
  assign n8697 = ~n8680 & n8696;
  assign n8698 = n8679 & ~n8697;
  assign n8713 = n8712 ^ n8701;
  assign n8766 = n8698 & ~n8713;
  assign n8780 = n8779 ^ n8769;
  assign n8997 = ~n8766 & ~n8780;
  assign n8998 = n8937 ^ n8934;
  assign n8999 = n8997 & ~n8998;
  assign n9000 = n8940 ^ n8932;
  assign n9001 = n8999 & ~n9000;
  assign n9065 = n9002 ^ n9001;
  assign n9066 = n9065 ^ x337;
  assign n9067 = n9000 ^ n8999;
  assign n9068 = n9067 ^ x338;
  assign n9069 = n8998 ^ n8997;
  assign n9070 = n9069 ^ x339;
  assign n8781 = n8780 ^ n8766;
  assign n9071 = n8781 ^ x340;
  assign n8714 = n8713 ^ n8698;
  assign n8715 = n8714 ^ x341;
  assign n8716 = n8697 ^ n8679;
  assign n8717 = n8716 ^ x342;
  assign n8718 = n8696 ^ n8680;
  assign n8719 = n8718 ^ x343;
  assign n8720 = n8695 ^ n8681;
  assign n8721 = n8720 ^ x344;
  assign n8722 = n8694 ^ n8682;
  assign n8723 = n8722 ^ x345;
  assign n8724 = n8693 ^ n8692;
  assign n8725 = n8724 ^ x346;
  assign n8726 = n8691 ^ n8683;
  assign n8727 = n8726 ^ x347;
  assign n8728 = n8690 ^ n8689;
  assign n8729 = n8728 ^ x348;
  assign n8730 = n8688 ^ n8686;
  assign n8731 = n8730 ^ x349;
  assign n8732 = x351 & ~n8684;
  assign n8733 = n8732 ^ x350;
  assign n8734 = n8685 ^ n8684;
  assign n8735 = n8734 ^ n8732;
  assign n8736 = n8733 & ~n8735;
  assign n8737 = n8736 ^ x350;
  assign n8738 = n8737 ^ n8730;
  assign n8739 = n8731 & ~n8738;
  assign n8740 = n8739 ^ x349;
  assign n8741 = n8740 ^ n8728;
  assign n8742 = ~n8729 & n8741;
  assign n8743 = n8742 ^ x348;
  assign n8744 = n8743 ^ n8726;
  assign n8745 = n8727 & ~n8744;
  assign n8746 = n8745 ^ x347;
  assign n8747 = n8746 ^ n8724;
  assign n8748 = ~n8725 & n8747;
  assign n8749 = n8748 ^ x346;
  assign n8750 = n8749 ^ n8722;
  assign n8751 = n8723 & ~n8750;
  assign n8752 = n8751 ^ x345;
  assign n8753 = n8752 ^ n8720;
  assign n8754 = n8721 & ~n8753;
  assign n8755 = n8754 ^ x344;
  assign n8756 = n8755 ^ n8718;
  assign n8757 = n8719 & ~n8756;
  assign n8758 = n8757 ^ x343;
  assign n8759 = n8758 ^ n8716;
  assign n8760 = ~n8717 & n8759;
  assign n8761 = n8760 ^ x342;
  assign n8762 = n8761 ^ n8714;
  assign n8763 = ~n8715 & n8762;
  assign n8764 = n8763 ^ x341;
  assign n9072 = n8781 ^ n8764;
  assign n9073 = ~n9071 & n9072;
  assign n9074 = n9073 ^ x340;
  assign n9075 = n9074 ^ n9069;
  assign n9076 = n9070 & ~n9075;
  assign n9077 = n9076 ^ x339;
  assign n9078 = n9077 ^ n9067;
  assign n9079 = n9068 & ~n9078;
  assign n9080 = n9079 ^ x338;
  assign n9081 = n9080 ^ n9065;
  assign n9082 = n9066 & ~n9081;
  assign n9083 = n9082 ^ x337;
  assign n9410 = n9083 ^ x336;
  assign n9003 = n9001 & ~n9002;
  assign n8944 = n8943 ^ n8929;
  assign n8945 = ~n8930 & n8944;
  assign n8946 = n8945 ^ n6290;
  assign n8867 = n8866 ^ n8841;
  assign n8868 = ~n8845 & n8867;
  assign n8869 = n8868 ^ n8844;
  assign n8836 = n7618 ^ n6756;
  assign n8837 = n7970 & ~n8836;
  assign n8838 = n8837 ^ n6756;
  assign n8926 = n8869 ^ n8838;
  assign n8835 = n8504 ^ n8466;
  assign n8927 = n8926 ^ n8835;
  assign n8928 = n8927 ^ n6284;
  assign n8996 = n8946 ^ n8928;
  assign n9063 = n9003 ^ n8996;
  assign n9411 = n9410 ^ n9063;
  assign n9415 = n9414 ^ n9411;
  assign n8791 = n8533 ^ x300;
  assign n8792 = n8791 ^ n8449;
  assign n9417 = n7931 ^ n7689;
  assign n9418 = ~n8792 & ~n9417;
  assign n9419 = n9418 ^ n7689;
  assign n9416 = n9080 ^ n9066;
  assign n9420 = n9419 ^ n9416;
  assign n8797 = n8530 ^ n8452;
  assign n9423 = n7937 ^ n7671;
  assign n9424 = n8797 & ~n9423;
  assign n9425 = n9424 ^ n7671;
  assign n9421 = n9077 ^ x338;
  assign n9422 = n9421 ^ n9067;
  assign n9426 = n9425 ^ n9422;
  assign n9430 = n9074 ^ n9070;
  assign n8802 = n8527 ^ x302;
  assign n8803 = n8802 ^ n8453;
  assign n9427 = n7948 ^ n7651;
  assign n9428 = n8803 & n9427;
  assign n9429 = n9428 ^ n7651;
  assign n9431 = n9430 ^ n9429;
  assign n8808 = n8524 ^ x303;
  assign n9432 = n7953 ^ n7638;
  assign n9433 = ~n8808 & ~n9432;
  assign n9434 = n9433 ^ n7638;
  assign n8765 = n8764 ^ x340;
  assign n8782 = n8781 ^ n8765;
  assign n9435 = n9434 ^ n8782;
  assign n8813 = n8520 ^ x304;
  assign n8814 = n8813 ^ n8456;
  assign n9436 = n7959 ^ n7618;
  assign n9437 = n8814 & n9436;
  assign n9438 = n9437 ^ n7618;
  assign n9336 = n8761 ^ n8715;
  assign n9439 = n9438 ^ n9336;
  assign n8819 = n8517 ^ n8459;
  assign n9440 = n7964 ^ n7570;
  assign n9441 = ~n8819 & n9440;
  assign n9442 = n9441 ^ n7570;
  assign n9343 = n8758 ^ n8717;
  assign n9443 = n9442 ^ n9343;
  assign n8783 = n8514 ^ x306;
  assign n8784 = n8783 ^ n8460;
  assign n9444 = n7970 ^ n7489;
  assign n9445 = n8784 & ~n9444;
  assign n9446 = n9445 ^ n7489;
  assign n9351 = n8755 ^ x343;
  assign n9352 = n9351 ^ n8718;
  assign n9447 = n9446 ^ n9352;
  assign n8828 = n8511 ^ n8463;
  assign n9448 = n7975 ^ n7383;
  assign n9449 = n8828 & ~n9448;
  assign n9450 = n9449 ^ n7383;
  assign n9358 = n8752 ^ x344;
  assign n9359 = n9358 ^ n8720;
  assign n9451 = n9450 ^ n9359;
  assign n8830 = n8508 ^ x308;
  assign n9453 = n7978 ^ n7389;
  assign n9454 = ~n8830 & n9453;
  assign n9455 = n9454 ^ n7389;
  assign n9452 = n8749 ^ n8723;
  assign n9456 = n9455 ^ n9452;
  assign n9457 = n7986 ^ n7391;
  assign n9458 = n8835 & ~n9457;
  assign n9459 = n9458 ^ n7391;
  assign n9365 = n8746 ^ x346;
  assign n9366 = n9365 ^ n8724;
  assign n9460 = n9459 ^ n9366;
  assign n9462 = n7989 ^ n7400;
  assign n9463 = n8841 & ~n9462;
  assign n9464 = n9463 ^ n7400;
  assign n9461 = n8743 ^ n8727;
  assign n9465 = n9464 ^ n9461;
  assign n9468 = n7994 ^ n7405;
  assign n9469 = n8847 & n9468;
  assign n9470 = n9469 ^ n7405;
  assign n9466 = n8740 ^ x348;
  assign n9467 = n9466 ^ n8728;
  assign n9471 = n9470 ^ n9467;
  assign n9474 = n8002 ^ n7376;
  assign n9475 = n8856 & n9474;
  assign n9476 = n9475 ^ n7376;
  assign n9472 = n8737 ^ x349;
  assign n9473 = n9472 ^ n8730;
  assign n9477 = n9476 ^ n9473;
  assign n9327 = n8734 ^ n8733;
  assign n9324 = n8005 ^ n7415;
  assign n9325 = n8776 & n9324;
  assign n9326 = n9325 ^ n7415;
  assign n9328 = n9327 ^ n9326;
  assign n9286 = n8684 ^ x351;
  assign n9283 = n7421 ^ n7375;
  assign n9284 = ~n8709 & n9283;
  assign n9285 = n9284 ^ n7421;
  assign n9287 = n9286 ^ n9285;
  assign n9269 = n7899 ^ n7423;
  assign n9270 = n8675 & ~n9269;
  assign n9271 = n9270 ^ n7423;
  assign n9173 = n7263 ^ n6667;
  assign n9174 = n7883 & n9173;
  assign n9175 = n9174 ^ n6667;
  assign n9138 = n8545 ^ x296;
  assign n9139 = n9138 ^ n8441;
  assign n9134 = n7212 ^ n6672;
  assign n9135 = ~n7847 & n9134;
  assign n9136 = n9135 ^ n6672;
  assign n9168 = n9139 ^ n9136;
  assign n9037 = n8542 ^ n8444;
  assign n9033 = n7215 ^ n6677;
  assign n9034 = n7810 & ~n9033;
  assign n9035 = n9034 ^ n6677;
  assign n9130 = n9037 ^ n9035;
  assign n8900 = n7226 ^ n6687;
  assign n8901 = ~n8188 & ~n8900;
  assign n8902 = n8901 ^ n6687;
  assign n8987 = n8904 ^ n8902;
  assign n8788 = n7932 ^ n7244;
  assign n8789 = ~n7918 & n8788;
  assign n8790 = n8789 ^ n7244;
  assign n8793 = n8792 ^ n8790;
  assign n8794 = n7939 ^ n7052;
  assign n8795 = n7920 & ~n8794;
  assign n8796 = n8795 ^ n7052;
  assign n8798 = n8797 ^ n8796;
  assign n8799 = n7865 ^ n7035;
  assign n8800 = n7925 & ~n8799;
  assign n8801 = n8800 ^ n7035;
  assign n8804 = n8803 ^ n8801;
  assign n8805 = n7834 ^ n7021;
  assign n8806 = ~n7931 & n8805;
  assign n8807 = n8806 ^ n7021;
  assign n8809 = n8808 ^ n8807;
  assign n8810 = n7806 ^ n7008;
  assign n8811 = n7937 & ~n8810;
  assign n8812 = n8811 ^ n7008;
  assign n8815 = n8814 ^ n8812;
  assign n8816 = n7689 ^ n6991;
  assign n8817 = n7948 & ~n8816;
  assign n8818 = n8817 ^ n6991;
  assign n8820 = n8819 ^ n8818;
  assign n8821 = n7671 ^ n6973;
  assign n8822 = ~n7953 & n8821;
  assign n8823 = n8822 ^ n6973;
  assign n8824 = n8823 ^ n8784;
  assign n8825 = n7651 ^ n6958;
  assign n8826 = n7959 & ~n8825;
  assign n8827 = n8826 ^ n6958;
  assign n8829 = n8828 ^ n8827;
  assign n8831 = n7638 ^ n6885;
  assign n8832 = n7964 & n8831;
  assign n8833 = n8832 ^ n6885;
  assign n8834 = n8833 ^ n8830;
  assign n8839 = n8838 ^ n8835;
  assign n8870 = n8869 ^ n8835;
  assign n8871 = ~n8839 & n8870;
  assign n8872 = n8871 ^ n8838;
  assign n8873 = n8872 ^ n8830;
  assign n8874 = ~n8834 & ~n8873;
  assign n8875 = n8874 ^ n8833;
  assign n8876 = n8875 ^ n8828;
  assign n8877 = ~n8829 & ~n8876;
  assign n8878 = n8877 ^ n8827;
  assign n8879 = n8878 ^ n8784;
  assign n8880 = ~n8824 & n8879;
  assign n8881 = n8880 ^ n8823;
  assign n8882 = n8881 ^ n8819;
  assign n8883 = n8820 & ~n8882;
  assign n8884 = n8883 ^ n8818;
  assign n8885 = n8884 ^ n8814;
  assign n8886 = ~n8815 & n8885;
  assign n8887 = n8886 ^ n8812;
  assign n8888 = n8887 ^ n8808;
  assign n8889 = ~n8809 & ~n8888;
  assign n8890 = n8889 ^ n8807;
  assign n8891 = n8890 ^ n8803;
  assign n8892 = ~n8804 & ~n8891;
  assign n8893 = n8892 ^ n8801;
  assign n8894 = n8893 ^ n8797;
  assign n8895 = ~n8798 & n8894;
  assign n8896 = n8895 ^ n8796;
  assign n8897 = n8896 ^ n8792;
  assign n8898 = ~n8793 & ~n8897;
  assign n8899 = n8898 ^ n8790;
  assign n8988 = n8904 ^ n8899;
  assign n8989 = ~n8987 & ~n8988;
  assign n8990 = n8989 ^ n8902;
  assign n8984 = n8539 ^ x298;
  assign n8985 = n8984 ^ n8445;
  assign n9029 = n8990 ^ n8985;
  assign n8981 = n7220 ^ n6682;
  assign n8982 = n7915 & ~n8981;
  assign n8983 = n8982 ^ n6682;
  assign n9030 = n8990 ^ n8983;
  assign n9031 = n9029 & ~n9030;
  assign n9032 = n9031 ^ n8985;
  assign n9131 = n9037 ^ n9032;
  assign n9132 = n9130 & n9131;
  assign n9133 = n9132 ^ n9035;
  assign n9169 = n9139 ^ n9133;
  assign n9170 = n9168 & ~n9169;
  assign n9171 = n9170 ^ n9136;
  assign n9167 = n8548 ^ n8440;
  assign n9172 = n9171 ^ n9167;
  assign n9176 = n9175 ^ n9172;
  assign n9221 = n9176 ^ n5980;
  assign n9137 = n9136 ^ n9133;
  assign n9140 = n9139 ^ n9137;
  assign n9162 = n9140 ^ n5928;
  assign n9036 = n9035 ^ n9032;
  assign n9038 = n9037 ^ n9036;
  assign n9125 = n9038 ^ n5886;
  assign n8986 = n8985 ^ n8983;
  assign n8991 = n8990 ^ n8986;
  assign n9024 = n8991 ^ n5852;
  assign n8903 = n8902 ^ n8899;
  assign n8905 = n8904 ^ n8903;
  assign n8906 = n8905 ^ n5796;
  assign n8907 = n8896 ^ n8793;
  assign n8908 = n8907 ^ n6578;
  assign n8909 = n8893 ^ n8798;
  assign n8910 = n8909 ^ n6562;
  assign n8911 = n8890 ^ n8804;
  assign n8912 = n8911 ^ n6358;
  assign n8913 = n8887 ^ n8809;
  assign n8914 = n8913 ^ n6360;
  assign n8915 = n8884 ^ n8815;
  assign n8916 = n8915 ^ n6366;
  assign n8917 = n8881 ^ n8820;
  assign n8918 = n8917 ^ n6004;
  assign n8919 = n8878 ^ n8824;
  assign n8920 = n8919 ^ n6264;
  assign n8921 = n8875 ^ n8829;
  assign n8922 = n8921 ^ n6271;
  assign n8923 = n8872 ^ n8833;
  assign n8924 = n8923 ^ n8830;
  assign n8925 = n8924 ^ n6277;
  assign n8947 = n8946 ^ n8927;
  assign n8948 = n8928 & n8947;
  assign n8949 = n8948 ^ n6284;
  assign n8950 = n8949 ^ n8924;
  assign n8951 = ~n8925 & ~n8950;
  assign n8952 = n8951 ^ n6277;
  assign n8953 = n8952 ^ n8921;
  assign n8954 = ~n8922 & ~n8953;
  assign n8955 = n8954 ^ n6271;
  assign n8956 = n8955 ^ n8919;
  assign n8957 = n8920 & ~n8956;
  assign n8958 = n8957 ^ n6264;
  assign n8959 = n8958 ^ n8917;
  assign n8960 = ~n8918 & n8959;
  assign n8961 = n8960 ^ n6004;
  assign n8962 = n8961 ^ n8915;
  assign n8963 = ~n8916 & ~n8962;
  assign n8964 = n8963 ^ n6366;
  assign n8965 = n8964 ^ n8913;
  assign n8966 = ~n8914 & n8965;
  assign n8967 = n8966 ^ n6360;
  assign n8968 = n8967 ^ n8911;
  assign n8969 = n8912 & ~n8968;
  assign n8970 = n8969 ^ n6358;
  assign n8971 = n8970 ^ n8909;
  assign n8972 = ~n8910 & n8971;
  assign n8973 = n8972 ^ n6562;
  assign n8974 = n8973 ^ n8907;
  assign n8975 = ~n8908 & n8974;
  assign n8976 = n8975 ^ n6578;
  assign n8977 = n8976 ^ n8905;
  assign n8978 = n8906 & ~n8977;
  assign n8979 = n8978 ^ n5796;
  assign n9025 = n8991 ^ n8979;
  assign n9026 = n9024 & ~n9025;
  assign n9027 = n9026 ^ n5852;
  assign n9126 = n9038 ^ n9027;
  assign n9127 = n9125 & ~n9126;
  assign n9128 = n9127 ^ n5886;
  assign n9163 = n9140 ^ n9128;
  assign n9164 = n9162 & n9163;
  assign n9165 = n9164 ^ n5928;
  assign n9222 = n9176 ^ n9165;
  assign n9223 = n9221 & ~n9222;
  assign n9224 = n9223 ^ n5980;
  assign n9225 = n9224 ^ n6053;
  assign n9217 = n7267 ^ n6356;
  assign n9218 = n8070 & ~n9217;
  assign n9219 = n9218 ^ n6356;
  assign n9213 = n9175 ^ n9167;
  assign n9214 = n9172 & n9213;
  assign n9215 = n9214 ^ n9175;
  assign n9211 = n8551 ^ x294;
  assign n9212 = n9211 ^ n8437;
  assign n9216 = n9215 ^ n9212;
  assign n9220 = n9219 ^ n9216;
  assign n9226 = n9225 ^ n9220;
  assign n9166 = n9165 ^ n5980;
  assign n9177 = n9176 ^ n9166;
  assign n8980 = n8979 ^ n5852;
  assign n8992 = n8991 ^ n8980;
  assign n8993 = n8964 ^ n8914;
  assign n8994 = n8961 ^ n8916;
  assign n8995 = n8952 ^ n8922;
  assign n9004 = ~n8996 & ~n9003;
  assign n9005 = n8949 ^ n8925;
  assign n9006 = n9004 & ~n9005;
  assign n9007 = ~n8995 & ~n9006;
  assign n9008 = n8955 ^ n8920;
  assign n9009 = ~n9007 & n9008;
  assign n9010 = n8958 ^ n6004;
  assign n9011 = n9010 ^ n8917;
  assign n9012 = n9009 & ~n9011;
  assign n9013 = ~n8994 & n9012;
  assign n9014 = n8993 & n9013;
  assign n9015 = n8967 ^ n8912;
  assign n9016 = n9014 & ~n9015;
  assign n9017 = n8970 ^ n8910;
  assign n9018 = ~n9016 & ~n9017;
  assign n9019 = n8973 ^ n8908;
  assign n9020 = ~n9018 & n9019;
  assign n9021 = n8976 ^ n8906;
  assign n9022 = ~n9020 & n9021;
  assign n9023 = ~n8992 & ~n9022;
  assign n9028 = n9027 ^ n5886;
  assign n9039 = n9038 ^ n9028;
  assign n9124 = ~n9023 & n9039;
  assign n9129 = n9128 ^ n5928;
  assign n9141 = n9140 ^ n9129;
  assign n9178 = n9124 & n9141;
  assign n9210 = n9177 & ~n9178;
  assign n9227 = n9226 ^ n9210;
  assign n9263 = n9227 ^ x321;
  assign n9179 = n9178 ^ n9177;
  assign n9205 = n9179 ^ x322;
  assign n9142 = n9141 ^ n9124;
  assign n9143 = n9142 ^ x323;
  assign n9040 = n9039 ^ n9023;
  assign n9041 = n9040 ^ x324;
  assign n9042 = n9022 ^ n8992;
  assign n9043 = n9042 ^ x325;
  assign n9044 = n9021 ^ n9020;
  assign n9045 = n9044 ^ x326;
  assign n9046 = n9019 ^ n9018;
  assign n9047 = n9046 ^ x327;
  assign n9048 = n9017 ^ n9016;
  assign n9049 = n9048 ^ x328;
  assign n9050 = n9015 ^ n9014;
  assign n9051 = n9050 ^ x329;
  assign n9052 = n9013 ^ n8993;
  assign n9053 = n9052 ^ x330;
  assign n9054 = n9012 ^ n8994;
  assign n9055 = n9054 ^ x331;
  assign n9056 = n9011 ^ n9009;
  assign n9057 = n9056 ^ x332;
  assign n9058 = n9008 ^ n9007;
  assign n9059 = n9058 ^ x333;
  assign n9060 = n9006 ^ n8995;
  assign n9061 = n9060 ^ x334;
  assign n9064 = n9063 ^ x336;
  assign n9084 = n9083 ^ n9063;
  assign n9085 = n9064 & ~n9084;
  assign n9086 = n9085 ^ x336;
  assign n9062 = n9005 ^ n9004;
  assign n9087 = n9086 ^ n9062;
  assign n9088 = n9062 ^ x335;
  assign n9089 = n9087 & ~n9088;
  assign n9090 = n9089 ^ x335;
  assign n9091 = n9090 ^ n9060;
  assign n9092 = ~n9061 & n9091;
  assign n9093 = n9092 ^ x334;
  assign n9094 = n9093 ^ n9058;
  assign n9095 = ~n9059 & n9094;
  assign n9096 = n9095 ^ x333;
  assign n9097 = n9096 ^ n9056;
  assign n9098 = ~n9057 & n9097;
  assign n9099 = n9098 ^ x332;
  assign n9100 = n9099 ^ n9054;
  assign n9101 = ~n9055 & n9100;
  assign n9102 = n9101 ^ x331;
  assign n9103 = n9102 ^ n9052;
  assign n9104 = n9053 & ~n9103;
  assign n9105 = n9104 ^ x330;
  assign n9106 = n9105 ^ n9050;
  assign n9107 = ~n9051 & n9106;
  assign n9108 = n9107 ^ x329;
  assign n9109 = n9108 ^ n9048;
  assign n9110 = ~n9049 & n9109;
  assign n9111 = n9110 ^ x328;
  assign n9112 = n9111 ^ n9046;
  assign n9113 = ~n9047 & n9112;
  assign n9114 = n9113 ^ x327;
  assign n9115 = n9114 ^ n9044;
  assign n9116 = n9045 & ~n9115;
  assign n9117 = n9116 ^ x326;
  assign n9118 = n9117 ^ n9042;
  assign n9119 = n9043 & ~n9118;
  assign n9120 = n9119 ^ x325;
  assign n9121 = n9120 ^ n9040;
  assign n9122 = n9041 & ~n9121;
  assign n9123 = n9122 ^ x324;
  assign n9158 = n9142 ^ n9123;
  assign n9159 = ~n9143 & n9158;
  assign n9160 = n9159 ^ x323;
  assign n9206 = n9179 ^ n9160;
  assign n9207 = ~n9205 & n9206;
  assign n9208 = n9207 ^ x322;
  assign n9264 = n9227 ^ n9208;
  assign n9265 = n9263 & ~n9264;
  assign n9266 = n9265 ^ x321;
  assign n9267 = n9266 ^ x320;
  assign n9258 = n9220 ^ n6053;
  assign n9259 = n9224 ^ n9220;
  assign n9260 = ~n9258 & n9259;
  assign n9261 = n9260 ^ n6053;
  assign n9256 = ~n9210 & n9226;
  assign n9252 = n9219 ^ n9212;
  assign n9253 = ~n9216 & n9252;
  assign n9254 = n9253 ^ n9219;
  assign n9247 = n7306 ^ n6351;
  assign n9248 = n8100 & n9247;
  assign n9249 = n9248 ^ n6351;
  assign n9246 = n8554 ^ n8436;
  assign n9250 = n9249 ^ n9246;
  assign n9251 = n9250 ^ n6048;
  assign n9255 = n9254 ^ n9251;
  assign n9257 = n9256 ^ n9255;
  assign n9262 = n9261 ^ n9257;
  assign n9268 = n9267 ^ n9262;
  assign n9272 = n9271 ^ n9268;
  assign n9209 = n9208 ^ x321;
  assign n9228 = n9227 ^ n9209;
  assign n9201 = n7906 ^ n7432;
  assign n9202 = ~n8621 & ~n9201;
  assign n9203 = n9202 ^ n7432;
  assign n9242 = n9228 ^ n9203;
  assign n9181 = n8022 ^ n7434;
  assign n9182 = ~n7897 & n9181;
  assign n9183 = n9182 ^ n7434;
  assign n9161 = n9160 ^ x322;
  assign n9180 = n9179 ^ n9161;
  assign n9184 = n9183 ^ n9180;
  assign n9145 = n8028 ^ n7443;
  assign n9146 = n7903 & ~n9145;
  assign n9147 = n9146 ^ n7443;
  assign n9144 = n9143 ^ n9123;
  assign n9148 = n9147 ^ n9144;
  assign n9149 = n9120 ^ x324;
  assign n9150 = n9149 ^ n9040;
  assign n9151 = n8033 ^ n7370;
  assign n9152 = ~n7910 & ~n9151;
  assign n9153 = n9152 ^ n7370;
  assign n9154 = n9150 & ~n9153;
  assign n9155 = n9154 ^ n9144;
  assign n9156 = ~n9148 & ~n9155;
  assign n9157 = n9156 ^ n9154;
  assign n9198 = n9180 ^ n9157;
  assign n9199 = n9184 & n9198;
  assign n9200 = n9199 ^ n9183;
  assign n9243 = n9228 ^ n9200;
  assign n9244 = n9242 & n9243;
  assign n9245 = n9244 ^ n9203;
  assign n9280 = n9268 ^ n9245;
  assign n9281 = n9272 & ~n9280;
  assign n9282 = n9281 ^ n9271;
  assign n9321 = n9286 ^ n9282;
  assign n9322 = ~n9287 & n9321;
  assign n9323 = n9322 ^ n9285;
  assign n9478 = n9327 ^ n9323;
  assign n9479 = ~n9328 & ~n9478;
  assign n9480 = n9479 ^ n9326;
  assign n9481 = n9480 ^ n9473;
  assign n9482 = n9477 & n9481;
  assign n9483 = n9482 ^ n9476;
  assign n9484 = n9483 ^ n9467;
  assign n9485 = ~n9471 & n9484;
  assign n9486 = n9485 ^ n9470;
  assign n9487 = n9486 ^ n9461;
  assign n9488 = ~n9465 & ~n9487;
  assign n9489 = n9488 ^ n9464;
  assign n9490 = n9489 ^ n9366;
  assign n9491 = ~n9460 & ~n9490;
  assign n9492 = n9491 ^ n9459;
  assign n9493 = n9492 ^ n9452;
  assign n9494 = n9456 & ~n9493;
  assign n9495 = n9494 ^ n9455;
  assign n9496 = n9495 ^ n9359;
  assign n9497 = ~n9451 & ~n9496;
  assign n9498 = n9497 ^ n9450;
  assign n9499 = n9498 ^ n9352;
  assign n9500 = ~n9447 & n9499;
  assign n9501 = n9500 ^ n9446;
  assign n9502 = n9501 ^ n9343;
  assign n9503 = ~n9443 & ~n9502;
  assign n9504 = n9503 ^ n9442;
  assign n9505 = n9504 ^ n9336;
  assign n9506 = ~n9439 & n9505;
  assign n9507 = n9506 ^ n9438;
  assign n9508 = n9507 ^ n8782;
  assign n9509 = ~n9435 & n9508;
  assign n9510 = n9509 ^ n9434;
  assign n9511 = n9510 ^ n9430;
  assign n9512 = n9431 & ~n9511;
  assign n9513 = n9512 ^ n9429;
  assign n9514 = n9513 ^ n9422;
  assign n9515 = ~n9426 & ~n9514;
  assign n9516 = n9515 ^ n9425;
  assign n9517 = n9516 ^ n9416;
  assign n9518 = n9420 & n9517;
  assign n9519 = n9518 ^ n9419;
  assign n9520 = n9519 ^ n9411;
  assign n9521 = n9415 & ~n9520;
  assign n9522 = n9521 ^ n9414;
  assign n9409 = n9087 ^ x335;
  assign n9523 = n9522 ^ n9409;
  assign n9524 = n7920 ^ n7834;
  assign n9525 = ~n8985 & n9524;
  assign n9526 = n9525 ^ n7834;
  assign n9527 = n9526 ^ n9409;
  assign n9528 = n9523 & ~n9527;
  assign n9529 = n9528 ^ n9526;
  assign n9405 = n7918 ^ n7865;
  assign n9406 = n9037 & ~n9405;
  assign n9407 = n9406 ^ n7865;
  assign n9403 = n9090 ^ x334;
  assign n9404 = n9403 ^ n9060;
  assign n9408 = n9407 ^ n9404;
  assign n9593 = n9529 ^ n9408;
  assign n9594 = n9593 ^ n7035;
  assign n9595 = n9526 ^ n9523;
  assign n9596 = n9595 ^ n7021;
  assign n9597 = n9519 ^ n9414;
  assign n9598 = n9597 ^ n9411;
  assign n9599 = n9598 ^ n7008;
  assign n9600 = n9516 ^ n9420;
  assign n9601 = n9600 ^ n6991;
  assign n9602 = n9513 ^ n9426;
  assign n9603 = n9602 ^ n6973;
  assign n9604 = n9510 ^ n9431;
  assign n9605 = n9604 ^ n6958;
  assign n9606 = n9507 ^ n9435;
  assign n9607 = n9606 ^ n6885;
  assign n9608 = n9504 ^ n9438;
  assign n9609 = n9608 ^ n9336;
  assign n9610 = n9609 ^ n6756;
  assign n9611 = n9501 ^ n9443;
  assign n9612 = n9611 ^ n6261;
  assign n9613 = n9498 ^ n9446;
  assign n9614 = n9613 ^ n9352;
  assign n9615 = n9614 ^ n6269;
  assign n9616 = n9495 ^ n9451;
  assign n9617 = n9616 ^ n6275;
  assign n9618 = n9492 ^ n9455;
  assign n9619 = n9618 ^ n9452;
  assign n9620 = n9619 ^ n6282;
  assign n9621 = n9489 ^ n9460;
  assign n9622 = n9621 ^ n6288;
  assign n9623 = n9486 ^ n9464;
  assign n9624 = n9623 ^ n9461;
  assign n9625 = n9624 ^ n6295;
  assign n9626 = n9483 ^ n9470;
  assign n9627 = n9626 ^ n9467;
  assign n9628 = n9627 ^ n6301;
  assign n9629 = n9480 ^ n9476;
  assign n9630 = n9629 ^ n9473;
  assign n9631 = n9630 ^ n6307;
  assign n9329 = n9328 ^ n9323;
  assign n9330 = n9329 ^ n6314;
  assign n9288 = n9287 ^ n9282;
  assign n9289 = n9288 ^ n6322;
  assign n9273 = n9272 ^ n9245;
  assign n9274 = n9273 ^ n6324;
  assign n9204 = n9203 ^ n9200;
  assign n9229 = n9228 ^ n9204;
  assign n9230 = n9229 ^ n6330;
  assign n9185 = n9184 ^ n9157;
  assign n9186 = n9185 ^ n5990;
  assign n9187 = n9153 ^ n9150;
  assign n9188 = ~n6343 & ~n9187;
  assign n9189 = n9188 ^ n5997;
  assign n9190 = n9154 ^ n9147;
  assign n9191 = n9190 ^ n9144;
  assign n9192 = n9191 ^ n9188;
  assign n9193 = n9189 & ~n9192;
  assign n9194 = n9193 ^ n5997;
  assign n9195 = n9194 ^ n9185;
  assign n9196 = n9186 & ~n9195;
  assign n9197 = n9196 ^ n5990;
  assign n9239 = n9229 ^ n9197;
  assign n9240 = ~n9230 & n9239;
  assign n9241 = n9240 ^ n6330;
  assign n9277 = n9273 ^ n9241;
  assign n9278 = ~n9274 & ~n9277;
  assign n9279 = n9278 ^ n6324;
  assign n9318 = n9288 ^ n9279;
  assign n9319 = n9289 & ~n9318;
  assign n9320 = n9319 ^ n6322;
  assign n9632 = n9329 ^ n9320;
  assign n9633 = n9330 & ~n9632;
  assign n9634 = n9633 ^ n6314;
  assign n9635 = n9634 ^ n9630;
  assign n9636 = ~n9631 & ~n9635;
  assign n9637 = n9636 ^ n6307;
  assign n9638 = n9637 ^ n9627;
  assign n9639 = ~n9628 & n9638;
  assign n9640 = n9639 ^ n6301;
  assign n9641 = n9640 ^ n9624;
  assign n9642 = ~n9625 & n9641;
  assign n9643 = n9642 ^ n6295;
  assign n9644 = n9643 ^ n9621;
  assign n9645 = n9622 & ~n9644;
  assign n9646 = n9645 ^ n6288;
  assign n9647 = n9646 ^ n9619;
  assign n9648 = ~n9620 & ~n9647;
  assign n9649 = n9648 ^ n6282;
  assign n9650 = n9649 ^ n9616;
  assign n9651 = ~n9617 & ~n9650;
  assign n9652 = n9651 ^ n6275;
  assign n9653 = n9652 ^ n9614;
  assign n9654 = ~n9615 & ~n9653;
  assign n9655 = n9654 ^ n6269;
  assign n9656 = n9655 ^ n9611;
  assign n9657 = ~n9612 & n9656;
  assign n9658 = n9657 ^ n6261;
  assign n9659 = n9658 ^ n9609;
  assign n9660 = n9610 & ~n9659;
  assign n9661 = n9660 ^ n6756;
  assign n9662 = n9661 ^ n9606;
  assign n9663 = ~n9607 & ~n9662;
  assign n9664 = n9663 ^ n6885;
  assign n9665 = n9664 ^ n9604;
  assign n9666 = ~n9605 & ~n9665;
  assign n9667 = n9666 ^ n6958;
  assign n9668 = n9667 ^ n9602;
  assign n9669 = n9603 & ~n9668;
  assign n9670 = n9669 ^ n6973;
  assign n9671 = n9670 ^ n9600;
  assign n9672 = n9601 & ~n9671;
  assign n9673 = n9672 ^ n6991;
  assign n9674 = n9673 ^ n9598;
  assign n9675 = ~n9599 & n9674;
  assign n9676 = n9675 ^ n7008;
  assign n9677 = n9676 ^ n9595;
  assign n9678 = ~n9596 & ~n9677;
  assign n9679 = n9678 ^ n7021;
  assign n9680 = n9679 ^ n9593;
  assign n9681 = n9594 & n9680;
  assign n9682 = n9681 ^ n7035;
  assign n9534 = n8188 ^ n7939;
  assign n9535 = n9139 & ~n9534;
  assign n9536 = n9535 ^ n7939;
  assign n9530 = n9529 ^ n9407;
  assign n9531 = ~n9408 & ~n9530;
  assign n9532 = n9531 ^ n9404;
  assign n9402 = n9093 ^ n9059;
  assign n9533 = n9532 ^ n9402;
  assign n9592 = n9536 ^ n9533;
  assign n9683 = n9682 ^ n9592;
  assign n9684 = n9592 ^ n7052;
  assign n9685 = n9683 & ~n9684;
  assign n9686 = n9685 ^ n7052;
  assign n9541 = n7932 ^ n7915;
  assign n9542 = ~n9167 & n9541;
  assign n9543 = n9542 ^ n7932;
  assign n9400 = n9096 ^ x332;
  assign n9401 = n9400 ^ n9056;
  assign n9589 = n9543 ^ n9401;
  assign n9537 = n9536 ^ n9402;
  assign n9538 = ~n9533 & ~n9537;
  assign n9539 = n9538 ^ n9536;
  assign n9590 = n9589 ^ n9539;
  assign n9591 = n9590 ^ n7244;
  assign n9746 = n9686 ^ n9591;
  assign n9709 = n9683 ^ n7052;
  assign n9710 = n9676 ^ n9596;
  assign n9711 = n9673 ^ n9599;
  assign n9712 = n9667 ^ n9603;
  assign n9713 = n9655 ^ n9612;
  assign n9714 = n9649 ^ n9617;
  assign n9715 = n9640 ^ n9625;
  assign n9716 = n9634 ^ n9631;
  assign n9231 = n9230 ^ n9197;
  assign n9232 = n9194 ^ n5990;
  assign n9233 = n9232 ^ n9185;
  assign n9234 = n9187 ^ n6343;
  assign n9235 = n9191 ^ n9189;
  assign n9236 = n9234 & n9235;
  assign n9237 = n9233 & n9236;
  assign n9238 = n9231 & ~n9237;
  assign n9275 = n9274 ^ n9241;
  assign n9276 = n9238 & n9275;
  assign n9290 = n9289 ^ n9279;
  assign n9317 = ~n9276 & ~n9290;
  assign n9331 = n9330 ^ n9320;
  assign n9717 = n9317 & ~n9331;
  assign n9718 = ~n9716 & ~n9717;
  assign n9719 = n9637 ^ n9628;
  assign n9720 = n9718 & n9719;
  assign n9721 = ~n9715 & ~n9720;
  assign n9722 = n9643 ^ n6288;
  assign n9723 = n9722 ^ n9621;
  assign n9724 = n9721 & n9723;
  assign n9725 = n9646 ^ n9620;
  assign n9726 = ~n9724 & n9725;
  assign n9727 = ~n9714 & n9726;
  assign n9728 = n9652 ^ n6269;
  assign n9729 = n9728 ^ n9614;
  assign n9730 = n9727 & n9729;
  assign n9731 = ~n9713 & n9730;
  assign n9732 = n9658 ^ n9610;
  assign n9733 = ~n9731 & ~n9732;
  assign n9734 = n9661 ^ n9607;
  assign n9735 = n9733 & n9734;
  assign n9736 = n9664 ^ n9605;
  assign n9737 = ~n9735 & n9736;
  assign n9738 = ~n9712 & ~n9737;
  assign n9739 = n9670 ^ n9601;
  assign n9740 = n9738 & ~n9739;
  assign n9741 = n9711 & n9740;
  assign n9742 = n9710 & n9741;
  assign n9743 = n9679 ^ n9594;
  assign n9744 = n9742 & n9743;
  assign n9745 = ~n9709 & ~n9744;
  assign n9780 = n9746 ^ n9745;
  assign n9781 = n9780 ^ x359;
  assign n9782 = n9744 ^ n9709;
  assign n9783 = n9782 ^ x360;
  assign n9784 = n9743 ^ n9742;
  assign n9785 = n9784 ^ x361;
  assign n9786 = n9741 ^ n9710;
  assign n9787 = n9786 ^ x362;
  assign n9788 = n9740 ^ n9711;
  assign n9789 = n9788 ^ x363;
  assign n9790 = n9739 ^ n9738;
  assign n9791 = n9790 ^ x364;
  assign n9792 = n9737 ^ n9712;
  assign n9793 = n9792 ^ x365;
  assign n9794 = n9736 ^ n9735;
  assign n9795 = n9794 ^ x366;
  assign n9797 = n9732 ^ n9731;
  assign n9798 = n9797 ^ x368;
  assign n9799 = n9730 ^ n9713;
  assign n9800 = n9799 ^ x369;
  assign n9801 = n9729 ^ n9727;
  assign n9802 = n9801 ^ x370;
  assign n9803 = n9726 ^ n9714;
  assign n9804 = n9803 ^ x371;
  assign n9805 = n9725 ^ n9724;
  assign n9806 = n9805 ^ x372;
  assign n9807 = n9723 ^ n9721;
  assign n9808 = n9807 ^ x373;
  assign n9809 = n9720 ^ n9715;
  assign n9810 = n9809 ^ x374;
  assign n9811 = n9719 ^ n9718;
  assign n9812 = n9811 ^ x375;
  assign n9813 = n9717 ^ n9716;
  assign n9814 = n9813 ^ x376;
  assign n9332 = n9331 ^ n9317;
  assign n9333 = n9332 ^ x377;
  assign n9291 = n9290 ^ n9276;
  assign n9292 = n9291 ^ x378;
  assign n9293 = n9275 ^ n9238;
  assign n9294 = n9293 ^ x379;
  assign n9295 = n9237 ^ n9231;
  assign n9296 = n9295 ^ x380;
  assign n9297 = n9236 ^ n9233;
  assign n9298 = n9297 ^ x381;
  assign n9299 = x383 & ~n9234;
  assign n9300 = n9299 ^ x382;
  assign n9301 = n9235 ^ n9234;
  assign n9302 = n9301 ^ n9299;
  assign n9303 = n9300 & ~n9302;
  assign n9304 = n9303 ^ x382;
  assign n9305 = n9304 ^ n9297;
  assign n9306 = n9298 & ~n9305;
  assign n9307 = n9306 ^ x381;
  assign n9308 = n9307 ^ n9295;
  assign n9309 = n9296 & ~n9308;
  assign n9310 = n9309 ^ x380;
  assign n9311 = n9310 ^ n9293;
  assign n9312 = ~n9294 & n9311;
  assign n9313 = n9312 ^ x379;
  assign n9314 = n9313 ^ n9291;
  assign n9315 = n9292 & ~n9314;
  assign n9316 = n9315 ^ x378;
  assign n9815 = n9332 ^ n9316;
  assign n9816 = ~n9333 & n9815;
  assign n9817 = n9816 ^ x377;
  assign n9818 = n9817 ^ n9813;
  assign n9819 = ~n9814 & n9818;
  assign n9820 = n9819 ^ x376;
  assign n9821 = n9820 ^ n9811;
  assign n9822 = ~n9812 & n9821;
  assign n9823 = n9822 ^ x375;
  assign n9824 = n9823 ^ n9809;
  assign n9825 = n9810 & ~n9824;
  assign n9826 = n9825 ^ x374;
  assign n9827 = n9826 ^ n9807;
  assign n9828 = n9808 & ~n9827;
  assign n9829 = n9828 ^ x373;
  assign n9830 = n9829 ^ n9805;
  assign n9831 = n9806 & ~n9830;
  assign n9832 = n9831 ^ x372;
  assign n9833 = n9832 ^ n9803;
  assign n9834 = n9804 & ~n9833;
  assign n9835 = n9834 ^ x371;
  assign n9836 = n9835 ^ n9801;
  assign n9837 = ~n9802 & n9836;
  assign n9838 = n9837 ^ x370;
  assign n9839 = n9838 ^ n9799;
  assign n9840 = n9800 & ~n9839;
  assign n9841 = n9840 ^ x369;
  assign n9842 = n9841 ^ n9797;
  assign n9843 = n9798 & ~n9842;
  assign n9844 = n9843 ^ x368;
  assign n9796 = n9734 ^ n9733;
  assign n9845 = n9844 ^ n9796;
  assign n9846 = n9796 ^ x367;
  assign n9847 = ~n9845 & n9846;
  assign n9848 = n9847 ^ x367;
  assign n9849 = n9848 ^ n9794;
  assign n9850 = n9795 & ~n9849;
  assign n9851 = n9850 ^ x366;
  assign n9852 = n9851 ^ n9792;
  assign n9853 = n9793 & ~n9852;
  assign n9854 = n9853 ^ x365;
  assign n9855 = n9854 ^ n9790;
  assign n9856 = ~n9791 & n9855;
  assign n9857 = n9856 ^ x364;
  assign n9858 = n9857 ^ n9788;
  assign n9859 = n9789 & ~n9858;
  assign n9860 = n9859 ^ x363;
  assign n9861 = n9860 ^ n9786;
  assign n9862 = n9787 & ~n9861;
  assign n9863 = n9862 ^ x362;
  assign n9864 = n9863 ^ n9784;
  assign n9865 = n9785 & ~n9864;
  assign n9866 = n9865 ^ x361;
  assign n9867 = n9866 ^ n9782;
  assign n9868 = ~n9783 & n9867;
  assign n9869 = n9868 ^ x360;
  assign n9870 = n9869 ^ n9780;
  assign n9871 = ~n9781 & n9870;
  assign n9872 = n9871 ^ x359;
  assign n9687 = n9686 ^ n9590;
  assign n9688 = ~n9591 & ~n9687;
  assign n9689 = n9688 ^ n7244;
  assign n9540 = n9539 ^ n9401;
  assign n9544 = n9543 ^ n9539;
  assign n9545 = ~n9540 & ~n9544;
  assign n9546 = n9545 ^ n9401;
  assign n9396 = n7810 ^ n7226;
  assign n9397 = ~n9212 & n9396;
  assign n9398 = n9397 ^ n7226;
  assign n9586 = n9546 ^ n9398;
  assign n9395 = n9099 ^ n9055;
  assign n9587 = n9586 ^ n9395;
  assign n9588 = n9587 ^ n6687;
  assign n9748 = n9689 ^ n9588;
  assign n9747 = ~n9745 & n9746;
  assign n9778 = n9748 ^ n9747;
  assign n9779 = n9778 ^ x358;
  assign n10256 = n9872 ^ n9779;
  assign n11098 = n9150 ^ n8594;
  assign n11099 = n10256 & ~n11098;
  assign n11100 = n11099 ^ n8594;
  assign n10261 = n9869 ^ n9781;
  assign n9374 = n9117 ^ n9043;
  assign n11086 = n9374 ^ n9246;
  assign n11087 = ~n10261 & ~n11086;
  assign n11088 = n11087 ^ n9246;
  assign n10309 = n8797 ^ n7953;
  assign n10310 = ~n9409 & ~n10309;
  assign n10311 = n10310 ^ n7953;
  assign n10216 = n9829 ^ x372;
  assign n10217 = n10216 ^ n9805;
  assign n10312 = n10311 ^ n10217;
  assign n10313 = n8803 ^ n7959;
  assign n10314 = n9411 & n10313;
  assign n10315 = n10314 ^ n7959;
  assign n10224 = n9826 ^ n9808;
  assign n10316 = n10315 ^ n10224;
  assign n10153 = n9823 ^ n9810;
  assign n10150 = n8808 ^ n7964;
  assign n10151 = n9416 & ~n10150;
  assign n10152 = n10151 ^ n7964;
  assign n10154 = n10153 ^ n10152;
  assign n10040 = n9820 ^ x375;
  assign n10041 = n10040 ^ n9811;
  assign n10036 = n8814 ^ n7970;
  assign n10037 = n9422 & n10036;
  assign n10038 = n10037 ^ n7970;
  assign n10146 = n10041 ^ n10038;
  assign n9961 = n8819 ^ n7975;
  assign n9962 = n9430 & ~n9961;
  assign n9963 = n9962 ^ n7975;
  assign n9959 = n9817 ^ x376;
  assign n9960 = n9959 ^ n9813;
  assign n9964 = n9963 ^ n9960;
  assign n9334 = n9333 ^ n9316;
  assign n8785 = n8784 ^ n7978;
  assign n8786 = ~n8782 & n8785;
  assign n8787 = n8786 ^ n7978;
  assign n9335 = n9334 ^ n8787;
  assign n9340 = n9313 ^ x378;
  assign n9341 = n9340 ^ n9291;
  assign n9337 = n8828 ^ n7986;
  assign n9338 = ~n9336 & ~n9337;
  assign n9339 = n9338 ^ n7986;
  assign n9342 = n9341 ^ n9339;
  assign n9347 = n9310 ^ n9294;
  assign n9344 = n8830 ^ n7989;
  assign n9345 = ~n9343 & ~n9344;
  assign n9346 = n9345 ^ n7989;
  assign n9348 = n9347 ^ n9346;
  assign n9353 = n8835 ^ n7994;
  assign n9354 = n9352 & n9353;
  assign n9355 = n9354 ^ n7994;
  assign n9349 = n9307 ^ x380;
  assign n9350 = n9349 ^ n9295;
  assign n9356 = n9355 ^ n9350;
  assign n9360 = n8841 ^ n8002;
  assign n9361 = n9359 & n9360;
  assign n9362 = n9361 ^ n8002;
  assign n9357 = n9304 ^ n9298;
  assign n9363 = n9362 ^ n9357;
  assign n9936 = n9301 ^ n9300;
  assign n9367 = n8856 ^ n7375;
  assign n9368 = ~n9366 & n9367;
  assign n9369 = n9368 ^ n7375;
  assign n9364 = n9234 ^ x383;
  assign n9370 = n9369 ^ n9364;
  assign n9893 = n8776 ^ n7899;
  assign n9894 = n9461 & ~n9893;
  assign n9895 = n9894 ^ n7899;
  assign n9560 = n8100 ^ n7263;
  assign n9561 = ~n8583 & ~n9560;
  assign n9562 = n9561 ^ n7263;
  assign n9380 = n8070 ^ n7212;
  assign n9381 = ~n8591 & n9380;
  assign n9382 = n9381 ^ n7212;
  assign n9378 = n9108 ^ x328;
  assign n9379 = n9378 ^ n9048;
  assign n9383 = n9382 ^ n9379;
  assign n9385 = n7883 ^ n7215;
  assign n9386 = ~n8594 & ~n9385;
  assign n9387 = n9386 ^ n7215;
  assign n9384 = n9105 ^ n9051;
  assign n9388 = n9387 ^ n9384;
  assign n9391 = n7847 ^ n7220;
  assign n9392 = ~n9246 & ~n9391;
  assign n9393 = n9392 ^ n7220;
  assign n9389 = n9102 ^ x330;
  assign n9390 = n9389 ^ n9052;
  assign n9394 = n9393 ^ n9390;
  assign n9399 = n9398 ^ n9395;
  assign n9547 = n9546 ^ n9395;
  assign n9548 = ~n9399 & ~n9547;
  assign n9549 = n9548 ^ n9398;
  assign n9550 = n9549 ^ n9390;
  assign n9551 = n9394 & ~n9550;
  assign n9552 = n9551 ^ n9393;
  assign n9553 = n9552 ^ n9384;
  assign n9554 = n9388 & n9553;
  assign n9555 = n9554 ^ n9387;
  assign n9556 = n9555 ^ n9379;
  assign n9557 = ~n9383 & ~n9556;
  assign n9558 = n9557 ^ n9382;
  assign n9377 = n9111 ^ n9047;
  assign n9559 = n9558 ^ n9377;
  assign n9576 = n9562 ^ n9559;
  assign n9755 = n9576 ^ n6667;
  assign n9577 = n9555 ^ n9382;
  assign n9578 = n9577 ^ n9379;
  assign n9579 = n9578 ^ n6672;
  assign n9580 = n9552 ^ n9387;
  assign n9581 = n9580 ^ n9384;
  assign n9582 = n9581 ^ n6677;
  assign n9583 = n9549 ^ n9393;
  assign n9584 = n9583 ^ n9390;
  assign n9585 = n9584 ^ n6682;
  assign n9690 = n9689 ^ n9587;
  assign n9691 = ~n9588 & ~n9690;
  assign n9692 = n9691 ^ n6687;
  assign n9693 = n9692 ^ n9584;
  assign n9694 = ~n9585 & n9693;
  assign n9695 = n9694 ^ n6682;
  assign n9696 = n9695 ^ n9581;
  assign n9697 = n9582 & n9696;
  assign n9698 = n9697 ^ n6677;
  assign n9699 = n9698 ^ n9578;
  assign n9700 = n9579 & ~n9699;
  assign n9701 = n9700 ^ n6672;
  assign n9756 = n9701 ^ n9576;
  assign n9757 = ~n9755 & ~n9756;
  assign n9758 = n9757 ^ n6667;
  assign n9759 = n9758 ^ n6356;
  assign n9569 = n8039 ^ n7267;
  assign n9570 = n8578 & n9569;
  assign n9571 = n9570 ^ n7267;
  assign n9566 = n9114 ^ x326;
  assign n9567 = n9566 ^ n9044;
  assign n9563 = n9562 ^ n9377;
  assign n9564 = n9559 & n9563;
  assign n9565 = n9564 ^ n9562;
  assign n9568 = n9567 ^ n9565;
  assign n9754 = n9571 ^ n9568;
  assign n9760 = n9759 ^ n9754;
  assign n9702 = n9701 ^ n6667;
  assign n9703 = n9702 ^ n9576;
  assign n9704 = n9698 ^ n6672;
  assign n9705 = n9704 ^ n9578;
  assign n9706 = n9695 ^ n6677;
  assign n9707 = n9706 ^ n9581;
  assign n9708 = n9692 ^ n9585;
  assign n9749 = ~n9747 & n9748;
  assign n9750 = n9708 & ~n9749;
  assign n9751 = n9707 & ~n9750;
  assign n9752 = ~n9705 & n9751;
  assign n9753 = ~n9703 & ~n9752;
  assign n9768 = n9760 ^ n9753;
  assign n9769 = n9768 ^ x353;
  assign n9770 = n9752 ^ n9703;
  assign n9771 = n9770 ^ x354;
  assign n9772 = n9751 ^ n9705;
  assign n9773 = n9772 ^ x355;
  assign n9774 = n9750 ^ n9707;
  assign n9775 = n9774 ^ x356;
  assign n9776 = n9749 ^ n9708;
  assign n9777 = n9776 ^ x357;
  assign n9873 = n9872 ^ n9778;
  assign n9874 = n9779 & ~n9873;
  assign n9875 = n9874 ^ x358;
  assign n9876 = n9875 ^ n9776;
  assign n9877 = ~n9777 & n9876;
  assign n9878 = n9877 ^ x357;
  assign n9879 = n9878 ^ n9774;
  assign n9880 = n9775 & ~n9879;
  assign n9881 = n9880 ^ x356;
  assign n9882 = n9881 ^ n9772;
  assign n9883 = n9773 & ~n9882;
  assign n9884 = n9883 ^ x355;
  assign n9885 = n9884 ^ n9770;
  assign n9886 = n9771 & ~n9885;
  assign n9887 = n9886 ^ x354;
  assign n9888 = n9887 ^ n9768;
  assign n9889 = n9769 & ~n9888;
  assign n9890 = n9889 ^ x353;
  assign n9891 = n9890 ^ x352;
  assign n9763 = n9754 ^ n6356;
  assign n9764 = n9758 ^ n9754;
  assign n9765 = n9763 & ~n9764;
  assign n9766 = n9765 ^ n6356;
  assign n9761 = ~n9753 & n9760;
  assign n9572 = n9571 ^ n9567;
  assign n9573 = n9568 & n9572;
  assign n9574 = n9573 ^ n9571;
  assign n9371 = n8038 ^ n7306;
  assign n9372 = n8572 & ~n9371;
  assign n9373 = n9372 ^ n7306;
  assign n9375 = n9374 ^ n9373;
  assign n9376 = n9375 ^ n6351;
  assign n9575 = n9574 ^ n9376;
  assign n9762 = n9761 ^ n9575;
  assign n9767 = n9766 ^ n9762;
  assign n9892 = n9891 ^ n9767;
  assign n9896 = n9895 ^ n9892;
  assign n9899 = n8709 ^ n7906;
  assign n9900 = ~n9467 & n9899;
  assign n9901 = n9900 ^ n7906;
  assign n9897 = n9887 ^ x353;
  assign n9898 = n9897 ^ n9768;
  assign n9902 = n9901 ^ n9898;
  assign n9908 = n8621 ^ n8028;
  assign n9909 = n9327 & ~n9908;
  assign n9910 = n9909 ^ n8028;
  assign n9906 = n9881 ^ x355;
  assign n9907 = n9906 ^ n9772;
  assign n9911 = n9910 ^ n9907;
  assign n9912 = n8033 ^ n7897;
  assign n9913 = ~n9286 & ~n9912;
  assign n9914 = n9913 ^ n8033;
  assign n9915 = n9878 ^ x356;
  assign n9916 = n9915 ^ n9774;
  assign n9917 = n9914 & n9916;
  assign n9918 = n9917 ^ n9907;
  assign n9919 = ~n9911 & n9918;
  assign n9920 = n9919 ^ n9917;
  assign n9903 = n8675 ^ n8022;
  assign n9904 = n9473 & ~n9903;
  assign n9905 = n9904 ^ n8022;
  assign n9921 = n9920 ^ n9905;
  assign n9922 = n9884 ^ x354;
  assign n9923 = n9922 ^ n9770;
  assign n9924 = n9923 ^ n9920;
  assign n9925 = ~n9921 & ~n9924;
  assign n9926 = n9925 ^ n9905;
  assign n9927 = n9926 ^ n9898;
  assign n9928 = ~n9902 & n9927;
  assign n9929 = n9928 ^ n9901;
  assign n9930 = n9929 ^ n9892;
  assign n9931 = ~n9896 & n9930;
  assign n9932 = n9931 ^ n9895;
  assign n9933 = n9932 ^ n9364;
  assign n9934 = ~n9370 & ~n9933;
  assign n9935 = n9934 ^ n9369;
  assign n9937 = n9936 ^ n9935;
  assign n9938 = n8847 ^ n8005;
  assign n9939 = n9452 & ~n9938;
  assign n9940 = n9939 ^ n8005;
  assign n9941 = n9940 ^ n9936;
  assign n9942 = ~n9937 & ~n9941;
  assign n9943 = n9942 ^ n9940;
  assign n9944 = n9943 ^ n9357;
  assign n9945 = n9363 & n9944;
  assign n9946 = n9945 ^ n9362;
  assign n9947 = n9946 ^ n9350;
  assign n9948 = n9356 & ~n9947;
  assign n9949 = n9948 ^ n9355;
  assign n9950 = n9949 ^ n9347;
  assign n9951 = ~n9348 & n9950;
  assign n9952 = n9951 ^ n9346;
  assign n9953 = n9952 ^ n9341;
  assign n9954 = ~n9342 & ~n9953;
  assign n9955 = n9954 ^ n9339;
  assign n9956 = n9955 ^ n9334;
  assign n9957 = ~n9335 & ~n9956;
  assign n9958 = n9957 ^ n8787;
  assign n10033 = n9960 ^ n9958;
  assign n10034 = ~n9964 & n10033;
  assign n10035 = n10034 ^ n9963;
  assign n10147 = n10041 ^ n10035;
  assign n10148 = ~n10146 & n10147;
  assign n10149 = n10148 ^ n10038;
  assign n10317 = n10153 ^ n10149;
  assign n10318 = n10154 & ~n10317;
  assign n10319 = n10318 ^ n10152;
  assign n10320 = n10319 ^ n10224;
  assign n10321 = n10316 & ~n10320;
  assign n10322 = n10321 ^ n10315;
  assign n10323 = n10322 ^ n10217;
  assign n10324 = ~n10312 & ~n10323;
  assign n10325 = n10324 ^ n10311;
  assign n10305 = n8792 ^ n7948;
  assign n10306 = ~n9404 & ~n10305;
  assign n10307 = n10306 ^ n7948;
  assign n10413 = n10325 ^ n10307;
  assign n10209 = n9832 ^ n9804;
  assign n10414 = n10413 ^ n10209;
  assign n10415 = n10414 ^ n7651;
  assign n10416 = n10322 ^ n10312;
  assign n10417 = n10416 ^ n7638;
  assign n10418 = n10319 ^ n10315;
  assign n10419 = n10418 ^ n10224;
  assign n10420 = n10419 ^ n7618;
  assign n10155 = n10154 ^ n10149;
  assign n10156 = n10155 ^ n7570;
  assign n10039 = n10038 ^ n10035;
  assign n10042 = n10041 ^ n10039;
  assign n10043 = n10042 ^ n7489;
  assign n9965 = n9964 ^ n9958;
  assign n9966 = n9965 ^ n7383;
  assign n9967 = n9955 ^ n8787;
  assign n9968 = n9967 ^ n9334;
  assign n9969 = n9968 ^ n7389;
  assign n9970 = n9952 ^ n9342;
  assign n9971 = n9970 ^ n7391;
  assign n9972 = n9949 ^ n9346;
  assign n9973 = n9972 ^ n9347;
  assign n9974 = n9973 ^ n7400;
  assign n9975 = n9946 ^ n9356;
  assign n9976 = n9975 ^ n7405;
  assign n9977 = n9943 ^ n9362;
  assign n9978 = n9977 ^ n9357;
  assign n9979 = n9978 ^ n7376;
  assign n9980 = n9940 ^ n9937;
  assign n9981 = n9980 ^ n7415;
  assign n9982 = n9932 ^ n9369;
  assign n9983 = n9982 ^ n9364;
  assign n9984 = n9983 ^ n7421;
  assign n9985 = n9929 ^ n9895;
  assign n9986 = n9985 ^ n9892;
  assign n9987 = n9986 ^ n7423;
  assign n9988 = n9926 ^ n9902;
  assign n9989 = n9988 ^ n7432;
  assign n9990 = n9923 ^ n9921;
  assign n9991 = n9990 ^ n7434;
  assign n9992 = n9916 ^ n9914;
  assign n9993 = ~n7370 & n9992;
  assign n9994 = n9993 ^ n7443;
  assign n9995 = n9917 ^ n9910;
  assign n9996 = n9995 ^ n9907;
  assign n9997 = n9996 ^ n9993;
  assign n9998 = ~n9994 & ~n9997;
  assign n9999 = n9998 ^ n7443;
  assign n10000 = n9999 ^ n9990;
  assign n10001 = n9991 & ~n10000;
  assign n10002 = n10001 ^ n7434;
  assign n10003 = n10002 ^ n9988;
  assign n10004 = n9989 & n10003;
  assign n10005 = n10004 ^ n7432;
  assign n10006 = n10005 ^ n9986;
  assign n10007 = n9987 & ~n10006;
  assign n10008 = n10007 ^ n7423;
  assign n10009 = n10008 ^ n9983;
  assign n10010 = n9984 & ~n10009;
  assign n10011 = n10010 ^ n7421;
  assign n10012 = n10011 ^ n9980;
  assign n10013 = n9981 & n10012;
  assign n10014 = n10013 ^ n7415;
  assign n10015 = n10014 ^ n9978;
  assign n10016 = ~n9979 & ~n10015;
  assign n10017 = n10016 ^ n7376;
  assign n10018 = n10017 ^ n9975;
  assign n10019 = n9976 & ~n10018;
  assign n10020 = n10019 ^ n7405;
  assign n10021 = n10020 ^ n9973;
  assign n10022 = n9974 & n10021;
  assign n10023 = n10022 ^ n7400;
  assign n10024 = n10023 ^ n9970;
  assign n10025 = ~n9971 & ~n10024;
  assign n10026 = n10025 ^ n7391;
  assign n10027 = n10026 ^ n9968;
  assign n10028 = n9969 & ~n10027;
  assign n10029 = n10028 ^ n7389;
  assign n10030 = n10029 ^ n9965;
  assign n10031 = n9966 & n10030;
  assign n10032 = n10031 ^ n7383;
  assign n10143 = n10042 ^ n10032;
  assign n10144 = n10043 & ~n10143;
  assign n10145 = n10144 ^ n7489;
  assign n10421 = n10155 ^ n10145;
  assign n10422 = n10156 & n10421;
  assign n10423 = n10422 ^ n7570;
  assign n10424 = n10423 ^ n10419;
  assign n10425 = n10420 & ~n10424;
  assign n10426 = n10425 ^ n7618;
  assign n10427 = n10426 ^ n10416;
  assign n10428 = ~n10417 & n10427;
  assign n10429 = n10428 ^ n7638;
  assign n10430 = n10429 ^ n10414;
  assign n10431 = ~n10415 & n10430;
  assign n10432 = n10431 ^ n7651;
  assign n10308 = n10307 ^ n10209;
  assign n10326 = n10325 ^ n10209;
  assign n10327 = n10308 & n10326;
  assign n10328 = n10327 ^ n10307;
  assign n10301 = n8904 ^ n7937;
  assign n10302 = ~n9402 & n10301;
  assign n10303 = n10302 ^ n7937;
  assign n10410 = n10328 ^ n10303;
  assign n10201 = n9835 ^ x370;
  assign n10202 = n10201 ^ n9801;
  assign n10411 = n10410 ^ n10202;
  assign n10412 = n10411 ^ n7671;
  assign n10486 = n10432 ^ n10412;
  assign n10479 = n10429 ^ n10415;
  assign n10480 = n10423 ^ n10420;
  assign n10044 = n10043 ^ n10032;
  assign n10045 = n10029 ^ n9966;
  assign n10046 = n10026 ^ n9969;
  assign n10047 = n10023 ^ n9971;
  assign n10048 = n10014 ^ n9979;
  assign n10049 = n10002 ^ n7432;
  assign n10050 = n10049 ^ n9988;
  assign n10051 = n9999 ^ n7434;
  assign n10052 = n10051 ^ n9990;
  assign n10053 = n9992 ^ n7370;
  assign n10054 = n9996 ^ n9994;
  assign n10055 = ~n10053 & ~n10054;
  assign n10056 = ~n10052 & n10055;
  assign n10057 = n10050 & ~n10056;
  assign n10058 = n10005 ^ n7423;
  assign n10059 = n10058 ^ n9986;
  assign n10060 = n10057 & ~n10059;
  assign n10061 = n10008 ^ n7421;
  assign n10062 = n10061 ^ n9983;
  assign n10063 = ~n10060 & n10062;
  assign n10064 = n10011 ^ n7415;
  assign n10065 = n10064 ^ n9980;
  assign n10066 = n10063 & n10065;
  assign n10067 = ~n10048 & ~n10066;
  assign n10068 = n10017 ^ n9976;
  assign n10069 = n10067 & ~n10068;
  assign n10070 = n10020 ^ n7400;
  assign n10071 = n10070 ^ n9973;
  assign n10072 = ~n10069 & n10071;
  assign n10073 = n10047 & n10072;
  assign n10074 = ~n10046 & ~n10073;
  assign n10075 = ~n10045 & n10074;
  assign n10142 = n10044 & n10075;
  assign n10157 = n10156 ^ n10145;
  assign n10481 = n10142 & n10157;
  assign n10482 = n10480 & ~n10481;
  assign n10483 = n10426 ^ n10417;
  assign n10484 = n10482 & ~n10483;
  assign n10485 = n10479 & ~n10484;
  assign n10537 = n10486 ^ n10485;
  assign n10538 = n10537 ^ x397;
  assign n10539 = n10484 ^ n10479;
  assign n10540 = n10539 ^ x398;
  assign n10542 = n10481 ^ n10480;
  assign n10543 = n10542 ^ x400;
  assign n10158 = n10157 ^ n10142;
  assign n10159 = n10158 ^ x401;
  assign n10076 = n10075 ^ n10044;
  assign n10077 = n10076 ^ x402;
  assign n10078 = n10074 ^ n10045;
  assign n10079 = n10078 ^ x403;
  assign n10080 = n10073 ^ n10046;
  assign n10081 = n10080 ^ x404;
  assign n10082 = n10072 ^ n10047;
  assign n10083 = n10082 ^ x405;
  assign n10084 = n10071 ^ n10069;
  assign n10085 = n10084 ^ x406;
  assign n10086 = n10068 ^ n10067;
  assign n10087 = n10086 ^ x407;
  assign n10088 = n10066 ^ n10048;
  assign n10089 = n10088 ^ x408;
  assign n10090 = n10065 ^ n10063;
  assign n10091 = n10090 ^ x409;
  assign n10092 = n10062 ^ n10060;
  assign n10093 = n10092 ^ x410;
  assign n10094 = n10059 ^ n10057;
  assign n10095 = n10094 ^ x411;
  assign n10096 = n10056 ^ n10050;
  assign n10097 = n10096 ^ x412;
  assign n10098 = n10055 ^ n10052;
  assign n10099 = n10098 ^ x413;
  assign n10100 = x415 & n10053;
  assign n10101 = n10100 ^ x414;
  assign n10102 = n10054 ^ n10053;
  assign n10103 = n10102 ^ n10100;
  assign n10104 = n10101 & ~n10103;
  assign n10105 = n10104 ^ x414;
  assign n10106 = n10105 ^ n10098;
  assign n10107 = ~n10099 & n10106;
  assign n10108 = n10107 ^ x413;
  assign n10109 = n10108 ^ n10096;
  assign n10110 = n10097 & ~n10109;
  assign n10111 = n10110 ^ x412;
  assign n10112 = n10111 ^ n10094;
  assign n10113 = n10095 & ~n10112;
  assign n10114 = n10113 ^ x411;
  assign n10115 = n10114 ^ n10092;
  assign n10116 = ~n10093 & n10115;
  assign n10117 = n10116 ^ x410;
  assign n10118 = n10117 ^ n10090;
  assign n10119 = n10091 & ~n10118;
  assign n10120 = n10119 ^ x409;
  assign n10121 = n10120 ^ n10088;
  assign n10122 = ~n10089 & n10121;
  assign n10123 = n10122 ^ x408;
  assign n10124 = n10123 ^ n10086;
  assign n10125 = n10087 & ~n10124;
  assign n10126 = n10125 ^ x407;
  assign n10127 = n10126 ^ n10084;
  assign n10128 = ~n10085 & n10127;
  assign n10129 = n10128 ^ x406;
  assign n10130 = n10129 ^ n10082;
  assign n10131 = n10083 & ~n10130;
  assign n10132 = n10131 ^ x405;
  assign n10133 = n10132 ^ n10080;
  assign n10134 = ~n10081 & n10133;
  assign n10135 = n10134 ^ x404;
  assign n10136 = n10135 ^ n10078;
  assign n10137 = n10079 & ~n10136;
  assign n10138 = n10137 ^ x403;
  assign n10139 = n10138 ^ n10076;
  assign n10140 = ~n10077 & n10139;
  assign n10141 = n10140 ^ x402;
  assign n10544 = n10158 ^ n10141;
  assign n10545 = ~n10159 & n10544;
  assign n10546 = n10545 ^ x401;
  assign n10547 = n10546 ^ n10542;
  assign n10548 = ~n10543 & n10547;
  assign n10549 = n10548 ^ x400;
  assign n10541 = n10483 ^ n10482;
  assign n10550 = n10549 ^ n10541;
  assign n10551 = n10541 ^ x399;
  assign n10552 = n10550 & ~n10551;
  assign n10553 = n10552 ^ x399;
  assign n10554 = n10553 ^ n10539;
  assign n10555 = n10540 & ~n10554;
  assign n10556 = n10555 ^ x398;
  assign n10557 = n10556 ^ n10537;
  assign n10558 = ~n10538 & n10557;
  assign n10559 = n10558 ^ x397;
  assign n11084 = n10559 ^ x396;
  assign n10433 = n10432 ^ n10411;
  assign n10434 = n10412 & n10433;
  assign n10435 = n10434 ^ n7671;
  assign n10488 = n10435 ^ n7689;
  assign n10304 = n10303 ^ n10202;
  assign n10329 = n10328 ^ n10202;
  assign n10330 = ~n10304 & n10329;
  assign n10331 = n10330 ^ n10303;
  assign n10297 = n8985 ^ n7931;
  assign n10298 = ~n9401 & n10297;
  assign n10299 = n10298 ^ n7931;
  assign n10407 = n10331 ^ n10299;
  assign n10194 = n9838 ^ n9800;
  assign n10408 = n10407 ^ n10194;
  assign n10489 = n10488 ^ n10408;
  assign n10487 = ~n10485 & n10486;
  assign n10535 = n10489 ^ n10487;
  assign n11085 = n11084 ^ n10535;
  assign n11089 = n11088 ^ n11085;
  assign n10262 = n9866 ^ x360;
  assign n10263 = n10262 ^ n9782;
  assign n10994 = n9567 ^ n9212;
  assign n10995 = ~n10263 & ~n10994;
  assign n10996 = n10995 ^ n9212;
  assign n10993 = n10556 ^ n10538;
  assign n11090 = n10996 ^ n10993;
  assign n10276 = n9860 ^ x362;
  assign n10277 = n10276 ^ n9786;
  assign n10807 = n9379 ^ n9139;
  assign n10808 = n10277 & ~n10807;
  assign n10809 = n10808 ^ n9139;
  assign n10806 = n10550 ^ x399;
  assign n10810 = n10809 ^ n10806;
  assign n10692 = n10546 ^ x400;
  assign n10693 = n10692 ^ n10542;
  assign n10282 = n9857 ^ x363;
  assign n10283 = n10282 ^ n9788;
  assign n10689 = n9384 ^ n9037;
  assign n10690 = n10283 & ~n10689;
  assign n10691 = n10690 ^ n9037;
  assign n10694 = n10693 ^ n10691;
  assign n10161 = n9854 ^ x364;
  assign n10162 = n10161 ^ n9790;
  assign n10163 = n9390 ^ n8985;
  assign n10164 = ~n10162 & ~n10163;
  assign n10165 = n10164 ^ n8985;
  assign n10160 = n10159 ^ n10141;
  assign n10166 = n10165 ^ n10160;
  assign n10171 = n10138 ^ x402;
  assign n10172 = n10171 ^ n10076;
  assign n10167 = n9851 ^ n9793;
  assign n10168 = n9395 ^ n8904;
  assign n10169 = n10167 & ~n10168;
  assign n10170 = n10169 ^ n8904;
  assign n10173 = n10172 ^ n10170;
  assign n10178 = n10135 ^ n10079;
  assign n10174 = n9848 ^ n9795;
  assign n10175 = n9401 ^ n8792;
  assign n10176 = n10174 & n10175;
  assign n10177 = n10176 ^ n8792;
  assign n10179 = n10178 ^ n10177;
  assign n10184 = n10132 ^ x404;
  assign n10185 = n10184 ^ n10080;
  assign n10180 = n9845 ^ x367;
  assign n10181 = n9402 ^ n8797;
  assign n10182 = n10180 & ~n10181;
  assign n10183 = n10182 ^ n8797;
  assign n10186 = n10185 ^ n10183;
  assign n10192 = n10129 ^ n10083;
  assign n10187 = n9841 ^ x368;
  assign n10188 = n10187 ^ n9797;
  assign n10189 = n9404 ^ n8803;
  assign n10190 = n10188 & ~n10189;
  assign n10191 = n10190 ^ n8803;
  assign n10193 = n10192 ^ n10191;
  assign n10198 = n10126 ^ n10085;
  assign n10195 = n9409 ^ n8808;
  assign n10196 = n10194 & n10195;
  assign n10197 = n10196 ^ n8808;
  assign n10199 = n10198 ^ n10197;
  assign n10203 = n9411 ^ n8814;
  assign n10204 = ~n10202 & n10203;
  assign n10205 = n10204 ^ n8814;
  assign n10200 = n10123 ^ n10087;
  assign n10206 = n10205 ^ n10200;
  assign n10210 = n9416 ^ n8819;
  assign n10211 = n10209 & ~n10210;
  assign n10212 = n10211 ^ n8819;
  assign n10207 = n10120 ^ x408;
  assign n10208 = n10207 ^ n10088;
  assign n10213 = n10212 ^ n10208;
  assign n10218 = n9422 ^ n8784;
  assign n10219 = n10217 & n10218;
  assign n10220 = n10219 ^ n8784;
  assign n10214 = n10117 ^ x409;
  assign n10215 = n10214 ^ n10090;
  assign n10221 = n10220 ^ n10215;
  assign n10225 = n9430 ^ n8828;
  assign n10226 = n10224 & n10225;
  assign n10227 = n10226 ^ n8828;
  assign n10222 = n10114 ^ x410;
  assign n10223 = n10222 ^ n10092;
  assign n10228 = n10227 ^ n10223;
  assign n10232 = n10111 ^ n10095;
  assign n10229 = n8830 ^ n8782;
  assign n10230 = n10153 & n10229;
  assign n10231 = n10230 ^ n8830;
  assign n10233 = n10232 ^ n10231;
  assign n10237 = n10108 ^ x412;
  assign n10238 = n10237 ^ n10096;
  assign n10234 = n9336 ^ n8835;
  assign n10235 = ~n10041 & ~n10234;
  assign n10236 = n10235 ^ n8835;
  assign n10239 = n10238 ^ n10236;
  assign n10645 = n10105 ^ n10099;
  assign n10243 = n10102 ^ n10101;
  assign n10240 = n9352 ^ n8847;
  assign n10241 = ~n9334 & n10240;
  assign n10242 = n10241 ^ n8847;
  assign n10244 = n10243 ^ n10242;
  assign n10246 = n9359 ^ n8856;
  assign n10247 = n9341 & n10246;
  assign n10248 = n10247 ^ n8856;
  assign n10245 = n10053 ^ x415;
  assign n10249 = n10248 ^ n10245;
  assign n10599 = n9452 ^ n8776;
  assign n10600 = ~n9347 & n10599;
  assign n10601 = n10600 ^ n8776;
  assign n10271 = n9863 ^ n9785;
  assign n10268 = n8583 ^ n7883;
  assign n10269 = n9150 & ~n10268;
  assign n10270 = n10269 ^ n7883;
  assign n10272 = n10271 ^ n10270;
  assign n10273 = n8591 ^ n7847;
  assign n10274 = n9374 & n10273;
  assign n10275 = n10274 ^ n7847;
  assign n10278 = n10277 ^ n10275;
  assign n10279 = n8594 ^ n7810;
  assign n10280 = n9567 & ~n10279;
  assign n10281 = n10280 ^ n7810;
  assign n10284 = n10283 ^ n10281;
  assign n10285 = n9246 ^ n7915;
  assign n10286 = ~n9377 & ~n10285;
  assign n10287 = n10286 ^ n7915;
  assign n10288 = n10287 ^ n10162;
  assign n10289 = n9212 ^ n8188;
  assign n10290 = ~n9379 & n10289;
  assign n10291 = n10290 ^ n8188;
  assign n10292 = n10291 ^ n10167;
  assign n10293 = n9037 ^ n7925;
  assign n10294 = ~n9395 & n10293;
  assign n10295 = n10294 ^ n7925;
  assign n10296 = n10295 ^ n10188;
  assign n10300 = n10299 ^ n10194;
  assign n10332 = n10331 ^ n10194;
  assign n10333 = ~n10300 & ~n10332;
  assign n10334 = n10333 ^ n10299;
  assign n10335 = n10334 ^ n10188;
  assign n10336 = n10296 & n10335;
  assign n10337 = n10336 ^ n10295;
  assign n10338 = n10337 ^ n10180;
  assign n10339 = n9139 ^ n7920;
  assign n10340 = n9390 & n10339;
  assign n10341 = n10340 ^ n7920;
  assign n10342 = n10341 ^ n10180;
  assign n10343 = ~n10338 & n10342;
  assign n10344 = n10343 ^ n10341;
  assign n10345 = n10344 ^ n10174;
  assign n10346 = n9167 ^ n7918;
  assign n10347 = ~n9384 & n10346;
  assign n10348 = n10347 ^ n7918;
  assign n10349 = n10348 ^ n10174;
  assign n10350 = ~n10345 & ~n10349;
  assign n10351 = n10350 ^ n10348;
  assign n10352 = n10351 ^ n10167;
  assign n10353 = ~n10292 & n10352;
  assign n10354 = n10353 ^ n10291;
  assign n10355 = n10354 ^ n10162;
  assign n10356 = ~n10288 & ~n10355;
  assign n10357 = n10356 ^ n10287;
  assign n10358 = n10357 ^ n10283;
  assign n10359 = n10284 & ~n10358;
  assign n10360 = n10359 ^ n10281;
  assign n10361 = n10360 ^ n10277;
  assign n10362 = ~n10278 & ~n10361;
  assign n10363 = n10362 ^ n10275;
  assign n10364 = n10363 ^ n10271;
  assign n10365 = n10272 & n10364;
  assign n10366 = n10365 ^ n10270;
  assign n10264 = n8578 ^ n8070;
  assign n10265 = ~n9144 & n10264;
  assign n10266 = n10265 ^ n8070;
  assign n10384 = n10366 ^ n10266;
  assign n10385 = n10384 ^ n10263;
  assign n10386 = n10385 ^ n7212;
  assign n10387 = n10363 ^ n10270;
  assign n10388 = n10387 ^ n10271;
  assign n10389 = n10388 ^ n7215;
  assign n10390 = n10360 ^ n10275;
  assign n10391 = n10390 ^ n10277;
  assign n10392 = n10391 ^ n7220;
  assign n10393 = n10357 ^ n10281;
  assign n10394 = n10393 ^ n10283;
  assign n10395 = n10394 ^ n7226;
  assign n10396 = n10354 ^ n10288;
  assign n10397 = n10396 ^ n7932;
  assign n10398 = n10351 ^ n10291;
  assign n10399 = n10398 ^ n10167;
  assign n10400 = n10399 ^ n7939;
  assign n10401 = n10348 ^ n10345;
  assign n10402 = n10401 ^ n7865;
  assign n10403 = n10341 ^ n10338;
  assign n10404 = n10403 ^ n7834;
  assign n10405 = n10334 ^ n10296;
  assign n10406 = n10405 ^ n7806;
  assign n10409 = n10408 ^ n7689;
  assign n10436 = n10435 ^ n10408;
  assign n10437 = ~n10409 & ~n10436;
  assign n10438 = n10437 ^ n7689;
  assign n10439 = n10438 ^ n10405;
  assign n10440 = ~n10406 & n10439;
  assign n10441 = n10440 ^ n7806;
  assign n10442 = n10441 ^ n10403;
  assign n10443 = n10404 & ~n10442;
  assign n10444 = n10443 ^ n7834;
  assign n10445 = n10444 ^ n10401;
  assign n10446 = ~n10402 & n10445;
  assign n10447 = n10446 ^ n7865;
  assign n10448 = n10447 ^ n10399;
  assign n10449 = n10400 & ~n10448;
  assign n10450 = n10449 ^ n7939;
  assign n10451 = n10450 ^ n10396;
  assign n10452 = n10397 & ~n10451;
  assign n10453 = n10452 ^ n7932;
  assign n10454 = n10453 ^ n10394;
  assign n10455 = n10395 & ~n10454;
  assign n10456 = n10455 ^ n7226;
  assign n10457 = n10456 ^ n10391;
  assign n10458 = ~n10392 & n10457;
  assign n10459 = n10458 ^ n7220;
  assign n10460 = n10459 ^ n10388;
  assign n10461 = n10389 & n10460;
  assign n10462 = n10461 ^ n7215;
  assign n10463 = n10462 ^ n10385;
  assign n10464 = ~n10386 & ~n10463;
  assign n10465 = n10464 ^ n7212;
  assign n10471 = n10465 ^ n7263;
  assign n10371 = n8572 ^ n8100;
  assign n10372 = ~n9180 & n10371;
  assign n10373 = n10372 ^ n8100;
  assign n10267 = n10266 ^ n10263;
  assign n10367 = n10366 ^ n10263;
  assign n10368 = ~n10267 & n10367;
  assign n10369 = n10368 ^ n10266;
  assign n10370 = n10369 ^ n10261;
  assign n10382 = n10373 ^ n10370;
  assign n10472 = n10471 ^ n10382;
  assign n10473 = n10462 ^ n7212;
  assign n10474 = n10473 ^ n10385;
  assign n10475 = n10459 ^ n7215;
  assign n10476 = n10475 ^ n10388;
  assign n10477 = n10450 ^ n10397;
  assign n10478 = n10444 ^ n10402;
  assign n10490 = n10487 & n10489;
  assign n10491 = n10438 ^ n10406;
  assign n10492 = n10490 & ~n10491;
  assign n10493 = n10441 ^ n10404;
  assign n10494 = n10492 & n10493;
  assign n10495 = ~n10478 & n10494;
  assign n10496 = n10447 ^ n7939;
  assign n10497 = n10496 ^ n10399;
  assign n10498 = ~n10495 & ~n10497;
  assign n10499 = n10477 & ~n10498;
  assign n10500 = n10453 ^ n10395;
  assign n10501 = ~n10499 & ~n10500;
  assign n10502 = n10456 ^ n10392;
  assign n10503 = ~n10501 & ~n10502;
  assign n10504 = ~n10476 & ~n10503;
  assign n10505 = ~n10474 & n10504;
  assign n10506 = n10472 & ~n10505;
  assign n10383 = n10382 ^ n7263;
  assign n10466 = n10465 ^ n10382;
  assign n10467 = n10383 & n10466;
  assign n10468 = n10467 ^ n7263;
  assign n10469 = n10468 ^ n7267;
  assign n10374 = n10373 ^ n10261;
  assign n10375 = n10370 & ~n10374;
  assign n10376 = n10375 ^ n10373;
  assign n10257 = n8039 ^ n7910;
  assign n10258 = n9228 & ~n10257;
  assign n10259 = n10258 ^ n8039;
  assign n10260 = n10259 ^ n10256;
  assign n10381 = n10376 ^ n10260;
  assign n10470 = n10469 ^ n10381;
  assign n10514 = n10506 ^ n10470;
  assign n10515 = n10514 ^ x385;
  assign n10516 = n10505 ^ n10472;
  assign n10517 = n10516 ^ x386;
  assign n10518 = n10504 ^ n10474;
  assign n10519 = n10518 ^ x387;
  assign n10520 = n10503 ^ n10476;
  assign n10521 = n10520 ^ x388;
  assign n10522 = n10502 ^ n10501;
  assign n10523 = n10522 ^ x389;
  assign n10524 = n10500 ^ n10499;
  assign n10525 = n10524 ^ x390;
  assign n10527 = n10497 ^ n10495;
  assign n10528 = n10527 ^ x392;
  assign n10529 = n10494 ^ n10478;
  assign n10530 = n10529 ^ x393;
  assign n10531 = n10493 ^ n10492;
  assign n10532 = n10531 ^ x394;
  assign n10533 = n10491 ^ n10490;
  assign n10534 = n10533 ^ x395;
  assign n10536 = n10535 ^ x396;
  assign n10560 = n10559 ^ n10535;
  assign n10561 = n10536 & ~n10560;
  assign n10562 = n10561 ^ x396;
  assign n10563 = n10562 ^ n10533;
  assign n10564 = ~n10534 & n10563;
  assign n10565 = n10564 ^ x395;
  assign n10566 = n10565 ^ n10531;
  assign n10567 = n10532 & ~n10566;
  assign n10568 = n10567 ^ x394;
  assign n10569 = n10568 ^ n10529;
  assign n10570 = ~n10530 & n10569;
  assign n10571 = n10570 ^ x393;
  assign n10572 = n10571 ^ n10527;
  assign n10573 = ~n10528 & n10572;
  assign n10574 = n10573 ^ x392;
  assign n10526 = n10498 ^ n10477;
  assign n10575 = n10574 ^ n10526;
  assign n10576 = n10526 ^ x391;
  assign n10577 = n10575 & ~n10576;
  assign n10578 = n10577 ^ x391;
  assign n10579 = n10578 ^ n10524;
  assign n10580 = ~n10525 & n10579;
  assign n10581 = n10580 ^ x390;
  assign n10582 = n10581 ^ n10522;
  assign n10583 = n10523 & ~n10582;
  assign n10584 = n10583 ^ x389;
  assign n10585 = n10584 ^ n10520;
  assign n10586 = ~n10521 & n10585;
  assign n10587 = n10586 ^ x388;
  assign n10588 = n10587 ^ n10518;
  assign n10589 = n10519 & ~n10588;
  assign n10590 = n10589 ^ x387;
  assign n10591 = n10590 ^ n10516;
  assign n10592 = ~n10517 & n10591;
  assign n10593 = n10592 ^ x386;
  assign n10594 = n10593 ^ n10514;
  assign n10595 = n10515 & ~n10594;
  assign n10596 = n10595 ^ x385;
  assign n10597 = n10596 ^ x384;
  assign n10509 = n10381 ^ n7267;
  assign n10510 = n10468 ^ n10381;
  assign n10511 = n10509 & n10510;
  assign n10512 = n10511 ^ n7267;
  assign n10507 = n10470 & ~n10506;
  assign n10377 = n10376 ^ n10256;
  assign n10378 = n10260 & ~n10377;
  assign n10379 = n10378 ^ n10259;
  assign n10251 = n8038 ^ n7903;
  assign n10252 = n9268 & n10251;
  assign n10253 = n10252 ^ n8038;
  assign n10250 = n9875 ^ n9777;
  assign n10254 = n10253 ^ n10250;
  assign n10255 = n10254 ^ n7306;
  assign n10380 = n10379 ^ n10255;
  assign n10508 = n10507 ^ n10380;
  assign n10513 = n10512 ^ n10508;
  assign n10598 = n10597 ^ n10513;
  assign n10602 = n10601 ^ n10598;
  assign n10605 = n9366 ^ n8709;
  assign n10606 = n9350 & n10605;
  assign n10607 = n10606 ^ n8709;
  assign n10603 = n10593 ^ x385;
  assign n10604 = n10603 ^ n10514;
  assign n10608 = n10607 ^ n10604;
  assign n10614 = n9467 ^ n8621;
  assign n10615 = n9936 & n10614;
  assign n10616 = n10615 ^ n8621;
  assign n10612 = n10587 ^ x387;
  assign n10613 = n10612 ^ n10518;
  assign n10617 = n10616 ^ n10613;
  assign n10618 = n10584 ^ x388;
  assign n10619 = n10618 ^ n10520;
  assign n10620 = n9473 ^ n7897;
  assign n10621 = ~n9364 & ~n10620;
  assign n10622 = n10621 ^ n7897;
  assign n10623 = ~n10619 & ~n10622;
  assign n10624 = n10623 ^ n10613;
  assign n10625 = n10617 & n10624;
  assign n10626 = n10625 ^ n10623;
  assign n10609 = n9461 ^ n8675;
  assign n10610 = n9357 & n10609;
  assign n10611 = n10610 ^ n8675;
  assign n10627 = n10626 ^ n10611;
  assign n10628 = n10590 ^ x386;
  assign n10629 = n10628 ^ n10516;
  assign n10630 = n10629 ^ n10626;
  assign n10631 = n10627 & n10630;
  assign n10632 = n10631 ^ n10611;
  assign n10633 = n10632 ^ n10604;
  assign n10634 = ~n10608 & ~n10633;
  assign n10635 = n10634 ^ n10607;
  assign n10636 = n10635 ^ n10598;
  assign n10637 = ~n10602 & ~n10636;
  assign n10638 = n10637 ^ n10601;
  assign n10639 = n10638 ^ n10245;
  assign n10640 = n10249 & ~n10639;
  assign n10641 = n10640 ^ n10248;
  assign n10642 = n10641 ^ n10243;
  assign n10643 = n10244 & ~n10642;
  assign n10644 = n10643 ^ n10242;
  assign n10646 = n10645 ^ n10644;
  assign n10647 = n9343 ^ n8841;
  assign n10648 = ~n9960 & ~n10647;
  assign n10649 = n10648 ^ n8841;
  assign n10650 = n10649 ^ n10644;
  assign n10651 = ~n10646 & ~n10650;
  assign n10652 = n10651 ^ n10645;
  assign n10653 = n10652 ^ n10238;
  assign n10654 = n10239 & n10653;
  assign n10655 = n10654 ^ n10236;
  assign n10656 = n10655 ^ n10232;
  assign n10657 = ~n10233 & ~n10656;
  assign n10658 = n10657 ^ n10231;
  assign n10659 = n10658 ^ n10223;
  assign n10660 = ~n10228 & ~n10659;
  assign n10661 = n10660 ^ n10227;
  assign n10662 = n10661 ^ n10215;
  assign n10663 = n10221 & ~n10662;
  assign n10664 = n10663 ^ n10220;
  assign n10665 = n10664 ^ n10208;
  assign n10666 = n10213 & n10665;
  assign n10667 = n10666 ^ n10212;
  assign n10668 = n10667 ^ n10200;
  assign n10669 = n10206 & n10668;
  assign n10670 = n10669 ^ n10205;
  assign n10671 = n10670 ^ n10198;
  assign n10672 = n10199 & n10671;
  assign n10673 = n10672 ^ n10197;
  assign n10674 = n10673 ^ n10192;
  assign n10675 = n10193 & n10674;
  assign n10676 = n10675 ^ n10191;
  assign n10677 = n10676 ^ n10185;
  assign n10678 = ~n10186 & n10677;
  assign n10679 = n10678 ^ n10183;
  assign n10680 = n10679 ^ n10178;
  assign n10681 = ~n10179 & ~n10680;
  assign n10682 = n10681 ^ n10177;
  assign n10683 = n10682 ^ n10172;
  assign n10684 = ~n10173 & ~n10683;
  assign n10685 = n10684 ^ n10170;
  assign n10686 = n10685 ^ n10160;
  assign n10687 = n10166 & n10686;
  assign n10688 = n10687 ^ n10165;
  assign n10803 = n10693 ^ n10688;
  assign n10804 = ~n10694 & ~n10803;
  assign n10805 = n10804 ^ n10691;
  assign n10870 = n10806 ^ n10805;
  assign n10871 = ~n10810 & n10870;
  assign n10872 = n10871 ^ n10809;
  assign n10868 = n10553 ^ x398;
  assign n10869 = n10868 ^ n10539;
  assign n10873 = n10872 ^ n10869;
  assign n10865 = n9377 ^ n9167;
  assign n10866 = n10271 & n10865;
  assign n10867 = n10866 ^ n9167;
  assign n10997 = n10869 ^ n10867;
  assign n10998 = ~n10873 & ~n10997;
  assign n10999 = n10998 ^ n10867;
  assign n11091 = n10999 ^ n10993;
  assign n11092 = n11090 & ~n11091;
  assign n11093 = n11092 ^ n10996;
  assign n11094 = n11093 ^ n11085;
  assign n11095 = ~n11089 & n11094;
  assign n11096 = n11095 ^ n11088;
  assign n11083 = n10562 ^ n10534;
  assign n11097 = n11096 ^ n11083;
  assign n11136 = n11100 ^ n11097;
  assign n11137 = n11136 ^ n7810;
  assign n11138 = n11093 ^ n11089;
  assign n11139 = n11138 ^ n7915;
  assign n11000 = n10999 ^ n10996;
  assign n11001 = n11000 ^ n10993;
  assign n11140 = n11001 ^ n8188;
  assign n10874 = n10873 ^ n10867;
  assign n10875 = n10874 ^ n7918;
  assign n10811 = n10810 ^ n10805;
  assign n10812 = n10811 ^ n7920;
  assign n10695 = n10694 ^ n10688;
  assign n10696 = n10695 ^ n7925;
  assign n10697 = n10685 ^ n10166;
  assign n10698 = n10697 ^ n7931;
  assign n10699 = n10682 ^ n10173;
  assign n10700 = n10699 ^ n7937;
  assign n10701 = n10679 ^ n10179;
  assign n10702 = n10701 ^ n7948;
  assign n10703 = n10676 ^ n10183;
  assign n10704 = n10703 ^ n10185;
  assign n10705 = n10704 ^ n7953;
  assign n10706 = n10673 ^ n10193;
  assign n10707 = n10706 ^ n7959;
  assign n10708 = n10670 ^ n10199;
  assign n10709 = n10708 ^ n7964;
  assign n10710 = n10667 ^ n10206;
  assign n10711 = n10710 ^ n7970;
  assign n10712 = n10664 ^ n10213;
  assign n10713 = n10712 ^ n7975;
  assign n10714 = n10661 ^ n10221;
  assign n10715 = n10714 ^ n7978;
  assign n10716 = n10658 ^ n10228;
  assign n10717 = n10716 ^ n7986;
  assign n10718 = n10655 ^ n10233;
  assign n10719 = n10718 ^ n7989;
  assign n10720 = n10652 ^ n10239;
  assign n10721 = n10720 ^ n7994;
  assign n10722 = n10641 ^ n10244;
  assign n10723 = n10722 ^ n8005;
  assign n10724 = n10638 ^ n10248;
  assign n10725 = n10724 ^ n10245;
  assign n10726 = n10725 ^ n7375;
  assign n10727 = n10635 ^ n10601;
  assign n10728 = n10727 ^ n10598;
  assign n10729 = n10728 ^ n7899;
  assign n10730 = n10632 ^ n10607;
  assign n10731 = n10730 ^ n10604;
  assign n10732 = n10731 ^ n7906;
  assign n10733 = n10629 ^ n10627;
  assign n10734 = n10733 ^ n8022;
  assign n10735 = n10622 ^ n10619;
  assign n10736 = n8033 & n10735;
  assign n10737 = n10736 ^ n8028;
  assign n10738 = n10623 ^ n10616;
  assign n10739 = n10738 ^ n10613;
  assign n10740 = n10739 ^ n10736;
  assign n10741 = n10737 & n10740;
  assign n10742 = n10741 ^ n8028;
  assign n10743 = n10742 ^ n10733;
  assign n10744 = n10734 & n10743;
  assign n10745 = n10744 ^ n8022;
  assign n10746 = n10745 ^ n10731;
  assign n10747 = n10732 & ~n10746;
  assign n10748 = n10747 ^ n7906;
  assign n10749 = n10748 ^ n10728;
  assign n10750 = ~n10729 & n10749;
  assign n10751 = n10750 ^ n7899;
  assign n10752 = n10751 ^ n10725;
  assign n10753 = n10726 & n10752;
  assign n10754 = n10753 ^ n7375;
  assign n10755 = n10754 ^ n10722;
  assign n10756 = ~n10723 & ~n10755;
  assign n10757 = n10756 ^ n8005;
  assign n10758 = n10757 ^ n8002;
  assign n10759 = n10649 ^ n10645;
  assign n10760 = n10759 ^ n10644;
  assign n10761 = n10760 ^ n10757;
  assign n10762 = ~n10758 & ~n10761;
  assign n10763 = n10762 ^ n8002;
  assign n10764 = n10763 ^ n10720;
  assign n10765 = ~n10721 & n10764;
  assign n10766 = n10765 ^ n7994;
  assign n10767 = n10766 ^ n10718;
  assign n10768 = ~n10719 & n10767;
  assign n10769 = n10768 ^ n7989;
  assign n10770 = n10769 ^ n10716;
  assign n10771 = ~n10717 & ~n10770;
  assign n10772 = n10771 ^ n7986;
  assign n10773 = n10772 ^ n10714;
  assign n10774 = n10715 & n10773;
  assign n10775 = n10774 ^ n7978;
  assign n10776 = n10775 ^ n10712;
  assign n10777 = n10713 & ~n10776;
  assign n10778 = n10777 ^ n7975;
  assign n10779 = n10778 ^ n10710;
  assign n10780 = ~n10711 & n10779;
  assign n10781 = n10780 ^ n7970;
  assign n10782 = n10781 ^ n10708;
  assign n10783 = n10709 & ~n10782;
  assign n10784 = n10783 ^ n7964;
  assign n10785 = n10784 ^ n10706;
  assign n10786 = ~n10707 & n10785;
  assign n10787 = n10786 ^ n7959;
  assign n10788 = n10787 ^ n10704;
  assign n10789 = n10705 & n10788;
  assign n10790 = n10789 ^ n7953;
  assign n10791 = n10790 ^ n10701;
  assign n10792 = ~n10702 & ~n10791;
  assign n10793 = n10792 ^ n7948;
  assign n10794 = n10793 ^ n10699;
  assign n10795 = n10700 & ~n10794;
  assign n10796 = n10795 ^ n7937;
  assign n10797 = n10796 ^ n10697;
  assign n10798 = ~n10698 & ~n10797;
  assign n10799 = n10798 ^ n7931;
  assign n10800 = n10799 ^ n10695;
  assign n10801 = n10696 & n10800;
  assign n10802 = n10801 ^ n7925;
  assign n10862 = n10811 ^ n10802;
  assign n10863 = ~n10812 & n10862;
  assign n10864 = n10863 ^ n7920;
  assign n10989 = n10874 ^ n10864;
  assign n10990 = n10875 & n10989;
  assign n10991 = n10990 ^ n7918;
  assign n11141 = n11001 ^ n10991;
  assign n11142 = n11140 & ~n11141;
  assign n11143 = n11142 ^ n8188;
  assign n11144 = n11143 ^ n11138;
  assign n11145 = n11139 & n11144;
  assign n11146 = n11145 ^ n7915;
  assign n11147 = n11146 ^ n11136;
  assign n11148 = ~n11137 & n11147;
  assign n11149 = n11148 ^ n7810;
  assign n11101 = n11100 ^ n11083;
  assign n11102 = ~n11097 & n11101;
  assign n11103 = n11102 ^ n11100;
  assign n11079 = n9144 ^ n8591;
  assign n11080 = ~n10250 & n11079;
  assign n11081 = n11080 ^ n8591;
  assign n11133 = n11103 ^ n11081;
  assign n11077 = n10565 ^ x394;
  assign n11078 = n11077 ^ n10531;
  assign n11134 = n11133 ^ n11078;
  assign n11135 = n11134 ^ n7847;
  assign n11165 = n11149 ^ n11135;
  assign n11160 = n11143 ^ n11139;
  assign n10992 = n10991 ^ n8188;
  assign n11002 = n11001 ^ n10992;
  assign n10813 = n10812 ^ n10802;
  assign n10814 = n10784 ^ n10707;
  assign n10815 = n10781 ^ n10709;
  assign n10816 = n10778 ^ n10711;
  assign n10817 = n10775 ^ n10713;
  assign n10818 = n10769 ^ n10717;
  assign n10819 = n10766 ^ n10719;
  assign n10820 = n10763 ^ n10721;
  assign n10821 = n10754 ^ n10723;
  assign n10822 = n10751 ^ n7375;
  assign n10823 = n10822 ^ n10725;
  assign n10824 = n10748 ^ n7899;
  assign n10825 = n10824 ^ n10728;
  assign n10826 = n10735 ^ n8033;
  assign n10827 = n10739 ^ n10737;
  assign n10828 = n10826 & ~n10827;
  assign n10829 = n10742 ^ n8022;
  assign n10830 = n10829 ^ n10733;
  assign n10831 = n10828 & n10830;
  assign n10832 = n10745 ^ n7906;
  assign n10833 = n10832 ^ n10731;
  assign n10834 = ~n10831 & n10833;
  assign n10835 = ~n10825 & n10834;
  assign n10836 = ~n10823 & ~n10835;
  assign n10837 = ~n10821 & n10836;
  assign n10838 = n10760 ^ n8002;
  assign n10839 = n10838 ^ n10757;
  assign n10840 = ~n10837 & ~n10839;
  assign n10841 = n10820 & n10840;
  assign n10842 = ~n10819 & ~n10841;
  assign n10843 = ~n10818 & n10842;
  assign n10844 = n10772 ^ n10715;
  assign n10845 = ~n10843 & n10844;
  assign n10846 = ~n10817 & n10845;
  assign n10847 = n10816 & n10846;
  assign n10848 = ~n10815 & n10847;
  assign n10849 = ~n10814 & ~n10848;
  assign n10850 = n10787 ^ n10705;
  assign n10851 = n10849 & n10850;
  assign n10852 = n10790 ^ n10702;
  assign n10853 = ~n10851 & ~n10852;
  assign n10854 = n10793 ^ n10700;
  assign n10855 = ~n10853 & n10854;
  assign n10856 = n10796 ^ n7931;
  assign n10857 = n10856 ^ n10697;
  assign n10858 = n10855 & ~n10857;
  assign n10859 = n10799 ^ n10696;
  assign n10860 = n10858 & ~n10859;
  assign n10861 = ~n10813 & n10860;
  assign n10876 = n10875 ^ n10864;
  assign n11003 = n10861 & n10876;
  assign n11161 = n11002 & ~n11003;
  assign n11162 = ~n11160 & ~n11161;
  assign n11163 = n11146 ^ n11137;
  assign n11164 = ~n11162 & n11163;
  assign n11199 = n11165 ^ n11164;
  assign n11200 = n11199 ^ x421;
  assign n11201 = n11163 ^ n11162;
  assign n11202 = n11201 ^ x422;
  assign n11203 = n11161 ^ n11160;
  assign n11204 = n11203 ^ x423;
  assign n11004 = n11003 ^ n11002;
  assign n11205 = n11004 ^ x424;
  assign n10877 = n10876 ^ n10861;
  assign n10878 = n10877 ^ x425;
  assign n10879 = n10860 ^ n10813;
  assign n10880 = n10879 ^ x426;
  assign n10881 = n10859 ^ n10858;
  assign n10882 = n10881 ^ x427;
  assign n10883 = n10857 ^ n10855;
  assign n10884 = n10883 ^ x428;
  assign n10885 = n10854 ^ n10853;
  assign n10886 = n10885 ^ x429;
  assign n10887 = n10852 ^ n10851;
  assign n10888 = n10887 ^ x430;
  assign n10890 = n10848 ^ n10814;
  assign n10891 = n10890 ^ x432;
  assign n10892 = n10847 ^ n10815;
  assign n10893 = n10892 ^ x433;
  assign n10894 = n10846 ^ n10816;
  assign n10895 = n10894 ^ x434;
  assign n10896 = n10845 ^ n10817;
  assign n10897 = n10896 ^ x435;
  assign n10898 = n10844 ^ n10843;
  assign n10899 = n10898 ^ x436;
  assign n10900 = n10842 ^ n10818;
  assign n10901 = n10900 ^ x437;
  assign n10902 = n10841 ^ n10819;
  assign n10903 = n10902 ^ x438;
  assign n10904 = n10840 ^ n10820;
  assign n10905 = n10904 ^ x439;
  assign n10906 = n10836 ^ n10821;
  assign n10907 = n10906 ^ x441;
  assign n10908 = n10835 ^ n10823;
  assign n10909 = n10908 ^ x442;
  assign n10910 = n10834 ^ n10825;
  assign n10911 = n10910 ^ x443;
  assign n10912 = n10833 ^ n10831;
  assign n10913 = n10912 ^ x444;
  assign n10914 = n10830 ^ n10828;
  assign n10915 = n10914 ^ x445;
  assign n10916 = x447 & ~n10826;
  assign n10917 = n10916 ^ x446;
  assign n10918 = n10827 ^ n10826;
  assign n10919 = n10918 ^ n10916;
  assign n10920 = n10917 & n10919;
  assign n10921 = n10920 ^ x446;
  assign n10922 = n10921 ^ n10914;
  assign n10923 = n10915 & ~n10922;
  assign n10924 = n10923 ^ x445;
  assign n10925 = n10924 ^ n10912;
  assign n10926 = n10913 & ~n10925;
  assign n10927 = n10926 ^ x444;
  assign n10928 = n10927 ^ n10910;
  assign n10929 = n10911 & ~n10928;
  assign n10930 = n10929 ^ x443;
  assign n10931 = n10930 ^ n10908;
  assign n10932 = n10909 & ~n10931;
  assign n10933 = n10932 ^ x442;
  assign n10934 = n10933 ^ n10906;
  assign n10935 = ~n10907 & n10934;
  assign n10936 = n10935 ^ x441;
  assign n10937 = n10936 ^ x440;
  assign n10938 = n10839 ^ n10837;
  assign n10939 = n10938 ^ n10936;
  assign n10940 = n10937 & n10939;
  assign n10941 = n10940 ^ x440;
  assign n10942 = n10941 ^ n10904;
  assign n10943 = ~n10905 & n10942;
  assign n10944 = n10943 ^ x439;
  assign n10945 = n10944 ^ n10902;
  assign n10946 = n10903 & ~n10945;
  assign n10947 = n10946 ^ x438;
  assign n10948 = n10947 ^ n10900;
  assign n10949 = ~n10901 & n10948;
  assign n10950 = n10949 ^ x437;
  assign n10951 = n10950 ^ n10898;
  assign n10952 = n10899 & ~n10951;
  assign n10953 = n10952 ^ x436;
  assign n10954 = n10953 ^ n10896;
  assign n10955 = n10897 & ~n10954;
  assign n10956 = n10955 ^ x435;
  assign n10957 = n10956 ^ n10894;
  assign n10958 = ~n10895 & n10957;
  assign n10959 = n10958 ^ x434;
  assign n10960 = n10959 ^ n10892;
  assign n10961 = n10893 & ~n10960;
  assign n10962 = n10961 ^ x433;
  assign n10963 = n10962 ^ n10890;
  assign n10964 = n10891 & ~n10963;
  assign n10965 = n10964 ^ x432;
  assign n10889 = n10850 ^ n10849;
  assign n10966 = n10965 ^ n10889;
  assign n10967 = n10889 ^ x431;
  assign n10968 = ~n10966 & n10967;
  assign n10969 = n10968 ^ x431;
  assign n10970 = n10969 ^ n10887;
  assign n10971 = ~n10888 & n10970;
  assign n10972 = n10971 ^ x430;
  assign n10973 = n10972 ^ n10885;
  assign n10974 = ~n10886 & n10973;
  assign n10975 = n10974 ^ x429;
  assign n10976 = n10975 ^ n10883;
  assign n10977 = ~n10884 & n10976;
  assign n10978 = n10977 ^ x428;
  assign n10979 = n10978 ^ n10881;
  assign n10980 = ~n10882 & n10979;
  assign n10981 = n10980 ^ x427;
  assign n10982 = n10981 ^ n10879;
  assign n10983 = ~n10880 & n10982;
  assign n10984 = n10983 ^ x426;
  assign n10985 = n10984 ^ n10877;
  assign n10986 = n10878 & ~n10985;
  assign n10987 = n10986 ^ x425;
  assign n11206 = n11004 ^ n10987;
  assign n11207 = n11205 & ~n11206;
  assign n11208 = n11207 ^ x424;
  assign n11209 = n11208 ^ n11203;
  assign n11210 = n11204 & ~n11209;
  assign n11211 = n11210 ^ x423;
  assign n11212 = n11211 ^ n11201;
  assign n11213 = n11202 & ~n11212;
  assign n11214 = n11213 ^ x422;
  assign n11215 = n11214 ^ n11199;
  assign n11216 = n11200 & ~n11215;
  assign n11217 = n11216 ^ x421;
  assign n11254 = n11217 ^ x420;
  assign n11166 = ~n11164 & ~n11165;
  assign n11150 = n11149 ^ n11134;
  assign n11151 = ~n11135 & ~n11150;
  assign n11152 = n11151 ^ n7847;
  assign n11158 = n11152 ^ n7883;
  assign n11082 = n11081 ^ n11078;
  assign n11104 = n11103 ^ n11078;
  assign n11105 = ~n11082 & n11104;
  assign n11106 = n11105 ^ n11081;
  assign n11073 = n9180 ^ n8583;
  assign n11074 = n9916 & n11073;
  assign n11075 = n11074 ^ n8583;
  assign n11130 = n11106 ^ n11075;
  assign n11071 = n10568 ^ x393;
  assign n11072 = n11071 ^ n10529;
  assign n11131 = n11130 ^ n11072;
  assign n11159 = n11158 ^ n11131;
  assign n11197 = n11166 ^ n11159;
  assign n11255 = n11254 ^ n11197;
  assign n11251 = n9473 ^ n9357;
  assign n11252 = n10245 & n11251;
  assign n11253 = n11252 ^ n9473;
  assign n11333 = n11255 ^ n11253;
  assign n11397 = n11333 ^ n7897;
  assign n11667 = n11397 ^ x479;
  assign n11046 = n10921 ^ n10915;
  assign n12632 = n11046 ^ n10645;
  assign n12633 = ~n11667 & ~n12632;
  assign n12634 = n12633 ^ n10645;
  assign n11547 = n10956 ^ x434;
  assign n11548 = n11547 ^ n10894;
  assign n11544 = n10283 ^ n9395;
  assign n11545 = ~n10993 & ~n11544;
  assign n11546 = n11545 ^ n9395;
  assign n11549 = n11548 ^ n11546;
  assign n11447 = n10953 ^ n10897;
  assign n11444 = n10162 ^ n9401;
  assign n11445 = n10869 & n11444;
  assign n11446 = n11445 ^ n9401;
  assign n11448 = n11447 ^ n11446;
  assign n11431 = n10950 ^ x436;
  assign n11432 = n11431 ^ n10898;
  assign n11428 = n10167 ^ n9402;
  assign n11429 = ~n10806 & ~n11428;
  assign n11430 = n11429 ^ n9402;
  assign n11433 = n11432 ^ n11430;
  assign n11386 = n10947 ^ n10901;
  assign n11383 = n10174 ^ n9404;
  assign n11384 = ~n10693 & ~n11383;
  assign n11385 = n11384 ^ n9404;
  assign n11387 = n11386 ^ n11385;
  assign n11302 = n10944 ^ n10903;
  assign n11299 = n10180 ^ n9409;
  assign n11300 = ~n10160 & ~n11299;
  assign n11301 = n11300 ^ n9409;
  assign n11303 = n11302 ^ n11301;
  assign n11014 = n10941 ^ n10905;
  assign n11011 = n10188 ^ n9411;
  assign n11012 = ~n10172 & n11011;
  assign n11013 = n11012 ^ n9411;
  assign n11015 = n11014 ^ n11013;
  assign n11019 = n10938 ^ n10937;
  assign n11016 = n10194 ^ n9416;
  assign n11017 = n10178 & n11016;
  assign n11018 = n11017 ^ n9416;
  assign n11020 = n11019 ^ n11018;
  assign n11024 = n10933 ^ n10907;
  assign n11021 = n10202 ^ n9422;
  assign n11022 = ~n10185 & ~n11021;
  assign n11023 = n11022 ^ n9422;
  assign n11025 = n11024 ^ n11023;
  assign n11029 = n10930 ^ x442;
  assign n11030 = n11029 ^ n10908;
  assign n11026 = n10209 ^ n9430;
  assign n11027 = n10192 & n11026;
  assign n11028 = n11027 ^ n9430;
  assign n11031 = n11030 ^ n11028;
  assign n11035 = n10927 ^ n10911;
  assign n11032 = n10217 ^ n8782;
  assign n11033 = ~n10198 & ~n11032;
  assign n11034 = n11033 ^ n8782;
  assign n11036 = n11035 ^ n11034;
  assign n11039 = n10224 ^ n9336;
  assign n11040 = n10200 & ~n11039;
  assign n11041 = n11040 ^ n9336;
  assign n11037 = n10924 ^ x444;
  assign n11038 = n11037 ^ n10912;
  assign n11042 = n11041 ^ n11038;
  assign n11043 = n10153 ^ n9343;
  assign n11044 = ~n10208 & ~n11043;
  assign n11045 = n11044 ^ n9343;
  assign n11047 = n11046 ^ n11045;
  assign n11051 = n10918 ^ n10917;
  assign n11048 = n10041 ^ n9352;
  assign n11049 = n10215 & ~n11048;
  assign n11050 = n11049 ^ n9352;
  assign n11052 = n11051 ^ n11050;
  assign n11054 = n9960 ^ n9359;
  assign n11055 = ~n10223 & ~n11054;
  assign n11056 = n11055 ^ n9359;
  assign n11053 = n10826 ^ x447;
  assign n11057 = n11056 ^ n11053;
  assign n11232 = n9452 ^ n9334;
  assign n11233 = n10232 & ~n11232;
  assign n11234 = n11233 ^ n9452;
  assign n11114 = n9268 ^ n8572;
  assign n11115 = n9923 & n11114;
  assign n11116 = n11115 ^ n8572;
  assign n11067 = n9228 ^ n8578;
  assign n11068 = n9907 & n11067;
  assign n11069 = n11068 ^ n8578;
  assign n11065 = n10571 ^ x392;
  assign n11066 = n11065 ^ n10527;
  assign n11070 = n11069 ^ n11066;
  assign n11076 = n11075 ^ n11072;
  assign n11107 = n11106 ^ n11072;
  assign n11108 = n11076 & ~n11107;
  assign n11109 = n11108 ^ n11075;
  assign n11110 = n11109 ^ n11066;
  assign n11111 = ~n11070 & ~n11110;
  assign n11112 = n11111 ^ n11069;
  assign n11064 = n10575 ^ x391;
  assign n11113 = n11112 ^ n11064;
  assign n11169 = n11116 ^ n11113;
  assign n11178 = n11169 ^ n8100;
  assign n11128 = n11109 ^ n11069;
  assign n11129 = n11128 ^ n11066;
  assign n11170 = n11129 ^ n8070;
  assign n11132 = n11131 ^ n7883;
  assign n11153 = n11152 ^ n11131;
  assign n11154 = ~n11132 & ~n11153;
  assign n11155 = n11154 ^ n7883;
  assign n11171 = n11155 ^ n11129;
  assign n11172 = n11170 & ~n11171;
  assign n11173 = n11172 ^ n8070;
  assign n11179 = n11173 ^ n11169;
  assign n11180 = ~n11178 & n11179;
  assign n11181 = n11180 ^ n8100;
  assign n11182 = n11181 ^ n8039;
  assign n11121 = n9286 ^ n7910;
  assign n11122 = n9898 & n11121;
  assign n11123 = n11122 ^ n7910;
  assign n11117 = n11116 ^ n11064;
  assign n11118 = n11113 & ~n11117;
  assign n11119 = n11118 ^ n11116;
  assign n11006 = n10578 ^ x390;
  assign n11007 = n11006 ^ n10524;
  assign n11120 = n11119 ^ n11007;
  assign n11177 = n11123 ^ n11120;
  assign n11183 = n11182 ^ n11177;
  assign n11156 = n11155 ^ n8070;
  assign n11157 = n11156 ^ n11129;
  assign n11167 = ~n11159 & ~n11166;
  assign n11168 = ~n11157 & n11167;
  assign n11174 = n11173 ^ n8100;
  assign n11175 = n11174 ^ n11169;
  assign n11176 = ~n11168 & ~n11175;
  assign n11191 = n11183 ^ n11176;
  assign n11192 = n11191 ^ x417;
  assign n11193 = n11175 ^ n11168;
  assign n11194 = n11193 ^ x418;
  assign n11195 = n11167 ^ n11157;
  assign n11196 = n11195 ^ x419;
  assign n11198 = n11197 ^ x420;
  assign n11218 = n11217 ^ n11197;
  assign n11219 = ~n11198 & n11218;
  assign n11220 = n11219 ^ x420;
  assign n11221 = n11220 ^ n11195;
  assign n11222 = n11196 & ~n11221;
  assign n11223 = n11222 ^ x419;
  assign n11224 = n11223 ^ n11193;
  assign n11225 = n11194 & ~n11224;
  assign n11226 = n11225 ^ x418;
  assign n11227 = n11226 ^ n11191;
  assign n11228 = ~n11192 & n11227;
  assign n11229 = n11228 ^ x417;
  assign n11230 = n11229 ^ x416;
  assign n11186 = n11177 ^ n8039;
  assign n11187 = n11181 ^ n11177;
  assign n11188 = n11186 & ~n11187;
  assign n11189 = n11188 ^ n8039;
  assign n11184 = ~n11176 & ~n11183;
  assign n11124 = n11123 ^ n11007;
  assign n11125 = n11120 & n11124;
  assign n11126 = n11125 ^ n11123;
  assign n11061 = n10581 ^ n10523;
  assign n11058 = n9327 ^ n7903;
  assign n11059 = n9892 & n11058;
  assign n11060 = n11059 ^ n7903;
  assign n11062 = n11061 ^ n11060;
  assign n11063 = n11062 ^ n8038;
  assign n11127 = n11126 ^ n11063;
  assign n11185 = n11184 ^ n11127;
  assign n11190 = n11189 ^ n11185;
  assign n11231 = n11230 ^ n11190;
  assign n11235 = n11234 ^ n11231;
  assign n11238 = n9366 ^ n9341;
  assign n11239 = n10238 & ~n11238;
  assign n11240 = n11239 ^ n9366;
  assign n11236 = n11226 ^ x417;
  assign n11237 = n11236 ^ n11191;
  assign n11241 = n11240 ^ n11237;
  assign n11247 = n9467 ^ n9350;
  assign n11248 = n10243 & ~n11247;
  assign n11249 = n11248 ^ n9467;
  assign n11245 = n11220 ^ x419;
  assign n11246 = n11245 ^ n11195;
  assign n11250 = n11249 ^ n11246;
  assign n11256 = n11253 & ~n11255;
  assign n11257 = n11256 ^ n11246;
  assign n11258 = n11250 & n11257;
  assign n11259 = n11258 ^ n11256;
  assign n11242 = n9461 ^ n9347;
  assign n11243 = ~n10645 & ~n11242;
  assign n11244 = n11243 ^ n9461;
  assign n11260 = n11259 ^ n11244;
  assign n11261 = n11223 ^ x418;
  assign n11262 = n11261 ^ n11193;
  assign n11263 = n11262 ^ n11259;
  assign n11264 = n11260 & ~n11263;
  assign n11265 = n11264 ^ n11244;
  assign n11266 = n11265 ^ n11237;
  assign n11267 = n11241 & n11266;
  assign n11268 = n11267 ^ n11240;
  assign n11269 = n11268 ^ n11231;
  assign n11270 = n11235 & n11269;
  assign n11271 = n11270 ^ n11234;
  assign n11272 = n11271 ^ n11053;
  assign n11273 = ~n11057 & n11272;
  assign n11274 = n11273 ^ n11056;
  assign n11275 = n11274 ^ n11051;
  assign n11276 = ~n11052 & n11275;
  assign n11277 = n11276 ^ n11050;
  assign n11278 = n11277 ^ n11046;
  assign n11279 = ~n11047 & ~n11278;
  assign n11280 = n11279 ^ n11045;
  assign n11281 = n11280 ^ n11038;
  assign n11282 = ~n11042 & n11281;
  assign n11283 = n11282 ^ n11041;
  assign n11284 = n11283 ^ n11035;
  assign n11285 = ~n11036 & n11284;
  assign n11286 = n11285 ^ n11034;
  assign n11287 = n11286 ^ n11030;
  assign n11288 = n11031 & n11287;
  assign n11289 = n11288 ^ n11028;
  assign n11290 = n11289 ^ n11024;
  assign n11291 = ~n11025 & n11290;
  assign n11292 = n11291 ^ n11023;
  assign n11293 = n11292 ^ n11019;
  assign n11294 = ~n11020 & n11293;
  assign n11295 = n11294 ^ n11018;
  assign n11296 = n11295 ^ n11014;
  assign n11297 = ~n11015 & n11296;
  assign n11298 = n11297 ^ n11013;
  assign n11380 = n11302 ^ n11298;
  assign n11381 = ~n11303 & ~n11380;
  assign n11382 = n11381 ^ n11301;
  assign n11425 = n11386 ^ n11382;
  assign n11426 = n11387 & ~n11425;
  assign n11427 = n11426 ^ n11385;
  assign n11441 = n11432 ^ n11427;
  assign n11442 = ~n11433 & n11441;
  assign n11443 = n11442 ^ n11430;
  assign n11541 = n11447 ^ n11443;
  assign n11542 = ~n11448 & n11541;
  assign n11543 = n11542 ^ n11446;
  assign n11550 = n11549 ^ n11543;
  assign n11551 = n11550 ^ n8904;
  assign n11449 = n11448 ^ n11443;
  assign n11450 = n11449 ^ n8792;
  assign n11434 = n11433 ^ n11427;
  assign n11435 = n11434 ^ n8797;
  assign n11388 = n11387 ^ n11382;
  assign n11389 = n11388 ^ n8803;
  assign n11304 = n11303 ^ n11298;
  assign n11305 = n11304 ^ n8808;
  assign n11306 = n11295 ^ n11015;
  assign n11307 = n11306 ^ n8814;
  assign n11308 = n11292 ^ n11020;
  assign n11309 = n11308 ^ n8819;
  assign n11310 = n11289 ^ n11025;
  assign n11311 = n11310 ^ n8784;
  assign n11312 = n11286 ^ n11031;
  assign n11313 = n11312 ^ n8828;
  assign n11314 = n11283 ^ n11036;
  assign n11315 = n11314 ^ n8830;
  assign n11316 = n11280 ^ n11042;
  assign n11317 = n11316 ^ n8835;
  assign n11318 = n11277 ^ n11047;
  assign n11319 = n11318 ^ n8841;
  assign n11320 = n11274 ^ n11052;
  assign n11321 = n11320 ^ n8847;
  assign n11322 = n11271 ^ n11056;
  assign n11323 = n11322 ^ n11053;
  assign n11324 = n11323 ^ n8856;
  assign n11325 = n11268 ^ n11234;
  assign n11326 = n11325 ^ n11231;
  assign n11327 = n11326 ^ n8776;
  assign n11328 = n11265 ^ n11240;
  assign n11329 = n11328 ^ n11237;
  assign n11330 = n11329 ^ n8709;
  assign n11331 = n11262 ^ n11260;
  assign n11332 = n11331 ^ n8675;
  assign n11334 = ~n7897 & ~n11333;
  assign n11335 = n11334 ^ n8621;
  assign n11336 = n11256 ^ n11249;
  assign n11337 = n11336 ^ n11246;
  assign n11338 = n11337 ^ n11334;
  assign n11339 = ~n11335 & n11338;
  assign n11340 = n11339 ^ n8621;
  assign n11341 = n11340 ^ n11331;
  assign n11342 = n11332 & n11341;
  assign n11343 = n11342 ^ n8675;
  assign n11344 = n11343 ^ n11329;
  assign n11345 = ~n11330 & ~n11344;
  assign n11346 = n11345 ^ n8709;
  assign n11347 = n11346 ^ n11326;
  assign n11348 = ~n11327 & ~n11347;
  assign n11349 = n11348 ^ n8776;
  assign n11350 = n11349 ^ n11323;
  assign n11351 = ~n11324 & n11350;
  assign n11352 = n11351 ^ n8856;
  assign n11353 = n11352 ^ n11320;
  assign n11354 = ~n11321 & n11353;
  assign n11355 = n11354 ^ n8847;
  assign n11356 = n11355 ^ n11318;
  assign n11357 = ~n11319 & n11356;
  assign n11358 = n11357 ^ n8841;
  assign n11359 = n11358 ^ n11316;
  assign n11360 = n11317 & ~n11359;
  assign n11361 = n11360 ^ n8835;
  assign n11362 = n11361 ^ n11314;
  assign n11363 = ~n11315 & ~n11362;
  assign n11364 = n11363 ^ n8830;
  assign n11365 = n11364 ^ n11312;
  assign n11366 = ~n11313 & ~n11365;
  assign n11367 = n11366 ^ n8828;
  assign n11368 = n11367 ^ n11310;
  assign n11369 = ~n11311 & n11368;
  assign n11370 = n11369 ^ n8784;
  assign n11371 = n11370 ^ n11308;
  assign n11372 = n11309 & n11371;
  assign n11373 = n11372 ^ n8819;
  assign n11374 = n11373 ^ n11306;
  assign n11375 = ~n11307 & ~n11374;
  assign n11376 = n11375 ^ n8814;
  assign n11377 = n11376 ^ n11304;
  assign n11378 = n11305 & n11377;
  assign n11379 = n11378 ^ n8808;
  assign n11422 = n11388 ^ n11379;
  assign n11423 = ~n11389 & ~n11422;
  assign n11424 = n11423 ^ n8803;
  assign n11438 = n11434 ^ n11424;
  assign n11439 = n11435 & ~n11438;
  assign n11440 = n11439 ^ n8797;
  assign n11538 = n11449 ^ n11440;
  assign n11539 = ~n11450 & ~n11538;
  assign n11540 = n11539 ^ n8792;
  assign n11794 = n11550 ^ n11540;
  assign n11795 = ~n11551 & ~n11794;
  assign n11796 = n11795 ^ n8904;
  assign n11714 = n11548 ^ n11543;
  assign n11715 = n11549 & ~n11714;
  assign n11716 = n11715 ^ n11546;
  assign n11710 = n10277 ^ n9390;
  assign n11711 = n11085 & n11710;
  assign n11712 = n11711 ^ n9390;
  assign n11615 = n10959 ^ n10893;
  assign n11713 = n11712 ^ n11615;
  assign n11792 = n11716 ^ n11713;
  assign n11793 = n11792 ^ n8985;
  assign n11838 = n11796 ^ n11793;
  assign n11552 = n11551 ^ n11540;
  assign n11390 = n11389 ^ n11379;
  assign n11391 = n11376 ^ n11305;
  assign n11392 = n11370 ^ n11309;
  assign n11393 = n11367 ^ n11311;
  assign n11394 = n11358 ^ n11317;
  assign n11395 = n11340 ^ n8675;
  assign n11396 = n11395 ^ n11331;
  assign n11398 = n11337 ^ n11335;
  assign n11399 = n11397 & n11398;
  assign n11400 = ~n11396 & n11399;
  assign n11401 = n11343 ^ n11330;
  assign n11402 = ~n11400 & n11401;
  assign n11403 = n11346 ^ n11327;
  assign n11404 = n11402 & ~n11403;
  assign n11405 = n11349 ^ n11324;
  assign n11406 = ~n11404 & ~n11405;
  assign n11407 = n11352 ^ n11321;
  assign n11408 = n11406 & ~n11407;
  assign n11409 = n11355 ^ n11319;
  assign n11410 = ~n11408 & n11409;
  assign n11411 = ~n11394 & n11410;
  assign n11412 = n11361 ^ n11315;
  assign n11413 = ~n11411 & ~n11412;
  assign n11414 = n11364 ^ n11313;
  assign n11415 = n11413 & n11414;
  assign n11416 = n11393 & ~n11415;
  assign n11417 = ~n11392 & n11416;
  assign n11418 = n11373 ^ n11307;
  assign n11419 = n11417 & ~n11418;
  assign n11420 = ~n11391 & n11419;
  assign n11421 = n11390 & ~n11420;
  assign n11436 = n11435 ^ n11424;
  assign n11437 = n11421 & n11436;
  assign n11451 = n11450 ^ n11440;
  assign n11553 = ~n11437 & n11451;
  assign n11837 = n11552 & ~n11553;
  assign n11885 = n11838 ^ n11837;
  assign n11886 = n11885 ^ x460;
  assign n11554 = n11553 ^ n11552;
  assign n11555 = n11554 ^ x461;
  assign n11452 = n11451 ^ n11437;
  assign n11453 = n11452 ^ x462;
  assign n11455 = n11420 ^ n11390;
  assign n11456 = n11455 ^ x464;
  assign n11457 = n11419 ^ n11391;
  assign n11458 = n11457 ^ x465;
  assign n11459 = n11418 ^ n11417;
  assign n11460 = n11459 ^ x466;
  assign n11461 = n11416 ^ n11392;
  assign n11462 = n11461 ^ x467;
  assign n11463 = n11415 ^ n11393;
  assign n11464 = n11463 ^ x468;
  assign n11465 = n11414 ^ n11413;
  assign n11466 = n11465 ^ x469;
  assign n11467 = n11412 ^ n11411;
  assign n11468 = n11467 ^ x470;
  assign n11469 = n11410 ^ n11394;
  assign n11470 = n11469 ^ x471;
  assign n11471 = n11409 ^ n11408;
  assign n11472 = n11471 ^ x472;
  assign n11473 = n11407 ^ n11406;
  assign n11474 = n11473 ^ x473;
  assign n11475 = n11405 ^ n11404;
  assign n11476 = n11475 ^ x474;
  assign n11477 = n11403 ^ n11402;
  assign n11478 = n11477 ^ x475;
  assign n11479 = n11401 ^ n11400;
  assign n11480 = n11479 ^ x476;
  assign n11481 = n11399 ^ n11396;
  assign n11482 = n11481 ^ x477;
  assign n11483 = x479 & ~n11397;
  assign n11484 = n11483 ^ x478;
  assign n11485 = n11398 ^ n11397;
  assign n11486 = n11485 ^ n11483;
  assign n11487 = n11484 & ~n11486;
  assign n11488 = n11487 ^ x478;
  assign n11489 = n11488 ^ n11481;
  assign n11490 = ~n11482 & n11489;
  assign n11491 = n11490 ^ x477;
  assign n11492 = n11491 ^ n11479;
  assign n11493 = n11480 & ~n11492;
  assign n11494 = n11493 ^ x476;
  assign n11495 = n11494 ^ n11477;
  assign n11496 = n11478 & ~n11495;
  assign n11497 = n11496 ^ x475;
  assign n11498 = n11497 ^ n11475;
  assign n11499 = n11476 & ~n11498;
  assign n11500 = n11499 ^ x474;
  assign n11501 = n11500 ^ n11473;
  assign n11502 = ~n11474 & n11501;
  assign n11503 = n11502 ^ x473;
  assign n11504 = n11503 ^ n11471;
  assign n11505 = n11472 & ~n11504;
  assign n11506 = n11505 ^ x472;
  assign n11507 = n11506 ^ n11469;
  assign n11508 = n11470 & ~n11507;
  assign n11509 = n11508 ^ x471;
  assign n11510 = n11509 ^ n11467;
  assign n11511 = n11468 & ~n11510;
  assign n11512 = n11511 ^ x470;
  assign n11513 = n11512 ^ n11465;
  assign n11514 = n11466 & ~n11513;
  assign n11515 = n11514 ^ x469;
  assign n11516 = n11515 ^ n11463;
  assign n11517 = n11464 & ~n11516;
  assign n11518 = n11517 ^ x468;
  assign n11519 = n11518 ^ n11461;
  assign n11520 = n11462 & ~n11519;
  assign n11521 = n11520 ^ x467;
  assign n11522 = n11521 ^ n11459;
  assign n11523 = n11460 & ~n11522;
  assign n11524 = n11523 ^ x466;
  assign n11525 = n11524 ^ n11457;
  assign n11526 = n11458 & ~n11525;
  assign n11527 = n11526 ^ x465;
  assign n11528 = n11527 ^ n11455;
  assign n11529 = ~n11456 & n11528;
  assign n11530 = n11529 ^ x464;
  assign n11454 = n11436 ^ n11421;
  assign n11531 = n11530 ^ n11454;
  assign n11532 = n11454 ^ x463;
  assign n11533 = ~n11531 & n11532;
  assign n11534 = n11533 ^ x463;
  assign n11535 = n11534 ^ n11452;
  assign n11536 = n11453 & ~n11535;
  assign n11537 = n11536 ^ x462;
  assign n11887 = n11554 ^ n11537;
  assign n11888 = ~n11555 & n11887;
  assign n11889 = n11888 ^ x461;
  assign n11890 = n11889 ^ n11885;
  assign n11891 = n11886 & ~n11890;
  assign n11892 = n11891 ^ x460;
  assign n11839 = n11837 & n11838;
  assign n11797 = n11796 ^ n11792;
  assign n11798 = n11793 & n11797;
  assign n11799 = n11798 ^ n8985;
  assign n11717 = n11716 ^ n11615;
  assign n11718 = n11713 & n11717;
  assign n11719 = n11718 ^ n11712;
  assign n11706 = n10271 ^ n9384;
  assign n11707 = ~n11083 & ~n11706;
  assign n11708 = n11707 ^ n9384;
  assign n11608 = n10962 ^ x432;
  assign n11609 = n11608 ^ n10890;
  assign n11709 = n11708 ^ n11609;
  assign n11790 = n11719 ^ n11709;
  assign n11791 = n11790 ^ n9037;
  assign n11836 = n11799 ^ n11791;
  assign n11883 = n11839 ^ n11836;
  assign n11884 = n11883 ^ x459;
  assign n12165 = n11892 ^ n11884;
  assign n11675 = n11211 ^ x422;
  assign n11676 = n11675 ^ n11201;
  assign n12162 = n10619 ^ n9916;
  assign n12163 = n11676 & ~n12162;
  assign n12164 = n12163 ^ n9916;
  assign n12166 = n12165 ^ n12164;
  assign n12028 = n11889 ^ x460;
  assign n12029 = n12028 ^ n11885;
  assign n11677 = n11208 ^ n11204;
  assign n12025 = n11061 ^ n10250;
  assign n12026 = n11677 & ~n12025;
  assign n12027 = n12026 ^ n10250;
  assign n12030 = n12029 ^ n12027;
  assign n11556 = n11555 ^ n11537;
  assign n10988 = n10987 ^ x424;
  assign n11005 = n11004 ^ n10988;
  assign n11008 = n11007 ^ n10256;
  assign n11009 = n11005 & ~n11008;
  assign n11010 = n11009 ^ n10256;
  assign n11557 = n11556 ^ n11010;
  assign n11562 = n11534 ^ x462;
  assign n11563 = n11562 ^ n11452;
  assign n11558 = n10984 ^ n10878;
  assign n11559 = n11064 ^ n10261;
  assign n11560 = n11558 & n11559;
  assign n11561 = n11560 ^ n10261;
  assign n11564 = n11563 ^ n11561;
  assign n11570 = n11531 ^ x463;
  assign n11565 = n10981 ^ x426;
  assign n11566 = n11565 ^ n10879;
  assign n11567 = n11066 ^ n10263;
  assign n11568 = ~n11566 & n11567;
  assign n11569 = n11568 ^ n10263;
  assign n11571 = n11570 ^ n11569;
  assign n11576 = n11527 ^ x464;
  assign n11577 = n11576 ^ n11455;
  assign n11572 = n10978 ^ n10882;
  assign n11573 = n11072 ^ n10271;
  assign n11574 = ~n11572 & ~n11573;
  assign n11575 = n11574 ^ n10271;
  assign n11578 = n11577 ^ n11575;
  assign n11584 = n11524 ^ n11458;
  assign n11579 = n10975 ^ x428;
  assign n11580 = n11579 ^ n10883;
  assign n11581 = n11078 ^ n10277;
  assign n11582 = ~n11580 & n11581;
  assign n11583 = n11582 ^ n10277;
  assign n11585 = n11584 ^ n11583;
  assign n11590 = n11521 ^ x466;
  assign n11591 = n11590 ^ n11459;
  assign n11586 = n10972 ^ n10886;
  assign n11587 = n11083 ^ n10283;
  assign n11588 = ~n11586 & ~n11587;
  assign n11589 = n11588 ^ n10283;
  assign n11592 = n11591 ^ n11589;
  assign n11598 = n11518 ^ n11462;
  assign n11593 = n10969 ^ x430;
  assign n11594 = n11593 ^ n10887;
  assign n11595 = n11085 ^ n10162;
  assign n11596 = ~n11594 & ~n11595;
  assign n11597 = n11596 ^ n10162;
  assign n11599 = n11598 ^ n11597;
  assign n11602 = n10966 ^ x431;
  assign n11603 = n10993 ^ n10167;
  assign n11604 = n11602 & ~n11603;
  assign n11605 = n11604 ^ n10167;
  assign n11600 = n11515 ^ x468;
  assign n11601 = n11600 ^ n11463;
  assign n11606 = n11605 ^ n11601;
  assign n11610 = n10869 ^ n10174;
  assign n11611 = n11609 & n11610;
  assign n11612 = n11611 ^ n10174;
  assign n11607 = n11512 ^ n11466;
  assign n11613 = n11612 ^ n11607;
  assign n11616 = n10806 ^ n10180;
  assign n11617 = n11615 & ~n11616;
  assign n11618 = n11617 ^ n10180;
  assign n11614 = n11509 ^ n11468;
  assign n11619 = n11618 ^ n11614;
  assign n11622 = n10693 ^ n10188;
  assign n11623 = ~n11548 & ~n11622;
  assign n11624 = n11623 ^ n10188;
  assign n11620 = n11506 ^ x471;
  assign n11621 = n11620 ^ n11469;
  assign n11625 = n11624 ^ n11621;
  assign n11628 = n10194 ^ n10160;
  assign n11629 = n11447 & ~n11628;
  assign n11630 = n11629 ^ n10194;
  assign n11626 = n11503 ^ x472;
  assign n11627 = n11626 ^ n11471;
  assign n11631 = n11630 ^ n11627;
  assign n11633 = n10202 ^ n10172;
  assign n11634 = n11432 & n11633;
  assign n11635 = n11634 ^ n10202;
  assign n11632 = n11500 ^ n11474;
  assign n11636 = n11635 ^ n11632;
  assign n11639 = n10209 ^ n10178;
  assign n11640 = ~n11386 & n11639;
  assign n11641 = n11640 ^ n10209;
  assign n11637 = n11497 ^ x474;
  assign n11638 = n11637 ^ n11475;
  assign n11642 = n11641 ^ n11638;
  assign n11644 = n10217 ^ n10185;
  assign n11645 = n11302 & ~n11644;
  assign n11646 = n11645 ^ n10217;
  assign n11643 = n11494 ^ n11478;
  assign n11647 = n11646 ^ n11643;
  assign n11650 = n10224 ^ n10192;
  assign n11651 = ~n11014 & n11650;
  assign n11652 = n11651 ^ n10224;
  assign n11648 = n11491 ^ x476;
  assign n11649 = n11648 ^ n11479;
  assign n11653 = n11652 ^ n11649;
  assign n11655 = n10198 ^ n10153;
  assign n11656 = ~n11019 & ~n11655;
  assign n11657 = n11656 ^ n10153;
  assign n11654 = n11488 ^ n11482;
  assign n11658 = n11657 ^ n11654;
  assign n11662 = n11485 ^ n11484;
  assign n11659 = n10200 ^ n10041;
  assign n11660 = ~n11024 & ~n11659;
  assign n11661 = n11660 ^ n10041;
  assign n11663 = n11662 ^ n11661;
  assign n11664 = n10208 ^ n9960;
  assign n11665 = n11030 & n11664;
  assign n11666 = n11665 ^ n9960;
  assign n11668 = n11667 ^ n11666;
  assign n11928 = n10215 ^ n9334;
  assign n11929 = n11035 & ~n11928;
  assign n11930 = n11929 ^ n9334;
  assign n11698 = n10256 ^ n9567;
  assign n11699 = ~n11066 & n11698;
  assign n11700 = n11699 ^ n9567;
  assign n11701 = n11700 ^ n11586;
  assign n11702 = n10263 ^ n9379;
  assign n11703 = n11078 & n11702;
  assign n11704 = n11703 ^ n9379;
  assign n11705 = n11704 ^ n11602;
  assign n11720 = n11719 ^ n11609;
  assign n11721 = ~n11709 & ~n11720;
  assign n11722 = n11721 ^ n11708;
  assign n11723 = n11722 ^ n11602;
  assign n11724 = ~n11705 & n11723;
  assign n11725 = n11724 ^ n11704;
  assign n11726 = n11725 ^ n11594;
  assign n11727 = n10261 ^ n9377;
  assign n11728 = ~n11072 & n11727;
  assign n11729 = n11728 ^ n9377;
  assign n11730 = n11729 ^ n11594;
  assign n11731 = ~n11726 & n11730;
  assign n11732 = n11731 ^ n11729;
  assign n11733 = n11732 ^ n11586;
  assign n11734 = ~n11701 & ~n11733;
  assign n11735 = n11734 ^ n11700;
  assign n11694 = n10250 ^ n9374;
  assign n11695 = ~n11064 & ~n11694;
  assign n11696 = n11695 ^ n9374;
  assign n11697 = n11696 ^ n11580;
  assign n11781 = n11735 ^ n11697;
  assign n11782 = n11781 ^ n9246;
  assign n11783 = n11732 ^ n11700;
  assign n11784 = n11783 ^ n11586;
  assign n11785 = n11784 ^ n9212;
  assign n11786 = n11729 ^ n11726;
  assign n11787 = n11786 ^ n9167;
  assign n11788 = n11722 ^ n11705;
  assign n11789 = n11788 ^ n9139;
  assign n11800 = n11799 ^ n11790;
  assign n11801 = ~n11791 & ~n11800;
  assign n11802 = n11801 ^ n9037;
  assign n11803 = n11802 ^ n11788;
  assign n11804 = n11789 & ~n11803;
  assign n11805 = n11804 ^ n9139;
  assign n11806 = n11805 ^ n11786;
  assign n11807 = n11787 & n11806;
  assign n11808 = n11807 ^ n9167;
  assign n11809 = n11808 ^ n11784;
  assign n11810 = ~n11785 & n11809;
  assign n11811 = n11810 ^ n9212;
  assign n11812 = n11811 ^ n11781;
  assign n11813 = n11782 & ~n11812;
  assign n11814 = n11813 ^ n9246;
  assign n11736 = n11735 ^ n11580;
  assign n11737 = ~n11697 & n11736;
  assign n11738 = n11737 ^ n11696;
  assign n11690 = n9916 ^ n9150;
  assign n11691 = ~n11007 & n11690;
  assign n11692 = n11691 ^ n9150;
  assign n11778 = n11738 ^ n11692;
  assign n11779 = n11778 ^ n11572;
  assign n11780 = n11779 ^ n8594;
  assign n11832 = n11814 ^ n11780;
  assign n11833 = n11811 ^ n11782;
  assign n11834 = n11808 ^ n9212;
  assign n11835 = n11834 ^ n11784;
  assign n11840 = n11836 & n11839;
  assign n11841 = n11802 ^ n11789;
  assign n11842 = n11840 & n11841;
  assign n11843 = n11805 ^ n11787;
  assign n11844 = n11842 & n11843;
  assign n11845 = ~n11835 & ~n11844;
  assign n11846 = ~n11833 & ~n11845;
  assign n11847 = n11832 & ~n11846;
  assign n11815 = n11814 ^ n11779;
  assign n11816 = n11780 & ~n11815;
  assign n11817 = n11816 ^ n8594;
  assign n11693 = n11692 ^ n11572;
  assign n11739 = n11738 ^ n11572;
  assign n11740 = ~n11693 & n11739;
  assign n11741 = n11740 ^ n11692;
  assign n11686 = n9907 ^ n9144;
  assign n11687 = n11061 & ~n11686;
  assign n11688 = n11687 ^ n9144;
  assign n11775 = n11741 ^ n11688;
  assign n11776 = n11775 ^ n11566;
  assign n11777 = n11776 ^ n8591;
  assign n11848 = n11817 ^ n11777;
  assign n11849 = ~n11847 & n11848;
  assign n11818 = n11817 ^ n11776;
  assign n11819 = ~n11777 & n11818;
  assign n11820 = n11819 ^ n8591;
  assign n11689 = n11688 ^ n11566;
  assign n11742 = n11741 ^ n11566;
  assign n11743 = n11689 & n11742;
  assign n11744 = n11743 ^ n11688;
  assign n11682 = n9923 ^ n9180;
  assign n11683 = ~n10619 & ~n11682;
  assign n11684 = n11683 ^ n9180;
  assign n11772 = n11744 ^ n11684;
  assign n11773 = n11772 ^ n11558;
  assign n11774 = n11773 ^ n8583;
  assign n11850 = n11820 ^ n11774;
  assign n11851 = ~n11849 & ~n11850;
  assign n11821 = n11820 ^ n11773;
  assign n11822 = ~n11774 & n11821;
  assign n11823 = n11822 ^ n8583;
  assign n11685 = n11684 ^ n11558;
  assign n11745 = n11744 ^ n11558;
  assign n11746 = ~n11685 & n11745;
  assign n11747 = n11746 ^ n11684;
  assign n11678 = n9898 ^ n9228;
  assign n11679 = n10613 & n11678;
  assign n11680 = n11679 ^ n9228;
  assign n11769 = n11747 ^ n11680;
  assign n11770 = n11769 ^ n11005;
  assign n11771 = n11770 ^ n8578;
  assign n11852 = n11823 ^ n11771;
  assign n11853 = n11851 & ~n11852;
  assign n11824 = n11823 ^ n11770;
  assign n11825 = ~n11771 & ~n11824;
  assign n11826 = n11825 ^ n8578;
  assign n11752 = n9892 ^ n9268;
  assign n11753 = ~n10629 & n11752;
  assign n11754 = n11753 ^ n9268;
  assign n11681 = n11680 ^ n11005;
  assign n11748 = n11747 ^ n11005;
  assign n11749 = n11681 & n11748;
  assign n11750 = n11749 ^ n11680;
  assign n11751 = n11750 ^ n11677;
  assign n11767 = n11754 ^ n11751;
  assign n11768 = n11767 ^ n8572;
  assign n11854 = n11826 ^ n11768;
  assign n11855 = ~n11853 & n11854;
  assign n11827 = n11826 ^ n11767;
  assign n11828 = n11768 & ~n11827;
  assign n11829 = n11828 ^ n8572;
  assign n11830 = n11829 ^ n7910;
  assign n11759 = n9364 ^ n9286;
  assign n11760 = n10604 & n11759;
  assign n11761 = n11760 ^ n9286;
  assign n11755 = n11754 ^ n11677;
  assign n11756 = ~n11751 & n11755;
  assign n11757 = n11756 ^ n11754;
  assign n11758 = n11757 ^ n11676;
  assign n11766 = n11761 ^ n11758;
  assign n11831 = n11830 ^ n11766;
  assign n11863 = n11855 ^ n11831;
  assign n11864 = n11863 ^ x449;
  assign n11865 = n11854 ^ n11853;
  assign n11866 = n11865 ^ x450;
  assign n11867 = n11852 ^ n11851;
  assign n11868 = n11867 ^ x451;
  assign n11869 = n11850 ^ n11849;
  assign n11870 = n11869 ^ x452;
  assign n11871 = n11848 ^ n11847;
  assign n11872 = n11871 ^ x453;
  assign n11873 = n11846 ^ n11832;
  assign n11874 = n11873 ^ x454;
  assign n11875 = n11845 ^ n11833;
  assign n11876 = n11875 ^ x455;
  assign n11877 = n11844 ^ n11835;
  assign n11878 = n11877 ^ x456;
  assign n11879 = n11843 ^ n11842;
  assign n11880 = n11879 ^ x457;
  assign n11881 = n11841 ^ n11840;
  assign n11882 = n11881 ^ x458;
  assign n11893 = n11892 ^ n11883;
  assign n11894 = n11884 & ~n11893;
  assign n11895 = n11894 ^ x459;
  assign n11896 = n11895 ^ n11881;
  assign n11897 = n11882 & ~n11896;
  assign n11898 = n11897 ^ x458;
  assign n11899 = n11898 ^ n11879;
  assign n11900 = n11880 & ~n11899;
  assign n11901 = n11900 ^ x457;
  assign n11902 = n11901 ^ n11877;
  assign n11903 = ~n11878 & n11902;
  assign n11904 = n11903 ^ x456;
  assign n11905 = n11904 ^ n11875;
  assign n11906 = n11876 & ~n11905;
  assign n11907 = n11906 ^ x455;
  assign n11908 = n11907 ^ n11873;
  assign n11909 = n11874 & ~n11908;
  assign n11910 = n11909 ^ x454;
  assign n11911 = n11910 ^ n11871;
  assign n11912 = ~n11872 & n11911;
  assign n11913 = n11912 ^ x453;
  assign n11914 = n11913 ^ n11869;
  assign n11915 = ~n11870 & n11914;
  assign n11916 = n11915 ^ x452;
  assign n11917 = n11916 ^ n11867;
  assign n11918 = n11868 & ~n11917;
  assign n11919 = n11918 ^ x451;
  assign n11920 = n11919 ^ n11865;
  assign n11921 = ~n11866 & n11920;
  assign n11922 = n11921 ^ x450;
  assign n11923 = n11922 ^ n11863;
  assign n11924 = ~n11864 & n11923;
  assign n11925 = n11924 ^ x449;
  assign n11926 = n11925 ^ x448;
  assign n11858 = n11766 ^ n7910;
  assign n11859 = n11829 ^ n11766;
  assign n11860 = n11858 & n11859;
  assign n11861 = n11860 ^ n7910;
  assign n11856 = ~n11831 & ~n11855;
  assign n11762 = n11761 ^ n11676;
  assign n11763 = ~n11758 & ~n11762;
  assign n11764 = n11763 ^ n11761;
  assign n11670 = n9936 ^ n9327;
  assign n11671 = ~n10598 & n11670;
  assign n11672 = n11671 ^ n9327;
  assign n11669 = n11214 ^ n11200;
  assign n11673 = n11672 ^ n11669;
  assign n11674 = n11673 ^ n7903;
  assign n11765 = n11764 ^ n11674;
  assign n11857 = n11856 ^ n11765;
  assign n11862 = n11861 ^ n11857;
  assign n11927 = n11926 ^ n11862;
  assign n11931 = n11930 ^ n11927;
  assign n11938 = n11919 ^ x450;
  assign n11939 = n11938 ^ n11865;
  assign n11935 = n10232 ^ n9347;
  assign n11936 = n11046 & ~n11935;
  assign n11937 = n11936 ^ n9347;
  assign n11940 = n11939 ^ n11937;
  assign n11944 = n11916 ^ x451;
  assign n11945 = n11944 ^ n11867;
  assign n11941 = n10238 ^ n9350;
  assign n11942 = ~n11051 & n11941;
  assign n11943 = n11942 ^ n9350;
  assign n11946 = n11945 ^ n11943;
  assign n11947 = n11913 ^ x452;
  assign n11948 = n11947 ^ n11869;
  assign n11949 = n10645 ^ n9357;
  assign n11950 = ~n11053 & ~n11949;
  assign n11951 = n11950 ^ n9357;
  assign n11952 = ~n11948 & n11951;
  assign n11953 = n11952 ^ n11945;
  assign n11954 = ~n11946 & n11953;
  assign n11955 = n11954 ^ n11952;
  assign n11956 = n11955 ^ n11939;
  assign n11957 = n11940 & n11956;
  assign n11958 = n11957 ^ n11937;
  assign n11932 = n10223 ^ n9341;
  assign n11933 = n11038 & ~n11932;
  assign n11934 = n11933 ^ n9341;
  assign n11959 = n11958 ^ n11934;
  assign n11960 = n11922 ^ x449;
  assign n11961 = n11960 ^ n11863;
  assign n11962 = n11961 ^ n11958;
  assign n11963 = ~n11959 & ~n11962;
  assign n11964 = n11963 ^ n11934;
  assign n11965 = n11964 ^ n11927;
  assign n11966 = n11931 & n11965;
  assign n11967 = n11966 ^ n11930;
  assign n11968 = n11967 ^ n11667;
  assign n11969 = n11668 & ~n11968;
  assign n11970 = n11969 ^ n11666;
  assign n11971 = n11970 ^ n11662;
  assign n11972 = ~n11663 & n11971;
  assign n11973 = n11972 ^ n11661;
  assign n11974 = n11973 ^ n11654;
  assign n11975 = ~n11658 & ~n11974;
  assign n11976 = n11975 ^ n11657;
  assign n11977 = n11976 ^ n11649;
  assign n11978 = n11653 & ~n11977;
  assign n11979 = n11978 ^ n11652;
  assign n11980 = n11979 ^ n11643;
  assign n11981 = n11647 & ~n11980;
  assign n11982 = n11981 ^ n11646;
  assign n11983 = n11982 ^ n11638;
  assign n11984 = n11642 & ~n11983;
  assign n11985 = n11984 ^ n11641;
  assign n11986 = n11985 ^ n11632;
  assign n11987 = n11636 & n11986;
  assign n11988 = n11987 ^ n11635;
  assign n11989 = n11988 ^ n11627;
  assign n11990 = n11631 & n11989;
  assign n11991 = n11990 ^ n11630;
  assign n11992 = n11991 ^ n11621;
  assign n11993 = n11625 & ~n11992;
  assign n11994 = n11993 ^ n11624;
  assign n11995 = n11994 ^ n11614;
  assign n11996 = n11619 & ~n11995;
  assign n11997 = n11996 ^ n11618;
  assign n11998 = n11997 ^ n11607;
  assign n11999 = n11613 & ~n11998;
  assign n12000 = n11999 ^ n11612;
  assign n12001 = n12000 ^ n11601;
  assign n12002 = n11606 & ~n12001;
  assign n12003 = n12002 ^ n11605;
  assign n12004 = n12003 ^ n11598;
  assign n12005 = ~n11599 & ~n12004;
  assign n12006 = n12005 ^ n11597;
  assign n12007 = n12006 ^ n11591;
  assign n12008 = n11592 & n12007;
  assign n12009 = n12008 ^ n11589;
  assign n12010 = n12009 ^ n11584;
  assign n12011 = n11585 & ~n12010;
  assign n12012 = n12011 ^ n11583;
  assign n12013 = n12012 ^ n11577;
  assign n12014 = ~n11578 & n12013;
  assign n12015 = n12014 ^ n11575;
  assign n12016 = n12015 ^ n11570;
  assign n12017 = ~n11571 & ~n12016;
  assign n12018 = n12017 ^ n11569;
  assign n12019 = n12018 ^ n11563;
  assign n12020 = ~n11564 & n12019;
  assign n12021 = n12020 ^ n11561;
  assign n12022 = n12021 ^ n11556;
  assign n12023 = ~n11557 & ~n12022;
  assign n12024 = n12023 ^ n11010;
  assign n12159 = n12029 ^ n12024;
  assign n12160 = ~n12030 & ~n12159;
  assign n12161 = n12160 ^ n12027;
  assign n12167 = n12166 ^ n12161;
  assign n12168 = n12167 ^ n9150;
  assign n12031 = n12030 ^ n12024;
  assign n12032 = n12031 ^ n9374;
  assign n12033 = n12021 ^ n11557;
  assign n12034 = n12033 ^ n9567;
  assign n12035 = n12018 ^ n11564;
  assign n12036 = n12035 ^ n9377;
  assign n12037 = n12015 ^ n11571;
  assign n12038 = n12037 ^ n9379;
  assign n12039 = n12012 ^ n11575;
  assign n12040 = n12039 ^ n11577;
  assign n12041 = n12040 ^ n9384;
  assign n12042 = n12009 ^ n11583;
  assign n12043 = n12042 ^ n11584;
  assign n12044 = n12043 ^ n9390;
  assign n12045 = n12006 ^ n11589;
  assign n12046 = n12045 ^ n11591;
  assign n12047 = n12046 ^ n9395;
  assign n12048 = n12003 ^ n11597;
  assign n12049 = n12048 ^ n11598;
  assign n12050 = n12049 ^ n9401;
  assign n12051 = n12000 ^ n11606;
  assign n12052 = n12051 ^ n9402;
  assign n12053 = n11997 ^ n11613;
  assign n12054 = n12053 ^ n9404;
  assign n12055 = n11994 ^ n11619;
  assign n12056 = n12055 ^ n9409;
  assign n12057 = n11991 ^ n11625;
  assign n12058 = n12057 ^ n9411;
  assign n12059 = n11988 ^ n11631;
  assign n12060 = n12059 ^ n9416;
  assign n12061 = n11985 ^ n11636;
  assign n12062 = n12061 ^ n9422;
  assign n12063 = n11982 ^ n11642;
  assign n12064 = n12063 ^ n9430;
  assign n12065 = n11979 ^ n11647;
  assign n12066 = n12065 ^ n8782;
  assign n12067 = n11976 ^ n11653;
  assign n12068 = n12067 ^ n9336;
  assign n12069 = n11973 ^ n11658;
  assign n12070 = n12069 ^ n9343;
  assign n12071 = n11970 ^ n11663;
  assign n12072 = n12071 ^ n9352;
  assign n12073 = n11967 ^ n11668;
  assign n12074 = n12073 ^ n9359;
  assign n12075 = n11964 ^ n11931;
  assign n12076 = n12075 ^ n9452;
  assign n12077 = n11961 ^ n11959;
  assign n12078 = n12077 ^ n9366;
  assign n12079 = n11955 ^ n11937;
  assign n12080 = n12079 ^ n11939;
  assign n12081 = n12080 ^ n9461;
  assign n12082 = n11951 ^ n11948;
  assign n12083 = n9473 & ~n12082;
  assign n12084 = n12083 ^ n9467;
  assign n12085 = n11952 ^ n11943;
  assign n12086 = n12085 ^ n11945;
  assign n12087 = n12086 ^ n12083;
  assign n12088 = ~n12084 & ~n12087;
  assign n12089 = n12088 ^ n9467;
  assign n12090 = n12089 ^ n12080;
  assign n12091 = n12081 & n12090;
  assign n12092 = n12091 ^ n9461;
  assign n12093 = n12092 ^ n12077;
  assign n12094 = ~n12078 & ~n12093;
  assign n12095 = n12094 ^ n9366;
  assign n12096 = n12095 ^ n12075;
  assign n12097 = n12076 & n12096;
  assign n12098 = n12097 ^ n9452;
  assign n12099 = n12098 ^ n12073;
  assign n12100 = ~n12074 & n12099;
  assign n12101 = n12100 ^ n9359;
  assign n12102 = n12101 ^ n12071;
  assign n12103 = n12072 & ~n12102;
  assign n12104 = n12103 ^ n9352;
  assign n12105 = n12104 ^ n12069;
  assign n12106 = ~n12070 & ~n12105;
  assign n12107 = n12106 ^ n9343;
  assign n12108 = n12107 ^ n12067;
  assign n12109 = ~n12068 & n12108;
  assign n12110 = n12109 ^ n9336;
  assign n12111 = n12110 ^ n12065;
  assign n12112 = ~n12066 & n12111;
  assign n12113 = n12112 ^ n8782;
  assign n12114 = n12113 ^ n12063;
  assign n12115 = n12064 & n12114;
  assign n12116 = n12115 ^ n9430;
  assign n12117 = n12116 ^ n12061;
  assign n12118 = n12062 & ~n12117;
  assign n12119 = n12118 ^ n9422;
  assign n12120 = n12119 ^ n12059;
  assign n12121 = ~n12060 & n12120;
  assign n12122 = n12121 ^ n9416;
  assign n12123 = n12122 ^ n12057;
  assign n12124 = n12058 & ~n12123;
  assign n12125 = n12124 ^ n9411;
  assign n12126 = n12125 ^ n12055;
  assign n12127 = ~n12056 & ~n12126;
  assign n12128 = n12127 ^ n9409;
  assign n12129 = n12128 ^ n12053;
  assign n12130 = ~n12054 & n12129;
  assign n12131 = n12130 ^ n9404;
  assign n12132 = n12131 ^ n12051;
  assign n12133 = ~n12052 & n12132;
  assign n12134 = n12133 ^ n9402;
  assign n12135 = n12134 ^ n12049;
  assign n12136 = n12050 & ~n12135;
  assign n12137 = n12136 ^ n9401;
  assign n12138 = n12137 ^ n12046;
  assign n12139 = n12047 & ~n12138;
  assign n12140 = n12139 ^ n9395;
  assign n12141 = n12140 ^ n12043;
  assign n12142 = n12044 & n12141;
  assign n12143 = n12142 ^ n9390;
  assign n12144 = n12143 ^ n12040;
  assign n12145 = n12041 & n12144;
  assign n12146 = n12145 ^ n9384;
  assign n12147 = n12146 ^ n12037;
  assign n12148 = n12038 & ~n12147;
  assign n12149 = n12148 ^ n9379;
  assign n12150 = n12149 ^ n12035;
  assign n12151 = ~n12036 & n12150;
  assign n12152 = n12151 ^ n9377;
  assign n12153 = n12152 ^ n12033;
  assign n12154 = n12034 & n12153;
  assign n12155 = n12154 ^ n9567;
  assign n12156 = n12155 ^ n12031;
  assign n12157 = ~n12032 & n12156;
  assign n12158 = n12157 ^ n9374;
  assign n12169 = n12168 ^ n12158;
  assign n12170 = n12149 ^ n12036;
  assign n12171 = n12143 ^ n12041;
  assign n12172 = n12134 ^ n12050;
  assign n12173 = n12131 ^ n12052;
  assign n12174 = n12128 ^ n12054;
  assign n12175 = n12122 ^ n12058;
  assign n12176 = n12119 ^ n12060;
  assign n12177 = n12116 ^ n12062;
  assign n12178 = n12113 ^ n12064;
  assign n12179 = n12104 ^ n12070;
  assign n12180 = n12101 ^ n12072;
  assign n12181 = n12098 ^ n12074;
  assign n12182 = n12089 ^ n12081;
  assign n12183 = n12082 ^ n9473;
  assign n12184 = n12086 ^ n12084;
  assign n12185 = ~n12183 & ~n12184;
  assign n12186 = ~n12182 & n12185;
  assign n12187 = n12092 ^ n12078;
  assign n12188 = ~n12186 & n12187;
  assign n12189 = n12095 ^ n12076;
  assign n12190 = n12188 & n12189;
  assign n12191 = ~n12181 & ~n12190;
  assign n12192 = n12180 & n12191;
  assign n12193 = n12179 & ~n12192;
  assign n12194 = n12107 ^ n12068;
  assign n12195 = n12193 & ~n12194;
  assign n12196 = n12110 ^ n12066;
  assign n12197 = ~n12195 & n12196;
  assign n12198 = ~n12178 & n12197;
  assign n12199 = ~n12177 & ~n12198;
  assign n12200 = n12176 & n12199;
  assign n12201 = ~n12175 & n12200;
  assign n12202 = n12125 ^ n12056;
  assign n12203 = n12201 & n12202;
  assign n12204 = n12174 & ~n12203;
  assign n12205 = n12173 & n12204;
  assign n12206 = n12172 & ~n12205;
  assign n12207 = n12137 ^ n12047;
  assign n12208 = ~n12206 & ~n12207;
  assign n12209 = n12140 ^ n12044;
  assign n12210 = n12208 & ~n12209;
  assign n12211 = n12171 & n12210;
  assign n12212 = n12146 ^ n12038;
  assign n12213 = n12211 & ~n12212;
  assign n12214 = n12170 & n12213;
  assign n12215 = n12152 ^ n12034;
  assign n12216 = ~n12214 & n12215;
  assign n12217 = n12155 ^ n12032;
  assign n12218 = ~n12216 & ~n12217;
  assign n12360 = n12169 & ~n12218;
  assign n12354 = n11895 ^ x458;
  assign n12355 = n12354 ^ n11881;
  assign n12351 = n10613 ^ n9907;
  assign n12352 = n11669 & n12351;
  assign n12353 = n12352 ^ n9907;
  assign n12356 = n12355 ^ n12353;
  assign n12348 = n12165 ^ n12161;
  assign n12349 = n12166 & n12348;
  assign n12350 = n12349 ^ n12164;
  assign n12357 = n12356 ^ n12350;
  assign n12358 = n12357 ^ n9144;
  assign n12345 = n12167 ^ n12158;
  assign n12346 = ~n12168 & n12345;
  assign n12347 = n12346 ^ n9150;
  assign n12359 = n12358 ^ n12347;
  assign n12361 = n12360 ^ n12359;
  assign n12362 = n12361 ^ x485;
  assign n12219 = n12218 ^ n12169;
  assign n12220 = n12219 ^ x486;
  assign n12221 = n12217 ^ n12216;
  assign n12222 = n12221 ^ x487;
  assign n12223 = n12215 ^ n12214;
  assign n12224 = n12223 ^ x488;
  assign n12225 = n12213 ^ n12170;
  assign n12226 = n12225 ^ x489;
  assign n12227 = n12212 ^ n12211;
  assign n12228 = n12227 ^ x490;
  assign n12229 = n12210 ^ n12171;
  assign n12230 = n12229 ^ x491;
  assign n12231 = n12209 ^ n12208;
  assign n12232 = n12231 ^ x492;
  assign n12233 = n12207 ^ n12206;
  assign n12234 = n12233 ^ x493;
  assign n12235 = n12205 ^ n12172;
  assign n12236 = n12235 ^ x494;
  assign n12238 = n12203 ^ n12174;
  assign n12239 = n12238 ^ x496;
  assign n12240 = n12202 ^ n12201;
  assign n12241 = n12240 ^ x497;
  assign n12242 = n12200 ^ n12175;
  assign n12243 = n12242 ^ x498;
  assign n12244 = n12199 ^ n12176;
  assign n12245 = n12244 ^ x499;
  assign n12246 = n12198 ^ n12177;
  assign n12247 = n12246 ^ x500;
  assign n12248 = n12197 ^ n12178;
  assign n12249 = n12248 ^ x501;
  assign n12250 = n12196 ^ n12195;
  assign n12251 = n12250 ^ x502;
  assign n12252 = n12194 ^ n12193;
  assign n12253 = n12252 ^ x503;
  assign n12254 = n12192 ^ n12179;
  assign n12255 = n12254 ^ x504;
  assign n12256 = n12191 ^ n12180;
  assign n12257 = n12256 ^ x505;
  assign n12258 = n12190 ^ n12181;
  assign n12259 = n12258 ^ x506;
  assign n12260 = n12189 ^ n12188;
  assign n12261 = n12260 ^ x507;
  assign n12262 = n12187 ^ n12186;
  assign n12263 = n12262 ^ x508;
  assign n12264 = n12185 ^ n12182;
  assign n12265 = n12264 ^ x509;
  assign n12266 = x511 & n12183;
  assign n12267 = n12266 ^ x510;
  assign n12268 = n12184 ^ n12183;
  assign n12269 = n12268 ^ n12266;
  assign n12270 = n12267 & ~n12269;
  assign n12271 = n12270 ^ x510;
  assign n12272 = n12271 ^ n12264;
  assign n12273 = ~n12265 & n12272;
  assign n12274 = n12273 ^ x509;
  assign n12275 = n12274 ^ n12262;
  assign n12276 = n12263 & ~n12275;
  assign n12277 = n12276 ^ x508;
  assign n12278 = n12277 ^ n12260;
  assign n12279 = ~n12261 & n12278;
  assign n12280 = n12279 ^ x507;
  assign n12281 = n12280 ^ n12258;
  assign n12282 = n12259 & ~n12281;
  assign n12283 = n12282 ^ x506;
  assign n12284 = n12283 ^ n12256;
  assign n12285 = n12257 & ~n12284;
  assign n12286 = n12285 ^ x505;
  assign n12287 = n12286 ^ n12254;
  assign n12288 = n12255 & ~n12287;
  assign n12289 = n12288 ^ x504;
  assign n12290 = n12289 ^ n12252;
  assign n12291 = n12253 & ~n12290;
  assign n12292 = n12291 ^ x503;
  assign n12293 = n12292 ^ n12250;
  assign n12294 = ~n12251 & n12293;
  assign n12295 = n12294 ^ x502;
  assign n12296 = n12295 ^ n12248;
  assign n12297 = ~n12249 & n12296;
  assign n12298 = n12297 ^ x501;
  assign n12299 = n12298 ^ n12246;
  assign n12300 = ~n12247 & n12299;
  assign n12301 = n12300 ^ x500;
  assign n12302 = n12301 ^ n12244;
  assign n12303 = ~n12245 & n12302;
  assign n12304 = n12303 ^ x499;
  assign n12305 = n12304 ^ n12242;
  assign n12306 = n12243 & ~n12305;
  assign n12307 = n12306 ^ x498;
  assign n12308 = n12307 ^ n12240;
  assign n12309 = ~n12241 & n12308;
  assign n12310 = n12309 ^ x497;
  assign n12311 = n12310 ^ n12238;
  assign n12312 = ~n12239 & n12311;
  assign n12313 = n12312 ^ x496;
  assign n12237 = n12204 ^ n12173;
  assign n12314 = n12313 ^ n12237;
  assign n12315 = n12237 ^ x495;
  assign n12316 = ~n12314 & n12315;
  assign n12317 = n12316 ^ x495;
  assign n12318 = n12317 ^ n12235;
  assign n12319 = n12236 & ~n12318;
  assign n12320 = n12319 ^ x494;
  assign n12321 = n12320 ^ n12233;
  assign n12322 = n12234 & ~n12321;
  assign n12323 = n12322 ^ x493;
  assign n12324 = n12323 ^ n12231;
  assign n12325 = ~n12232 & n12324;
  assign n12326 = n12325 ^ x492;
  assign n12327 = n12326 ^ n12229;
  assign n12328 = n12230 & ~n12327;
  assign n12329 = n12328 ^ x491;
  assign n12330 = n12329 ^ n12227;
  assign n12331 = ~n12228 & n12330;
  assign n12332 = n12331 ^ x490;
  assign n12333 = n12332 ^ n12225;
  assign n12334 = n12226 & ~n12333;
  assign n12335 = n12334 ^ x489;
  assign n12336 = n12335 ^ n12223;
  assign n12337 = n12224 & ~n12336;
  assign n12338 = n12337 ^ x488;
  assign n12339 = n12338 ^ n12221;
  assign n12340 = n12222 & ~n12339;
  assign n12341 = n12340 ^ x487;
  assign n12342 = n12341 ^ n12219;
  assign n12343 = n12220 & ~n12342;
  assign n12344 = n12343 ^ x486;
  assign n12592 = n12361 ^ n12344;
  assign n12593 = n12362 & ~n12592;
  assign n12594 = n12593 ^ x485;
  assign n12630 = n12594 ^ x484;
  assign n12561 = ~n12359 & ~n12360;
  assign n12553 = n12357 ^ n12347;
  assign n12554 = ~n12358 & ~n12553;
  assign n12555 = n12554 ^ n9144;
  assign n12525 = n12355 ^ n12350;
  assign n12526 = n12356 & ~n12525;
  assign n12527 = n12526 ^ n12353;
  assign n12521 = n10629 ^ n9923;
  assign n12522 = ~n11255 & ~n12521;
  assign n12523 = n12522 ^ n9923;
  assign n12412 = n11898 ^ n11880;
  assign n12524 = n12523 ^ n12412;
  assign n12551 = n12527 ^ n12524;
  assign n12552 = n12551 ^ n9180;
  assign n12560 = n12555 ^ n12552;
  assign n12590 = n12561 ^ n12560;
  assign n12631 = n12630 ^ n12590;
  assign n12798 = n12634 ^ n12631;
  assign n12907 = n12798 ^ n9357;
  assign n13006 = n2358 & ~n12907;
  assign n13007 = n13006 ^ n3242;
  assign n12635 = ~n12631 & ~n12634;
  assign n12626 = n11038 ^ n10238;
  assign n12627 = n11662 & n12626;
  assign n12628 = n12627 ^ n10238;
  assign n12801 = n12635 ^ n12628;
  assign n12591 = n12590 ^ x484;
  assign n12595 = n12594 ^ n12590;
  assign n12596 = ~n12591 & n12595;
  assign n12597 = n12596 ^ x484;
  assign n12562 = ~n12560 & ~n12561;
  assign n12556 = n12555 ^ n12551;
  assign n12557 = ~n12552 & n12556;
  assign n12558 = n12557 ^ n9180;
  assign n12528 = n12527 ^ n12412;
  assign n12529 = n12524 & ~n12528;
  assign n12530 = n12529 ^ n12523;
  assign n12517 = n10604 ^ n9898;
  assign n12518 = n11246 & n12517;
  assign n12519 = n12518 ^ n9898;
  assign n12405 = n11901 ^ x456;
  assign n12406 = n12405 ^ n11877;
  assign n12520 = n12519 ^ n12406;
  assign n12549 = n12530 ^ n12520;
  assign n12550 = n12549 ^ n9228;
  assign n12559 = n12558 ^ n12550;
  assign n12588 = n12562 ^ n12559;
  assign n12589 = n12588 ^ x483;
  assign n12625 = n12597 ^ n12589;
  assign n12802 = n12801 ^ n12625;
  assign n12799 = n9357 & n12798;
  assign n12800 = n12799 ^ n9350;
  assign n12908 = n12802 ^ n12800;
  assign n13008 = n12908 ^ n12907;
  assign n13009 = n13008 ^ n13006;
  assign n13010 = n13007 & ~n13009;
  assign n13011 = n13010 ^ n3242;
  assign n12909 = n12907 & n12908;
  assign n12803 = n12802 ^ n12799;
  assign n12804 = n12800 & ~n12803;
  assign n12805 = n12804 ^ n9350;
  assign n12629 = n12628 ^ n12625;
  assign n12636 = n12635 ^ n12625;
  assign n12637 = ~n12629 & n12636;
  assign n12638 = n12637 ^ n12635;
  assign n12598 = n12597 ^ n12588;
  assign n12599 = n12589 & ~n12598;
  assign n12600 = n12599 ^ x483;
  assign n12622 = n12600 ^ x482;
  assign n12566 = n12558 ^ n12549;
  assign n12567 = ~n12550 & ~n12566;
  assign n12568 = n12567 ^ n9228;
  assign n12535 = n10598 ^ n9892;
  assign n12536 = n11262 & ~n12535;
  assign n12537 = n12536 ^ n9892;
  assign n12531 = n12530 ^ n12406;
  assign n12532 = ~n12520 & n12531;
  assign n12533 = n12532 ^ n12519;
  assign n12398 = n11904 ^ n11876;
  assign n12534 = n12533 ^ n12398;
  assign n12564 = n12537 ^ n12534;
  assign n12565 = n12564 ^ n9268;
  assign n12569 = n12568 ^ n12565;
  assign n12563 = ~n12559 & n12562;
  assign n12586 = n12569 ^ n12563;
  assign n12623 = n12622 ^ n12586;
  assign n12619 = n11035 ^ n10232;
  assign n12620 = ~n11654 & n12619;
  assign n12621 = n12620 ^ n10232;
  assign n12624 = n12623 ^ n12621;
  assign n12796 = n12638 ^ n12624;
  assign n12797 = n12796 ^ n9347;
  assign n12906 = n12805 ^ n12797;
  assign n13004 = n12909 ^ n12906;
  assign n13005 = n13004 ^ n541;
  assign n13197 = n13011 ^ n13005;
  assign n12471 = n12286 ^ x504;
  assign n12472 = n12471 ^ n12254;
  assign n13194 = n11614 ^ n11302;
  assign n13195 = n12472 & n13194;
  assign n13196 = n13195 ^ n11302;
  assign n13198 = n13197 ^ n13196;
  assign n13203 = n12907 ^ n2358;
  assign n12479 = n12280 ^ x506;
  assign n12480 = n12479 ^ n12258;
  assign n13200 = n11627 ^ n11019;
  assign n13201 = n12480 & ~n13200;
  assign n13202 = n13201 ^ n11019;
  assign n13204 = n13203 ^ n13202;
  assign n12488 = n12277 ^ n12261;
  assign n13205 = n11632 ^ n11024;
  assign n13206 = ~n12488 & n13205;
  assign n13207 = n13206 ^ n11024;
  assign n12379 = n11262 ^ n10629;
  assign n12380 = ~n11948 & ~n12379;
  assign n12381 = n12380 ^ n10629;
  assign n12378 = n12332 ^ n12226;
  assign n12382 = n12381 ^ n12378;
  assign n12385 = n11910 ^ n11872;
  assign n12386 = n11246 ^ n10613;
  assign n12387 = ~n12385 & n12386;
  assign n12388 = n12387 ^ n10613;
  assign n12383 = n12329 ^ x490;
  assign n12384 = n12383 ^ n12227;
  assign n12389 = n12388 ^ n12384;
  assign n12395 = n12326 ^ x491;
  assign n12396 = n12395 ^ n12229;
  assign n12390 = n11907 ^ x454;
  assign n12391 = n12390 ^ n11873;
  assign n12392 = n11255 ^ n10619;
  assign n12393 = n12391 & n12392;
  assign n12394 = n12393 ^ n10619;
  assign n12397 = n12396 ^ n12394;
  assign n12402 = n12323 ^ x492;
  assign n12403 = n12402 ^ n12231;
  assign n12399 = n11669 ^ n11061;
  assign n12400 = n12398 & n12399;
  assign n12401 = n12400 ^ n11061;
  assign n12404 = n12403 ^ n12401;
  assign n12410 = n12320 ^ n12234;
  assign n12407 = n11676 ^ n11007;
  assign n12408 = ~n12406 & ~n12407;
  assign n12409 = n12408 ^ n11007;
  assign n12411 = n12410 ^ n12409;
  assign n12416 = n12317 ^ x494;
  assign n12417 = n12416 ^ n12235;
  assign n12413 = n11677 ^ n11064;
  assign n12414 = n12412 & ~n12413;
  assign n12415 = n12414 ^ n11064;
  assign n12418 = n12417 ^ n12415;
  assign n12422 = n12314 ^ x495;
  assign n12419 = n11066 ^ n11005;
  assign n12420 = n12355 & ~n12419;
  assign n12421 = n12420 ^ n11066;
  assign n12423 = n12422 ^ n12421;
  assign n12427 = n12310 ^ x496;
  assign n12428 = n12427 ^ n12238;
  assign n12424 = n11558 ^ n11072;
  assign n12425 = n12165 & ~n12424;
  assign n12426 = n12425 ^ n11072;
  assign n12429 = n12428 ^ n12426;
  assign n12433 = n12307 ^ n12241;
  assign n12430 = n11566 ^ n11078;
  assign n12431 = n12029 & ~n12430;
  assign n12432 = n12431 ^ n11078;
  assign n12434 = n12433 ^ n12432;
  assign n12438 = n12304 ^ x498;
  assign n12439 = n12438 ^ n12242;
  assign n12435 = n11572 ^ n11083;
  assign n12436 = ~n11556 & n12435;
  assign n12437 = n12436 ^ n11083;
  assign n12440 = n12439 ^ n12437;
  assign n12444 = n12301 ^ n12245;
  assign n12441 = n11580 ^ n11085;
  assign n12442 = n11563 & ~n12441;
  assign n12443 = n12442 ^ n11085;
  assign n12445 = n12444 ^ n12443;
  assign n12448 = n11586 ^ n10993;
  assign n12449 = n11570 & n12448;
  assign n12450 = n12449 ^ n10993;
  assign n12446 = n12298 ^ x500;
  assign n12447 = n12446 ^ n12246;
  assign n12451 = n12450 ^ n12447;
  assign n12455 = n12295 ^ n12249;
  assign n12452 = n11594 ^ n10869;
  assign n12453 = ~n11577 & ~n12452;
  assign n12454 = n12453 ^ n10869;
  assign n12456 = n12455 ^ n12454;
  assign n12460 = n12292 ^ n12251;
  assign n12457 = n11602 ^ n10806;
  assign n12458 = n11584 & ~n12457;
  assign n12459 = n12458 ^ n10806;
  assign n12461 = n12460 ^ n12459;
  assign n12465 = n12289 ^ x503;
  assign n12466 = n12465 ^ n12252;
  assign n12462 = n11609 ^ n10693;
  assign n12463 = n11591 & ~n12462;
  assign n12464 = n12463 ^ n10693;
  assign n12467 = n12466 ^ n12464;
  assign n12468 = n11615 ^ n10160;
  assign n12469 = n11598 & ~n12468;
  assign n12470 = n12469 ^ n10160;
  assign n12473 = n12472 ^ n12470;
  assign n12475 = n11548 ^ n10172;
  assign n12476 = n11601 & n12475;
  assign n12477 = n12476 ^ n10172;
  assign n12474 = n12283 ^ n12257;
  assign n12478 = n12477 ^ n12474;
  assign n12481 = n11447 ^ n10178;
  assign n12482 = n11607 & n12481;
  assign n12483 = n12482 ^ n10178;
  assign n12484 = n12483 ^ n12480;
  assign n12485 = n11432 ^ n10185;
  assign n12486 = n11614 & ~n12485;
  assign n12487 = n12486 ^ n10185;
  assign n12489 = n12488 ^ n12487;
  assign n12493 = n12274 ^ x508;
  assign n12494 = n12493 ^ n12262;
  assign n12490 = n11386 ^ n10192;
  assign n12491 = n11621 & ~n12490;
  assign n12492 = n12491 ^ n10192;
  assign n12495 = n12494 ^ n12492;
  assign n12499 = n12271 ^ x509;
  assign n12500 = n12499 ^ n12264;
  assign n12496 = n11302 ^ n10198;
  assign n12497 = n11627 & ~n12496;
  assign n12498 = n12497 ^ n10198;
  assign n12501 = n12500 ^ n12498;
  assign n12503 = n11014 ^ n10200;
  assign n12504 = ~n11632 & ~n12503;
  assign n12505 = n12504 ^ n10200;
  assign n12502 = n12268 ^ n12267;
  assign n12506 = n12505 ^ n12502;
  assign n12508 = n11019 ^ n10208;
  assign n12509 = n11638 & n12508;
  assign n12510 = n12509 ^ n10208;
  assign n12507 = n12183 ^ x511;
  assign n12511 = n12510 ^ n12507;
  assign n12609 = n11024 ^ n10215;
  assign n12610 = n11643 & ~n12609;
  assign n12611 = n12610 ^ n10215;
  assign n12572 = n12568 ^ n12564;
  assign n12573 = n12565 & ~n12572;
  assign n12574 = n12573 ^ n9268;
  assign n12575 = n12574 ^ n9286;
  assign n12542 = n10245 ^ n9364;
  assign n12543 = ~n11237 & ~n12542;
  assign n12544 = n12543 ^ n9364;
  assign n12538 = n12537 ^ n12398;
  assign n12539 = ~n12534 & n12538;
  assign n12540 = n12539 ^ n12537;
  assign n12541 = n12540 ^ n12391;
  assign n12571 = n12544 ^ n12541;
  assign n12576 = n12575 ^ n12571;
  assign n12570 = ~n12563 & n12569;
  assign n12584 = n12576 ^ n12570;
  assign n12585 = n12584 ^ x481;
  assign n12587 = n12586 ^ x482;
  assign n12601 = n12600 ^ n12586;
  assign n12602 = ~n12587 & n12601;
  assign n12603 = n12602 ^ x482;
  assign n12604 = n12603 ^ n12584;
  assign n12605 = ~n12585 & n12604;
  assign n12606 = n12605 ^ x481;
  assign n12607 = n12606 ^ x480;
  assign n12579 = n12571 ^ n9286;
  assign n12580 = n12574 ^ n12571;
  assign n12581 = n12579 & n12580;
  assign n12582 = n12581 ^ n9286;
  assign n12577 = ~n12570 & ~n12576;
  assign n12545 = n12544 ^ n12391;
  assign n12546 = ~n12541 & ~n12545;
  assign n12547 = n12546 ^ n12544;
  assign n12512 = n10243 ^ n9936;
  assign n12513 = n11231 & n12512;
  assign n12514 = n12513 ^ n9936;
  assign n12515 = n12514 ^ n12385;
  assign n12516 = n12515 ^ n9327;
  assign n12548 = n12547 ^ n12516;
  assign n12578 = n12577 ^ n12548;
  assign n12583 = n12582 ^ n12578;
  assign n12608 = n12607 ^ n12583;
  assign n12612 = n12611 ^ n12608;
  assign n12615 = n11030 ^ n10223;
  assign n12616 = n11649 & ~n12615;
  assign n12617 = n12616 ^ n10223;
  assign n12613 = n12603 ^ x481;
  assign n12614 = n12613 ^ n12584;
  assign n12618 = n12617 ^ n12614;
  assign n12639 = n12638 ^ n12623;
  assign n12640 = ~n12624 & n12639;
  assign n12641 = n12640 ^ n12621;
  assign n12642 = n12641 ^ n12614;
  assign n12643 = n12618 & n12642;
  assign n12644 = n12643 ^ n12617;
  assign n12645 = n12644 ^ n12608;
  assign n12646 = n12612 & n12645;
  assign n12647 = n12646 ^ n12611;
  assign n12648 = n12647 ^ n12507;
  assign n12649 = ~n12511 & ~n12648;
  assign n12650 = n12649 ^ n12510;
  assign n12651 = n12650 ^ n12502;
  assign n12652 = n12506 & n12651;
  assign n12653 = n12652 ^ n12505;
  assign n12654 = n12653 ^ n12500;
  assign n12655 = n12501 & n12654;
  assign n12656 = n12655 ^ n12498;
  assign n12657 = n12656 ^ n12494;
  assign n12658 = n12495 & n12657;
  assign n12659 = n12658 ^ n12492;
  assign n12660 = n12659 ^ n12488;
  assign n12661 = n12489 & n12660;
  assign n12662 = n12661 ^ n12487;
  assign n12663 = n12662 ^ n12480;
  assign n12664 = n12484 & n12663;
  assign n12665 = n12664 ^ n12483;
  assign n12666 = n12665 ^ n12474;
  assign n12667 = ~n12478 & ~n12666;
  assign n12668 = n12667 ^ n12477;
  assign n12669 = n12668 ^ n12472;
  assign n12670 = ~n12473 & n12669;
  assign n12671 = n12670 ^ n12470;
  assign n12672 = n12671 ^ n12466;
  assign n12673 = ~n12467 & n12672;
  assign n12674 = n12673 ^ n12464;
  assign n12675 = n12674 ^ n12460;
  assign n12676 = n12461 & ~n12675;
  assign n12677 = n12676 ^ n12459;
  assign n12678 = n12677 ^ n12455;
  assign n12679 = ~n12456 & ~n12678;
  assign n12680 = n12679 ^ n12454;
  assign n12681 = n12680 ^ n12447;
  assign n12682 = n12451 & n12681;
  assign n12683 = n12682 ^ n12450;
  assign n12684 = n12683 ^ n12444;
  assign n12685 = ~n12445 & ~n12684;
  assign n12686 = n12685 ^ n12443;
  assign n12687 = n12686 ^ n12439;
  assign n12688 = ~n12440 & ~n12687;
  assign n12689 = n12688 ^ n12437;
  assign n12690 = n12689 ^ n12433;
  assign n12691 = ~n12434 & ~n12690;
  assign n12692 = n12691 ^ n12432;
  assign n12693 = n12692 ^ n12428;
  assign n12694 = n12429 & n12693;
  assign n12695 = n12694 ^ n12426;
  assign n12696 = n12695 ^ n12422;
  assign n12697 = ~n12423 & n12696;
  assign n12698 = n12697 ^ n12421;
  assign n12699 = n12698 ^ n12417;
  assign n12700 = ~n12418 & n12699;
  assign n12701 = n12700 ^ n12415;
  assign n12702 = n12701 ^ n12410;
  assign n12703 = ~n12411 & n12702;
  assign n12704 = n12703 ^ n12409;
  assign n12705 = n12704 ^ n12403;
  assign n12706 = ~n12404 & ~n12705;
  assign n12707 = n12706 ^ n12401;
  assign n12708 = n12707 ^ n12396;
  assign n12709 = ~n12397 & ~n12708;
  assign n12710 = n12709 ^ n12394;
  assign n12711 = n12710 ^ n12384;
  assign n12712 = ~n12389 & ~n12711;
  assign n12713 = n12712 ^ n12388;
  assign n12714 = n12713 ^ n12378;
  assign n12715 = ~n12382 & ~n12714;
  assign n12716 = n12715 ^ n12381;
  assign n12374 = n11237 ^ n10604;
  assign n12375 = n11945 & ~n12374;
  assign n12376 = n12375 ^ n10604;
  assign n12738 = n12716 ^ n12376;
  assign n12372 = n12335 ^ x488;
  assign n12373 = n12372 ^ n12223;
  assign n12739 = n12738 ^ n12373;
  assign n12740 = n12739 ^ n9898;
  assign n12741 = n12713 ^ n12381;
  assign n12742 = n12741 ^ n12378;
  assign n12743 = n12742 ^ n9923;
  assign n12744 = n12710 ^ n12388;
  assign n12745 = n12744 ^ n12384;
  assign n12746 = n12745 ^ n9907;
  assign n12747 = n12707 ^ n12397;
  assign n12748 = n12747 ^ n9916;
  assign n12749 = n12704 ^ n12404;
  assign n12750 = n12749 ^ n10250;
  assign n12751 = n12701 ^ n12411;
  assign n12752 = n12751 ^ n10256;
  assign n12753 = n12698 ^ n12418;
  assign n12754 = n12753 ^ n10261;
  assign n12755 = n12695 ^ n12423;
  assign n12756 = n12755 ^ n10263;
  assign n12757 = n12692 ^ n12429;
  assign n12758 = n12757 ^ n10271;
  assign n12759 = n12689 ^ n12434;
  assign n12760 = n12759 ^ n10277;
  assign n12761 = n12686 ^ n12440;
  assign n12762 = n12761 ^ n10283;
  assign n12763 = n12683 ^ n12443;
  assign n12764 = n12763 ^ n12444;
  assign n12765 = n12764 ^ n10162;
  assign n12766 = n12680 ^ n12450;
  assign n12767 = n12766 ^ n12447;
  assign n12768 = n12767 ^ n10167;
  assign n12769 = n12677 ^ n12454;
  assign n12770 = n12769 ^ n12455;
  assign n12771 = n12770 ^ n10174;
  assign n12772 = n12674 ^ n12461;
  assign n12773 = n12772 ^ n10180;
  assign n12774 = n12671 ^ n12467;
  assign n12775 = n12774 ^ n10188;
  assign n12776 = n12668 ^ n12473;
  assign n12777 = n12776 ^ n10194;
  assign n12778 = n12665 ^ n12478;
  assign n12779 = n12778 ^ n10202;
  assign n12780 = n12662 ^ n12484;
  assign n12781 = n12780 ^ n10209;
  assign n12782 = n12659 ^ n12489;
  assign n12783 = n12782 ^ n10217;
  assign n12784 = n12656 ^ n12495;
  assign n12785 = n12784 ^ n10224;
  assign n12786 = n12653 ^ n12501;
  assign n12787 = n12786 ^ n10153;
  assign n12788 = n12650 ^ n12506;
  assign n12789 = n12788 ^ n10041;
  assign n12790 = n12647 ^ n12511;
  assign n12791 = n12790 ^ n9960;
  assign n12792 = n12644 ^ n12612;
  assign n12793 = n12792 ^ n9334;
  assign n12794 = n12641 ^ n12618;
  assign n12795 = n12794 ^ n9341;
  assign n12806 = n12805 ^ n12796;
  assign n12807 = n12797 & n12806;
  assign n12808 = n12807 ^ n9347;
  assign n12809 = n12808 ^ n12794;
  assign n12810 = n12795 & n12809;
  assign n12811 = n12810 ^ n9341;
  assign n12812 = n12811 ^ n12792;
  assign n12813 = n12793 & n12812;
  assign n12814 = n12813 ^ n9334;
  assign n12815 = n12814 ^ n12790;
  assign n12816 = n12791 & ~n12815;
  assign n12817 = n12816 ^ n9960;
  assign n12818 = n12817 ^ n12788;
  assign n12819 = n12789 & ~n12818;
  assign n12820 = n12819 ^ n10041;
  assign n12821 = n12820 ^ n12786;
  assign n12822 = n12787 & n12821;
  assign n12823 = n12822 ^ n10153;
  assign n12824 = n12823 ^ n12784;
  assign n12825 = ~n12785 & n12824;
  assign n12826 = n12825 ^ n10224;
  assign n12827 = n12826 ^ n12782;
  assign n12828 = n12783 & ~n12827;
  assign n12829 = n12828 ^ n10217;
  assign n12830 = n12829 ^ n12780;
  assign n12831 = ~n12781 & n12830;
  assign n12832 = n12831 ^ n10209;
  assign n12833 = n12832 ^ n12778;
  assign n12834 = n12779 & n12833;
  assign n12835 = n12834 ^ n10202;
  assign n12836 = n12835 ^ n12776;
  assign n12837 = n12777 & n12836;
  assign n12838 = n12837 ^ n10194;
  assign n12839 = n12838 ^ n12774;
  assign n12840 = n12775 & ~n12839;
  assign n12841 = n12840 ^ n10188;
  assign n12842 = n12841 ^ n12772;
  assign n12843 = ~n12773 & n12842;
  assign n12844 = n12843 ^ n10180;
  assign n12845 = n12844 ^ n12770;
  assign n12846 = n12771 & ~n12845;
  assign n12847 = n12846 ^ n10174;
  assign n12848 = n12847 ^ n12767;
  assign n12849 = n12768 & ~n12848;
  assign n12850 = n12849 ^ n10167;
  assign n12851 = n12850 ^ n12764;
  assign n12852 = ~n12765 & ~n12851;
  assign n12853 = n12852 ^ n10162;
  assign n12854 = n12853 ^ n12761;
  assign n12855 = ~n12762 & ~n12854;
  assign n12856 = n12855 ^ n10283;
  assign n12857 = n12856 ^ n12759;
  assign n12858 = n12760 & ~n12857;
  assign n12859 = n12858 ^ n10277;
  assign n12860 = n12859 ^ n12757;
  assign n12861 = n12758 & ~n12860;
  assign n12862 = n12861 ^ n10271;
  assign n12863 = n12862 ^ n12755;
  assign n12864 = ~n12756 & ~n12863;
  assign n12865 = n12864 ^ n10263;
  assign n12866 = n12865 ^ n12753;
  assign n12867 = ~n12754 & n12866;
  assign n12868 = n12867 ^ n10261;
  assign n12869 = n12868 ^ n12751;
  assign n12870 = n12752 & n12869;
  assign n12871 = n12870 ^ n10256;
  assign n12872 = n12871 ^ n12749;
  assign n12873 = ~n12750 & ~n12872;
  assign n12874 = n12873 ^ n10250;
  assign n12875 = n12874 ^ n12747;
  assign n12876 = ~n12748 & ~n12875;
  assign n12877 = n12876 ^ n9916;
  assign n12878 = n12877 ^ n12745;
  assign n12879 = n12746 & ~n12878;
  assign n12880 = n12879 ^ n9907;
  assign n12881 = n12880 ^ n12742;
  assign n12882 = ~n12743 & n12881;
  assign n12883 = n12882 ^ n9923;
  assign n12884 = n12883 ^ n12739;
  assign n12885 = ~n12740 & n12884;
  assign n12886 = n12885 ^ n9898;
  assign n12721 = n11231 ^ n10598;
  assign n12722 = ~n11939 & ~n12721;
  assign n12723 = n12722 ^ n10598;
  assign n12377 = n12376 ^ n12373;
  assign n12717 = n12716 ^ n12373;
  assign n12718 = n12377 & n12717;
  assign n12719 = n12718 ^ n12376;
  assign n12371 = n12338 ^ n12222;
  assign n12720 = n12719 ^ n12371;
  assign n12736 = n12723 ^ n12720;
  assign n12737 = n12736 ^ n9892;
  assign n12949 = n12886 ^ n12737;
  assign n12892 = n12877 ^ n12746;
  assign n12893 = n12874 ^ n12748;
  assign n12894 = n12868 ^ n12752;
  assign n12895 = n12862 ^ n12756;
  assign n12896 = n12859 ^ n12758;
  assign n12897 = n12853 ^ n12762;
  assign n12898 = n12850 ^ n12765;
  assign n12899 = n12841 ^ n12773;
  assign n12900 = n12835 ^ n12777;
  assign n12901 = n12829 ^ n12781;
  assign n12902 = n12826 ^ n12783;
  assign n12903 = n12817 ^ n12789;
  assign n12904 = n12811 ^ n12793;
  assign n12905 = n12808 ^ n12795;
  assign n12910 = n12906 & n12909;
  assign n12911 = n12905 & ~n12910;
  assign n12912 = ~n12904 & n12911;
  assign n12913 = n12814 ^ n12791;
  assign n12914 = ~n12912 & ~n12913;
  assign n12915 = ~n12903 & n12914;
  assign n12916 = n12820 ^ n12787;
  assign n12917 = ~n12915 & n12916;
  assign n12918 = n12823 ^ n12785;
  assign n12919 = n12917 & n12918;
  assign n12920 = n12902 & ~n12919;
  assign n12921 = ~n12901 & n12920;
  assign n12922 = n12832 ^ n12779;
  assign n12923 = ~n12921 & ~n12922;
  assign n12924 = n12900 & n12923;
  assign n12925 = n12838 ^ n12775;
  assign n12926 = n12924 & ~n12925;
  assign n12927 = n12899 & n12926;
  assign n12928 = n12844 ^ n12771;
  assign n12929 = ~n12927 & n12928;
  assign n12930 = n12847 ^ n12768;
  assign n12931 = n12929 & n12930;
  assign n12932 = n12898 & ~n12931;
  assign n12933 = n12897 & ~n12932;
  assign n12934 = n12856 ^ n12760;
  assign n12935 = n12933 & n12934;
  assign n12936 = n12896 & n12935;
  assign n12937 = ~n12895 & n12936;
  assign n12938 = n12865 ^ n12754;
  assign n12939 = n12937 & n12938;
  assign n12940 = n12894 & ~n12939;
  assign n12941 = n12871 ^ n12750;
  assign n12942 = ~n12940 & ~n12941;
  assign n12943 = ~n12893 & ~n12942;
  assign n12944 = n12892 & ~n12943;
  assign n12945 = n12880 ^ n12743;
  assign n12946 = ~n12944 & n12945;
  assign n12947 = n12883 ^ n12740;
  assign n12948 = n12946 & n12947;
  assign n12959 = n12949 ^ n12948;
  assign n12960 = n12959 ^ n678;
  assign n12961 = n12947 ^ n12946;
  assign n12962 = n12961 ^ n1949;
  assign n12963 = n12945 ^ n12944;
  assign n12964 = n12963 ^ n1805;
  assign n12966 = n12942 ^ n12893;
  assign n12967 = n12966 ^ n1701;
  assign n12968 = n12941 ^ n12940;
  assign n12969 = n12968 ^ n1651;
  assign n12970 = n12939 ^ n12894;
  assign n12971 = n12970 ^ n1641;
  assign n12973 = n12936 ^ n12895;
  assign n12974 = n12973 ^ n2899;
  assign n12976 = n12934 ^ n12933;
  assign n12977 = n12976 ^ n1562;
  assign n12978 = n12932 ^ n12897;
  assign n12979 = n12978 ^ n2632;
  assign n12980 = n12931 ^ n12898;
  assign n12981 = n12980 ^ n1515;
  assign n12983 = n12928 ^ n12927;
  assign n2456 = x433 ^ x81;
  assign n2457 = n2456 ^ x273;
  assign n2458 = n2457 ^ x17;
  assign n12984 = n12983 ^ n2458;
  assign n12986 = n12925 ^ n12924;
  assign n12987 = n12986 ^ n1299;
  assign n12989 = n12922 ^ n12921;
  assign n1112 = x437 ^ x85;
  assign n1113 = n1112 ^ x277;
  assign n1114 = n1113 ^ x21;
  assign n12990 = n12989 ^ n1114;
  assign n12992 = n12919 ^ n12902;
  assign n12993 = n12992 ^ n973;
  assign n12995 = n12916 ^ n12915;
  assign n12996 = n12995 ^ n958;
  assign n12997 = n12914 ^ n12903;
  assign n12998 = n12997 ^ n608;
  assign n12999 = n12913 ^ n12912;
  assign n13000 = n12999 ^ n647;
  assign n13001 = n12911 ^ n12904;
  assign n13002 = n13001 ^ n567;
  assign n13012 = n13011 ^ n13004;
  assign n13013 = n13005 & ~n13012;
  assign n13014 = n13013 ^ n541;
  assign n13003 = n12910 ^ n12905;
  assign n13015 = n13014 ^ n13003;
  assign n13016 = n13003 ^ n547;
  assign n13017 = ~n13015 & n13016;
  assign n13018 = n13017 ^ n547;
  assign n13019 = n13018 ^ n13001;
  assign n13020 = n13002 & ~n13019;
  assign n13021 = n13020 ^ n567;
  assign n13022 = n13021 ^ n12999;
  assign n13023 = n13000 & ~n13022;
  assign n13024 = n13023 ^ n647;
  assign n13025 = n13024 ^ n12997;
  assign n13026 = ~n12998 & n13025;
  assign n13027 = n13026 ^ n608;
  assign n13028 = n13027 ^ n12995;
  assign n13029 = n12996 & ~n13028;
  assign n13030 = n13029 ^ n958;
  assign n12994 = n12918 ^ n12917;
  assign n13031 = n13030 ^ n12994;
  assign n13032 = n12994 ^ n791;
  assign n13033 = n13031 & ~n13032;
  assign n13034 = n13033 ^ n791;
  assign n13035 = n13034 ^ n12992;
  assign n13036 = ~n12993 & n13035;
  assign n13037 = n13036 ^ n973;
  assign n12991 = n12920 ^ n12901;
  assign n13038 = n13037 ^ n12991;
  assign n13039 = n12991 ^ n992;
  assign n13040 = n13038 & ~n13039;
  assign n13041 = n13040 ^ n992;
  assign n13042 = n13041 ^ n12989;
  assign n13043 = ~n12990 & n13042;
  assign n13044 = n13043 ^ n1114;
  assign n12988 = n12923 ^ n12900;
  assign n13045 = n13044 ^ n12988;
  assign n13046 = n12988 ^ n1287;
  assign n13047 = n13045 & ~n13046;
  assign n13048 = n13047 ^ n1287;
  assign n13049 = n13048 ^ n12986;
  assign n13050 = n12987 & ~n13049;
  assign n13051 = n13050 ^ n1299;
  assign n12985 = n12926 ^ n12899;
  assign n13052 = n13051 ^ n12985;
  assign n13053 = n12985 ^ n2477;
  assign n13054 = n13052 & ~n13053;
  assign n13055 = n13054 ^ n2477;
  assign n13056 = n13055 ^ n12983;
  assign n13057 = ~n12984 & n13056;
  assign n13058 = n13057 ^ n2458;
  assign n12982 = n12930 ^ n12929;
  assign n13059 = n13058 ^ n12982;
  assign n13060 = n12982 ^ n2464;
  assign n13061 = ~n13059 & n13060;
  assign n13062 = n13061 ^ n2464;
  assign n13063 = n13062 ^ n12980;
  assign n13064 = n12981 & ~n13063;
  assign n13065 = n13064 ^ n1515;
  assign n13066 = n13065 ^ n12978;
  assign n13067 = ~n12979 & n13066;
  assign n13068 = n13067 ^ n2632;
  assign n13069 = n13068 ^ n12976;
  assign n13070 = n12977 & ~n13069;
  assign n13071 = n13070 ^ n1562;
  assign n12975 = n12935 ^ n12896;
  assign n13072 = n13071 ^ n12975;
  assign n13073 = n12975 ^ n2744;
  assign n13074 = ~n13072 & n13073;
  assign n13075 = n13074 ^ n2744;
  assign n13076 = n13075 ^ n12973;
  assign n13077 = ~n12974 & n13076;
  assign n13078 = n13077 ^ n2899;
  assign n12972 = n12938 ^ n12937;
  assign n13079 = n13078 ^ n12972;
  assign n13080 = n12972 ^ n1635;
  assign n13081 = ~n13079 & n13080;
  assign n13082 = n13081 ^ n1635;
  assign n13083 = n13082 ^ n12970;
  assign n13084 = n12971 & ~n13083;
  assign n13085 = n13084 ^ n1641;
  assign n13086 = n13085 ^ n12968;
  assign n13087 = n12969 & ~n13086;
  assign n13088 = n13087 ^ n1651;
  assign n13089 = n13088 ^ n12966;
  assign n13090 = ~n12967 & n13089;
  assign n13091 = n13090 ^ n1701;
  assign n12965 = n12943 ^ n12892;
  assign n13092 = n13091 ^ n12965;
  assign n13093 = n12965 ^ n1808;
  assign n13094 = n13092 & ~n13093;
  assign n13095 = n13094 ^ n1808;
  assign n13096 = n13095 ^ n12963;
  assign n13097 = n12964 & ~n13096;
  assign n13098 = n13097 ^ n1805;
  assign n13099 = n13098 ^ n12961;
  assign n13100 = ~n12962 & n13099;
  assign n13101 = n13100 ^ n1949;
  assign n13102 = n13101 ^ n12959;
  assign n13103 = n12960 & ~n13102;
  assign n13104 = n13103 ^ n678;
  assign n12950 = ~n12948 & ~n12949;
  assign n12887 = n12886 ^ n12736;
  assign n12888 = ~n12737 & n12887;
  assign n12889 = n12888 ^ n9892;
  assign n12890 = n12889 ^ n9364;
  assign n12728 = n11053 ^ n10245;
  assign n12729 = ~n11961 & ~n12728;
  assign n12730 = n12729 ^ n10245;
  assign n12724 = n12723 ^ n12371;
  assign n12725 = ~n12720 & ~n12724;
  assign n12726 = n12725 ^ n12723;
  assign n12369 = n12341 ^ x486;
  assign n12370 = n12369 ^ n12219;
  assign n12727 = n12726 ^ n12370;
  assign n12735 = n12730 ^ n12727;
  assign n12891 = n12890 ^ n12735;
  assign n12958 = n12950 ^ n12891;
  assign n13105 = n13104 ^ n12958;
  assign n2127 = x418 ^ x66;
  assign n2128 = n2127 ^ x258;
  assign n2129 = n2128 ^ x2;
  assign n13106 = n12958 ^ n2129;
  assign n13107 = n13105 & ~n13106;
  assign n13108 = n13107 ^ n2129;
  assign n13109 = n13108 ^ n2342;
  assign n12953 = n12735 ^ n9364;
  assign n12954 = n12889 ^ n12735;
  assign n12955 = n12953 & n12954;
  assign n12956 = n12955 ^ n9364;
  assign n12951 = ~n12891 & ~n12950;
  assign n12731 = n12730 ^ n12370;
  assign n12732 = n12727 & n12731;
  assign n12733 = n12732 ^ n12730;
  assign n12364 = n11051 ^ n10243;
  assign n12365 = ~n11927 & ~n12364;
  assign n12366 = n12365 ^ n10243;
  assign n12363 = n12362 ^ n12344;
  assign n12367 = n12366 ^ n12363;
  assign n12368 = n12367 ^ n9936;
  assign n12734 = n12733 ^ n12368;
  assign n12952 = n12951 ^ n12734;
  assign n12957 = n12956 ^ n12952;
  assign n13110 = n13109 ^ n12957;
  assign n13208 = n13207 ^ n13110;
  assign n13210 = n11638 ^ n11030;
  assign n13211 = n12494 & n13210;
  assign n13212 = n13211 ^ n11030;
  assign n13209 = n13105 ^ n2129;
  assign n13213 = n13212 ^ n13209;
  assign n13227 = n11643 ^ n11035;
  assign n13228 = ~n12500 & n13227;
  assign n13229 = n13228 ^ n11035;
  assign n13215 = n11649 ^ n11038;
  assign n13216 = n12502 & n13215;
  assign n13217 = n13216 ^ n11038;
  assign n13214 = n13098 ^ n12962;
  assign n13218 = n13217 ^ n13214;
  assign n13219 = n13095 ^ n12964;
  assign n13220 = n11654 ^ n11046;
  assign n13221 = n12507 & ~n13220;
  assign n13222 = n13221 ^ n11046;
  assign n13223 = n13219 & n13222;
  assign n13224 = n13223 ^ n13214;
  assign n13225 = n13218 & ~n13224;
  assign n13226 = n13225 ^ n13223;
  assign n13230 = n13229 ^ n13226;
  assign n13231 = n13101 ^ n12960;
  assign n13232 = n13231 ^ n13226;
  assign n13233 = n13230 & ~n13232;
  assign n13234 = n13233 ^ n13229;
  assign n13235 = n13234 ^ n13209;
  assign n13236 = ~n13213 & n13235;
  assign n13237 = n13236 ^ n13212;
  assign n13238 = n13237 ^ n13110;
  assign n13239 = ~n13208 & ~n13238;
  assign n13240 = n13239 ^ n13207;
  assign n13241 = n13240 ^ n13203;
  assign n13242 = n13204 & ~n13241;
  assign n13243 = n13242 ^ n13202;
  assign n13199 = n13008 ^ n13007;
  assign n13244 = n13243 ^ n13199;
  assign n13245 = n11621 ^ n11014;
  assign n13246 = n12474 & ~n13245;
  assign n13247 = n13246 ^ n11014;
  assign n13248 = n13247 ^ n13199;
  assign n13249 = n13244 & ~n13248;
  assign n13250 = n13249 ^ n13247;
  assign n13251 = n13250 ^ n13197;
  assign n13252 = n13198 & n13251;
  assign n13253 = n13252 ^ n13196;
  assign n13189 = n11607 ^ n11386;
  assign n13190 = n12466 & ~n13189;
  assign n13191 = n13190 ^ n11386;
  assign n13354 = n13253 ^ n13191;
  assign n13192 = n13015 ^ n547;
  assign n13355 = n13354 ^ n13192;
  assign n13356 = n13355 ^ n10192;
  assign n13357 = n13250 ^ n13196;
  assign n13358 = n13357 ^ n13197;
  assign n13359 = n13358 ^ n10198;
  assign n13360 = n13247 ^ n13244;
  assign n13361 = n13360 ^ n10200;
  assign n13362 = n13240 ^ n13202;
  assign n13363 = n13362 ^ n13203;
  assign n13364 = n13363 ^ n10208;
  assign n13365 = n13237 ^ n13207;
  assign n13366 = n13365 ^ n13110;
  assign n13367 = n13366 ^ n10215;
  assign n13368 = n13234 ^ n13213;
  assign n13369 = n13368 ^ n10223;
  assign n13370 = n13231 ^ n13229;
  assign n13371 = n13370 ^ n13226;
  assign n13372 = n13371 ^ n10232;
  assign n13373 = n13222 ^ n13219;
  assign n13374 = ~n10645 & n13373;
  assign n13375 = n13374 ^ n10238;
  assign n13376 = n13223 ^ n13217;
  assign n13377 = n13376 ^ n13214;
  assign n13378 = n13377 ^ n13374;
  assign n13379 = n13375 & n13378;
  assign n13380 = n13379 ^ n10238;
  assign n13381 = n13380 ^ n13371;
  assign n13382 = n13372 & ~n13381;
  assign n13383 = n13382 ^ n10232;
  assign n13384 = n13383 ^ n13368;
  assign n13385 = n13369 & n13384;
  assign n13386 = n13385 ^ n10223;
  assign n13387 = n13386 ^ n13366;
  assign n13388 = ~n13367 & ~n13387;
  assign n13389 = n13388 ^ n10215;
  assign n13390 = n13389 ^ n13363;
  assign n13391 = n13364 & n13390;
  assign n13392 = n13391 ^ n10208;
  assign n13393 = n13392 ^ n13360;
  assign n13394 = n13361 & n13393;
  assign n13395 = n13394 ^ n10200;
  assign n13396 = n13395 ^ n13358;
  assign n13397 = n13359 & n13396;
  assign n13398 = n13397 ^ n10198;
  assign n13399 = n13398 ^ n13355;
  assign n13400 = ~n13356 & ~n13399;
  assign n13401 = n13400 ^ n10192;
  assign n13193 = n13192 ^ n13191;
  assign n13254 = n13253 ^ n13192;
  assign n13255 = ~n13193 & ~n13254;
  assign n13256 = n13255 ^ n13191;
  assign n13185 = n11601 ^ n11432;
  assign n13186 = ~n12460 & n13185;
  assign n13187 = n13186 ^ n11432;
  assign n13351 = n13256 ^ n13187;
  assign n13184 = n13018 ^ n13002;
  assign n13352 = n13351 ^ n13184;
  assign n13353 = n13352 ^ n10185;
  assign n13477 = n13401 ^ n13353;
  assign n13478 = n13389 ^ n13364;
  assign n13479 = n13386 ^ n13367;
  assign n13480 = n13380 ^ n13372;
  assign n13481 = n13373 ^ n10645;
  assign n13482 = n13377 ^ n13375;
  assign n13483 = ~n13481 & ~n13482;
  assign n13484 = n13480 & n13483;
  assign n13485 = n13383 ^ n13369;
  assign n13486 = ~n13484 & ~n13485;
  assign n13487 = ~n13479 & n13486;
  assign n13488 = n13478 & ~n13487;
  assign n13489 = n13392 ^ n13361;
  assign n13490 = n13488 & ~n13489;
  assign n13491 = n13395 ^ n13359;
  assign n13492 = ~n13490 & ~n13491;
  assign n13493 = n13398 ^ n13356;
  assign n13494 = n13492 & ~n13493;
  assign n13495 = n13477 & ~n13494;
  assign n13402 = n13401 ^ n13352;
  assign n13403 = n13353 & n13402;
  assign n13404 = n13403 ^ n10185;
  assign n13188 = n13187 ^ n13184;
  assign n13257 = n13256 ^ n13184;
  assign n13258 = n13188 & n13257;
  assign n13259 = n13258 ^ n13187;
  assign n13180 = n11598 ^ n11447;
  assign n13181 = ~n12455 & n13180;
  assign n13182 = n13181 ^ n11447;
  assign n13348 = n13259 ^ n13182;
  assign n13179 = n13021 ^ n13000;
  assign n13349 = n13348 ^ n13179;
  assign n13350 = n13349 ^ n10178;
  assign n13496 = n13404 ^ n13350;
  assign n13497 = n13495 & ~n13496;
  assign n13265 = n11591 ^ n11548;
  assign n13266 = ~n12447 & ~n13265;
  assign n13267 = n13266 ^ n11548;
  assign n13263 = n13024 ^ n12998;
  assign n13409 = n13267 ^ n13263;
  assign n13183 = n13182 ^ n13179;
  assign n13260 = n13259 ^ n13179;
  assign n13261 = n13183 & ~n13260;
  assign n13262 = n13261 ^ n13182;
  assign n13410 = n13409 ^ n13262;
  assign n13475 = n13410 ^ n10172;
  assign n13405 = n13404 ^ n13349;
  assign n13406 = n13350 & n13405;
  assign n13407 = n13406 ^ n10178;
  assign n13476 = n13475 ^ n13407;
  assign n13544 = n13497 ^ n13476;
  assign n1234 = x469 ^ x117;
  assign n1235 = n1234 ^ x309;
  assign n1236 = n1235 ^ x53;
  assign n13545 = n13544 ^ n1236;
  assign n13547 = n13494 ^ n13477;
  assign n13548 = n13547 ^ n862;
  assign n13550 = n13491 ^ n13490;
  assign n13551 = n13550 ^ n755;
  assign n13552 = n13489 ^ n13488;
  assign n13553 = n13552 ^ n658;
  assign n13554 = n13487 ^ n13478;
  assign n13555 = n13554 ^ n599;
  assign n13556 = n13486 ^ n13479;
  assign n13557 = n13556 ^ n593;
  assign n13559 = n13483 ^ n13480;
  assign n13563 = n13562 ^ n13559;
  assign n13567 = n13481 & n13566;
  assign n13568 = n13567 ^ n672;
  assign n13569 = n13482 ^ n13481;
  assign n13570 = n13569 ^ n13567;
  assign n13571 = n13568 & ~n13570;
  assign n13572 = n13571 ^ n672;
  assign n13573 = n13572 ^ n13559;
  assign n13574 = n13563 & ~n13573;
  assign n13575 = n13574 ^ n13562;
  assign n13558 = n13485 ^ n13484;
  assign n13576 = n13575 ^ n13558;
  assign n13577 = n13558 ^ n3252;
  assign n13578 = n13576 & ~n13577;
  assign n13579 = n13578 ^ n3252;
  assign n13580 = n13579 ^ n13556;
  assign n13581 = n13557 & ~n13580;
  assign n13582 = n13581 ^ n593;
  assign n13583 = n13582 ^ n13554;
  assign n13584 = ~n13555 & n13583;
  assign n13585 = n13584 ^ n599;
  assign n13586 = n13585 ^ n13552;
  assign n13587 = ~n13553 & n13586;
  assign n13588 = n13587 ^ n658;
  assign n13589 = n13588 ^ n13550;
  assign n13590 = ~n13551 & n13589;
  assign n13591 = n13590 ^ n755;
  assign n13549 = n13493 ^ n13492;
  assign n13592 = n13591 ^ n13549;
  assign n13593 = n13549 ^ n856;
  assign n13594 = ~n13592 & n13593;
  assign n13595 = n13594 ^ n856;
  assign n13596 = n13595 ^ n13547;
  assign n13597 = ~n13548 & n13596;
  assign n13598 = n13597 ^ n862;
  assign n13546 = n13496 ^ n13495;
  assign n13599 = n13598 ^ n13546;
  assign n997 = x470 ^ x118;
  assign n998 = n997 ^ x310;
  assign n999 = n998 ^ x54;
  assign n13600 = n13546 ^ n999;
  assign n13601 = n13599 & ~n13600;
  assign n13602 = n13601 ^ n999;
  assign n13603 = n13602 ^ n13544;
  assign n13604 = n13545 & ~n13603;
  assign n13605 = n13604 ^ n1236;
  assign n13408 = n13407 ^ n10172;
  assign n13411 = n13410 ^ n13407;
  assign n13412 = ~n13408 & ~n13411;
  assign n13413 = n13412 ^ n10172;
  assign n13264 = n13263 ^ n13262;
  assign n13268 = n13267 ^ n13262;
  assign n13269 = ~n13264 & n13268;
  assign n13270 = n13269 ^ n13263;
  assign n13175 = n11615 ^ n11584;
  assign n13176 = ~n12444 & n13175;
  assign n13177 = n13176 ^ n11615;
  assign n13345 = n13270 ^ n13177;
  assign n13174 = n13027 ^ n12996;
  assign n13346 = n13345 ^ n13174;
  assign n13347 = n13346 ^ n10160;
  assign n13499 = n13413 ^ n13347;
  assign n13498 = n13476 & ~n13497;
  assign n13543 = n13499 ^ n13498;
  assign n13606 = n13605 ^ n13543;
  assign n1170 = x468 ^ x116;
  assign n1171 = n1170 ^ x308;
  assign n1172 = n1171 ^ x52;
  assign n13607 = n13543 ^ n1172;
  assign n13608 = n13606 & ~n13607;
  assign n13609 = n13608 ^ n1172;
  assign n13414 = n13413 ^ n13346;
  assign n13415 = n13347 & ~n13414;
  assign n13416 = n13415 ^ n10160;
  assign n13178 = n13177 ^ n13174;
  assign n13271 = n13270 ^ n13174;
  assign n13272 = n13178 & n13271;
  assign n13273 = n13272 ^ n13177;
  assign n13170 = n11609 ^ n11577;
  assign n13171 = n12439 & ~n13170;
  assign n13172 = n13171 ^ n11609;
  assign n13169 = n13031 ^ n791;
  assign n13173 = n13172 ^ n13169;
  assign n13343 = n13273 ^ n13173;
  assign n13344 = n13343 ^ n10693;
  assign n13501 = n13416 ^ n13344;
  assign n13500 = n13498 & n13499;
  assign n13541 = n13501 ^ n13500;
  assign n1416 = x467 ^ x115;
  assign n1417 = n1416 ^ x307;
  assign n1418 = n1417 ^ x51;
  assign n13542 = n13541 ^ n1418;
  assign n13715 = n13609 ^ n13542;
  assign n13144 = n13048 ^ n12987;
  assign n15100 = n13715 ^ n13144;
  assign n13773 = n13572 ^ n13563;
  assign n13770 = n12460 ^ n11614;
  assign n13771 = n13174 & ~n13770;
  assign n13772 = n13771 ^ n11614;
  assign n13774 = n13773 ^ n13772;
  assign n13777 = n12472 ^ n11627;
  assign n13778 = n13179 & n13777;
  assign n13779 = n13778 ^ n11627;
  assign n13776 = n13566 ^ n13481;
  assign n13780 = n13779 ^ n13776;
  assign n13864 = n12480 ^ n11638;
  assign n13865 = n13192 & n13864;
  assign n13866 = n13865 ^ n11638;
  assign n13818 = n11927 ^ n11231;
  assign n13819 = ~n12623 & ~n13818;
  assign n13820 = n13819 ^ n11231;
  assign n13795 = n11961 ^ n11237;
  assign n13796 = n12625 & n13795;
  assign n13797 = n13796 ^ n11237;
  assign n13688 = n13082 ^ n12971;
  assign n13813 = n13797 ^ n13688;
  assign n13784 = n11939 ^ n11262;
  assign n13785 = ~n12631 & ~n13784;
  assign n13786 = n13785 ^ n11262;
  assign n13694 = n13079 ^ n1635;
  assign n13787 = n13786 ^ n13694;
  assign n13464 = n13075 ^ n12974;
  assign n13460 = n11945 ^ n11246;
  assign n13461 = n12363 & n13460;
  assign n13462 = n13461 ^ n11246;
  assign n13788 = n13464 ^ n13462;
  assign n13314 = n13072 ^ n2744;
  assign n13310 = n11948 ^ n11255;
  assign n13311 = n12370 & n13310;
  assign n13312 = n13311 ^ n11255;
  assign n13456 = n13314 ^ n13312;
  assign n13117 = n13068 ^ n12977;
  assign n13114 = n12385 ^ n11669;
  assign n13115 = n12371 & ~n13114;
  assign n13116 = n13115 ^ n11669;
  assign n13118 = n13117 ^ n13116;
  assign n13122 = n13065 ^ n12979;
  assign n13119 = n12391 ^ n11676;
  assign n13120 = n12373 & n13119;
  assign n13121 = n13120 ^ n11676;
  assign n13123 = n13122 ^ n13121;
  assign n13127 = n13062 ^ n12981;
  assign n13124 = n12398 ^ n11677;
  assign n13125 = n12378 & n13124;
  assign n13126 = n13125 ^ n11677;
  assign n13128 = n13127 ^ n13126;
  assign n13132 = n13059 ^ n2464;
  assign n13129 = n12406 ^ n11005;
  assign n13130 = ~n12384 & ~n13129;
  assign n13131 = n13130 ^ n11005;
  assign n13133 = n13132 ^ n13131;
  assign n13135 = n12412 ^ n11558;
  assign n13136 = n12396 & n13135;
  assign n13137 = n13136 ^ n11558;
  assign n13134 = n13055 ^ n12984;
  assign n13138 = n13137 ^ n13134;
  assign n13140 = n12355 ^ n11566;
  assign n13141 = ~n12403 & ~n13140;
  assign n13142 = n13141 ^ n11566;
  assign n13139 = n13052 ^ n2477;
  assign n13143 = n13142 ^ n13139;
  assign n13145 = n12165 ^ n11572;
  assign n13146 = n12410 & ~n13145;
  assign n13147 = n13146 ^ n11572;
  assign n13148 = n13147 ^ n13144;
  assign n13150 = n12029 ^ n11580;
  assign n13151 = n12417 & ~n13150;
  assign n13152 = n13151 ^ n11580;
  assign n13149 = n13045 ^ n1287;
  assign n13153 = n13152 ^ n13149;
  assign n13155 = n11586 ^ n11556;
  assign n13156 = n12422 & n13155;
  assign n13157 = n13156 ^ n11586;
  assign n13154 = n13041 ^ n12990;
  assign n13158 = n13157 ^ n13154;
  assign n13160 = n11594 ^ n11563;
  assign n13161 = ~n12428 & ~n13160;
  assign n13162 = n13161 ^ n11594;
  assign n13159 = n13038 ^ n992;
  assign n13163 = n13162 ^ n13159;
  assign n13165 = n11602 ^ n11570;
  assign n13166 = ~n12433 & n13165;
  assign n13167 = n13166 ^ n11602;
  assign n13164 = n13034 ^ n12993;
  assign n13168 = n13167 ^ n13164;
  assign n13274 = n13273 ^ n13169;
  assign n13275 = ~n13173 & n13274;
  assign n13276 = n13275 ^ n13172;
  assign n13277 = n13276 ^ n13164;
  assign n13278 = ~n13168 & n13277;
  assign n13279 = n13278 ^ n13167;
  assign n13280 = n13279 ^ n13159;
  assign n13281 = n13163 & n13280;
  assign n13282 = n13281 ^ n13162;
  assign n13283 = n13282 ^ n13154;
  assign n13284 = n13158 & ~n13283;
  assign n13285 = n13284 ^ n13157;
  assign n13286 = n13285 ^ n13149;
  assign n13287 = n13153 & ~n13286;
  assign n13288 = n13287 ^ n13152;
  assign n13289 = n13288 ^ n13144;
  assign n13290 = ~n13148 & n13289;
  assign n13291 = n13290 ^ n13147;
  assign n13292 = n13291 ^ n13139;
  assign n13293 = n13143 & ~n13292;
  assign n13294 = n13293 ^ n13142;
  assign n13295 = n13294 ^ n13134;
  assign n13296 = ~n13138 & ~n13295;
  assign n13297 = n13296 ^ n13137;
  assign n13298 = n13297 ^ n13132;
  assign n13299 = n13133 & ~n13298;
  assign n13300 = n13299 ^ n13131;
  assign n13301 = n13300 ^ n13127;
  assign n13302 = n13128 & ~n13301;
  assign n13303 = n13302 ^ n13126;
  assign n13304 = n13303 ^ n13122;
  assign n13305 = ~n13123 & n13304;
  assign n13306 = n13305 ^ n13121;
  assign n13307 = n13306 ^ n13117;
  assign n13308 = n13118 & ~n13307;
  assign n13309 = n13308 ^ n13116;
  assign n13457 = n13314 ^ n13309;
  assign n13458 = ~n13456 & ~n13457;
  assign n13459 = n13458 ^ n13312;
  assign n13789 = n13464 ^ n13459;
  assign n13790 = ~n13788 & ~n13789;
  assign n13791 = n13790 ^ n13462;
  assign n13792 = n13791 ^ n13694;
  assign n13793 = n13787 & ~n13792;
  assign n13794 = n13793 ^ n13786;
  assign n13814 = n13794 ^ n13688;
  assign n13815 = ~n13813 & ~n13814;
  assign n13816 = n13815 ^ n13797;
  assign n13682 = n13085 ^ n12969;
  assign n13817 = n13816 ^ n13682;
  assign n13821 = n13820 ^ n13817;
  assign n13822 = n13821 ^ n10598;
  assign n13798 = n13797 ^ n13794;
  assign n13799 = n13798 ^ n13688;
  assign n13800 = n13799 ^ n10604;
  assign n13801 = n13791 ^ n13786;
  assign n13802 = n13801 ^ n13694;
  assign n13803 = n13802 ^ n10629;
  assign n13463 = n13462 ^ n13459;
  assign n13465 = n13464 ^ n13463;
  assign n13466 = n13465 ^ n10613;
  assign n13313 = n13312 ^ n13309;
  assign n13315 = n13314 ^ n13313;
  assign n13316 = n13315 ^ n10619;
  assign n13317 = n13306 ^ n13118;
  assign n13318 = n13317 ^ n11061;
  assign n13319 = n13303 ^ n13123;
  assign n13320 = n13319 ^ n11007;
  assign n13321 = n13300 ^ n13128;
  assign n13322 = n13321 ^ n11064;
  assign n13323 = n13297 ^ n13133;
  assign n13324 = n13323 ^ n11066;
  assign n13325 = n13294 ^ n13137;
  assign n13326 = n13325 ^ n13134;
  assign n13327 = n13326 ^ n11072;
  assign n13328 = n13291 ^ n13143;
  assign n13329 = n13328 ^ n11078;
  assign n13330 = n13288 ^ n13148;
  assign n13331 = n13330 ^ n11083;
  assign n13332 = n13285 ^ n13152;
  assign n13333 = n13332 ^ n13149;
  assign n13334 = n13333 ^ n11085;
  assign n13335 = n13282 ^ n13157;
  assign n13336 = n13335 ^ n13154;
  assign n13337 = n13336 ^ n10993;
  assign n13338 = n13279 ^ n13162;
  assign n13339 = n13338 ^ n13159;
  assign n13340 = n13339 ^ n10869;
  assign n13341 = n13276 ^ n13168;
  assign n13342 = n13341 ^ n10806;
  assign n13417 = n13416 ^ n13343;
  assign n13418 = n13344 & ~n13417;
  assign n13419 = n13418 ^ n10693;
  assign n13420 = n13419 ^ n13341;
  assign n13421 = n13342 & ~n13420;
  assign n13422 = n13421 ^ n10806;
  assign n13423 = n13422 ^ n13339;
  assign n13424 = n13340 & n13423;
  assign n13425 = n13424 ^ n10869;
  assign n13426 = n13425 ^ n13336;
  assign n13427 = n13337 & n13426;
  assign n13428 = n13427 ^ n10993;
  assign n13429 = n13428 ^ n13333;
  assign n13430 = ~n13334 & ~n13429;
  assign n13431 = n13430 ^ n11085;
  assign n13432 = n13431 ^ n13330;
  assign n13433 = ~n13331 & ~n13432;
  assign n13434 = n13433 ^ n11083;
  assign n13435 = n13434 ^ n13328;
  assign n13436 = ~n13329 & ~n13435;
  assign n13437 = n13436 ^ n11078;
  assign n13438 = n13437 ^ n13326;
  assign n13439 = ~n13327 & ~n13438;
  assign n13440 = n13439 ^ n11072;
  assign n13441 = n13440 ^ n13323;
  assign n13442 = ~n13324 & n13441;
  assign n13443 = n13442 ^ n11066;
  assign n13444 = n13443 ^ n13321;
  assign n13445 = ~n13322 & n13444;
  assign n13446 = n13445 ^ n11064;
  assign n13447 = n13446 ^ n13319;
  assign n13448 = n13320 & ~n13447;
  assign n13449 = n13448 ^ n11007;
  assign n13450 = n13449 ^ n13317;
  assign n13451 = n13318 & n13450;
  assign n13452 = n13451 ^ n11061;
  assign n13453 = n13452 ^ n13315;
  assign n13454 = n13316 & n13453;
  assign n13455 = n13454 ^ n10619;
  assign n13804 = n13465 ^ n13455;
  assign n13805 = n13466 & n13804;
  assign n13806 = n13805 ^ n10613;
  assign n13807 = n13806 ^ n13802;
  assign n13808 = ~n13803 & ~n13807;
  assign n13809 = n13808 ^ n10629;
  assign n13810 = n13809 ^ n13799;
  assign n13811 = ~n13800 & ~n13810;
  assign n13812 = n13811 ^ n10604;
  assign n13856 = n13821 ^ n13812;
  assign n13857 = n13822 & n13856;
  assign n13858 = n13857 ^ n10598;
  assign n13859 = n13858 ^ n10245;
  assign n13852 = n11667 ^ n11053;
  assign n13853 = ~n12614 & n13852;
  assign n13854 = n13853 ^ n11053;
  assign n13848 = n13820 ^ n13682;
  assign n13849 = n13817 & n13848;
  assign n13850 = n13849 ^ n13820;
  assign n13676 = n13088 ^ n12967;
  assign n13851 = n13850 ^ n13676;
  assign n13855 = n13854 ^ n13851;
  assign n13860 = n13859 ^ n13855;
  assign n13823 = n13822 ^ n13812;
  assign n13824 = n13809 ^ n13800;
  assign n13467 = n13466 ^ n13455;
  assign n13468 = n13452 ^ n13316;
  assign n13469 = n13449 ^ n13318;
  assign n13470 = n13446 ^ n11007;
  assign n13471 = n13470 ^ n13319;
  assign n13472 = n13443 ^ n13322;
  assign n13473 = n13431 ^ n13331;
  assign n13474 = n13419 ^ n13342;
  assign n13502 = n13500 & n13501;
  assign n13503 = n13474 & n13502;
  assign n13504 = n13422 ^ n13340;
  assign n13505 = ~n13503 & ~n13504;
  assign n13506 = n13425 ^ n13337;
  assign n13507 = n13505 & n13506;
  assign n13508 = n13428 ^ n13334;
  assign n13509 = ~n13507 & ~n13508;
  assign n13510 = ~n13473 & ~n13509;
  assign n13511 = n13434 ^ n13329;
  assign n13512 = n13510 & n13511;
  assign n13513 = n13437 ^ n13327;
  assign n13514 = n13512 & ~n13513;
  assign n13515 = n13440 ^ n13324;
  assign n13516 = n13514 & n13515;
  assign n13517 = n13472 & n13516;
  assign n13518 = n13471 & ~n13517;
  assign n13519 = ~n13469 & ~n13518;
  assign n13520 = ~n13468 & ~n13519;
  assign n13825 = ~n13467 & ~n13520;
  assign n13826 = n13806 ^ n13803;
  assign n13827 = ~n13825 & n13826;
  assign n13828 = ~n13824 & n13827;
  assign n13847 = n13823 & ~n13828;
  assign n13861 = n13860 ^ n13847;
  assign n13862 = n13861 ^ n2213;
  assign n13829 = n13828 ^ n13823;
  assign n13830 = n13829 ^ n2028;
  assign n13832 = n13826 ^ n13825;
  assign n13833 = n13832 ^ n1890;
  assign n13522 = n13519 ^ n13468;
  assign n13523 = n13522 ^ n1772;
  assign n13524 = n13518 ^ n13469;
  assign n13525 = n13524 ^ n1780;
  assign n13526 = n13517 ^ n13471;
  assign n13527 = n13526 ^ n1604;
  assign n13529 = n13515 ^ n13514;
  assign n13530 = n13529 ^ n1511;
  assign n13532 = n13511 ^ n13510;
  assign n13533 = n13532 ^ n1490;
  assign n13534 = n13509 ^ n13473;
  assign n13535 = n13534 ^ n2600;
  assign n13538 = n13504 ^ n13503;
  assign n13539 = n13538 ^ n2432;
  assign n13610 = n13609 ^ n13541;
  assign n13611 = ~n13542 & n13610;
  assign n13612 = n13611 ^ n1418;
  assign n13540 = n13502 ^ n13474;
  assign n13613 = n13612 ^ n13540;
  assign n13614 = n13540 ^ n1434;
  assign n13615 = n13613 & ~n13614;
  assign n13616 = n13615 ^ n1434;
  assign n13617 = n13616 ^ n13538;
  assign n13618 = n13539 & ~n13617;
  assign n13619 = n13618 ^ n2432;
  assign n13537 = n13506 ^ n13505;
  assign n13620 = n13619 ^ n13537;
  assign n13621 = n13537 ^ n2606;
  assign n13622 = ~n13620 & n13621;
  assign n13623 = n13622 ^ n2606;
  assign n13536 = n13508 ^ n13507;
  assign n13624 = n13623 ^ n13536;
  assign n13625 = n13536 ^ n2594;
  assign n13626 = n13624 & ~n13625;
  assign n13627 = n13626 ^ n2594;
  assign n13628 = n13627 ^ n13534;
  assign n13629 = n13535 & ~n13628;
  assign n13630 = n13629 ^ n2600;
  assign n13631 = n13630 ^ n13532;
  assign n13632 = n13533 & ~n13631;
  assign n13633 = n13632 ^ n1490;
  assign n13531 = n13513 ^ n13512;
  assign n13634 = n13633 ^ n13531;
  assign n13635 = n13531 ^ n1573;
  assign n13636 = n13634 & ~n13635;
  assign n13637 = n13636 ^ n1573;
  assign n13638 = n13637 ^ n13529;
  assign n13639 = n13530 & ~n13638;
  assign n13640 = n13639 ^ n1511;
  assign n13528 = n13516 ^ n13472;
  assign n13641 = n13640 ^ n13528;
  assign n13642 = n13528 ^ n2944;
  assign n13643 = ~n13641 & n13642;
  assign n13644 = n13643 ^ n2944;
  assign n13645 = n13644 ^ n13526;
  assign n13646 = n13527 & ~n13645;
  assign n13647 = n13646 ^ n1604;
  assign n13648 = n13647 ^ n13524;
  assign n13649 = n13525 & ~n13648;
  assign n13650 = n13649 ^ n1780;
  assign n13651 = n13650 ^ n13522;
  assign n13652 = ~n13523 & n13651;
  assign n13653 = n13652 ^ n1772;
  assign n13521 = n13520 ^ n13467;
  assign n13654 = n13653 ^ n13521;
  assign n13834 = n13521 ^ n1792;
  assign n13835 = ~n13654 & n13834;
  assign n13836 = n13835 ^ n1792;
  assign n13837 = n13836 ^ n13832;
  assign n13838 = n13833 & ~n13837;
  assign n13839 = n13838 ^ n1890;
  assign n13831 = n13827 ^ n13824;
  assign n13840 = n13839 ^ n13831;
  assign n13841 = n13831 ^ n1902;
  assign n13842 = ~n13840 & n13841;
  assign n13843 = n13842 ^ n1902;
  assign n13844 = n13843 ^ n13829;
  assign n13845 = ~n13830 & n13844;
  assign n13846 = n13845 ^ n2028;
  assign n13863 = n13862 ^ n13846;
  assign n13867 = n13866 ^ n13863;
  assign n13869 = n12488 ^ n11643;
  assign n13870 = n13197 & ~n13869;
  assign n13871 = n13870 ^ n11643;
  assign n13868 = n13843 ^ n13830;
  assign n13872 = n13871 ^ n13868;
  assign n13874 = n12494 ^ n11649;
  assign n13875 = n13199 & n13874;
  assign n13876 = n13875 ^ n11649;
  assign n13873 = n13840 ^ n1902;
  assign n13877 = n13876 ^ n13873;
  assign n13878 = n12500 ^ n11654;
  assign n13879 = ~n13203 & n13878;
  assign n13880 = n13879 ^ n11654;
  assign n13881 = n13836 ^ n13833;
  assign n13882 = ~n13880 & n13881;
  assign n13883 = n13882 ^ n13873;
  assign n13884 = ~n13877 & n13883;
  assign n13885 = n13884 ^ n13882;
  assign n13886 = n13885 ^ n13868;
  assign n13887 = ~n13872 & n13886;
  assign n13888 = n13887 ^ n13871;
  assign n13889 = n13888 ^ n13863;
  assign n13890 = n13867 & ~n13889;
  assign n13891 = n13890 ^ n13866;
  assign n13781 = n12474 ^ n11632;
  assign n13782 = n13184 & ~n13781;
  assign n13783 = n13782 ^ n11632;
  assign n13892 = n13891 ^ n13783;
  assign n13909 = n13861 ^ n13846;
  assign n13910 = n13862 & ~n13909;
  assign n13911 = n13910 ^ n2213;
  assign n13912 = n13911 ^ n518;
  assign n13904 = n13855 ^ n10245;
  assign n13905 = n13858 ^ n13855;
  assign n13906 = n13904 & n13905;
  assign n13907 = n13906 ^ n10245;
  assign n13902 = ~n13847 & n13860;
  assign n13898 = n13854 ^ n13676;
  assign n13899 = n13851 & n13898;
  assign n13900 = n13899 ^ n13854;
  assign n13893 = n11662 ^ n11051;
  assign n13894 = n12608 & ~n13893;
  assign n13895 = n13894 ^ n11051;
  assign n13670 = n13092 ^ n1808;
  assign n13896 = n13895 ^ n13670;
  assign n13897 = n13896 ^ n10243;
  assign n13901 = n13900 ^ n13897;
  assign n13903 = n13902 ^ n13901;
  assign n13908 = n13907 ^ n13903;
  assign n13913 = n13912 ^ n13908;
  assign n13914 = n13913 ^ n13891;
  assign n13915 = ~n13892 & ~n13914;
  assign n13916 = n13915 ^ n13783;
  assign n13917 = n13916 ^ n13776;
  assign n13918 = n13780 & n13917;
  assign n13919 = n13918 ^ n13779;
  assign n13775 = n13569 ^ n13568;
  assign n13920 = n13919 ^ n13775;
  assign n13921 = n12466 ^ n11621;
  assign n13922 = ~n13263 & n13921;
  assign n13923 = n13922 ^ n11621;
  assign n13924 = n13923 ^ n13775;
  assign n13925 = ~n13920 & n13924;
  assign n13926 = n13925 ^ n13923;
  assign n13927 = n13926 ^ n13773;
  assign n13928 = n13774 & ~n13927;
  assign n13929 = n13928 ^ n13772;
  assign n13765 = n12455 ^ n11607;
  assign n13766 = ~n13169 & ~n13765;
  assign n13767 = n13766 ^ n11607;
  assign n14056 = n13929 ^ n13767;
  assign n13768 = n13576 ^ n3252;
  assign n14057 = n14056 ^ n13768;
  assign n14058 = n14057 ^ n11386;
  assign n14059 = n13926 ^ n13774;
  assign n14060 = n14059 ^ n11302;
  assign n14061 = n13923 ^ n13920;
  assign n14062 = n14061 ^ n11014;
  assign n14065 = n13913 ^ n13892;
  assign n14066 = n14065 ^ n11024;
  assign n14067 = n13888 ^ n13867;
  assign n14068 = n14067 ^ n11030;
  assign n14069 = n13885 ^ n13872;
  assign n14070 = n14069 ^ n11035;
  assign n14071 = n13881 ^ n13880;
  assign n14072 = n11046 & ~n14071;
  assign n14073 = n14072 ^ n11038;
  assign n14074 = n13882 ^ n13876;
  assign n14075 = n14074 ^ n13873;
  assign n14076 = n14075 ^ n14072;
  assign n14077 = n14073 & ~n14076;
  assign n14078 = n14077 ^ n11038;
  assign n14079 = n14078 ^ n14069;
  assign n14080 = ~n14070 & n14079;
  assign n14081 = n14080 ^ n11035;
  assign n14082 = n14081 ^ n14067;
  assign n14083 = n14068 & ~n14082;
  assign n14084 = n14083 ^ n11030;
  assign n14085 = n14084 ^ n14065;
  assign n14086 = n14066 & n14085;
  assign n14087 = n14086 ^ n11024;
  assign n14063 = n13916 ^ n13779;
  assign n14064 = n14063 ^ n13776;
  assign n14088 = n14087 ^ n14064;
  assign n14089 = n14064 ^ n11019;
  assign n14090 = ~n14088 & n14089;
  assign n14091 = n14090 ^ n11019;
  assign n14092 = n14091 ^ n14061;
  assign n14093 = ~n14062 & n14092;
  assign n14094 = n14093 ^ n11014;
  assign n14095 = n14094 ^ n14059;
  assign n14096 = n14060 & n14095;
  assign n14097 = n14096 ^ n11302;
  assign n14098 = n14097 ^ n14057;
  assign n14099 = n14058 & n14098;
  assign n14100 = n14099 ^ n11386;
  assign n13769 = n13768 ^ n13767;
  assign n13930 = n13929 ^ n13768;
  assign n13931 = ~n13769 & n13930;
  assign n13932 = n13931 ^ n13767;
  assign n13760 = n12447 ^ n11601;
  assign n13761 = ~n13164 & ~n13760;
  assign n13762 = n13761 ^ n11601;
  assign n14053 = n13932 ^ n13762;
  assign n13763 = n13579 ^ n13557;
  assign n14054 = n14053 ^ n13763;
  assign n14055 = n14054 ^ n11432;
  assign n14196 = n14100 ^ n14055;
  assign n14179 = n14091 ^ n14062;
  assign n14180 = n14084 ^ n14066;
  assign n14181 = n14081 ^ n14068;
  assign n14182 = n14071 ^ n11046;
  assign n14183 = n14075 ^ n14073;
  assign n14184 = ~n14182 & n14183;
  assign n14185 = n14078 ^ n14070;
  assign n14186 = n14184 & ~n14185;
  assign n14187 = ~n14181 & ~n14186;
  assign n14188 = ~n14180 & n14187;
  assign n14189 = n14088 ^ n11019;
  assign n14190 = ~n14188 & ~n14189;
  assign n14191 = n14179 & n14190;
  assign n14192 = n14094 ^ n14060;
  assign n14193 = ~n14191 & n14192;
  assign n14194 = n14097 ^ n14058;
  assign n14195 = n14193 & ~n14194;
  assign n14264 = n14196 ^ n14195;
  assign n14265 = n14264 ^ n934;
  assign n14267 = n14192 ^ n14191;
  assign n14268 = n14267 ^ n826;
  assign n14269 = n14190 ^ n14179;
  assign n14270 = n14269 ^ n820;
  assign n14271 = n14189 ^ n14188;
  assign n14272 = n14271 ^ n717;
  assign n14273 = n14187 ^ n14180;
  assign n14277 = n14276 ^ n14273;
  assign n14279 = n14185 ^ n14184;
  assign n14280 = n14279 ^ n635;
  assign n14281 = n2303 & n14182;
  assign n14282 = n14281 ^ n528;
  assign n14283 = n14183 ^ n14182;
  assign n14284 = n14283 ^ n14281;
  assign n14285 = n14282 & n14284;
  assign n14286 = n14285 ^ n528;
  assign n14287 = n14286 ^ n14279;
  assign n14288 = ~n14280 & n14287;
  assign n14289 = n14288 ^ n635;
  assign n14278 = n14186 ^ n14181;
  assign n14290 = n14289 ^ n14278;
  assign n14291 = n14278 ^ n515;
  assign n14292 = n14290 & ~n14291;
  assign n14293 = n14292 ^ n515;
  assign n14294 = n14293 ^ n14273;
  assign n14295 = n14277 & ~n14294;
  assign n14296 = n14295 ^ n14276;
  assign n14297 = n14296 ^ n14271;
  assign n14298 = n14272 & ~n14297;
  assign n14299 = n14298 ^ n717;
  assign n14300 = n14299 ^ n14269;
  assign n14301 = n14270 & ~n14300;
  assign n14302 = n14301 ^ n820;
  assign n14303 = n14302 ^ n14267;
  assign n14304 = n14268 & ~n14303;
  assign n14305 = n14304 ^ n826;
  assign n14266 = n14194 ^ n14193;
  assign n14306 = n14305 ^ n14266;
  assign n14307 = n14266 ^ n838;
  assign n14308 = ~n14306 & n14307;
  assign n14309 = n14308 ^ n838;
  assign n14310 = n14309 ^ n14264;
  assign n14311 = n14265 & ~n14310;
  assign n14312 = n14311 ^ n934;
  assign n14197 = ~n14195 & ~n14196;
  assign n14101 = n14100 ^ n14054;
  assign n14102 = n14055 & n14101;
  assign n14103 = n14102 ^ n11432;
  assign n13764 = n13763 ^ n13762;
  assign n13933 = n13932 ^ n13763;
  assign n13934 = n13764 & ~n13933;
  assign n13935 = n13934 ^ n13762;
  assign n13756 = n12444 ^ n11598;
  assign n13757 = ~n13159 & ~n13756;
  assign n13758 = n13757 ^ n11598;
  assign n14050 = n13935 ^ n13758;
  assign n13755 = n13582 ^ n13555;
  assign n14051 = n14050 ^ n13755;
  assign n14052 = n14051 ^ n11447;
  assign n14178 = n14103 ^ n14052;
  assign n14263 = n14197 ^ n14178;
  assign n14313 = n14312 ^ n14263;
  assign n14314 = n14263 ^ n948;
  assign n14315 = n14313 & ~n14314;
  assign n14316 = n14315 ^ n948;
  assign n14198 = ~n14178 & n14197;
  assign n14104 = n14103 ^ n14051;
  assign n14105 = ~n14052 & n14104;
  assign n14106 = n14105 ^ n11447;
  assign n13759 = n13758 ^ n13755;
  assign n13936 = n13935 ^ n13755;
  assign n13937 = ~n13759 & n13936;
  assign n13938 = n13937 ^ n13758;
  assign n13753 = n13585 ^ n13553;
  assign n13750 = n12439 ^ n11591;
  assign n13751 = ~n13154 & n13750;
  assign n13752 = n13751 ^ n11591;
  assign n13754 = n13753 ^ n13752;
  assign n14048 = n13938 ^ n13754;
  assign n14049 = n14048 ^ n11548;
  assign n14177 = n14106 ^ n14049;
  assign n14261 = n14198 ^ n14177;
  assign n14262 = n14261 ^ n1094;
  assign n14582 = n14316 ^ n14262;
  assign n15101 = n15100 ^ n14582;
  assign n14398 = n13184 ^ n12488;
  assign n14399 = n13773 & ~n14398;
  assign n14400 = n14399 ^ n12488;
  assign n13686 = n13630 ^ n13533;
  assign n13683 = n12385 ^ n12363;
  assign n13684 = n13682 & ~n13683;
  assign n13685 = n13684 ^ n12385;
  assign n13687 = n13686 ^ n13685;
  assign n13692 = n13627 ^ n13535;
  assign n13689 = n12391 ^ n12370;
  assign n13690 = n13688 & n13689;
  assign n13691 = n13690 ^ n12391;
  assign n13693 = n13692 ^ n13691;
  assign n13698 = n13624 ^ n2594;
  assign n13695 = n12398 ^ n12371;
  assign n13696 = n13694 & n13695;
  assign n13697 = n13696 ^ n12398;
  assign n13699 = n13698 ^ n13697;
  assign n13703 = n13620 ^ n2606;
  assign n13700 = n12406 ^ n12373;
  assign n13701 = ~n13464 & ~n13700;
  assign n13702 = n13701 ^ n12406;
  assign n13704 = n13703 ^ n13702;
  assign n13708 = n13616 ^ n13539;
  assign n13705 = n12412 ^ n12378;
  assign n13706 = n13314 & n13705;
  assign n13707 = n13706 ^ n12412;
  assign n13709 = n13708 ^ n13707;
  assign n13713 = n13613 ^ n1434;
  assign n13710 = n12384 ^ n12355;
  assign n13711 = n13117 & ~n13710;
  assign n13712 = n13711 ^ n12355;
  assign n13714 = n13713 ^ n13712;
  assign n13716 = n12396 ^ n12165;
  assign n13717 = ~n13122 & n13716;
  assign n13718 = n13717 ^ n12165;
  assign n13719 = n13718 ^ n13715;
  assign n13721 = n12403 ^ n12029;
  assign n13722 = n13127 & ~n13721;
  assign n13723 = n13722 ^ n12029;
  assign n13720 = n13606 ^ n1172;
  assign n13724 = n13723 ^ n13720;
  assign n13726 = n12410 ^ n11556;
  assign n13727 = n13132 & ~n13726;
  assign n13728 = n13727 ^ n11556;
  assign n13725 = n13602 ^ n13545;
  assign n13729 = n13728 ^ n13725;
  assign n13733 = n13599 ^ n999;
  assign n13730 = n12417 ^ n11563;
  assign n13731 = ~n13134 & n13730;
  assign n13732 = n13731 ^ n11563;
  assign n13734 = n13733 ^ n13732;
  assign n13736 = n12422 ^ n11570;
  assign n13737 = ~n13139 & n13736;
  assign n13738 = n13737 ^ n11570;
  assign n13735 = n13595 ^ n13548;
  assign n13739 = n13738 ^ n13735;
  assign n13741 = n12428 ^ n11577;
  assign n13742 = n13144 & n13741;
  assign n13743 = n13742 ^ n11577;
  assign n13740 = n13592 ^ n856;
  assign n13744 = n13743 ^ n13740;
  assign n13748 = n13588 ^ n13551;
  assign n13745 = n12433 ^ n11584;
  assign n13746 = ~n13149 & ~n13745;
  assign n13747 = n13746 ^ n11584;
  assign n13749 = n13748 ^ n13747;
  assign n13939 = n13938 ^ n13753;
  assign n13940 = ~n13754 & n13939;
  assign n13941 = n13940 ^ n13752;
  assign n13942 = n13941 ^ n13748;
  assign n13943 = ~n13749 & n13942;
  assign n13944 = n13943 ^ n13747;
  assign n13945 = n13944 ^ n13740;
  assign n13946 = ~n13744 & ~n13945;
  assign n13947 = n13946 ^ n13743;
  assign n13948 = n13947 ^ n13735;
  assign n13949 = ~n13739 & ~n13948;
  assign n13950 = n13949 ^ n13738;
  assign n13951 = n13950 ^ n13733;
  assign n13952 = ~n13734 & n13951;
  assign n13953 = n13952 ^ n13732;
  assign n13954 = n13953 ^ n13725;
  assign n13955 = ~n13729 & ~n13954;
  assign n13956 = n13955 ^ n13728;
  assign n13957 = n13956 ^ n13720;
  assign n13958 = ~n13724 & ~n13957;
  assign n13959 = n13958 ^ n13723;
  assign n13960 = n13959 ^ n13715;
  assign n13961 = ~n13719 & n13960;
  assign n13962 = n13961 ^ n13718;
  assign n13963 = n13962 ^ n13713;
  assign n13964 = ~n13714 & n13963;
  assign n13965 = n13964 ^ n13712;
  assign n13966 = n13965 ^ n13708;
  assign n13967 = n13709 & ~n13966;
  assign n13968 = n13967 ^ n13707;
  assign n13969 = n13968 ^ n13703;
  assign n13970 = ~n13704 & ~n13969;
  assign n13971 = n13970 ^ n13702;
  assign n13972 = n13971 ^ n13698;
  assign n13973 = ~n13699 & ~n13972;
  assign n13974 = n13973 ^ n13697;
  assign n13975 = n13974 ^ n13692;
  assign n13976 = n13693 & ~n13975;
  assign n13977 = n13976 ^ n13691;
  assign n13978 = n13977 ^ n13686;
  assign n13979 = ~n13687 & ~n13978;
  assign n13980 = n13979 ^ n13685;
  assign n13680 = n13634 ^ n1573;
  assign n13677 = n12631 ^ n11948;
  assign n13678 = ~n13676 & n13677;
  assign n13679 = n13678 ^ n11948;
  assign n13681 = n13680 ^ n13679;
  assign n14019 = n13980 ^ n13681;
  assign n14020 = n14019 ^ n11255;
  assign n14021 = n13977 ^ n13687;
  assign n14022 = n14021 ^ n11669;
  assign n14023 = n13974 ^ n13693;
  assign n14024 = n14023 ^ n11676;
  assign n14025 = n13971 ^ n13699;
  assign n14026 = n14025 ^ n11677;
  assign n14027 = n13968 ^ n13704;
  assign n14028 = n14027 ^ n11005;
  assign n14029 = n13965 ^ n13709;
  assign n14030 = n14029 ^ n11558;
  assign n14031 = n13962 ^ n13714;
  assign n14032 = n14031 ^ n11566;
  assign n14033 = n13959 ^ n13719;
  assign n14034 = n14033 ^ n11572;
  assign n14035 = n13956 ^ n13724;
  assign n14036 = n14035 ^ n11580;
  assign n14037 = n13953 ^ n13729;
  assign n14038 = n14037 ^ n11586;
  assign n14039 = n13950 ^ n13732;
  assign n14040 = n14039 ^ n13733;
  assign n14041 = n14040 ^ n11594;
  assign n14042 = n13947 ^ n13739;
  assign n14043 = n14042 ^ n11602;
  assign n14044 = n13944 ^ n13744;
  assign n14045 = n14044 ^ n11609;
  assign n14046 = n13941 ^ n13749;
  assign n14047 = n14046 ^ n11615;
  assign n14107 = n14106 ^ n14048;
  assign n14108 = n14049 & n14107;
  assign n14109 = n14108 ^ n11548;
  assign n14110 = n14109 ^ n14046;
  assign n14111 = ~n14047 & ~n14110;
  assign n14112 = n14111 ^ n11615;
  assign n14113 = n14112 ^ n14044;
  assign n14114 = ~n14045 & n14113;
  assign n14115 = n14114 ^ n11609;
  assign n14116 = n14115 ^ n14042;
  assign n14117 = n14043 & ~n14116;
  assign n14118 = n14117 ^ n11602;
  assign n14119 = n14118 ^ n14040;
  assign n14120 = n14041 & n14119;
  assign n14121 = n14120 ^ n11594;
  assign n14122 = n14121 ^ n14037;
  assign n14123 = n14038 & ~n14122;
  assign n14124 = n14123 ^ n11586;
  assign n14125 = n14124 ^ n14035;
  assign n14126 = ~n14036 & n14125;
  assign n14127 = n14126 ^ n11580;
  assign n14128 = n14127 ^ n14033;
  assign n14129 = n14034 & ~n14128;
  assign n14130 = n14129 ^ n11572;
  assign n14131 = n14130 ^ n14031;
  assign n14132 = n14032 & ~n14131;
  assign n14133 = n14132 ^ n11566;
  assign n14134 = n14133 ^ n14029;
  assign n14135 = n14030 & n14134;
  assign n14136 = n14135 ^ n11558;
  assign n14137 = n14136 ^ n14027;
  assign n14138 = ~n14028 & n14137;
  assign n14139 = n14138 ^ n11005;
  assign n14140 = n14139 ^ n14025;
  assign n14141 = n14026 & ~n14140;
  assign n14142 = n14141 ^ n11677;
  assign n14143 = n14142 ^ n14023;
  assign n14144 = n14024 & ~n14143;
  assign n14145 = n14144 ^ n11676;
  assign n14146 = n14145 ^ n14021;
  assign n14147 = ~n14022 & n14146;
  assign n14148 = n14147 ^ n11669;
  assign n14149 = n14148 ^ n14019;
  assign n14150 = n14020 & n14149;
  assign n14151 = n14150 ^ n11255;
  assign n13981 = n13980 ^ n13680;
  assign n13982 = n13681 & ~n13981;
  assign n13983 = n13982 ^ n13679;
  assign n13674 = n13637 ^ n13530;
  assign n13671 = n12625 ^ n11945;
  assign n13672 = ~n13670 & n13671;
  assign n13673 = n13672 ^ n11945;
  assign n13675 = n13674 ^ n13673;
  assign n14017 = n13983 ^ n13675;
  assign n14018 = n14017 ^ n11246;
  assign n14168 = n14151 ^ n14018;
  assign n14169 = n14145 ^ n14022;
  assign n14170 = n14142 ^ n14024;
  assign n14171 = n14136 ^ n14028;
  assign n14172 = n14130 ^ n14032;
  assign n14173 = n14127 ^ n14034;
  assign n14174 = n14121 ^ n14038;
  assign n14175 = n14115 ^ n14043;
  assign n14176 = n14112 ^ n14045;
  assign n14199 = ~n14177 & ~n14198;
  assign n14200 = n14109 ^ n14047;
  assign n14201 = n14199 & ~n14200;
  assign n14202 = n14176 & n14201;
  assign n14203 = ~n14175 & n14202;
  assign n14204 = n14118 ^ n14041;
  assign n14205 = ~n14203 & n14204;
  assign n14206 = ~n14174 & n14205;
  assign n14207 = n14124 ^ n14036;
  assign n14208 = ~n14206 & ~n14207;
  assign n14209 = ~n14173 & ~n14208;
  assign n14210 = ~n14172 & n14209;
  assign n14211 = n14133 ^ n14030;
  assign n14212 = n14210 & ~n14211;
  assign n14213 = ~n14171 & n14212;
  assign n14214 = n14139 ^ n14026;
  assign n14215 = n14213 & n14214;
  assign n14216 = ~n14170 & ~n14215;
  assign n14217 = ~n14169 & ~n14216;
  assign n14218 = n14148 ^ n14020;
  assign n14219 = ~n14217 & ~n14218;
  assign n14220 = n14168 & ~n14219;
  assign n14152 = n14151 ^ n14017;
  assign n14153 = ~n14018 & ~n14152;
  assign n14154 = n14153 ^ n11246;
  assign n13984 = n13983 ^ n13674;
  assign n13985 = n13675 & n13984;
  assign n13986 = n13985 ^ n13673;
  assign n13666 = n12623 ^ n11939;
  assign n13667 = n13219 & n13666;
  assign n13668 = n13667 ^ n11939;
  assign n14014 = n13986 ^ n13668;
  assign n13665 = n13641 ^ n2944;
  assign n14015 = n14014 ^ n13665;
  assign n14016 = n14015 ^ n11262;
  assign n14167 = n14154 ^ n14016;
  assign n14236 = n14220 ^ n14167;
  assign n14237 = n14236 ^ n1814;
  assign n14239 = n14218 ^ n14217;
  assign n14240 = n14239 ^ n1719;
  assign n14241 = n14216 ^ n14169;
  assign n14242 = n14241 ^ n1627;
  assign n14243 = n14215 ^ n14170;
  assign n14244 = n14243 ^ n1621;
  assign n14246 = n14212 ^ n14171;
  assign n14247 = n14246 ^ n1500;
  assign n14249 = n14209 ^ n14172;
  assign n14250 = n14249 ^ n2627;
  assign n14251 = n14208 ^ n14173;
  assign n14252 = n14251 ^ n2772;
  assign n14255 = n14204 ^ n14203;
  assign n2468 = x497 ^ x145;
  assign n2469 = n2468 ^ x337;
  assign n2470 = n2469 ^ x81;
  assign n14256 = n14255 ^ n2470;
  assign n14258 = n14201 ^ n14176;
  assign n14259 = n14258 ^ n1279;
  assign n14317 = n14316 ^ n14261;
  assign n14318 = ~n14262 & n14317;
  assign n14319 = n14318 ^ n1094;
  assign n14260 = n14200 ^ n14199;
  assign n14320 = n14319 ^ n14260;
  assign n1271 = x500 ^ x148;
  assign n1272 = n1271 ^ x340;
  assign n1273 = n1272 ^ x84;
  assign n14321 = n14260 ^ n1273;
  assign n14322 = ~n14320 & n14321;
  assign n14323 = n14322 ^ n1273;
  assign n14324 = n14323 ^ n14258;
  assign n14325 = ~n14259 & n14324;
  assign n14326 = n14325 ^ n1279;
  assign n14257 = n14202 ^ n14175;
  assign n14327 = n14326 ^ n14257;
  assign n2421 = x498 ^ x146;
  assign n2422 = n2421 ^ x338;
  assign n2423 = n2422 ^ x82;
  assign n14328 = n14257 ^ n2423;
  assign n14329 = ~n14327 & n14328;
  assign n14330 = n14329 ^ n2423;
  assign n14331 = n14330 ^ n14255;
  assign n14332 = ~n14256 & n14331;
  assign n14333 = n14332 ^ n2470;
  assign n14254 = n14205 ^ n14174;
  assign n14334 = n14333 ^ n14254;
  assign n14335 = n14254 ^ n1550;
  assign n14336 = n14334 & ~n14335;
  assign n14337 = n14336 ^ n1550;
  assign n14253 = n14207 ^ n14206;
  assign n14338 = n14337 ^ n14253;
  assign n14339 = n14253 ^ n2535;
  assign n14340 = n14338 & ~n14339;
  assign n14341 = n14340 ^ n2535;
  assign n14342 = n14341 ^ n14251;
  assign n14343 = n14252 & ~n14342;
  assign n14344 = n14343 ^ n2772;
  assign n14345 = n14344 ^ n14249;
  assign n14346 = ~n14250 & n14345;
  assign n14347 = n14346 ^ n2627;
  assign n14248 = n14211 ^ n14210;
  assign n14348 = n14347 ^ n14248;
  assign n14349 = n14248 ^ n2786;
  assign n14350 = n14348 & ~n14349;
  assign n14351 = n14350 ^ n2786;
  assign n14352 = n14351 ^ n14246;
  assign n14353 = ~n14247 & n14352;
  assign n14354 = n14353 ^ n1500;
  assign n14245 = n14214 ^ n14213;
  assign n14355 = n14354 ^ n14245;
  assign n14356 = n14245 ^ n1537;
  assign n14357 = ~n14355 & n14356;
  assign n14358 = n14357 ^ n1537;
  assign n14359 = n14358 ^ n14243;
  assign n14360 = ~n14244 & n14359;
  assign n14361 = n14360 ^ n1621;
  assign n14362 = n14361 ^ n14241;
  assign n14363 = n14242 & ~n14362;
  assign n14364 = n14363 ^ n1627;
  assign n14365 = n14364 ^ n14239;
  assign n14366 = ~n14240 & n14365;
  assign n14367 = n14366 ^ n1719;
  assign n14238 = n14219 ^ n14168;
  assign n14368 = n14367 ^ n14238;
  assign n14369 = n14238 ^ n1996;
  assign n14370 = n14368 & ~n14369;
  assign n14371 = n14370 ^ n1996;
  assign n14372 = n14371 ^ n14236;
  assign n14373 = n14237 & ~n14372;
  assign n14374 = n14373 ^ n1814;
  assign n14221 = n14167 & ~n14220;
  assign n14155 = n14154 ^ n14015;
  assign n14156 = ~n14016 & n14155;
  assign n14157 = n14156 ^ n11262;
  assign n13669 = n13668 ^ n13665;
  assign n13987 = n13986 ^ n13665;
  assign n13988 = ~n13669 & ~n13987;
  assign n13989 = n13988 ^ n13668;
  assign n13660 = n12614 ^ n11961;
  assign n13661 = ~n13214 & n13660;
  assign n13662 = n13661 ^ n11961;
  assign n14011 = n13989 ^ n13662;
  assign n13663 = n13644 ^ n13527;
  assign n14012 = n14011 ^ n13663;
  assign n14013 = n14012 ^ n11237;
  assign n14166 = n14157 ^ n14013;
  assign n14235 = n14221 ^ n14166;
  assign n14375 = n14374 ^ n14235;
  assign n14376 = n14235 ^ n1989;
  assign n14377 = n14375 & ~n14376;
  assign n14378 = n14377 ^ n1989;
  assign n14158 = n14157 ^ n14012;
  assign n14159 = ~n14013 & ~n14158;
  assign n14160 = n14159 ^ n11237;
  assign n13994 = n12608 ^ n11927;
  assign n13995 = n13231 & ~n13994;
  assign n13996 = n13995 ^ n11927;
  assign n13664 = n13663 ^ n13662;
  assign n13990 = n13989 ^ n13663;
  assign n13991 = ~n13664 & n13990;
  assign n13992 = n13991 ^ n13662;
  assign n13659 = n13647 ^ n13525;
  assign n13993 = n13992 ^ n13659;
  assign n14009 = n13996 ^ n13993;
  assign n14010 = n14009 ^ n11231;
  assign n14223 = n14160 ^ n14010;
  assign n14222 = n14166 & n14221;
  assign n14233 = n14223 ^ n14222;
  assign n14234 = n14233 ^ n2021;
  assign n14397 = n14378 ^ n14234;
  assign n14401 = n14400 ^ n14397;
  assign n14405 = n14375 ^ n1989;
  assign n14402 = n13192 ^ n12494;
  assign n14403 = n13775 & n14402;
  assign n14404 = n14403 ^ n12494;
  assign n14406 = n14405 ^ n14404;
  assign n14407 = n14371 ^ n14237;
  assign n14408 = n13197 ^ n12500;
  assign n14409 = n13776 & ~n14408;
  assign n14410 = n14409 ^ n12500;
  assign n14411 = n14407 & ~n14410;
  assign n14412 = n14411 ^ n14405;
  assign n14413 = n14406 & ~n14412;
  assign n14414 = n14413 ^ n14411;
  assign n14415 = n14414 ^ n14397;
  assign n14416 = ~n14401 & ~n14415;
  assign n14417 = n14416 ^ n14400;
  assign n14393 = n13179 ^ n12480;
  assign n14394 = ~n13768 & n14393;
  assign n14395 = n14394 ^ n12480;
  assign n14379 = n14378 ^ n14233;
  assign n14380 = n14234 & ~n14379;
  assign n14381 = n14380 ^ n2021;
  assign n14224 = ~n14222 & ~n14223;
  assign n14161 = n14160 ^ n14009;
  assign n14162 = n14010 & n14161;
  assign n14163 = n14162 ^ n11231;
  assign n14164 = n14163 ^ n11053;
  assign n14001 = n12507 ^ n11667;
  assign n14002 = ~n13209 & ~n14001;
  assign n14003 = n14002 ^ n11667;
  assign n13997 = n13996 ^ n13659;
  assign n13998 = n13993 & ~n13997;
  assign n13999 = n13998 ^ n13996;
  assign n13658 = n13650 ^ n13523;
  assign n14000 = n13999 ^ n13658;
  assign n14008 = n14003 ^ n14000;
  assign n14165 = n14164 ^ n14008;
  assign n14232 = n14224 ^ n14165;
  assign n14382 = n14381 ^ n14232;
  assign n14392 = n14382 ^ n2149;
  assign n14396 = n14395 ^ n14392;
  assign n14423 = n14417 ^ n14396;
  assign n14424 = n14423 ^ n11638;
  assign n14425 = n14414 ^ n14401;
  assign n14426 = n14425 ^ n11643;
  assign n14427 = n14410 ^ n14407;
  assign n14428 = ~n11654 & ~n14427;
  assign n14429 = n14428 ^ n11649;
  assign n14430 = n14411 ^ n14404;
  assign n14431 = n14430 ^ n14405;
  assign n14432 = n14431 ^ n14428;
  assign n14433 = n14429 & n14432;
  assign n14434 = n14433 ^ n11649;
  assign n14435 = n14434 ^ n14425;
  assign n14436 = ~n14426 & n14435;
  assign n14437 = n14436 ^ n11643;
  assign n14438 = n14437 ^ n14423;
  assign n14439 = n14424 & ~n14438;
  assign n14440 = n14439 ^ n11638;
  assign n14418 = n14417 ^ n14392;
  assign n14419 = ~n14396 & ~n14418;
  assign n14420 = n14419 ^ n14395;
  assign n14388 = n13263 ^ n12474;
  assign n14389 = n13763 & ~n14388;
  assign n14390 = n14389 ^ n12474;
  assign n14383 = n14232 ^ n2149;
  assign n14384 = n14382 & ~n14383;
  assign n14385 = n14384 ^ n2149;
  assign n14386 = n14385 ^ n2308;
  assign n14227 = n14008 ^ n11053;
  assign n14228 = n14163 ^ n14008;
  assign n14229 = n14227 & n14228;
  assign n14230 = n14229 ^ n11053;
  assign n14225 = ~n14165 & ~n14224;
  assign n14004 = n14003 ^ n13658;
  assign n14005 = ~n14000 & n14004;
  assign n14006 = n14005 ^ n14003;
  assign n13655 = n13654 ^ n1792;
  assign n13111 = n12502 ^ n11662;
  assign n13112 = n13110 & n13111;
  assign n13113 = n13112 ^ n11662;
  assign n13656 = n13655 ^ n13113;
  assign n13657 = n13656 ^ n11051;
  assign n14007 = n14006 ^ n13657;
  assign n14226 = n14225 ^ n14007;
  assign n14231 = n14230 ^ n14226;
  assign n14387 = n14386 ^ n14231;
  assign n14391 = n14390 ^ n14387;
  assign n14421 = n14420 ^ n14391;
  assign n14422 = n14421 ^ n11632;
  assign n14463 = n14440 ^ n14422;
  assign n14456 = n14437 ^ n14424;
  assign n14457 = n14434 ^ n14426;
  assign n14458 = n14427 ^ n11654;
  assign n14459 = n14431 ^ n14429;
  assign n14460 = n14458 & ~n14459;
  assign n14461 = ~n14457 & n14460;
  assign n14462 = ~n14456 & ~n14461;
  assign n14467 = n14463 ^ n14462;
  assign n14468 = n14467 ^ n562;
  assign n14470 = n14460 ^ n14457;
  assign n14471 = n14470 ^ n3245;
  assign n14475 = ~n14458 & n14474;
  assign n14479 = n14478 ^ n14475;
  assign n14480 = n14459 ^ n14458;
  assign n14481 = n14480 ^ n14475;
  assign n14482 = n14479 & n14481;
  assign n14483 = n14482 ^ n14478;
  assign n14484 = n14483 ^ n14470;
  assign n14485 = ~n14471 & n14484;
  assign n14486 = n14485 ^ n3245;
  assign n14469 = n14461 ^ n14456;
  assign n14487 = n14486 ^ n14469;
  assign n14488 = n14469 ^ n556;
  assign n14489 = n14487 & ~n14488;
  assign n14490 = n14489 ^ n556;
  assign n14491 = n14490 ^ n14467;
  assign n14492 = ~n14468 & n14491;
  assign n14493 = n14492 ^ n562;
  assign n14464 = n14462 & n14463;
  assign n14451 = n14182 ^ n2303;
  assign n14448 = n13174 ^ n12472;
  assign n14449 = ~n13755 & n14448;
  assign n14450 = n14449 ^ n12472;
  assign n14452 = n14451 ^ n14450;
  assign n14444 = n14420 ^ n14390;
  assign n14445 = n14420 ^ n14387;
  assign n14446 = n14444 & ~n14445;
  assign n14447 = n14446 ^ n14390;
  assign n14453 = n14452 ^ n14447;
  assign n14454 = n14453 ^ n11627;
  assign n14441 = n14440 ^ n14421;
  assign n14442 = ~n14422 & ~n14441;
  assign n14443 = n14442 ^ n11632;
  assign n14455 = n14454 ^ n14443;
  assign n14465 = n14464 ^ n14455;
  assign n14466 = n14465 ^ n585;
  assign n14518 = n14493 ^ n14466;
  assign n14516 = n14313 ^ n948;
  assign n14515 = n13720 ^ n13149;
  assign n14517 = n14516 ^ n14515;
  assign n14519 = n14518 ^ n14517;
  assign n15065 = n14474 ^ n14458;
  assign n15040 = n13768 ^ n13192;
  assign n14506 = n14283 ^ n14282;
  assign n15041 = n15040 ^ n14506;
  assign n14684 = n14341 ^ n14252;
  assign n14676 = n14338 ^ n2535;
  assign n14555 = n13688 ^ n12373;
  assign n14556 = n13674 & n14555;
  assign n14557 = n14556 ^ n12373;
  assign n14554 = n14334 ^ n1550;
  assign n14558 = n14557 ^ n14554;
  assign n14560 = n13694 ^ n12378;
  assign n14561 = ~n13680 & n14560;
  assign n14562 = n14561 ^ n12378;
  assign n14559 = n14330 ^ n14256;
  assign n14563 = n14562 ^ n14559;
  assign n14567 = n14327 ^ n2423;
  assign n14564 = n13464 ^ n12384;
  assign n14565 = n13686 & n14564;
  assign n14566 = n14565 ^ n12384;
  assign n14568 = n14567 ^ n14566;
  assign n14570 = n13314 ^ n12396;
  assign n14571 = n13692 & n14570;
  assign n14572 = n14571 ^ n12396;
  assign n14569 = n14323 ^ n14259;
  assign n14573 = n14572 ^ n14569;
  assign n14577 = n14320 ^ n1273;
  assign n14574 = n13117 ^ n12403;
  assign n14575 = ~n13698 & ~n14574;
  assign n14576 = n14575 ^ n12403;
  assign n14578 = n14577 ^ n14576;
  assign n14579 = n13122 ^ n12410;
  assign n14580 = n13703 & ~n14579;
  assign n14581 = n14580 ^ n12410;
  assign n14583 = n14582 ^ n14581;
  assign n14584 = n13127 ^ n12417;
  assign n14585 = n13708 & n14584;
  assign n14586 = n14585 ^ n12417;
  assign n14587 = n14586 ^ n14516;
  assign n14591 = n14309 ^ n14265;
  assign n14588 = n13132 ^ n12422;
  assign n14589 = ~n13713 & n14588;
  assign n14590 = n14589 ^ n12422;
  assign n14592 = n14591 ^ n14590;
  assign n14596 = n14306 ^ n838;
  assign n14593 = n13134 ^ n12428;
  assign n14594 = ~n13715 & n14593;
  assign n14595 = n14594 ^ n12428;
  assign n14597 = n14596 ^ n14595;
  assign n14599 = n13139 ^ n12433;
  assign n14600 = ~n13720 & n14599;
  assign n14601 = n14600 ^ n12433;
  assign n14598 = n14302 ^ n14268;
  assign n14602 = n14601 ^ n14598;
  assign n14606 = n14299 ^ n14270;
  assign n14603 = n13144 ^ n12439;
  assign n14604 = n13725 & n14603;
  assign n14605 = n14604 ^ n12439;
  assign n14607 = n14606 ^ n14605;
  assign n14611 = n14296 ^ n14272;
  assign n14608 = n13149 ^ n12444;
  assign n14609 = ~n13733 & n14608;
  assign n14610 = n14609 ^ n12444;
  assign n14612 = n14611 ^ n14610;
  assign n14614 = n13154 ^ n12447;
  assign n14615 = ~n13735 & n14614;
  assign n14616 = n14615 ^ n12447;
  assign n14613 = n14293 ^ n14277;
  assign n14617 = n14616 ^ n14613;
  assign n14619 = n13159 ^ n12455;
  assign n14620 = n13740 & n14619;
  assign n14621 = n14620 ^ n12455;
  assign n14618 = n14290 ^ n515;
  assign n14622 = n14621 ^ n14618;
  assign n14626 = n14286 ^ n14280;
  assign n14623 = n13164 ^ n12460;
  assign n14624 = ~n13748 & n14623;
  assign n14625 = n14624 ^ n12460;
  assign n14627 = n14626 ^ n14625;
  assign n14503 = n13169 ^ n12466;
  assign n14504 = ~n13753 & ~n14503;
  assign n14505 = n14504 ^ n12466;
  assign n14507 = n14506 ^ n14505;
  assign n14500 = n14451 ^ n14447;
  assign n14501 = n14452 & ~n14500;
  assign n14502 = n14501 ^ n14450;
  assign n14628 = n14506 ^ n14502;
  assign n14629 = ~n14507 & n14628;
  assign n14630 = n14629 ^ n14505;
  assign n14631 = n14630 ^ n14626;
  assign n14632 = n14627 & n14631;
  assign n14633 = n14632 ^ n14625;
  assign n14634 = n14633 ^ n14618;
  assign n14635 = n14622 & ~n14634;
  assign n14636 = n14635 ^ n14621;
  assign n14637 = n14636 ^ n14613;
  assign n14638 = ~n14617 & n14637;
  assign n14639 = n14638 ^ n14616;
  assign n14640 = n14639 ^ n14611;
  assign n14641 = ~n14612 & n14640;
  assign n14642 = n14641 ^ n14610;
  assign n14643 = n14642 ^ n14606;
  assign n14644 = n14607 & n14643;
  assign n14645 = n14644 ^ n14605;
  assign n14646 = n14645 ^ n14598;
  assign n14647 = ~n14602 & ~n14646;
  assign n14648 = n14647 ^ n14601;
  assign n14649 = n14648 ^ n14596;
  assign n14650 = ~n14597 & n14649;
  assign n14651 = n14650 ^ n14595;
  assign n14652 = n14651 ^ n14591;
  assign n14653 = n14592 & n14652;
  assign n14654 = n14653 ^ n14590;
  assign n14655 = n14654 ^ n14516;
  assign n14656 = ~n14587 & n14655;
  assign n14657 = n14656 ^ n14586;
  assign n14658 = n14657 ^ n14582;
  assign n14659 = ~n14583 & n14658;
  assign n14660 = n14659 ^ n14581;
  assign n14661 = n14660 ^ n14577;
  assign n14662 = ~n14578 & ~n14661;
  assign n14663 = n14662 ^ n14576;
  assign n14664 = n14663 ^ n14569;
  assign n14665 = ~n14573 & ~n14664;
  assign n14666 = n14665 ^ n14572;
  assign n14667 = n14666 ^ n14567;
  assign n14668 = ~n14568 & ~n14667;
  assign n14669 = n14668 ^ n14566;
  assign n14670 = n14669 ^ n14559;
  assign n14671 = ~n14563 & ~n14670;
  assign n14672 = n14671 ^ n14562;
  assign n14673 = n14672 ^ n14554;
  assign n14674 = ~n14558 & n14673;
  assign n14675 = n14674 ^ n14557;
  assign n14677 = n14676 ^ n14675;
  assign n14678 = n13682 ^ n12371;
  assign n14679 = n13665 & n14678;
  assign n14680 = n14679 ^ n12371;
  assign n14681 = n14680 ^ n14676;
  assign n14682 = n14677 & ~n14681;
  assign n14683 = n14682 ^ n14680;
  assign n14685 = n14684 ^ n14683;
  assign n14686 = n13676 ^ n12370;
  assign n14687 = n13663 & ~n14686;
  assign n14688 = n14687 ^ n12370;
  assign n14689 = n14688 ^ n14683;
  assign n14690 = n14685 & ~n14689;
  assign n14691 = n14690 ^ n14684;
  assign n14550 = n13670 ^ n12363;
  assign n14551 = n13659 & ~n14550;
  assign n14552 = n14551 ^ n12363;
  assign n14549 = n14344 ^ n14250;
  assign n14553 = n14552 ^ n14549;
  assign n14738 = n14691 ^ n14553;
  assign n14739 = n14738 ^ n12385;
  assign n14740 = n14688 ^ n14684;
  assign n14741 = n14740 ^ n14683;
  assign n14742 = n14741 ^ n12391;
  assign n14743 = n14680 ^ n14677;
  assign n14744 = n14743 ^ n12398;
  assign n14745 = n14672 ^ n14558;
  assign n14746 = n14745 ^ n12406;
  assign n14747 = n14669 ^ n14563;
  assign n14748 = n14747 ^ n12412;
  assign n14749 = n14666 ^ n14568;
  assign n14750 = n14749 ^ n12355;
  assign n14751 = n14663 ^ n14572;
  assign n14752 = n14751 ^ n14569;
  assign n14753 = n14752 ^ n12165;
  assign n14754 = n14660 ^ n14578;
  assign n14755 = n14754 ^ n12029;
  assign n14756 = n14657 ^ n14583;
  assign n14757 = n14756 ^ n11556;
  assign n14758 = n14654 ^ n14587;
  assign n14759 = n14758 ^ n11563;
  assign n14760 = n14651 ^ n14592;
  assign n14761 = n14760 ^ n11570;
  assign n14762 = n14648 ^ n14595;
  assign n14763 = n14762 ^ n14596;
  assign n14764 = n14763 ^ n11577;
  assign n14765 = n14645 ^ n14602;
  assign n14766 = n14765 ^ n11584;
  assign n14767 = n14642 ^ n14605;
  assign n14768 = n14767 ^ n14606;
  assign n14769 = n14768 ^ n11591;
  assign n14770 = n14639 ^ n14612;
  assign n14771 = n14770 ^ n11598;
  assign n14772 = n14636 ^ n14617;
  assign n14773 = n14772 ^ n11601;
  assign n14774 = n14633 ^ n14622;
  assign n14775 = n14774 ^ n11607;
  assign n14776 = n14630 ^ n14627;
  assign n14777 = n14776 ^ n11614;
  assign n14508 = n14507 ^ n14502;
  assign n14509 = n14508 ^ n11621;
  assign n14497 = n14453 ^ n14443;
  assign n14498 = n14454 & n14497;
  assign n14499 = n14498 ^ n11627;
  assign n14778 = n14508 ^ n14499;
  assign n14779 = ~n14509 & n14778;
  assign n14780 = n14779 ^ n11621;
  assign n14781 = n14780 ^ n14776;
  assign n14782 = n14777 & ~n14781;
  assign n14783 = n14782 ^ n11614;
  assign n14784 = n14783 ^ n14774;
  assign n14785 = ~n14775 & n14784;
  assign n14786 = n14785 ^ n11607;
  assign n14787 = n14786 ^ n14772;
  assign n14788 = n14773 & ~n14787;
  assign n14789 = n14788 ^ n11601;
  assign n14790 = n14789 ^ n14770;
  assign n14791 = n14771 & ~n14790;
  assign n14792 = n14791 ^ n11598;
  assign n14793 = n14792 ^ n14768;
  assign n14794 = ~n14769 & n14793;
  assign n14795 = n14794 ^ n11591;
  assign n14796 = n14795 ^ n14765;
  assign n14797 = ~n14766 & n14796;
  assign n14798 = n14797 ^ n11584;
  assign n14799 = n14798 ^ n14763;
  assign n14800 = ~n14764 & ~n14799;
  assign n14801 = n14800 ^ n11577;
  assign n14802 = n14801 ^ n14760;
  assign n14803 = ~n14761 & ~n14802;
  assign n14804 = n14803 ^ n11570;
  assign n14805 = n14804 ^ n14758;
  assign n14806 = ~n14759 & n14805;
  assign n14807 = n14806 ^ n11563;
  assign n14808 = n14807 ^ n14756;
  assign n14809 = n14757 & n14808;
  assign n14810 = n14809 ^ n11556;
  assign n14811 = n14810 ^ n14754;
  assign n14812 = ~n14755 & ~n14811;
  assign n14813 = n14812 ^ n12029;
  assign n14814 = n14813 ^ n14752;
  assign n14815 = n14753 & ~n14814;
  assign n14816 = n14815 ^ n12165;
  assign n14817 = n14816 ^ n14749;
  assign n14818 = ~n14750 & n14817;
  assign n14819 = n14818 ^ n12355;
  assign n14820 = n14819 ^ n14747;
  assign n14821 = n14748 & ~n14820;
  assign n14822 = n14821 ^ n12412;
  assign n14823 = n14822 ^ n14745;
  assign n14824 = n14746 & n14823;
  assign n14825 = n14824 ^ n12406;
  assign n14826 = n14825 ^ n14743;
  assign n14827 = ~n14744 & ~n14826;
  assign n14828 = n14827 ^ n12398;
  assign n14829 = n14828 ^ n14741;
  assign n14830 = n14742 & ~n14829;
  assign n14831 = n14830 ^ n12391;
  assign n14832 = n14831 ^ n14738;
  assign n14833 = n14739 & n14832;
  assign n14834 = n14833 ^ n12385;
  assign n14692 = n14691 ^ n14549;
  assign n14693 = ~n14553 & n14692;
  assign n14694 = n14693 ^ n14552;
  assign n14545 = n13219 ^ n12631;
  assign n14546 = ~n13658 & ~n14545;
  assign n14547 = n14546 ^ n12631;
  assign n14736 = n14694 ^ n14547;
  assign n14544 = n14348 ^ n2786;
  assign n14737 = n14736 ^ n14544;
  assign n14835 = n14834 ^ n14737;
  assign n14887 = n14835 ^ n11948;
  assign n14849 = n14831 ^ n14739;
  assign n14850 = n14822 ^ n14746;
  assign n14851 = n14819 ^ n14748;
  assign n14852 = n14816 ^ n14750;
  assign n14853 = n14810 ^ n14755;
  assign n14854 = n14807 ^ n14757;
  assign n14855 = n14804 ^ n14759;
  assign n14856 = n14798 ^ n14764;
  assign n14857 = n14789 ^ n14771;
  assign n14858 = n14780 ^ n14777;
  assign n14510 = n14509 ^ n14499;
  assign n14511 = ~n14455 & ~n14464;
  assign n14859 = ~n14510 & n14511;
  assign n14860 = ~n14858 & ~n14859;
  assign n14861 = n14783 ^ n14775;
  assign n14862 = n14860 & n14861;
  assign n14863 = n14786 ^ n14773;
  assign n14864 = ~n14862 & n14863;
  assign n14865 = n14857 & n14864;
  assign n14866 = n14792 ^ n14769;
  assign n14867 = ~n14865 & n14866;
  assign n14868 = n14795 ^ n14766;
  assign n14869 = n14867 & n14868;
  assign n14870 = n14856 & n14869;
  assign n14871 = n14801 ^ n14761;
  assign n14872 = n14870 & ~n14871;
  assign n14873 = ~n14855 & ~n14872;
  assign n14874 = n14854 & n14873;
  assign n14875 = ~n14853 & ~n14874;
  assign n14876 = n14813 ^ n14753;
  assign n14877 = ~n14875 & n14876;
  assign n14878 = ~n14852 & n14877;
  assign n14879 = n14851 & n14878;
  assign n14880 = n14850 & n14879;
  assign n14881 = n14825 ^ n12398;
  assign n14882 = n14881 ^ n14743;
  assign n14883 = n14880 & n14882;
  assign n14884 = n14828 ^ n14742;
  assign n14885 = ~n14883 & ~n14884;
  assign n14886 = n14849 & ~n14885;
  assign n14915 = n14887 ^ n14886;
  assign n14916 = n14915 ^ n1693;
  assign n14917 = n14885 ^ n14849;
  assign n14918 = n14917 ^ n1683;
  assign n14919 = n14884 ^ n14883;
  assign n14920 = n14919 ^ n1677;
  assign n14922 = n14879 ^ n14850;
  assign n14923 = n14922 ^ n2808;
  assign n14925 = n14877 ^ n14852;
  assign n14926 = n14925 ^ n2689;
  assign n14927 = n14876 ^ n14875;
  assign n14928 = n14927 ^ n1518;
  assign n14931 = n14872 ^ n14855;
  assign n14932 = n14931 ^ n2510;
  assign n14934 = n14869 ^ n14856;
  assign n14935 = n14934 ^ n1395;
  assign n14937 = n14866 ^ n14865;
  assign n1074 = n992 ^ x181;
  assign n1075 = n1074 ^ x373;
  assign n1076 = n1075 ^ x117;
  assign n14938 = n14937 ^ n1076;
  assign n14940 = n14863 ^ n14862;
  assign n14941 = n14940 ^ n851;
  assign n14943 = n14859 ^ n14858;
  assign n14944 = n14943 ^ n744;
  assign n14512 = n14511 ^ n14510;
  assign n14513 = n14512 ^ n653;
  assign n14494 = n14493 ^ n14465;
  assign n14495 = n14466 & ~n14494;
  assign n14496 = n14495 ^ n585;
  assign n14945 = n14512 ^ n14496;
  assign n14946 = ~n14513 & n14945;
  assign n14947 = n14946 ^ n653;
  assign n14948 = n14947 ^ n14943;
  assign n14949 = ~n14944 & n14948;
  assign n14950 = n14949 ^ n744;
  assign n14942 = n14861 ^ n14860;
  assign n14951 = n14950 ^ n14942;
  assign n14952 = n14942 ^ n1043;
  assign n14953 = n14951 & ~n14952;
  assign n14954 = n14953 ^ n1043;
  assign n14955 = n14954 ^ n14940;
  assign n14956 = ~n14941 & n14955;
  assign n14957 = n14956 ^ n851;
  assign n14939 = n14864 ^ n14857;
  assign n14958 = n14957 ^ n14939;
  assign n1056 = n973 ^ x182;
  assign n1057 = n1056 ^ x374;
  assign n1058 = n1057 ^ x118;
  assign n14959 = n14939 ^ n1058;
  assign n14960 = ~n14958 & n14959;
  assign n14961 = n14960 ^ n1058;
  assign n14962 = n14961 ^ n14937;
  assign n14963 = n14938 & ~n14962;
  assign n14964 = n14963 ^ n1076;
  assign n14936 = n14868 ^ n14867;
  assign n14965 = n14964 ^ n14936;
  assign n1205 = n1114 ^ x180;
  assign n1206 = n1205 ^ x372;
  assign n1207 = n1206 ^ x116;
  assign n14966 = n14936 ^ n1207;
  assign n14967 = n14965 & ~n14966;
  assign n14968 = n14967 ^ n1207;
  assign n14969 = n14968 ^ n14934;
  assign n14970 = ~n14935 & n14969;
  assign n14971 = n14970 ^ n1395;
  assign n14933 = n14871 ^ n14870;
  assign n14972 = n14971 ^ n14933;
  assign n14973 = n14933 ^ n1407;
  assign n14974 = ~n14972 & n14973;
  assign n14975 = n14974 ^ n1407;
  assign n14976 = n14975 ^ n14931;
  assign n14977 = n14932 & ~n14976;
  assign n14978 = n14977 ^ n2510;
  assign n14930 = n14873 ^ n14854;
  assign n14979 = n14978 ^ n14930;
  assign n2515 = n2458 ^ x176;
  assign n2516 = n2515 ^ x368;
  assign n2517 = n2516 ^ x112;
  assign n14980 = n14930 ^ n2517;
  assign n14981 = ~n14979 & n14980;
  assign n14982 = n14981 ^ n2517;
  assign n14929 = n14874 ^ n14853;
  assign n14983 = n14982 ^ n14929;
  assign n14984 = n14929 ^ n2529;
  assign n14985 = n14983 & ~n14984;
  assign n14986 = n14985 ^ n2529;
  assign n14987 = n14986 ^ n14927;
  assign n14988 = ~n14928 & n14987;
  assign n14989 = n14988 ^ n1518;
  assign n14990 = n14989 ^ n14925;
  assign n14991 = ~n14926 & n14990;
  assign n14992 = n14991 ^ n2689;
  assign n14924 = n14878 ^ n14851;
  assign n14993 = n14992 ^ n14924;
  assign n14994 = n14924 ^ n1568;
  assign n14995 = ~n14993 & n14994;
  assign n14996 = n14995 ^ n1568;
  assign n14997 = n14996 ^ n14922;
  assign n14998 = n14923 & ~n14997;
  assign n14999 = n14998 ^ n2808;
  assign n14921 = n14882 ^ n14880;
  assign n15000 = n14999 ^ n14921;
  assign n15001 = n14921 ^ n2972;
  assign n15002 = ~n15000 & n15001;
  assign n15003 = n15002 ^ n2972;
  assign n15004 = n15003 ^ n14919;
  assign n15005 = ~n14920 & n15004;
  assign n15006 = n15005 ^ n1677;
  assign n15007 = n15006 ^ n14917;
  assign n15008 = ~n14918 & n15007;
  assign n15009 = n15008 ^ n1683;
  assign n15010 = n15009 ^ n14915;
  assign n15011 = ~n14916 & n15010;
  assign n15012 = n15011 ^ n1693;
  assign n14836 = n14737 ^ n11948;
  assign n14837 = n14835 & ~n14836;
  assign n14838 = n14837 ^ n11948;
  assign n14548 = n14547 ^ n14544;
  assign n14695 = n14694 ^ n14544;
  assign n14696 = n14548 & n14695;
  assign n14697 = n14696 ^ n14547;
  assign n14540 = n13214 ^ n12625;
  assign n14541 = n13655 & ~n14540;
  assign n14542 = n14541 ^ n12625;
  assign n14733 = n14697 ^ n14542;
  assign n14539 = n14351 ^ n14247;
  assign n14734 = n14733 ^ n14539;
  assign n14735 = n14734 ^ n11945;
  assign n14889 = n14838 ^ n14735;
  assign n14888 = ~n14886 & ~n14887;
  assign n14914 = n14889 ^ n14888;
  assign n15013 = n15012 ^ n14914;
  assign n15014 = n14914 ^ n1760;
  assign n15015 = ~n15013 & n15014;
  assign n15016 = n15015 ^ n1760;
  assign n14839 = n14838 ^ n14734;
  assign n14840 = n14735 & n14839;
  assign n14841 = n14840 ^ n11945;
  assign n14543 = n14542 ^ n14539;
  assign n14698 = n14697 ^ n14539;
  assign n14699 = ~n14543 & ~n14698;
  assign n14700 = n14699 ^ n14542;
  assign n14535 = n13231 ^ n12623;
  assign n14536 = n13881 & ~n14535;
  assign n14537 = n14536 ^ n12623;
  assign n14730 = n14700 ^ n14537;
  assign n14534 = n14355 ^ n1537;
  assign n14731 = n14730 ^ n14534;
  assign n14732 = n14731 ^ n11939;
  assign n14891 = n14841 ^ n14732;
  assign n14890 = ~n14888 & ~n14889;
  assign n14913 = n14891 ^ n14890;
  assign n15017 = n15016 ^ n14913;
  assign n15036 = n15017 ^ n1874;
  assign n15037 = n14451 ^ n13197;
  assign n15038 = n15037 ^ n13773;
  assign n15039 = ~n15036 & n15038;
  assign n15042 = n15041 ^ n15039;
  assign n15018 = n14913 ^ n1874;
  assign n15019 = n15017 & ~n15018;
  assign n15020 = n15019 ^ n1874;
  assign n14842 = n14841 ^ n14731;
  assign n14843 = n14732 & n14842;
  assign n14844 = n14843 ^ n11939;
  assign n14538 = n14537 ^ n14534;
  assign n14701 = n14700 ^ n14534;
  assign n14702 = ~n14538 & ~n14701;
  assign n14703 = n14702 ^ n14537;
  assign n14529 = n13209 ^ n12614;
  assign n14530 = n13873 & n14529;
  assign n14531 = n14530 ^ n12614;
  assign n14727 = n14703 ^ n14531;
  assign n14532 = n14358 ^ n14244;
  assign n14728 = n14727 ^ n14532;
  assign n14729 = n14728 ^ n11961;
  assign n14893 = n14844 ^ n14729;
  assign n14892 = ~n14890 & ~n14891;
  assign n14912 = n14893 ^ n14892;
  assign n15021 = n15020 ^ n14912;
  assign n15043 = n15021 ^ n1871;
  assign n15044 = n15043 ^ n15041;
  assign n15045 = n15042 & n15044;
  assign n15046 = n15045 ^ n15039;
  assign n15022 = n14912 ^ n1871;
  assign n15023 = n15021 & ~n15022;
  assign n15024 = n15023 ^ n1871;
  assign n14894 = n14892 & n14893;
  assign n14845 = n14844 ^ n14728;
  assign n14846 = n14729 & ~n14845;
  assign n14847 = n14846 ^ n11961;
  assign n14709 = n13110 ^ n12608;
  assign n14710 = ~n13868 & n14709;
  assign n14711 = n14710 ^ n12608;
  assign n14707 = n14361 ^ n14242;
  assign n14533 = n14532 ^ n14531;
  assign n14704 = n14703 ^ n14532;
  assign n14705 = n14533 & ~n14704;
  assign n14706 = n14705 ^ n14531;
  assign n14708 = n14707 ^ n14706;
  assign n14725 = n14711 ^ n14708;
  assign n14726 = n14725 ^ n11927;
  assign n14848 = n14847 ^ n14726;
  assign n14910 = n14894 ^ n14848;
  assign n14911 = n14910 ^ n2036;
  assign n15035 = n15024 ^ n14911;
  assign n15047 = n15046 ^ n15035;
  assign n15048 = n13763 ^ n13184;
  assign n15049 = n15048 ^ n14626;
  assign n15050 = n15049 ^ n15035;
  assign n15051 = ~n15047 & ~n15050;
  assign n15052 = n15051 ^ n15049;
  assign n15025 = n15024 ^ n14910;
  assign n15026 = n14911 & ~n15025;
  assign n15027 = n15026 ^ n2036;
  assign n14897 = n14847 ^ n14725;
  assign n14898 = n14726 & ~n14897;
  assign n14899 = n14898 ^ n11927;
  assign n14900 = n14899 ^ n11667;
  assign n14717 = n13203 ^ n12507;
  assign n14718 = n13863 & ~n14717;
  assign n14719 = n14718 ^ n12507;
  assign n14715 = n14364 ^ n14240;
  assign n14712 = n14711 ^ n14707;
  assign n14713 = n14708 & n14712;
  assign n14714 = n14713 ^ n14711;
  assign n14716 = n14715 ^ n14714;
  assign n14896 = n14719 ^ n14716;
  assign n14901 = n14900 ^ n14896;
  assign n14895 = ~n14848 & ~n14894;
  assign n14909 = n14901 ^ n14895;
  assign n15028 = n15027 ^ n14909;
  assign n15034 = n15028 ^ n681;
  assign n15053 = n15052 ^ n15034;
  assign n15054 = n13755 ^ n13179;
  assign n15055 = n15054 ^ n14618;
  assign n15056 = n15055 ^ n15034;
  assign n15057 = n15053 & n15056;
  assign n15058 = n15057 ^ n15055;
  assign n15029 = n14909 ^ n681;
  assign n15030 = ~n15028 & n15029;
  assign n15031 = n15030 ^ n681;
  assign n2223 = n2129 ^ x161;
  assign n2224 = n2223 ^ x353;
  assign n2225 = n2224 ^ x97;
  assign n15032 = n15031 ^ n2225;
  assign n14904 = n14896 ^ n11667;
  assign n14905 = n14899 ^ n14896;
  assign n14906 = n14904 & ~n14905;
  assign n14907 = n14906 ^ n11667;
  assign n14902 = ~n14895 & n14901;
  assign n14720 = n14719 ^ n14715;
  assign n14721 = n14716 & ~n14720;
  assign n14722 = n14721 ^ n14719;
  assign n14723 = n14722 ^ n11662;
  assign n14525 = n13199 ^ n12502;
  assign n14526 = n13913 & n14525;
  assign n14527 = n14526 ^ n12502;
  assign n14524 = n14368 ^ n1996;
  assign n14528 = n14527 ^ n14524;
  assign n14724 = n14723 ^ n14528;
  assign n14903 = n14902 ^ n14724;
  assign n14908 = n14907 ^ n14903;
  assign n15033 = n15032 ^ n14908;
  assign n15059 = n15058 ^ n15033;
  assign n15060 = n13753 ^ n13263;
  assign n15061 = n15060 ^ n14613;
  assign n15062 = n15061 ^ n15033;
  assign n15063 = n15059 & ~n15062;
  assign n15064 = n15063 ^ n15061;
  assign n15066 = n15065 ^ n15064;
  assign n15067 = n13748 ^ n13174;
  assign n15068 = n15067 ^ n14611;
  assign n15069 = n15068 ^ n15065;
  assign n15070 = n15066 & n15069;
  assign n15071 = n15070 ^ n15068;
  assign n14523 = n14480 ^ n14479;
  assign n15072 = n15071 ^ n14523;
  assign n15073 = n13740 ^ n13169;
  assign n15074 = n15073 ^ n14606;
  assign n15075 = n15074 ^ n14523;
  assign n15076 = ~n15072 & n15075;
  assign n15077 = n15076 ^ n15074;
  assign n14522 = n14483 ^ n14471;
  assign n15078 = n15077 ^ n14522;
  assign n15079 = n13735 ^ n13164;
  assign n15080 = n15079 ^ n14598;
  assign n15081 = n15080 ^ n14522;
  assign n15082 = ~n15078 & ~n15081;
  assign n15083 = n15082 ^ n15080;
  assign n14521 = n14487 ^ n556;
  assign n15084 = n15083 ^ n14521;
  assign n15085 = n13733 ^ n13159;
  assign n15086 = n15085 ^ n14596;
  assign n15087 = n15086 ^ n14521;
  assign n15088 = n15084 & ~n15087;
  assign n15089 = n15088 ^ n15086;
  assign n14520 = n14490 ^ n14468;
  assign n15090 = n15089 ^ n14520;
  assign n15091 = n13725 ^ n13154;
  assign n15092 = n15091 ^ n14591;
  assign n15093 = n15092 ^ n14520;
  assign n15094 = n15090 & n15093;
  assign n15095 = n15094 ^ n15092;
  assign n15096 = n15095 ^ n14518;
  assign n15097 = ~n14519 & n15096;
  assign n15098 = n15097 ^ n14517;
  assign n14514 = n14513 ^ n14496;
  assign n15099 = n15098 ^ n14514;
  assign n15111 = n15101 ^ n15099;
  assign n15112 = n15111 ^ n12439;
  assign n15113 = n15095 ^ n14519;
  assign n15114 = n15113 ^ n12444;
  assign n15115 = n15092 ^ n15090;
  assign n15116 = n15115 ^ n12447;
  assign n15117 = n15086 ^ n15084;
  assign n15118 = n15117 ^ n12455;
  assign n15119 = n15080 ^ n15078;
  assign n15120 = n15119 ^ n12460;
  assign n15121 = n15074 ^ n15072;
  assign n15122 = n15121 ^ n12466;
  assign n15123 = n15068 ^ n15066;
  assign n15124 = n15123 ^ n12472;
  assign n15125 = n15061 ^ n15059;
  assign n15126 = n15125 ^ n12474;
  assign n15127 = n15055 ^ n15053;
  assign n15128 = n15127 ^ n12480;
  assign n15129 = n15049 ^ n15047;
  assign n15130 = n15129 ^ n12488;
  assign n15131 = n15038 ^ n15036;
  assign n15132 = ~n12500 & ~n15131;
  assign n15133 = n15132 ^ n12494;
  assign n15134 = n15043 ^ n15042;
  assign n15135 = n15134 ^ n15132;
  assign n15136 = n15133 & n15135;
  assign n15137 = n15136 ^ n12494;
  assign n15138 = n15137 ^ n15129;
  assign n15139 = n15130 & n15138;
  assign n15140 = n15139 ^ n12488;
  assign n15141 = n15140 ^ n15127;
  assign n15142 = ~n15128 & ~n15141;
  assign n15143 = n15142 ^ n12480;
  assign n15144 = n15143 ^ n15125;
  assign n15145 = ~n15126 & n15144;
  assign n15146 = n15145 ^ n12474;
  assign n15147 = n15146 ^ n15123;
  assign n15148 = n15124 & ~n15147;
  assign n15149 = n15148 ^ n12472;
  assign n15150 = n15149 ^ n15121;
  assign n15151 = ~n15122 & n15150;
  assign n15152 = n15151 ^ n12466;
  assign n15153 = n15152 ^ n15119;
  assign n15154 = ~n15120 & ~n15153;
  assign n15155 = n15154 ^ n12460;
  assign n15156 = n15155 ^ n15117;
  assign n15157 = n15118 & ~n15156;
  assign n15158 = n15157 ^ n12455;
  assign n15159 = n15158 ^ n15115;
  assign n15160 = ~n15116 & n15159;
  assign n15161 = n15160 ^ n12447;
  assign n15162 = n15161 ^ n15113;
  assign n15163 = ~n15114 & n15162;
  assign n15164 = n15163 ^ n12444;
  assign n15165 = n15164 ^ n15111;
  assign n15166 = n15112 & n15165;
  assign n15167 = n15166 ^ n12439;
  assign n15106 = n13713 ^ n13139;
  assign n15107 = n15106 ^ n14577;
  assign n15105 = n14947 ^ n14944;
  assign n15108 = n15107 ^ n15105;
  assign n15102 = n15101 ^ n14514;
  assign n15103 = ~n15099 & ~n15102;
  assign n15104 = n15103 ^ n15101;
  assign n15109 = n15108 ^ n15104;
  assign n15110 = n15109 ^ n12433;
  assign n15181 = n15167 ^ n15110;
  assign n15182 = n15164 ^ n15112;
  assign n15183 = n15149 ^ n15122;
  assign n15184 = n15140 ^ n15128;
  assign n15185 = n15137 ^ n15130;
  assign n15186 = n15131 ^ n12500;
  assign n15187 = n15134 ^ n15133;
  assign n15188 = n15186 & ~n15187;
  assign n15189 = n15185 & n15188;
  assign n15190 = n15184 & n15189;
  assign n15191 = n15143 ^ n15126;
  assign n15192 = n15190 & ~n15191;
  assign n15193 = n15146 ^ n15124;
  assign n15194 = ~n15192 & ~n15193;
  assign n15195 = ~n15183 & ~n15194;
  assign n15196 = n15152 ^ n15120;
  assign n15197 = ~n15195 & n15196;
  assign n15198 = n15155 ^ n15118;
  assign n15199 = n15197 & n15198;
  assign n15200 = n15158 ^ n15116;
  assign n15201 = n15199 & ~n15200;
  assign n15202 = n15161 ^ n15114;
  assign n15203 = ~n15201 & n15202;
  assign n15204 = n15182 & ~n15203;
  assign n15205 = n15181 & ~n15204;
  assign n15174 = n15105 ^ n15104;
  assign n15175 = ~n15108 & n15174;
  assign n15176 = n15175 ^ n15107;
  assign n15173 = n14951 ^ n1043;
  assign n15177 = n15176 ^ n15173;
  assign n15171 = n13708 ^ n13134;
  assign n15172 = n15171 ^ n14569;
  assign n15178 = n15177 ^ n15172;
  assign n15179 = n15178 ^ n12428;
  assign n15168 = n15167 ^ n15109;
  assign n15169 = n15110 & n15168;
  assign n15170 = n15169 ^ n12433;
  assign n15180 = n15179 ^ n15170;
  assign n15221 = n15205 ^ n15180;
  assign n1266 = n1172 ^ x211;
  assign n1267 = n1266 ^ x403;
  assign n1268 = n1267 ^ x147;
  assign n15222 = n15221 ^ n1268;
  assign n15223 = n15204 ^ n15181;
  assign n1342 = n1236 ^ x212;
  assign n1343 = n1342 ^ x404;
  assign n1344 = n1343 ^ x148;
  assign n15224 = n15223 ^ n1344;
  assign n15225 = n15203 ^ n15182;
  assign n1081 = n999 ^ x213;
  assign n1082 = n1081 ^ x405;
  assign n1083 = n1082 ^ x149;
  assign n15226 = n15225 ^ n1083;
  assign n15228 = n15200 ^ n15199;
  assign n15229 = n15228 ^ n922;
  assign n15231 = n15196 ^ n15195;
  assign n15232 = n15231 ^ n667;
  assign n15233 = n15194 ^ n15183;
  assign n15234 = n15233 ^ n626;
  assign n15236 = n15191 ^ n15190;
  assign n15237 = n15236 ^ n3258;
  assign n15238 = n15189 ^ n15184;
  assign n15242 = n15241 ^ n15238;
  assign n15243 = n15188 ^ n15185;
  assign n15244 = n15243 ^ n675;
  assign n15245 = n521 & ~n15186;
  assign n15249 = n15248 ^ n15245;
  assign n15250 = n15187 ^ n15186;
  assign n15251 = n15250 ^ n15245;
  assign n15252 = n15249 & n15251;
  assign n15253 = n15252 ^ n15248;
  assign n15254 = n15253 ^ n15243;
  assign n15255 = n15244 & ~n15254;
  assign n15256 = n15255 ^ n675;
  assign n15257 = n15256 ^ n15238;
  assign n15258 = n15242 & ~n15257;
  assign n15259 = n15258 ^ n15241;
  assign n15260 = n15259 ^ n15236;
  assign n15261 = ~n15237 & n15260;
  assign n15262 = n15261 ^ n3258;
  assign n15235 = n15193 ^ n15192;
  assign n15263 = n15262 ^ n15235;
  assign n15264 = n15235 ^ n620;
  assign n15265 = n15263 & ~n15264;
  assign n15266 = n15265 ^ n620;
  assign n15267 = n15266 ^ n15233;
  assign n15268 = n15234 & ~n15267;
  assign n15269 = n15268 ^ n626;
  assign n15270 = n15269 ^ n15231;
  assign n15271 = n15232 & ~n15270;
  assign n15272 = n15271 ^ n667;
  assign n15230 = n15198 ^ n15197;
  assign n15273 = n15272 ^ n15230;
  assign n15274 = n15230 ^ n806;
  assign n15275 = n15273 & ~n15274;
  assign n15276 = n15275 ^ n806;
  assign n15277 = n15276 ^ n15228;
  assign n15278 = n15229 & ~n15277;
  assign n15279 = n15278 ^ n922;
  assign n15227 = n15202 ^ n15201;
  assign n15280 = n15279 ^ n15227;
  assign n15281 = n15227 ^ n928;
  assign n15282 = n15280 & ~n15281;
  assign n15283 = n15282 ^ n928;
  assign n15284 = n15283 ^ n15225;
  assign n15285 = n15226 & ~n15284;
  assign n15286 = n15285 ^ n1083;
  assign n15287 = n15286 ^ n15223;
  assign n15288 = ~n15224 & n15287;
  assign n15289 = n15288 ^ n1344;
  assign n15290 = n15289 ^ n15221;
  assign n15291 = n15222 & ~n15290;
  assign n15292 = n15291 ^ n1268;
  assign n15214 = n14567 ^ n13132;
  assign n15215 = n15214 ^ n13703;
  assign n15213 = n14954 ^ n14941;
  assign n15216 = n15215 ^ n15213;
  assign n15210 = n15173 ^ n15172;
  assign n15211 = n15177 & ~n15210;
  assign n15212 = n15211 ^ n15172;
  assign n15217 = n15216 ^ n15212;
  assign n15218 = n15217 ^ n12422;
  assign n15207 = n15178 ^ n15170;
  assign n15208 = n15179 & ~n15207;
  assign n15209 = n15208 ^ n12428;
  assign n15219 = n15218 ^ n15209;
  assign n15206 = n15180 & ~n15205;
  assign n15220 = n15219 ^ n15206;
  assign n15293 = n15292 ^ n15220;
  assign n2410 = n1418 ^ x210;
  assign n2411 = n2410 ^ x402;
  assign n2412 = n2411 ^ x146;
  assign n15602 = n15220 ^ n2412;
  assign n15603 = ~n15293 & n15602;
  assign n15604 = n15603 ^ n2412;
  assign n15472 = n15217 ^ n15209;
  assign n15473 = ~n15218 & ~n15472;
  assign n15474 = n15473 ^ n12422;
  assign n15369 = n13698 ^ n13127;
  assign n15370 = n15369 ^ n14559;
  assign n15365 = n15213 ^ n15212;
  assign n15366 = ~n15216 & n15365;
  assign n15367 = n15366 ^ n15215;
  assign n15325 = n14958 ^ n1058;
  assign n15368 = n15367 ^ n15325;
  assign n15470 = n15370 ^ n15368;
  assign n15471 = n15470 ^ n12417;
  assign n15527 = n15474 ^ n15471;
  assign n15526 = n15206 & ~n15219;
  assign n15600 = n15527 ^ n15526;
  assign n15601 = n15600 ^ n3026;
  assign n15761 = n15604 ^ n15601;
  assign n15296 = n14989 ^ n14926;
  assign n15295 = n14539 ^ n13674;
  assign n15297 = n15296 ^ n15295;
  assign n15294 = n15293 ^ n2412;
  assign n15298 = n15297 ^ n15294;
  assign n15303 = n15286 ^ n15224;
  assign n15301 = n14983 ^ n2529;
  assign n15300 = n14549 ^ n13686;
  assign n15302 = n15301 ^ n15300;
  assign n15304 = n15303 ^ n15302;
  assign n15307 = n14979 ^ n2517;
  assign n15306 = n14684 ^ n13692;
  assign n15308 = n15307 ^ n15306;
  assign n15305 = n15283 ^ n15226;
  assign n15309 = n15308 ^ n15305;
  assign n15314 = n15276 ^ n15229;
  assign n15312 = n14972 ^ n1407;
  assign n15311 = n14554 ^ n13703;
  assign n15313 = n15312 ^ n15311;
  assign n15315 = n15314 ^ n15313;
  assign n15320 = n15269 ^ n15232;
  assign n15318 = n14965 ^ n1207;
  assign n15317 = n14567 ^ n13713;
  assign n15319 = n15318 ^ n15317;
  assign n15321 = n15320 ^ n15319;
  assign n15324 = n14577 ^ n13720;
  assign n15326 = n15325 ^ n15324;
  assign n15323 = n15263 ^ n620;
  assign n15327 = n15326 ^ n15323;
  assign n15332 = n15256 ^ n15242;
  assign n15330 = n14516 ^ n13733;
  assign n15331 = n15330 ^ n15173;
  assign n15333 = n15332 ^ n15331;
  assign n15337 = n15250 ^ n15249;
  assign n15335 = n14596 ^ n13740;
  assign n15336 = n15335 ^ n14514;
  assign n15338 = n15337 ^ n15336;
  assign n15439 = n13913 ^ n13110;
  assign n15440 = n15439 ^ n14397;
  assign n15437 = n15006 ^ n14918;
  assign n15424 = n15000 ^ n2972;
  assign n15417 = n14996 ^ n14923;
  assign n15398 = n14986 ^ n14928;
  assign n15344 = n13682 ^ n13659;
  assign n15345 = n15344 ^ n14534;
  assign n15346 = n15345 ^ n15301;
  assign n15347 = n13688 ^ n13663;
  assign n15348 = n15347 ^ n14539;
  assign n15349 = n15348 ^ n15307;
  assign n15351 = n13694 ^ n13665;
  assign n15352 = n15351 ^ n14544;
  assign n15350 = n14975 ^ n14932;
  assign n15353 = n15352 ^ n15350;
  assign n15354 = n13674 ^ n13464;
  assign n15355 = n15354 ^ n14549;
  assign n15356 = n15355 ^ n15312;
  assign n15358 = n13686 ^ n13117;
  assign n15359 = n15358 ^ n14676;
  assign n15360 = n15359 ^ n15318;
  assign n15363 = n14961 ^ n14938;
  assign n15361 = n13692 ^ n13122;
  assign n15362 = n15361 ^ n14554;
  assign n15364 = n15363 ^ n15362;
  assign n15371 = n15370 ^ n15325;
  assign n15372 = ~n15368 & n15371;
  assign n15373 = n15372 ^ n15370;
  assign n15374 = n15373 ^ n15363;
  assign n15375 = n15364 & ~n15374;
  assign n15376 = n15375 ^ n15362;
  assign n15377 = n15376 ^ n15318;
  assign n15378 = n15360 & n15377;
  assign n15379 = n15378 ^ n15359;
  assign n15357 = n14968 ^ n14935;
  assign n15380 = n15379 ^ n15357;
  assign n15381 = n13680 ^ n13314;
  assign n15382 = n15381 ^ n14684;
  assign n15383 = n15382 ^ n15357;
  assign n15384 = ~n15380 & n15383;
  assign n15385 = n15384 ^ n15382;
  assign n15386 = n15385 ^ n15312;
  assign n15387 = n15356 & n15386;
  assign n15388 = n15387 ^ n15355;
  assign n15389 = n15388 ^ n15350;
  assign n15390 = ~n15353 & ~n15389;
  assign n15391 = n15390 ^ n15352;
  assign n15392 = n15391 ^ n15307;
  assign n15393 = ~n15349 & n15392;
  assign n15394 = n15393 ^ n15348;
  assign n15395 = n15394 ^ n15345;
  assign n15396 = ~n15346 & n15395;
  assign n15397 = n15396 ^ n15301;
  assign n15399 = n15398 ^ n15397;
  assign n15400 = n13676 ^ n13658;
  assign n15401 = n15400 ^ n14532;
  assign n15402 = n15401 ^ n15398;
  assign n15403 = ~n15399 & n15402;
  assign n15404 = n15403 ^ n15401;
  assign n15405 = n15404 ^ n15296;
  assign n15406 = n13670 ^ n13655;
  assign n15407 = n15406 ^ n14707;
  assign n15408 = n15407 ^ n15296;
  assign n15409 = ~n15405 & n15408;
  assign n15410 = n15409 ^ n15407;
  assign n15343 = n14993 ^ n1568;
  assign n15411 = n15410 ^ n15343;
  assign n15412 = n13881 ^ n13219;
  assign n15413 = n15412 ^ n14715;
  assign n15414 = n15413 ^ n15343;
  assign n15415 = n15411 & ~n15414;
  assign n15416 = n15415 ^ n15413;
  assign n15418 = n15417 ^ n15416;
  assign n15419 = n13873 ^ n13214;
  assign n15420 = n15419 ^ n14524;
  assign n15421 = n15420 ^ n15417;
  assign n15422 = n15418 & n15421;
  assign n15423 = n15422 ^ n15420;
  assign n15425 = n15424 ^ n15423;
  assign n15426 = n13868 ^ n13231;
  assign n15427 = n15426 ^ n14407;
  assign n15428 = n15427 ^ n15424;
  assign n15429 = ~n15425 & ~n15428;
  assign n15430 = n15429 ^ n15427;
  assign n15342 = n15003 ^ n14920;
  assign n15431 = n15430 ^ n15342;
  assign n15432 = n13863 ^ n13209;
  assign n15433 = n15432 ^ n14405;
  assign n15434 = n15433 ^ n15342;
  assign n15435 = ~n15431 & ~n15434;
  assign n15436 = n15435 ^ n15433;
  assign n15438 = n15437 ^ n15436;
  assign n15441 = n15440 ^ n15438;
  assign n15442 = n15441 ^ n12608;
  assign n15443 = n15433 ^ n15431;
  assign n15444 = n15443 ^ n12614;
  assign n15445 = n15427 ^ n15425;
  assign n15446 = n15445 ^ n12623;
  assign n15447 = n15420 ^ n15418;
  assign n15448 = n15447 ^ n12625;
  assign n15449 = n15413 ^ n15411;
  assign n15450 = n15449 ^ n12631;
  assign n15451 = n15407 ^ n15405;
  assign n15452 = n15451 ^ n12363;
  assign n15453 = n15401 ^ n15399;
  assign n15454 = n15453 ^ n12370;
  assign n15455 = n15394 ^ n15346;
  assign n15456 = n15455 ^ n12371;
  assign n15457 = n15391 ^ n15349;
  assign n15458 = n15457 ^ n12373;
  assign n15459 = n15388 ^ n15352;
  assign n15460 = n15459 ^ n15350;
  assign n15461 = n15460 ^ n12378;
  assign n15462 = n15385 ^ n15356;
  assign n15463 = n15462 ^ n12384;
  assign n15464 = n15382 ^ n15380;
  assign n15465 = n15464 ^ n12396;
  assign n15466 = n15376 ^ n15360;
  assign n15467 = n15466 ^ n12403;
  assign n15468 = n15373 ^ n15364;
  assign n15469 = n15468 ^ n12410;
  assign n15475 = n15474 ^ n15470;
  assign n15476 = n15471 & ~n15475;
  assign n15477 = n15476 ^ n12417;
  assign n15478 = n15477 ^ n15468;
  assign n15479 = n15469 & ~n15478;
  assign n15480 = n15479 ^ n12410;
  assign n15481 = n15480 ^ n15466;
  assign n15482 = ~n15467 & ~n15481;
  assign n15483 = n15482 ^ n12403;
  assign n15484 = n15483 ^ n15464;
  assign n15485 = ~n15465 & ~n15484;
  assign n15486 = n15485 ^ n12396;
  assign n15487 = n15486 ^ n15462;
  assign n15488 = n15463 & n15487;
  assign n15489 = n15488 ^ n12384;
  assign n15490 = n15489 ^ n15460;
  assign n15491 = ~n15461 & ~n15490;
  assign n15492 = n15491 ^ n12378;
  assign n15493 = n15492 ^ n15457;
  assign n15494 = n15458 & ~n15493;
  assign n15495 = n15494 ^ n12373;
  assign n15496 = n15495 ^ n15455;
  assign n15497 = n15456 & ~n15496;
  assign n15498 = n15497 ^ n12371;
  assign n15499 = n15498 ^ n15453;
  assign n15500 = ~n15454 & n15499;
  assign n15501 = n15500 ^ n12370;
  assign n15502 = n15501 ^ n15451;
  assign n15503 = ~n15452 & n15502;
  assign n15504 = n15503 ^ n12363;
  assign n15505 = n15504 ^ n15449;
  assign n15506 = ~n15450 & ~n15505;
  assign n15507 = n15506 ^ n12631;
  assign n15508 = n15507 ^ n15447;
  assign n15509 = ~n15448 & ~n15508;
  assign n15510 = n15509 ^ n12625;
  assign n15511 = n15510 ^ n15445;
  assign n15512 = n15446 & n15511;
  assign n15513 = n15512 ^ n12623;
  assign n15514 = n15513 ^ n15443;
  assign n15515 = ~n15444 & n15514;
  assign n15516 = n15515 ^ n12614;
  assign n15556 = n15516 ^ n15441;
  assign n15557 = ~n15442 & ~n15556;
  assign n15558 = n15557 ^ n12608;
  assign n15559 = n15558 ^ n12507;
  assign n15553 = n15009 ^ n14916;
  assign n15550 = n15440 ^ n15437;
  assign n15551 = n15438 & ~n15550;
  assign n15552 = n15551 ^ n15440;
  assign n15554 = n15553 ^ n15552;
  assign n15548 = n13776 ^ n13203;
  assign n15549 = n15548 ^ n14392;
  assign n15555 = n15554 ^ n15549;
  assign n15560 = n15559 ^ n15555;
  assign n15517 = n15516 ^ n15442;
  assign n15518 = n15513 ^ n15444;
  assign n15519 = n15510 ^ n15446;
  assign n15520 = n15501 ^ n15452;
  assign n15521 = n15498 ^ n15454;
  assign n15522 = n15495 ^ n15456;
  assign n15523 = n15489 ^ n15461;
  assign n15524 = n15480 ^ n15467;
  assign n15525 = n15477 ^ n15469;
  assign n15528 = n15526 & ~n15527;
  assign n15529 = ~n15525 & n15528;
  assign n15530 = ~n15524 & ~n15529;
  assign n15531 = n15483 ^ n15465;
  assign n15532 = n15530 & n15531;
  assign n15533 = n15486 ^ n15463;
  assign n15534 = ~n15532 & ~n15533;
  assign n15535 = ~n15523 & n15534;
  assign n15536 = n15492 ^ n15458;
  assign n15537 = ~n15535 & n15536;
  assign n15538 = ~n15522 & ~n15537;
  assign n15539 = n15521 & n15538;
  assign n15540 = ~n15520 & ~n15539;
  assign n15541 = n15504 ^ n15450;
  assign n15542 = ~n15540 & n15541;
  assign n15543 = n15507 ^ n15448;
  assign n15544 = n15542 & ~n15543;
  assign n15545 = ~n15519 & n15544;
  assign n15546 = n15518 & ~n15545;
  assign n15547 = ~n15517 & ~n15546;
  assign n15577 = n15560 ^ n15547;
  assign n15578 = n15577 ^ n2115;
  assign n15583 = n15541 ^ n15540;
  assign n15584 = n15583 ^ n1845;
  assign n15585 = n15539 ^ n15520;
  assign n15586 = n15585 ^ n1616;
  assign n15588 = n15537 ^ n15522;
  assign n15589 = n15588 ^ n1532;
  assign n15591 = n15534 ^ n15523;
  assign n15592 = n15591 ^ n1493;
  assign n15594 = n15531 ^ n15530;
  assign n15595 = n15594 ^ n2651;
  assign n15596 = n15529 ^ n15524;
  assign n15597 = n15596 ^ n2654;
  assign n15598 = n15528 ^ n15525;
  assign n15599 = n15598 ^ n2488;
  assign n15605 = n15604 ^ n15600;
  assign n15606 = n15601 & ~n15605;
  assign n15607 = n15606 ^ n3026;
  assign n15608 = n15607 ^ n15598;
  assign n15609 = n15599 & ~n15608;
  assign n15610 = n15609 ^ n2488;
  assign n15611 = n15610 ^ n15596;
  assign n15612 = n15597 & ~n15611;
  assign n15613 = n15612 ^ n2654;
  assign n15614 = n15613 ^ n15594;
  assign n15615 = n15595 & ~n15614;
  assign n15616 = n15615 ^ n2651;
  assign n15593 = n15533 ^ n15532;
  assign n15617 = n15616 ^ n15593;
  assign n15618 = n15593 ^ n2671;
  assign n15619 = n15617 & ~n15618;
  assign n15620 = n15619 ^ n2671;
  assign n15621 = n15620 ^ n15591;
  assign n15622 = n15592 & ~n15621;
  assign n15623 = n15622 ^ n1493;
  assign n15590 = n15536 ^ n15535;
  assign n15624 = n15623 ^ n15590;
  assign n15625 = n15590 ^ n1582;
  assign n15626 = n15624 & ~n15625;
  assign n15627 = n15626 ^ n1582;
  assign n15628 = n15627 ^ n15588;
  assign n15629 = ~n15589 & n15628;
  assign n15630 = n15629 ^ n1532;
  assign n15587 = n15538 ^ n15521;
  assign n15631 = n15630 ^ n15587;
  assign n15635 = n15634 ^ n15587;
  assign n15636 = n15631 & ~n15635;
  assign n15637 = n15636 ^ n15634;
  assign n15638 = n15637 ^ n15585;
  assign n15639 = n15586 & ~n15638;
  assign n15640 = n15639 ^ n1616;
  assign n15641 = n15640 ^ n15583;
  assign n15642 = n15584 & ~n15641;
  assign n15643 = n15642 ^ n1845;
  assign n15582 = n15543 ^ n15542;
  assign n15644 = n15643 ^ n15582;
  assign n15645 = n15582 ^ n1838;
  assign n15646 = ~n15644 & n15645;
  assign n15647 = n15646 ^ n1838;
  assign n15581 = n15544 ^ n15519;
  assign n15648 = n15647 ^ n15581;
  assign n15649 = n15581 ^ n1858;
  assign n15650 = ~n15648 & n15649;
  assign n15651 = n15650 ^ n1858;
  assign n15580 = n15545 ^ n15518;
  assign n15652 = n15651 ^ n15580;
  assign n15653 = n15580 ^ n1964;
  assign n15654 = n15652 & ~n15653;
  assign n15655 = n15654 ^ n1964;
  assign n15579 = n15546 ^ n15517;
  assign n15656 = n15655 ^ n15579;
  assign n15657 = n15579 ^ n1970;
  assign n15658 = n15656 & ~n15657;
  assign n15659 = n15658 ^ n1970;
  assign n15660 = n15659 ^ n15577;
  assign n15661 = ~n15578 & n15660;
  assign n15662 = n15661 ^ n2115;
  assign n15663 = n15662 ^ n2315;
  assign n15570 = n15555 ^ n12507;
  assign n15571 = n15558 ^ n15555;
  assign n15572 = ~n15570 & n15571;
  assign n15573 = n15572 ^ n12507;
  assign n15574 = n15573 ^ n12502;
  assign n15568 = n15013 ^ n1760;
  assign n15564 = n15553 ^ n15549;
  assign n15565 = n15554 & ~n15564;
  assign n15566 = n15565 ^ n15549;
  assign n15562 = n13775 ^ n13199;
  assign n15563 = n15562 ^ n14387;
  assign n15567 = n15566 ^ n15563;
  assign n15569 = n15568 ^ n15567;
  assign n15575 = n15574 ^ n15569;
  assign n15561 = n15547 & n15560;
  assign n15576 = n15575 ^ n15561;
  assign n15664 = n15663 ^ n15576;
  assign n15340 = n14606 ^ n13753;
  assign n15341 = n15340 ^ n14520;
  assign n15665 = n15664 ^ n15341;
  assign n15673 = n14618 ^ n13768;
  assign n15674 = n15673 ^ n14523;
  assign n15669 = n15648 ^ n1858;
  assign n15670 = n14626 ^ n13773;
  assign n15671 = n15670 ^ n15065;
  assign n15672 = n15669 & n15671;
  assign n15675 = n15674 ^ n15672;
  assign n15676 = n15652 ^ n1964;
  assign n15677 = n15676 ^ n15674;
  assign n15678 = ~n15675 & ~n15677;
  assign n15679 = n15678 ^ n15672;
  assign n15668 = n15656 ^ n1970;
  assign n15680 = n15679 ^ n15668;
  assign n15681 = n14522 ^ n13763;
  assign n15682 = n15681 ^ n14613;
  assign n15683 = n15682 ^ n15668;
  assign n15684 = n15680 & n15683;
  assign n15685 = n15684 ^ n15682;
  assign n15666 = n15659 ^ n2115;
  assign n15667 = n15666 ^ n15577;
  assign n15686 = n15685 ^ n15667;
  assign n15687 = n14611 ^ n13755;
  assign n15688 = n15687 ^ n14521;
  assign n15689 = n15688 ^ n15667;
  assign n15690 = ~n15686 & ~n15689;
  assign n15691 = n15690 ^ n15688;
  assign n15692 = n15691 ^ n15664;
  assign n15693 = ~n15665 & n15692;
  assign n15694 = n15693 ^ n15341;
  assign n15339 = n15186 ^ n521;
  assign n15695 = n15694 ^ n15339;
  assign n15696 = n14598 ^ n13748;
  assign n15697 = n15696 ^ n14518;
  assign n15698 = n15697 ^ n15339;
  assign n15699 = n15695 & n15698;
  assign n15700 = n15699 ^ n15697;
  assign n15701 = n15700 ^ n15337;
  assign n15702 = n15338 & ~n15701;
  assign n15703 = n15702 ^ n15336;
  assign n15334 = n15253 ^ n15244;
  assign n15704 = n15703 ^ n15334;
  assign n15705 = n14591 ^ n13735;
  assign n15706 = n15705 ^ n15105;
  assign n15707 = n15706 ^ n15334;
  assign n15708 = n15704 & n15707;
  assign n15709 = n15708 ^ n15706;
  assign n15710 = n15709 ^ n15332;
  assign n15711 = ~n15333 & ~n15710;
  assign n15712 = n15711 ^ n15331;
  assign n15328 = n15259 ^ n3258;
  assign n15329 = n15328 ^ n15236;
  assign n15713 = n15712 ^ n15329;
  assign n15714 = n14582 ^ n13725;
  assign n15715 = n15714 ^ n15213;
  assign n15716 = n15715 ^ n15329;
  assign n15717 = ~n15713 & ~n15716;
  assign n15718 = n15717 ^ n15715;
  assign n15719 = n15718 ^ n15323;
  assign n15720 = n15327 & n15719;
  assign n15721 = n15720 ^ n15326;
  assign n15322 = n15266 ^ n15234;
  assign n15722 = n15721 ^ n15322;
  assign n15723 = n14569 ^ n13715;
  assign n15724 = n15723 ^ n15363;
  assign n15725 = n15724 ^ n15322;
  assign n15726 = n15722 & n15725;
  assign n15727 = n15726 ^ n15724;
  assign n15728 = n15727 ^ n15320;
  assign n15729 = n15321 & ~n15728;
  assign n15730 = n15729 ^ n15319;
  assign n15316 = n15273 ^ n806;
  assign n15731 = n15730 ^ n15316;
  assign n15732 = n14559 ^ n13708;
  assign n15733 = n15732 ^ n15357;
  assign n15734 = n15733 ^ n15316;
  assign n15735 = n15731 & ~n15734;
  assign n15736 = n15735 ^ n15733;
  assign n15737 = n15736 ^ n15314;
  assign n15738 = ~n15315 & ~n15737;
  assign n15739 = n15738 ^ n15313;
  assign n15310 = n15280 ^ n928;
  assign n15740 = n15739 ^ n15310;
  assign n15741 = n14676 ^ n13698;
  assign n15742 = n15741 ^ n15350;
  assign n15743 = n15742 ^ n15310;
  assign n15744 = ~n15740 & ~n15743;
  assign n15745 = n15744 ^ n15742;
  assign n15746 = n15745 ^ n15305;
  assign n15747 = n15309 & ~n15746;
  assign n15748 = n15747 ^ n15308;
  assign n15749 = n15748 ^ n15303;
  assign n15750 = ~n15304 & n15749;
  assign n15751 = n15750 ^ n15302;
  assign n15299 = n15289 ^ n15222;
  assign n15752 = n15751 ^ n15299;
  assign n15753 = n14544 ^ n13680;
  assign n15754 = n15753 ^ n15398;
  assign n15755 = n15754 ^ n15299;
  assign n15756 = ~n15752 & ~n15755;
  assign n15757 = n15756 ^ n15754;
  assign n15758 = n15757 ^ n15294;
  assign n15759 = n15298 & n15758;
  assign n15760 = n15759 ^ n15297;
  assign n15762 = n15761 ^ n15760;
  assign n15763 = n14534 ^ n13665;
  assign n15764 = n15763 ^ n15343;
  assign n16064 = n15764 ^ n15761;
  assign n16065 = ~n15762 & n16064;
  assign n16066 = n16065 ^ n15764;
  assign n16062 = n15607 ^ n15599;
  assign n16060 = n14532 ^ n13663;
  assign n16061 = n16060 ^ n15417;
  assign n16063 = n16062 ^ n16061;
  assign n16098 = n16066 ^ n16063;
  assign n16099 = n16098 ^ n13688;
  assign n15765 = n15764 ^ n15762;
  assign n15766 = n15765 ^ n13694;
  assign n15767 = n15757 ^ n15298;
  assign n15768 = n15767 ^ n13464;
  assign n15769 = n15754 ^ n15752;
  assign n15770 = n15769 ^ n13314;
  assign n15771 = n15748 ^ n15304;
  assign n15772 = n15771 ^ n13117;
  assign n15773 = n15745 ^ n15309;
  assign n15774 = n15773 ^ n13122;
  assign n15775 = n15742 ^ n15740;
  assign n15776 = n15775 ^ n13127;
  assign n15777 = n15736 ^ n15315;
  assign n15778 = n15777 ^ n13132;
  assign n15779 = n15733 ^ n15731;
  assign n15780 = n15779 ^ n13134;
  assign n15781 = n15727 ^ n15321;
  assign n15782 = n15781 ^ n13139;
  assign n15783 = n15724 ^ n15722;
  assign n15784 = n15783 ^ n13144;
  assign n15785 = n15718 ^ n15327;
  assign n15786 = n15785 ^ n13149;
  assign n15787 = n15715 ^ n15713;
  assign n15788 = n15787 ^ n13154;
  assign n15789 = n15709 ^ n15333;
  assign n15790 = n15789 ^ n13159;
  assign n15791 = n15706 ^ n15704;
  assign n15792 = n15791 ^ n13164;
  assign n15793 = n15700 ^ n15338;
  assign n15794 = n15793 ^ n13169;
  assign n15795 = n15697 ^ n15695;
  assign n15796 = n15795 ^ n13174;
  assign n15797 = n15691 ^ n15665;
  assign n15798 = n15797 ^ n13263;
  assign n15799 = n15688 ^ n15686;
  assign n15800 = n15799 ^ n13179;
  assign n15801 = n15682 ^ n15680;
  assign n15802 = n15801 ^ n13184;
  assign n15803 = n15671 ^ n15669;
  assign n15804 = n13197 & n15803;
  assign n15805 = n15804 ^ n13192;
  assign n15806 = n15676 ^ n15675;
  assign n15807 = n15806 ^ n15804;
  assign n15808 = n15805 & ~n15807;
  assign n15809 = n15808 ^ n13192;
  assign n15810 = n15809 ^ n15801;
  assign n15811 = n15802 & ~n15810;
  assign n15812 = n15811 ^ n13184;
  assign n15813 = n15812 ^ n15799;
  assign n15814 = n15800 & ~n15813;
  assign n15815 = n15814 ^ n13179;
  assign n15816 = n15815 ^ n15797;
  assign n15817 = n15798 & n15816;
  assign n15818 = n15817 ^ n13263;
  assign n15819 = n15818 ^ n15795;
  assign n15820 = n15796 & n15819;
  assign n15821 = n15820 ^ n13174;
  assign n15822 = n15821 ^ n15793;
  assign n15823 = n15794 & n15822;
  assign n15824 = n15823 ^ n13169;
  assign n15825 = n15824 ^ n15791;
  assign n15826 = n15792 & ~n15825;
  assign n15827 = n15826 ^ n13164;
  assign n15828 = n15827 ^ n15789;
  assign n15829 = n15790 & ~n15828;
  assign n15830 = n15829 ^ n13159;
  assign n15831 = n15830 ^ n15787;
  assign n15832 = ~n15788 & n15831;
  assign n15833 = n15832 ^ n13154;
  assign n15834 = n15833 ^ n15785;
  assign n15835 = ~n15786 & n15834;
  assign n15836 = n15835 ^ n13149;
  assign n15837 = n15836 ^ n15783;
  assign n15838 = ~n15784 & ~n15837;
  assign n15839 = n15838 ^ n13144;
  assign n15840 = n15839 ^ n15781;
  assign n15841 = ~n15782 & ~n15840;
  assign n15842 = n15841 ^ n13139;
  assign n15843 = n15842 ^ n15779;
  assign n15844 = n15780 & ~n15843;
  assign n15845 = n15844 ^ n13134;
  assign n15846 = n15845 ^ n15777;
  assign n15847 = ~n15778 & ~n15846;
  assign n15848 = n15847 ^ n13132;
  assign n15849 = n15848 ^ n15775;
  assign n15850 = n15776 & ~n15849;
  assign n15851 = n15850 ^ n13127;
  assign n15852 = n15851 ^ n15773;
  assign n15853 = ~n15774 & ~n15852;
  assign n15854 = n15853 ^ n13122;
  assign n15855 = n15854 ^ n15771;
  assign n15856 = ~n15772 & ~n15855;
  assign n15857 = n15856 ^ n13117;
  assign n15858 = n15857 ^ n15769;
  assign n15859 = ~n15770 & n15858;
  assign n15860 = n15859 ^ n13314;
  assign n15861 = n15860 ^ n15767;
  assign n15862 = n15768 & n15861;
  assign n15863 = n15862 ^ n13464;
  assign n16100 = n15863 ^ n15765;
  assign n16101 = n15766 & n16100;
  assign n16102 = n16101 ^ n13694;
  assign n16103 = n16102 ^ n16098;
  assign n16104 = ~n16099 & n16103;
  assign n16105 = n16104 ^ n13688;
  assign n16067 = n16066 ^ n16062;
  assign n16068 = ~n16063 & ~n16067;
  assign n16069 = n16068 ^ n16061;
  assign n16058 = n15610 ^ n15597;
  assign n16056 = n14707 ^ n13659;
  assign n16057 = n16056 ^ n15424;
  assign n16059 = n16058 ^ n16057;
  assign n16096 = n16069 ^ n16059;
  assign n16097 = n16096 ^ n13682;
  assign n16123 = n16105 ^ n16097;
  assign n15864 = n15863 ^ n15766;
  assign n15865 = n15860 ^ n15768;
  assign n15866 = n15857 ^ n15770;
  assign n15867 = n15851 ^ n15774;
  assign n15868 = n15845 ^ n15778;
  assign n15869 = n15842 ^ n15780;
  assign n15870 = n15836 ^ n15784;
  assign n15871 = n15827 ^ n15790;
  assign n15872 = n15812 ^ n15800;
  assign n15873 = n15803 ^ n13197;
  assign n15874 = n15806 ^ n15805;
  assign n15875 = n15873 & n15874;
  assign n15876 = n15809 ^ n15802;
  assign n15877 = n15875 & n15876;
  assign n15878 = n15872 & n15877;
  assign n15879 = n15815 ^ n15798;
  assign n15880 = n15878 & n15879;
  assign n15881 = n15818 ^ n15796;
  assign n15882 = ~n15880 & n15881;
  assign n15883 = n15821 ^ n15794;
  assign n15884 = ~n15882 & n15883;
  assign n15885 = n15824 ^ n15792;
  assign n15886 = ~n15884 & n15885;
  assign n15887 = n15871 & n15886;
  assign n15888 = n15830 ^ n15788;
  assign n15889 = n15887 & ~n15888;
  assign n15890 = n15833 ^ n15786;
  assign n15891 = ~n15889 & n15890;
  assign n15892 = ~n15870 & ~n15891;
  assign n15893 = n15839 ^ n15782;
  assign n15894 = ~n15892 & ~n15893;
  assign n15895 = n15869 & ~n15894;
  assign n15896 = ~n15868 & n15895;
  assign n15897 = n15848 ^ n15776;
  assign n15898 = n15896 & ~n15897;
  assign n15899 = n15867 & n15898;
  assign n15900 = n15854 ^ n15772;
  assign n15901 = ~n15899 & n15900;
  assign n15902 = ~n15866 & n15901;
  assign n15903 = ~n15865 & ~n15902;
  assign n16120 = n15864 & n15903;
  assign n16121 = n16102 ^ n16099;
  assign n16122 = ~n16120 & ~n16121;
  assign n16196 = n16123 ^ n16122;
  assign n16197 = n16196 ^ n1506;
  assign n15904 = n15903 ^ n15864;
  assign n15905 = n15904 ^ n2684;
  assign n15907 = n15901 ^ n15866;
  assign n15908 = n15907 ^ n2576;
  assign n15909 = n15900 ^ n15899;
  assign n15910 = n15909 ^ n1553;
  assign n15911 = n15898 ^ n15867;
  assign n2498 = n2470 ^ x240;
  assign n2499 = n2498 ^ x432;
  assign n2500 = n2499 ^ x176;
  assign n15912 = n15911 ^ n2500;
  assign n15913 = n15897 ^ n15896;
  assign n2445 = n2423 ^ x241;
  assign n2446 = n2445 ^ x433;
  assign n2447 = n2446 ^ x177;
  assign n15914 = n15913 ^ n2447;
  assign n15916 = n15894 ^ n15869;
  assign n1379 = n1273 ^ x243;
  assign n1380 = n1379 ^ x435;
  assign n1381 = n1380 ^ x179;
  assign n15917 = n15916 ^ n1381;
  assign n15918 = n15893 ^ n15892;
  assign n15919 = n15918 ^ n1187;
  assign n15920 = n15891 ^ n15870;
  assign n1030 = n948 ^ x245;
  assign n1031 = n1030 ^ x437;
  assign n1032 = n1031 ^ x181;
  assign n15921 = n15920 ^ n1032;
  assign n15923 = n15888 ^ n15887;
  assign n15924 = n15923 ^ n904;
  assign n15926 = n15885 ^ n15884;
  assign n15927 = n15926 ^ n886;
  assign n15928 = n15883 ^ n15882;
  assign n15929 = n15928 ^ n726;
  assign n15931 = n15879 ^ n15878;
  assign n15932 = n15931 ^ n551;
  assign n15933 = n15877 ^ n15872;
  assign n15934 = n15933 ^ n638;
  assign n15935 = n15876 ^ n15875;
  assign n532 = n528 ^ x254;
  assign n533 = n532 ^ x446;
  assign n534 = n533 ^ x190;
  assign n15936 = n15935 ^ n534;
  assign n15940 = ~n15873 & n15939;
  assign n15941 = n15940 ^ n3275;
  assign n15942 = n15874 ^ n15873;
  assign n15943 = n15942 ^ n15940;
  assign n15944 = n15941 & ~n15943;
  assign n15945 = n15944 ^ n3275;
  assign n15946 = n15945 ^ n15935;
  assign n15947 = n15936 & ~n15946;
  assign n15948 = n15947 ^ n534;
  assign n15949 = n15948 ^ n15933;
  assign n15950 = n15934 & ~n15949;
  assign n15951 = n15950 ^ n638;
  assign n15952 = n15951 ^ n15931;
  assign n15953 = n15932 & ~n15952;
  assign n15954 = n15953 ^ n551;
  assign n15930 = n15881 ^ n15880;
  assign n15955 = n15954 ^ n15930;
  assign n15959 = n15958 ^ n15930;
  assign n15960 = ~n15955 & n15959;
  assign n15961 = n15960 ^ n15958;
  assign n15962 = n15961 ^ n15928;
  assign n15963 = ~n15929 & n15962;
  assign n15964 = n15963 ^ n726;
  assign n15965 = n15964 ^ n15926;
  assign n15966 = n15927 & ~n15965;
  assign n15967 = n15966 ^ n886;
  assign n15925 = n15886 ^ n15871;
  assign n15968 = n15967 ^ n15925;
  assign n15969 = n15925 ^ n892;
  assign n15970 = n15968 & ~n15969;
  assign n15971 = n15970 ^ n892;
  assign n15972 = n15971 ^ n15923;
  assign n15973 = n15924 & ~n15972;
  assign n15974 = n15973 ^ n904;
  assign n15922 = n15890 ^ n15889;
  assign n15975 = n15974 ^ n15922;
  assign n1018 = n934 ^ x246;
  assign n1019 = n1018 ^ x438;
  assign n1020 = n1019 ^ x182;
  assign n15976 = n15922 ^ n1020;
  assign n15977 = n15975 & ~n15976;
  assign n15978 = n15977 ^ n1020;
  assign n15979 = n15978 ^ n15920;
  assign n15980 = ~n15921 & n15979;
  assign n15981 = n15980 ^ n1032;
  assign n15982 = n15981 ^ n15918;
  assign n15983 = n15919 & ~n15982;
  assign n15984 = n15983 ^ n1187;
  assign n15985 = n15984 ^ n15916;
  assign n15986 = n15917 & ~n15985;
  assign n15987 = n15986 ^ n1381;
  assign n15915 = n15895 ^ n15868;
  assign n15988 = n15987 ^ n15915;
  assign n15989 = n15915 ^ n1387;
  assign n15990 = ~n15988 & n15989;
  assign n15991 = n15990 ^ n1387;
  assign n15992 = n15991 ^ n15913;
  assign n15993 = n15914 & ~n15992;
  assign n15994 = n15993 ^ n2447;
  assign n15995 = n15994 ^ n15911;
  assign n15996 = ~n15912 & n15995;
  assign n15997 = n15996 ^ n2500;
  assign n15998 = n15997 ^ n15909;
  assign n15999 = ~n15910 & n15998;
  assign n16000 = n15999 ^ n1553;
  assign n16001 = n16000 ^ n15907;
  assign n16002 = ~n15908 & n16001;
  assign n16003 = n16002 ^ n2576;
  assign n15906 = n15902 ^ n15865;
  assign n16004 = n16003 ^ n15906;
  assign n16005 = n15906 ^ n2838;
  assign n16006 = n16004 & ~n16005;
  assign n16007 = n16006 ^ n2838;
  assign n16199 = n16007 ^ n15904;
  assign n16200 = ~n15905 & n16199;
  assign n16201 = n16200 ^ n2684;
  assign n16198 = n16121 ^ n16120;
  assign n16202 = n16201 ^ n16198;
  assign n16203 = n16198 ^ n2852;
  assign n16204 = ~n16202 & n16203;
  assign n16205 = n16204 ^ n2852;
  assign n16206 = n16205 ^ n16196;
  assign n16207 = n16197 & ~n16206;
  assign n16208 = n16207 ^ n1506;
  assign n16106 = n16105 ^ n16096;
  assign n16107 = ~n16097 & n16106;
  assign n16108 = n16107 ^ n13682;
  assign n16074 = n15342 ^ n13658;
  assign n16075 = n16074 ^ n14715;
  assign n16070 = n16069 ^ n16058;
  assign n16071 = n16059 & n16070;
  assign n16072 = n16071 ^ n16057;
  assign n16032 = n15613 ^ n15595;
  assign n16073 = n16072 ^ n16032;
  assign n16094 = n16075 ^ n16073;
  assign n16095 = n16094 ^ n13676;
  assign n16125 = n16108 ^ n16095;
  assign n16124 = ~n16122 & n16123;
  assign n16195 = n16125 ^ n16124;
  assign n16209 = n16208 ^ n16195;
  assign n16765 = n16209 ^ n1546;
  assign n16762 = n15034 ^ n14392;
  assign n16763 = n16762 ^ n15676;
  assign n16598 = n16205 ^ n16197;
  assign n16595 = n15035 ^ n14397;
  assign n16596 = n16595 ^ n15669;
  assign n16758 = n16598 ^ n16596;
  assign n16401 = n16202 ^ n2852;
  assign n16398 = n15043 ^ n14405;
  assign n16267 = n15644 ^ n1838;
  assign n16399 = n16398 ^ n16267;
  assign n16591 = n16401 ^ n16399;
  assign n16010 = n15036 ^ n14407;
  assign n16009 = n15640 ^ n15584;
  assign n16011 = n16010 ^ n16009;
  assign n16008 = n16007 ^ n15905;
  assign n16012 = n16011 ^ n16008;
  assign n16016 = n15553 ^ n14715;
  assign n16015 = n15634 ^ n15631;
  assign n16017 = n16016 ^ n16015;
  assign n16014 = n16000 ^ n15908;
  assign n16018 = n16017 ^ n16014;
  assign n16021 = n15437 ^ n14707;
  assign n16020 = n15627 ^ n15589;
  assign n16022 = n16021 ^ n16020;
  assign n16019 = n15997 ^ n15910;
  assign n16023 = n16022 ^ n16019;
  assign n16026 = n15624 ^ n1582;
  assign n16025 = n15342 ^ n14532;
  assign n16027 = n16026 ^ n16025;
  assign n16024 = n15994 ^ n15912;
  assign n16028 = n16027 ^ n16024;
  assign n16373 = n15991 ^ n15914;
  assign n16031 = n15343 ^ n14544;
  assign n16033 = n16032 ^ n16031;
  assign n16030 = n15984 ^ n15917;
  assign n16034 = n16033 ^ n16030;
  assign n16345 = n15975 ^ n1020;
  assign n16338 = n15971 ^ n15924;
  assign n16331 = n15968 ^ n892;
  assign n16324 = n15964 ^ n15927;
  assign n16317 = n15961 ^ n15929;
  assign n16310 = n15958 ^ n15955;
  assign n16303 = n15951 ^ n15932;
  assign n16039 = n15948 ^ n15934;
  assign n16037 = n15325 ^ n14516;
  assign n16038 = n16037 ^ n15316;
  assign n16040 = n16039 ^ n16038;
  assign n16044 = n15942 ^ n15941;
  assign n16042 = n15173 ^ n14596;
  assign n16043 = n16042 ^ n15322;
  assign n16045 = n16044 ^ n16043;
  assign n16284 = n15939 ^ n15873;
  assign n16086 = n14405 ^ n13873;
  assign n16087 = n16086 ^ n15568;
  assign n16049 = n14407 ^ n13881;
  assign n16050 = n16049 ^ n15553;
  assign n16048 = n15620 ^ n15592;
  assign n16051 = n16050 ^ n16048;
  assign n16053 = n14524 ^ n13655;
  assign n16054 = n16053 ^ n15437;
  assign n16052 = n15617 ^ n2671;
  assign n16055 = n16054 ^ n16052;
  assign n16076 = n16075 ^ n16032;
  assign n16077 = ~n16073 & ~n16076;
  assign n16078 = n16077 ^ n16075;
  assign n16079 = n16078 ^ n16052;
  assign n16080 = ~n16055 & ~n16079;
  assign n16081 = n16080 ^ n16054;
  assign n16082 = n16081 ^ n16048;
  assign n16083 = ~n16051 & ~n16082;
  assign n16084 = n16083 ^ n16050;
  assign n16085 = n16084 ^ n16026;
  assign n16088 = n16087 ^ n16085;
  assign n16089 = n16088 ^ n13214;
  assign n16090 = n16081 ^ n16051;
  assign n16091 = n16090 ^ n13219;
  assign n16092 = n16078 ^ n16055;
  assign n16093 = n16092 ^ n13670;
  assign n16109 = n16108 ^ n16094;
  assign n16110 = n16095 & n16109;
  assign n16111 = n16110 ^ n13676;
  assign n16112 = n16111 ^ n16092;
  assign n16113 = ~n16093 & n16112;
  assign n16114 = n16113 ^ n13670;
  assign n16115 = n16114 ^ n16090;
  assign n16116 = ~n16091 & ~n16115;
  assign n16117 = n16116 ^ n13219;
  assign n16138 = n16117 ^ n16088;
  assign n16139 = n16089 & n16138;
  assign n16140 = n16139 ^ n13214;
  assign n16141 = n16140 ^ n13231;
  assign n16135 = n14397 ^ n13868;
  assign n16136 = n16135 ^ n15036;
  assign n16131 = n16087 ^ n16026;
  assign n16132 = ~n16085 & n16131;
  assign n16133 = n16132 ^ n16087;
  assign n16134 = n16133 ^ n16020;
  assign n16137 = n16136 ^ n16134;
  assign n16142 = n16141 ^ n16137;
  assign n16118 = n16117 ^ n16089;
  assign n16119 = n16114 ^ n16091;
  assign n16126 = n16124 & ~n16125;
  assign n16127 = n16111 ^ n16093;
  assign n16128 = ~n16126 & n16127;
  assign n16129 = ~n16119 & ~n16128;
  assign n16130 = ~n16118 & n16129;
  assign n16188 = n16142 ^ n16130;
  assign n16189 = n16188 ^ n2074;
  assign n16191 = n16128 ^ n16119;
  assign n16192 = n16191 ^ n1669;
  assign n16193 = n16127 ^ n16126;
  assign n16194 = n16193 ^ n1663;
  assign n16210 = n16195 ^ n1546;
  assign n16211 = ~n16209 & n16210;
  assign n16212 = n16211 ^ n1546;
  assign n16213 = n16212 ^ n16193;
  assign n16214 = ~n16194 & n16213;
  assign n16215 = n16214 ^ n1663;
  assign n16216 = n16215 ^ n16191;
  assign n16217 = ~n16192 & n16216;
  assign n16218 = n16217 ^ n1669;
  assign n16190 = n16129 ^ n16118;
  assign n16219 = n16218 ^ n16190;
  assign n16220 = n16190 ^ n1748;
  assign n16221 = ~n16219 & n16220;
  assign n16222 = n16221 ^ n1748;
  assign n16223 = n16222 ^ n16188;
  assign n16224 = ~n16189 & n16223;
  assign n16225 = n16224 ^ n2074;
  assign n16152 = n16137 ^ n13231;
  assign n16153 = n16140 ^ n16137;
  assign n16154 = n16152 & n16153;
  assign n16155 = n16154 ^ n13231;
  assign n16148 = n14392 ^ n13863;
  assign n16149 = n16148 ^ n15043;
  assign n16144 = n16136 ^ n16020;
  assign n16145 = ~n16134 & ~n16144;
  assign n16146 = n16145 ^ n16136;
  assign n16147 = n16146 ^ n16015;
  assign n16150 = n16149 ^ n16147;
  assign n16151 = n16150 ^ n13209;
  assign n16156 = n16155 ^ n16151;
  assign n16143 = n16130 & n16142;
  assign n16187 = n16156 ^ n16143;
  assign n16226 = n16225 ^ n16187;
  assign n16227 = n16187 ^ n1880;
  assign n16228 = n16226 & ~n16227;
  assign n16229 = n16228 ^ n1880;
  assign n16167 = n16155 ^ n16150;
  assign n16168 = n16151 & n16167;
  assign n16169 = n16168 ^ n13209;
  assign n16161 = n16149 ^ n16015;
  assign n16162 = n16147 & ~n16161;
  assign n16163 = n16162 ^ n16149;
  assign n16160 = n15637 ^ n15586;
  assign n16164 = n16163 ^ n16160;
  assign n16158 = n14387 ^ n13913;
  assign n16159 = n16158 ^ n15035;
  assign n16165 = n16164 ^ n16159;
  assign n16166 = n16165 ^ n13110;
  assign n16170 = n16169 ^ n16166;
  assign n16157 = ~n16143 & n16156;
  assign n16185 = n16170 ^ n16157;
  assign n16186 = n16185 ^ n2088;
  assign n16237 = n16229 ^ n16186;
  assign n16235 = n14613 ^ n14520;
  assign n16236 = n16235 ^ n15334;
  assign n16238 = n16237 ^ n16236;
  assign n16243 = n14618 ^ n14521;
  assign n16244 = n16243 ^ n15337;
  assign n16239 = n16222 ^ n16189;
  assign n16240 = n14626 ^ n14522;
  assign n16241 = n16240 ^ n15339;
  assign n16242 = ~n16239 & ~n16241;
  assign n16245 = n16244 ^ n16242;
  assign n16246 = n16226 ^ n1880;
  assign n16247 = n16246 ^ n16244;
  assign n16248 = ~n16245 & ~n16247;
  assign n16249 = n16248 ^ n16242;
  assign n16250 = n16249 ^ n16237;
  assign n16251 = ~n16238 & ~n16250;
  assign n16252 = n16251 ^ n16236;
  assign n16230 = n16229 ^ n16185;
  assign n16231 = n16186 & ~n16230;
  assign n16232 = n16231 ^ n2088;
  assign n16179 = n16169 ^ n16165;
  assign n16180 = n16166 & n16179;
  assign n16181 = n16180 ^ n13110;
  assign n16182 = n16181 ^ n13203;
  assign n16174 = n16160 ^ n16159;
  assign n16175 = ~n16164 & n16174;
  assign n16176 = n16175 ^ n16159;
  assign n16177 = n16176 ^ n16009;
  assign n16172 = n14451 ^ n13776;
  assign n16173 = n16172 ^ n15034;
  assign n16178 = n16177 ^ n16173;
  assign n16183 = n16182 ^ n16178;
  assign n16171 = ~n16157 & n16170;
  assign n16184 = n16183 ^ n16171;
  assign n16233 = n16232 ^ n16184;
  assign n16234 = n16233 ^ n2107;
  assign n16253 = n16252 ^ n16234;
  assign n16254 = n15332 ^ n14518;
  assign n16255 = n16254 ^ n14611;
  assign n16256 = n16255 ^ n16252;
  assign n16257 = ~n16253 & ~n16256;
  assign n16258 = n16257 ^ n16255;
  assign n16046 = n14606 ^ n14514;
  assign n16047 = n16046 ^ n15329;
  assign n16259 = n16258 ^ n16047;
  assign n16276 = n16184 ^ n2107;
  assign n16277 = n16233 & ~n16276;
  assign n16278 = n16277 ^ n2107;
  assign n16279 = n16278 ^ n2241;
  assign n16269 = n16178 ^ n13203;
  assign n16270 = n16181 ^ n16178;
  assign n16271 = ~n16269 & ~n16270;
  assign n16272 = n16271 ^ n13203;
  assign n16273 = n16272 ^ n13199;
  assign n16263 = n16173 ^ n16009;
  assign n16264 = ~n16177 & n16263;
  assign n16265 = n16264 ^ n16173;
  assign n16261 = n14506 ^ n13775;
  assign n16262 = n16261 ^ n15033;
  assign n16266 = n16265 ^ n16262;
  assign n16268 = n16267 ^ n16266;
  assign n16274 = n16273 ^ n16268;
  assign n16260 = n16171 & n16183;
  assign n16275 = n16274 ^ n16260;
  assign n16280 = n16279 ^ n16275;
  assign n16281 = n16280 ^ n16258;
  assign n16282 = n16259 & ~n16281;
  assign n16283 = n16282 ^ n16047;
  assign n16285 = n16284 ^ n16283;
  assign n16286 = n15105 ^ n14598;
  assign n16287 = n16286 ^ n15323;
  assign n16288 = n16287 ^ n16284;
  assign n16289 = n16285 & ~n16288;
  assign n16290 = n16289 ^ n16287;
  assign n16291 = n16290 ^ n16044;
  assign n16292 = ~n16045 & ~n16291;
  assign n16293 = n16292 ^ n16043;
  assign n16041 = n15945 ^ n15936;
  assign n16294 = n16293 ^ n16041;
  assign n16295 = n15213 ^ n14591;
  assign n16296 = n16295 ^ n15320;
  assign n16297 = n16296 ^ n16041;
  assign n16298 = n16294 & ~n16297;
  assign n16299 = n16298 ^ n16296;
  assign n16300 = n16299 ^ n16039;
  assign n16301 = n16040 & n16300;
  assign n16302 = n16301 ^ n16038;
  assign n16304 = n16303 ^ n16302;
  assign n16305 = n15363 ^ n14582;
  assign n16306 = n16305 ^ n15314;
  assign n16307 = n16306 ^ n16303;
  assign n16308 = ~n16304 & ~n16307;
  assign n16309 = n16308 ^ n16306;
  assign n16311 = n16310 ^ n16309;
  assign n16312 = n15318 ^ n14577;
  assign n16313 = n16312 ^ n15310;
  assign n16314 = n16313 ^ n16310;
  assign n16315 = n16311 & n16314;
  assign n16316 = n16315 ^ n16313;
  assign n16318 = n16317 ^ n16316;
  assign n16319 = n15357 ^ n14569;
  assign n16320 = n16319 ^ n15305;
  assign n16321 = n16320 ^ n16317;
  assign n16322 = n16318 & ~n16321;
  assign n16323 = n16322 ^ n16320;
  assign n16325 = n16324 ^ n16323;
  assign n16326 = n15312 ^ n14567;
  assign n16327 = n16326 ^ n15303;
  assign n16328 = n16327 ^ n16324;
  assign n16329 = ~n16325 & ~n16328;
  assign n16330 = n16329 ^ n16327;
  assign n16332 = n16331 ^ n16330;
  assign n16333 = n15350 ^ n14559;
  assign n16334 = n16333 ^ n15299;
  assign n16335 = n16334 ^ n16331;
  assign n16336 = ~n16332 & n16335;
  assign n16337 = n16336 ^ n16334;
  assign n16339 = n16338 ^ n16337;
  assign n16340 = n15307 ^ n14554;
  assign n16341 = n16340 ^ n15294;
  assign n16342 = n16341 ^ n16338;
  assign n16343 = n16339 & ~n16342;
  assign n16344 = n16343 ^ n16341;
  assign n16346 = n16345 ^ n16344;
  assign n16347 = n15761 ^ n15301;
  assign n16348 = n16347 ^ n14676;
  assign n16349 = n16348 ^ n16345;
  assign n16350 = ~n16346 & ~n16349;
  assign n16351 = n16350 ^ n16348;
  assign n16036 = n15978 ^ n15921;
  assign n16352 = n16351 ^ n16036;
  assign n16353 = n15398 ^ n14684;
  assign n16354 = n16353 ^ n16062;
  assign n16355 = n16354 ^ n16036;
  assign n16356 = n16352 & n16355;
  assign n16357 = n16356 ^ n16354;
  assign n16035 = n15981 ^ n15919;
  assign n16358 = n16357 ^ n16035;
  assign n16359 = n15296 ^ n14549;
  assign n16360 = n16359 ^ n16058;
  assign n16361 = n16360 ^ n16035;
  assign n16362 = n16358 & n16361;
  assign n16363 = n16362 ^ n16360;
  assign n16364 = n16363 ^ n16030;
  assign n16365 = ~n16034 & ~n16364;
  assign n16366 = n16365 ^ n16033;
  assign n16029 = n15988 ^ n1387;
  assign n16367 = n16366 ^ n16029;
  assign n16368 = n15417 ^ n14539;
  assign n16369 = n16368 ^ n16052;
  assign n16370 = n16369 ^ n16029;
  assign n16371 = n16367 & n16370;
  assign n16372 = n16371 ^ n16369;
  assign n16374 = n16373 ^ n16372;
  assign n16375 = n15424 ^ n14534;
  assign n16376 = n16375 ^ n16048;
  assign n16377 = n16376 ^ n16373;
  assign n16378 = ~n16374 & n16377;
  assign n16379 = n16378 ^ n16376;
  assign n16380 = n16379 ^ n16027;
  assign n16381 = n16028 & n16380;
  assign n16382 = n16381 ^ n16024;
  assign n16383 = n16382 ^ n16022;
  assign n16384 = ~n16023 & n16383;
  assign n16385 = n16384 ^ n16019;
  assign n16386 = n16385 ^ n16014;
  assign n16387 = n16018 & ~n16386;
  assign n16388 = n16387 ^ n16017;
  assign n16013 = n16004 ^ n2838;
  assign n16389 = n16388 ^ n16013;
  assign n16390 = n15568 ^ n14524;
  assign n16391 = n16390 ^ n16160;
  assign n16392 = n16391 ^ n16013;
  assign n16393 = ~n16389 & n16392;
  assign n16394 = n16393 ^ n16391;
  assign n16395 = n16394 ^ n16008;
  assign n16396 = n16012 & ~n16395;
  assign n16397 = n16396 ^ n16011;
  assign n16592 = n16401 ^ n16397;
  assign n16593 = n16591 & n16592;
  assign n16594 = n16593 ^ n16399;
  assign n16759 = n16598 ^ n16594;
  assign n16760 = n16758 & ~n16759;
  assign n16761 = n16760 ^ n16596;
  assign n16764 = n16763 ^ n16761;
  assign n16766 = n16765 ^ n16764;
  assign n16767 = n16766 ^ n13863;
  assign n16597 = n16596 ^ n16594;
  assign n16599 = n16598 ^ n16597;
  assign n16754 = n16599 ^ n13868;
  assign n16403 = n16394 ^ n16012;
  assign n16404 = n16403 ^ n13881;
  assign n16406 = n16385 ^ n16018;
  assign n16407 = n16406 ^ n13658;
  assign n16408 = n16382 ^ n16023;
  assign n16409 = n16408 ^ n13659;
  assign n16410 = n16379 ^ n16028;
  assign n16411 = n16410 ^ n13663;
  assign n16412 = n16376 ^ n16374;
  assign n16413 = n16412 ^ n13665;
  assign n16416 = n16360 ^ n16358;
  assign n16417 = n16416 ^ n13686;
  assign n16418 = n16354 ^ n16352;
  assign n16419 = n16418 ^ n13692;
  assign n16420 = n16348 ^ n16346;
  assign n16421 = n16420 ^ n13698;
  assign n16422 = n16341 ^ n16339;
  assign n16423 = n16422 ^ n13703;
  assign n16424 = n16334 ^ n16332;
  assign n16425 = n16424 ^ n13708;
  assign n16426 = n16327 ^ n16325;
  assign n16427 = n16426 ^ n13713;
  assign n16428 = n16320 ^ n16318;
  assign n16429 = n16428 ^ n13715;
  assign n16430 = n16313 ^ n16311;
  assign n16431 = n16430 ^ n13720;
  assign n16432 = n16306 ^ n16304;
  assign n16433 = n16432 ^ n13725;
  assign n16434 = n16299 ^ n16040;
  assign n16435 = n16434 ^ n13733;
  assign n16436 = n16296 ^ n16294;
  assign n16437 = n16436 ^ n13735;
  assign n16438 = n16290 ^ n16045;
  assign n16439 = n16438 ^ n13740;
  assign n16440 = n16287 ^ n16285;
  assign n16441 = n16440 ^ n13748;
  assign n16442 = n16280 ^ n16047;
  assign n16443 = n16442 ^ n16258;
  assign n16444 = n16443 ^ n13753;
  assign n16445 = n16255 ^ n16253;
  assign n16446 = n16445 ^ n13755;
  assign n16447 = n16249 ^ n16238;
  assign n16448 = n16447 ^ n13763;
  assign n16449 = n16241 ^ n16239;
  assign n16450 = n13773 & n16449;
  assign n16451 = n16450 ^ n13768;
  assign n16452 = n16246 ^ n16245;
  assign n16453 = n16452 ^ n16450;
  assign n16454 = ~n16451 & ~n16453;
  assign n16455 = n16454 ^ n13768;
  assign n16456 = n16455 ^ n16447;
  assign n16457 = ~n16448 & ~n16456;
  assign n16458 = n16457 ^ n13763;
  assign n16459 = n16458 ^ n16445;
  assign n16460 = ~n16446 & ~n16459;
  assign n16461 = n16460 ^ n13755;
  assign n16462 = n16461 ^ n16443;
  assign n16463 = ~n16444 & n16462;
  assign n16464 = n16463 ^ n13753;
  assign n16465 = n16464 ^ n16440;
  assign n16466 = n16441 & ~n16465;
  assign n16467 = n16466 ^ n13748;
  assign n16468 = n16467 ^ n16438;
  assign n16469 = ~n16439 & ~n16468;
  assign n16470 = n16469 ^ n13740;
  assign n16471 = n16470 ^ n16436;
  assign n16472 = ~n16437 & ~n16471;
  assign n16473 = n16472 ^ n13735;
  assign n16474 = n16473 ^ n16434;
  assign n16475 = n16435 & ~n16474;
  assign n16476 = n16475 ^ n13733;
  assign n16477 = n16476 ^ n16432;
  assign n16478 = ~n16433 & ~n16477;
  assign n16479 = n16478 ^ n13725;
  assign n16480 = n16479 ^ n16430;
  assign n16481 = n16431 & n16480;
  assign n16482 = n16481 ^ n13720;
  assign n16483 = n16482 ^ n16428;
  assign n16484 = n16429 & ~n16483;
  assign n16485 = n16484 ^ n13715;
  assign n16486 = n16485 ^ n16426;
  assign n16487 = n16427 & ~n16486;
  assign n16488 = n16487 ^ n13713;
  assign n16489 = n16488 ^ n16424;
  assign n16490 = ~n16425 & ~n16489;
  assign n16491 = n16490 ^ n13708;
  assign n16492 = n16491 ^ n16422;
  assign n16493 = n16423 & ~n16492;
  assign n16494 = n16493 ^ n13703;
  assign n16495 = n16494 ^ n16420;
  assign n16496 = ~n16421 & ~n16495;
  assign n16497 = n16496 ^ n13698;
  assign n16498 = n16497 ^ n16418;
  assign n16499 = n16419 & n16498;
  assign n16500 = n16499 ^ n13692;
  assign n16501 = n16500 ^ n16416;
  assign n16502 = ~n16417 & n16501;
  assign n16503 = n16502 ^ n13686;
  assign n16415 = n16363 ^ n16034;
  assign n16504 = n16503 ^ n16415;
  assign n16505 = n16415 ^ n13680;
  assign n16506 = n16504 & n16505;
  assign n16507 = n16506 ^ n13680;
  assign n16414 = n16369 ^ n16367;
  assign n16508 = n16507 ^ n16414;
  assign n16509 = n16414 ^ n13674;
  assign n16510 = ~n16508 & ~n16509;
  assign n16511 = n16510 ^ n13674;
  assign n16512 = n16511 ^ n16412;
  assign n16513 = n16413 & ~n16512;
  assign n16514 = n16513 ^ n13665;
  assign n16515 = n16514 ^ n16410;
  assign n16516 = n16411 & ~n16515;
  assign n16517 = n16516 ^ n13663;
  assign n16518 = n16517 ^ n16408;
  assign n16519 = n16409 & ~n16518;
  assign n16520 = n16519 ^ n13659;
  assign n16521 = n16520 ^ n16406;
  assign n16522 = n16407 & n16521;
  assign n16523 = n16522 ^ n13658;
  assign n16405 = n16391 ^ n16389;
  assign n16524 = n16523 ^ n16405;
  assign n16525 = n16405 ^ n13655;
  assign n16526 = ~n16524 & ~n16525;
  assign n16527 = n16526 ^ n13655;
  assign n16528 = n16527 ^ n16403;
  assign n16529 = ~n16404 & n16528;
  assign n16530 = n16529 ^ n13881;
  assign n16400 = n16399 ^ n16397;
  assign n16402 = n16401 ^ n16400;
  assign n16531 = n16530 ^ n16402;
  assign n16587 = n16402 ^ n13873;
  assign n16588 = n16531 & ~n16587;
  assign n16589 = n16588 ^ n13873;
  assign n16755 = n16599 ^ n16589;
  assign n16756 = ~n16754 & ~n16755;
  assign n16757 = n16756 ^ n13868;
  assign n16768 = n16767 ^ n16757;
  assign n16532 = n16531 ^ n13873;
  assign n16533 = n16520 ^ n16407;
  assign n16534 = n16517 ^ n16409;
  assign n16535 = n16514 ^ n16411;
  assign n16536 = n16511 ^ n16413;
  assign n16537 = n16508 ^ n13674;
  assign n16538 = n16500 ^ n16417;
  assign n16539 = n16497 ^ n16419;
  assign n16540 = n16494 ^ n13698;
  assign n16541 = n16540 ^ n16420;
  assign n16542 = n16491 ^ n16423;
  assign n16543 = n16482 ^ n16429;
  assign n16544 = n16479 ^ n16431;
  assign n16545 = n16476 ^ n16433;
  assign n16546 = n16473 ^ n16435;
  assign n16547 = n16470 ^ n16437;
  assign n16548 = n16458 ^ n16446;
  assign n16549 = n16449 ^ n13773;
  assign n16550 = n16452 ^ n16451;
  assign n16551 = n16549 & ~n16550;
  assign n16552 = n16455 ^ n16448;
  assign n16553 = n16551 & n16552;
  assign n16554 = ~n16548 & n16553;
  assign n16555 = n16461 ^ n16444;
  assign n16556 = n16554 & n16555;
  assign n16557 = n16464 ^ n16441;
  assign n16558 = ~n16556 & n16557;
  assign n16559 = n16467 ^ n16439;
  assign n16560 = ~n16558 & n16559;
  assign n16561 = n16547 & ~n16560;
  assign n16562 = n16546 & n16561;
  assign n16563 = ~n16545 & n16562;
  assign n16564 = n16544 & ~n16563;
  assign n16565 = n16543 & ~n16564;
  assign n16566 = n16485 ^ n16427;
  assign n16567 = ~n16565 & ~n16566;
  assign n16568 = n16488 ^ n16425;
  assign n16569 = ~n16567 & ~n16568;
  assign n16570 = ~n16542 & n16569;
  assign n16571 = n16541 & n16570;
  assign n16572 = n16539 & n16571;
  assign n16573 = ~n16538 & ~n16572;
  assign n16574 = n16504 ^ n13680;
  assign n16575 = n16573 & n16574;
  assign n16576 = ~n16537 & ~n16575;
  assign n16577 = ~n16536 & n16576;
  assign n16578 = n16535 & ~n16577;
  assign n16579 = ~n16534 & ~n16578;
  assign n16580 = ~n16533 & n16579;
  assign n16581 = n16524 ^ n13655;
  assign n16582 = ~n16580 & n16581;
  assign n16583 = n16527 ^ n13881;
  assign n16584 = n16583 ^ n16403;
  assign n16585 = ~n16582 & n16584;
  assign n16586 = n16532 & n16585;
  assign n16590 = n16589 ^ n13868;
  assign n16600 = n16599 ^ n16590;
  assign n16769 = n16586 & n16600;
  assign n16778 = ~n16768 & ~n16769;
  assign n16788 = n16766 ^ n16757;
  assign n16789 = n16767 & n16788;
  assign n16790 = n16789 ^ n13863;
  assign n16784 = n15033 ^ n14387;
  assign n16785 = n16784 ^ n15668;
  assign n16783 = n16212 ^ n16194;
  assign n16786 = n16785 ^ n16783;
  assign n16779 = n16765 ^ n16763;
  assign n16780 = n16765 ^ n16761;
  assign n16781 = n16779 & ~n16780;
  assign n16782 = n16781 ^ n16763;
  assign n16787 = n16786 ^ n16782;
  assign n16791 = n16790 ^ n16787;
  assign n16792 = n16791 ^ n13913;
  assign n16835 = ~n16778 & n16792;
  assign n16830 = n16215 ^ n16192;
  assign n16828 = n15667 ^ n14451;
  assign n16829 = n16828 ^ n15065;
  assign n16831 = n16830 ^ n16829;
  assign n16825 = n16783 ^ n16782;
  assign n16826 = ~n16786 & n16825;
  assign n16827 = n16826 ^ n16785;
  assign n16832 = n16831 ^ n16827;
  assign n16833 = n16832 ^ n13776;
  assign n16822 = n16787 ^ n13913;
  assign n16823 = n16791 & ~n16822;
  assign n16824 = n16823 ^ n13913;
  assign n16834 = n16833 ^ n16824;
  assign n16836 = n16835 ^ n16834;
  assign n16837 = n16836 ^ n2120;
  assign n16793 = n16792 ^ n16778;
  assign n16794 = n16793 ^ n1943;
  assign n16770 = n16769 ^ n16768;
  assign n16771 = n16770 ^ n1946;
  assign n16601 = n16600 ^ n16586;
  assign n16750 = n16601 ^ n1826;
  assign n16602 = n16585 ^ n16532;
  assign n16603 = n16602 ^ n1714;
  assign n16604 = n16584 ^ n16582;
  assign n16605 = n16604 ^ n1708;
  assign n16606 = n16581 ^ n16580;
  assign n16607 = n16606 ^ n1738;
  assign n16608 = n16579 ^ n16533;
  assign n16612 = n16611 ^ n16608;
  assign n16725 = n16578 ^ n16534;
  assign n16613 = n16577 ^ n16535;
  assign n16614 = n16613 ^ n1577;
  assign n16615 = n16576 ^ n16536;
  assign n16616 = n16615 ^ n2741;
  assign n16617 = n16575 ^ n16537;
  assign n16618 = n16617 ^ n1521;
  assign n16620 = n16572 ^ n16538;
  assign n2557 = n2517 ^ x271;
  assign n2558 = n2557 ^ x463;
  assign n2559 = n2558 ^ x207;
  assign n16621 = n16620 ^ n2559;
  assign n16622 = n16571 ^ n16539;
  assign n16623 = n16622 ^ n2552;
  assign n16624 = n16570 ^ n16541;
  assign n16625 = n16624 ^ n3161;
  assign n16626 = n16569 ^ n16542;
  assign n16627 = n16626 ^ n3014;
  assign n16628 = n16568 ^ n16567;
  assign n1313 = n1207 ^ x275;
  assign n1314 = n1313 ^ x467;
  assign n1315 = n1314 ^ x211;
  assign n16629 = n16628 ^ n1315;
  assign n16631 = n16564 ^ n16543;
  assign n1133 = n1058 ^ x277;
  assign n1134 = n1133 ^ x469;
  assign n1135 = n1134 ^ x213;
  assign n16632 = n16631 ^ n1135;
  assign n16634 = n16562 ^ n16545;
  assign n16635 = n16634 ^ n1143;
  assign n16637 = n16560 ^ n16547;
  assign n16638 = n16637 ^ n662;
  assign n16639 = n16559 ^ n16558;
  assign n16640 = n16639 ^ n612;
  assign n16642 = n16555 ^ n16554;
  assign n16643 = n16642 ^ n574;
  assign n16644 = n16553 ^ n16548;
  assign n16645 = n16644 ^ n3248;
  assign n16646 = n16552 ^ n16551;
  assign n16650 = n16649 ^ n16646;
  assign n2325 = n2225 ^ x256;
  assign n2326 = n2325 ^ x448;
  assign n2327 = n2326 ^ x192;
  assign n16651 = n2327 & ~n16549;
  assign n16655 = n16654 ^ n16651;
  assign n16656 = n16550 ^ n16549;
  assign n16657 = n16656 ^ n16651;
  assign n16658 = n16655 & n16657;
  assign n16659 = n16658 ^ n16654;
  assign n16660 = n16659 ^ n16646;
  assign n16661 = n16650 & ~n16660;
  assign n16662 = n16661 ^ n16649;
  assign n16663 = n16662 ^ n16644;
  assign n16664 = ~n16645 & n16663;
  assign n16665 = n16664 ^ n3248;
  assign n16666 = n16665 ^ n16642;
  assign n16667 = n16643 & ~n16666;
  assign n16668 = n16667 ^ n574;
  assign n16641 = n16557 ^ n16556;
  assign n16669 = n16668 ^ n16641;
  assign n16670 = n16641 ^ n580;
  assign n16671 = ~n16669 & n16670;
  assign n16672 = n16671 ^ n580;
  assign n16673 = n16672 ^ n16639;
  assign n16674 = ~n16640 & n16673;
  assign n16675 = n16674 ^ n612;
  assign n16676 = n16675 ^ n16637;
  assign n16677 = n16638 & ~n16676;
  assign n16678 = n16677 ^ n662;
  assign n16636 = n16561 ^ n16546;
  assign n16679 = n16678 ^ n16636;
  assign n16680 = n16636 ^ n795;
  assign n16681 = n16679 & ~n16680;
  assign n16682 = n16681 ^ n795;
  assign n16683 = n16682 ^ n16634;
  assign n16684 = n16635 & ~n16683;
  assign n16685 = n16684 ^ n1143;
  assign n16633 = n16563 ^ n16544;
  assign n16686 = n16685 ^ n16633;
  assign n16687 = n16633 ^ n917;
  assign n16688 = n16686 & ~n16687;
  assign n16689 = n16688 ^ n917;
  assign n16690 = n16689 ^ n16631;
  assign n16691 = n16632 & ~n16690;
  assign n16692 = n16691 ^ n1135;
  assign n16630 = n16566 ^ n16565;
  assign n16693 = n16692 ^ n16630;
  assign n1164 = n1076 ^ x276;
  assign n1165 = n1164 ^ x468;
  assign n1166 = n1165 ^ x212;
  assign n16694 = n16630 ^ n1166;
  assign n16695 = ~n16693 & n16694;
  assign n16696 = n16695 ^ n1166;
  assign n16697 = n16696 ^ n16628;
  assign n16698 = ~n16629 & n16697;
  assign n16699 = n16698 ^ n1315;
  assign n16700 = n16699 ^ n16626;
  assign n16701 = n16627 & ~n16700;
  assign n16702 = n16701 ^ n3014;
  assign n16703 = n16702 ^ n16624;
  assign n16704 = ~n16625 & n16703;
  assign n16705 = n16704 ^ n3161;
  assign n16706 = n16705 ^ n2552;
  assign n16707 = ~n16623 & ~n16706;
  assign n16708 = n16707 ^ n16622;
  assign n16709 = n16708 ^ n2559;
  assign n16710 = n16621 & n16709;
  assign n16711 = n16710 ^ n16620;
  assign n16619 = n16574 ^ n16573;
  assign n16712 = n16711 ^ n16619;
  assign n16713 = n16619 ^ n2571;
  assign n16714 = ~n16712 & n16713;
  assign n16715 = n16714 ^ n2571;
  assign n16716 = n16715 ^ n16617;
  assign n16717 = ~n16618 & n16716;
  assign n16718 = n16717 ^ n1521;
  assign n16719 = n16718 ^ n16615;
  assign n16720 = n16616 & ~n16719;
  assign n16721 = n16720 ^ n2741;
  assign n16722 = n16721 ^ n16613;
  assign n16723 = ~n16614 & n16722;
  assign n16724 = n16723 ^ n1577;
  assign n16726 = n16725 ^ n16724;
  assign n16727 = n16725 ^ n2873;
  assign n16728 = n16726 & ~n16727;
  assign n16729 = n16728 ^ n2873;
  assign n16730 = n16729 ^ n16608;
  assign n16731 = n16612 & ~n16730;
  assign n16732 = n16731 ^ n16611;
  assign n16733 = n16732 ^ n16606;
  assign n16734 = ~n16607 & n16733;
  assign n16735 = n16734 ^ n1738;
  assign n16736 = n16735 ^ n16604;
  assign n16737 = n16605 & ~n16736;
  assign n16738 = n16737 ^ n1708;
  assign n16739 = n16738 ^ n16602;
  assign n16740 = ~n16603 & n16739;
  assign n16741 = n16740 ^ n1714;
  assign n16751 = n16741 ^ n16601;
  assign n16752 = ~n16750 & n16751;
  assign n16753 = n16752 ^ n1826;
  assign n16795 = n16753 ^ n1946;
  assign n16796 = n16771 & ~n16795;
  assign n16797 = n16796 ^ n16770;
  assign n16819 = n16797 ^ n16793;
  assign n16820 = n16794 & ~n16819;
  assign n16821 = n16820 ^ n1943;
  assign n16838 = n16837 ^ n16821;
  assign n16816 = n15323 ^ n14518;
  assign n16817 = n16816 ^ n16039;
  assign n16776 = n16041 ^ n15329;
  assign n16777 = n16776 ^ n14520;
  assign n16747 = n15332 ^ n14521;
  assign n16748 = n16747 ^ n16044;
  assign n16742 = n16741 ^ n1826;
  assign n16743 = n16742 ^ n16601;
  assign n16744 = n16284 ^ n15334;
  assign n16745 = n16744 ^ n14522;
  assign n16746 = ~n16743 & n16745;
  assign n16749 = n16748 ^ n16746;
  assign n16772 = n16771 ^ n16753;
  assign n16773 = n16772 ^ n16748;
  assign n16774 = ~n16749 & n16773;
  assign n16775 = n16774 ^ n16746;
  assign n16812 = n16777 ^ n16775;
  assign n16798 = n16797 ^ n16794;
  assign n16813 = n16798 ^ n16775;
  assign n16814 = n16812 & ~n16813;
  assign n16815 = n16814 ^ n16777;
  assign n16818 = n16817 ^ n16815;
  assign n16839 = n16838 ^ n16818;
  assign n16840 = n16839 ^ n14611;
  assign n16799 = n16798 ^ n16777;
  assign n16800 = n16799 ^ n16775;
  assign n16801 = n16800 ^ n14613;
  assign n16802 = n16745 ^ n16743;
  assign n16803 = ~n14626 & ~n16802;
  assign n16804 = n16803 ^ n14618;
  assign n16805 = n16772 ^ n16749;
  assign n16806 = n16805 ^ n16803;
  assign n16807 = ~n16804 & n16806;
  assign n16808 = n16807 ^ n14618;
  assign n16809 = n16808 ^ n16800;
  assign n16810 = n16801 & n16809;
  assign n16811 = n16810 ^ n14613;
  assign n16841 = n16840 ^ n16811;
  assign n16842 = n16802 ^ n14626;
  assign n16843 = n16805 ^ n16804;
  assign n16844 = n16842 & n16843;
  assign n16845 = n16808 ^ n16801;
  assign n16846 = n16844 & ~n16845;
  assign n16847 = n16841 & n16846;
  assign n16875 = n16839 ^ n16811;
  assign n16876 = n16840 & ~n16875;
  assign n16877 = n16876 ^ n14611;
  assign n16871 = n15322 ^ n14514;
  assign n16872 = n16871 ^ n16303;
  assign n16867 = n16830 ^ n16827;
  assign n16868 = ~n16831 & n16867;
  assign n16869 = n16868 ^ n16829;
  assign n16863 = n16832 ^ n16824;
  assign n16864 = ~n16833 & n16863;
  assign n16865 = n16864 ^ n13776;
  assign n16859 = n16836 ^ n16821;
  assign n16860 = ~n16837 & n16859;
  assign n16861 = n16860 ^ n2120;
  assign n16857 = n16219 ^ n1748;
  assign n16852 = n16834 & n16835;
  assign n16853 = n16852 ^ n684;
  assign n16854 = n16853 ^ n16261;
  assign n16855 = n16854 ^ n15664;
  assign n16856 = n16855 ^ n14523;
  assign n16858 = n16857 ^ n16856;
  assign n16862 = n16861 ^ n16858;
  assign n16866 = n16865 ^ n16862;
  assign n16870 = n16869 ^ n16866;
  assign n16873 = n16872 ^ n16870;
  assign n16848 = n16838 ^ n16817;
  assign n16849 = n16838 ^ n16815;
  assign n16850 = n16848 & n16849;
  assign n16851 = n16850 ^ n16817;
  assign n16874 = n16873 ^ n16851;
  assign n16878 = n16877 ^ n16874;
  assign n16879 = n16878 ^ n14606;
  assign n16923 = n16847 & n16879;
  assign n16918 = n15320 ^ n15105;
  assign n16919 = n16918 ^ n16310;
  assign n16917 = n16549 ^ n2327;
  assign n16920 = n16919 ^ n16917;
  assign n16914 = n16872 ^ n16851;
  assign n16915 = ~n16873 & ~n16914;
  assign n16916 = n16915 ^ n16870;
  assign n16921 = n16920 ^ n16916;
  assign n16910 = n16874 ^ n14606;
  assign n16911 = ~n16878 & n16910;
  assign n16912 = n16911 ^ n14606;
  assign n16913 = n16912 ^ n14598;
  assign n16922 = n16921 ^ n16913;
  assign n16924 = n16923 ^ n16922;
  assign n16925 = n16924 ^ n3264;
  assign n16880 = n16879 ^ n16847;
  assign n16884 = n16883 ^ n16880;
  assign n16885 = n16846 ^ n16841;
  assign n16886 = n16885 ^ n699;
  assign n16896 = n15248 ^ x318;
  assign n16897 = n16896 ^ x510;
  assign n16898 = n16897 ^ x254;
  assign n16890 = ~n16842 & n16889;
  assign n522 = n521 ^ x319;
  assign n523 = n522 ^ x511;
  assign n524 = n523 ^ x255;
  assign n16891 = n16890 ^ n524;
  assign n16892 = n16843 ^ n16842;
  assign n16893 = n16892 ^ n16890;
  assign n16894 = n16891 & ~n16893;
  assign n16895 = n16894 ^ n524;
  assign n16899 = n16898 ^ n16895;
  assign n16900 = n16845 ^ n16844;
  assign n16901 = n16900 ^ n16895;
  assign n16902 = n16899 & n16901;
  assign n16903 = n16902 ^ n16898;
  assign n16904 = n16903 ^ n16885;
  assign n16905 = n16886 & ~n16904;
  assign n16906 = n16905 ^ n699;
  assign n16907 = n16906 ^ n16880;
  assign n16908 = n16884 & ~n16907;
  assign n16909 = n16908 ^ n16883;
  assign n17389 = n16924 ^ n16909;
  assign n17390 = ~n16925 & n17389;
  assign n17391 = n17390 ^ n3264;
  assign n17522 = n17391 ^ n767;
  assign n17271 = ~n16922 & ~n16923;
  assign n17178 = n16921 ^ n14598;
  assign n17179 = n16921 ^ n16912;
  assign n17180 = n17178 & ~n17179;
  assign n17181 = n17180 ^ n14598;
  assign n17269 = n17181 ^ n14596;
  assign n17041 = n16917 ^ n16916;
  assign n17042 = n16920 & n17041;
  assign n17043 = n17042 ^ n16919;
  assign n17038 = n15316 ^ n15173;
  assign n17039 = n17038 ^ n16317;
  assign n17175 = n17043 ^ n17039;
  assign n17037 = n16656 ^ n16655;
  assign n17176 = n17175 ^ n17037;
  assign n17270 = n17269 ^ n17176;
  assign n17387 = n17271 ^ n17270;
  assign n17523 = n17522 ^ n17387;
  assign n17520 = n16030 ^ n15299;
  assign n17007 = n16689 ^ n16632;
  assign n17521 = n17520 ^ n17007;
  assign n17524 = n17523 ^ n17521;
  assign n16928 = n16686 ^ n917;
  assign n16927 = n16035 ^ n15303;
  assign n16929 = n16928 ^ n16927;
  assign n16926 = n16925 ^ n16909;
  assign n16930 = n16929 ^ n16926;
  assign n16934 = n16906 ^ n16884;
  assign n16932 = n16682 ^ n16635;
  assign n16931 = n16036 ^ n15305;
  assign n16933 = n16932 ^ n16931;
  assign n16935 = n16934 ^ n16933;
  assign n16939 = n16903 ^ n16886;
  assign n16937 = n16679 ^ n795;
  assign n16936 = n16345 ^ n15310;
  assign n16938 = n16937 ^ n16936;
  assign n16940 = n16939 ^ n16938;
  assign n16944 = n16900 ^ n16899;
  assign n16942 = n16675 ^ n16638;
  assign n16941 = n16338 ^ n15314;
  assign n16943 = n16942 ^ n16941;
  assign n16945 = n16944 ^ n16943;
  assign n16949 = n16892 ^ n16891;
  assign n16947 = n16672 ^ n16640;
  assign n16946 = n16331 ^ n15316;
  assign n16948 = n16947 ^ n16946;
  assign n16950 = n16949 ^ n16948;
  assign n16954 = n16889 ^ n16842;
  assign n16952 = n16669 ^ n580;
  assign n16951 = n16324 ^ n15320;
  assign n16953 = n16952 ^ n16951;
  assign n16955 = n16954 ^ n16953;
  assign n16964 = n15667 ^ n15034;
  assign n16965 = n16964 ^ n16246;
  assign n16963 = n16729 ^ n16612;
  assign n16966 = n16965 ^ n16963;
  assign n16971 = n15676 ^ n15043;
  assign n16972 = n16971 ^ n16857;
  assign n16969 = n16721 ^ n1577;
  assign n16970 = n16969 ^ n16613;
  assign n16973 = n16972 ^ n16970;
  assign n16976 = n16718 ^ n2741;
  assign n16977 = n16976 ^ n16615;
  assign n16974 = n16830 ^ n15669;
  assign n16975 = n16974 ^ n15036;
  assign n16978 = n16977 ^ n16975;
  assign n17101 = n16715 ^ n16618;
  assign n16981 = n16712 ^ n2571;
  assign n16979 = n16009 ^ n15553;
  assign n16980 = n16979 ^ n16765;
  assign n16982 = n16981 ^ n16980;
  assign n16985 = n16708 ^ n16621;
  assign n16983 = n16160 ^ n15437;
  assign n16984 = n16983 ^ n16598;
  assign n16986 = n16985 ^ n16984;
  assign n16988 = n16015 ^ n15342;
  assign n16989 = n16988 ^ n16401;
  assign n16987 = n16705 ^ n16623;
  assign n16990 = n16989 ^ n16987;
  assign n16992 = n16020 ^ n15424;
  assign n16993 = n16992 ^ n16008;
  assign n16991 = n16702 ^ n16625;
  assign n16994 = n16993 ^ n16991;
  assign n16996 = n16026 ^ n15417;
  assign n16997 = n16996 ^ n16013;
  assign n16995 = n16699 ^ n16627;
  assign n16998 = n16997 ^ n16995;
  assign n17001 = n16696 ^ n16629;
  assign n16999 = n16048 ^ n15343;
  assign n17000 = n16999 ^ n16014;
  assign n17002 = n17001 ^ n17000;
  assign n17005 = n16693 ^ n1166;
  assign n17003 = n16052 ^ n15296;
  assign n17004 = n17003 ^ n16019;
  assign n17006 = n17005 ^ n17004;
  assign n17008 = n16032 ^ n15398;
  assign n17009 = n17008 ^ n16024;
  assign n17010 = n17009 ^ n17007;
  assign n17011 = n16058 ^ n15301;
  assign n17012 = n17011 ^ n16373;
  assign n17013 = n17012 ^ n16928;
  assign n17014 = n16062 ^ n15307;
  assign n17015 = n17014 ^ n16029;
  assign n17016 = n17015 ^ n16932;
  assign n17017 = n15761 ^ n15350;
  assign n17018 = n17017 ^ n16030;
  assign n17019 = n17018 ^ n16937;
  assign n17020 = n15312 ^ n15294;
  assign n17021 = n17020 ^ n16035;
  assign n17022 = n17021 ^ n16942;
  assign n17023 = n15318 ^ n15303;
  assign n17024 = n17023 ^ n16345;
  assign n17025 = n17024 ^ n16952;
  assign n17026 = n15363 ^ n15305;
  assign n17027 = n17026 ^ n16338;
  assign n16957 = n16665 ^ n16643;
  assign n17028 = n17027 ^ n16957;
  assign n17031 = n16662 ^ n16645;
  assign n17029 = n15325 ^ n15310;
  assign n17030 = n17029 ^ n16331;
  assign n17032 = n17031 ^ n17030;
  assign n17034 = n15314 ^ n15213;
  assign n17035 = n17034 ^ n16324;
  assign n17033 = n16659 ^ n16650;
  assign n17036 = n17035 ^ n17033;
  assign n17040 = n17039 ^ n17037;
  assign n17044 = n17043 ^ n17037;
  assign n17045 = n17040 & ~n17044;
  assign n17046 = n17045 ^ n17039;
  assign n17047 = n17046 ^ n17033;
  assign n17048 = ~n17036 & n17047;
  assign n17049 = n17048 ^ n17035;
  assign n17050 = n17049 ^ n17031;
  assign n17051 = ~n17032 & ~n17050;
  assign n17052 = n17051 ^ n17030;
  assign n17053 = n17052 ^ n16957;
  assign n17054 = n17028 & ~n17053;
  assign n17055 = n17054 ^ n17027;
  assign n17056 = n17055 ^ n16952;
  assign n17057 = ~n17025 & ~n17056;
  assign n17058 = n17057 ^ n17024;
  assign n17059 = n17058 ^ n16947;
  assign n17060 = n15357 ^ n15299;
  assign n17061 = n17060 ^ n16036;
  assign n17062 = n17061 ^ n16947;
  assign n17063 = ~n17059 & ~n17062;
  assign n17064 = n17063 ^ n17061;
  assign n17065 = n17064 ^ n16942;
  assign n17066 = n17022 & ~n17065;
  assign n17067 = n17066 ^ n17021;
  assign n17068 = n17067 ^ n16937;
  assign n17069 = ~n17019 & n17068;
  assign n17070 = n17069 ^ n17018;
  assign n17071 = n17070 ^ n16932;
  assign n17072 = n17016 & ~n17071;
  assign n17073 = n17072 ^ n17015;
  assign n17074 = n17073 ^ n16928;
  assign n17075 = n17013 & n17074;
  assign n17076 = n17075 ^ n17012;
  assign n17077 = n17076 ^ n17007;
  assign n17078 = n17010 & n17077;
  assign n17079 = n17078 ^ n17009;
  assign n17080 = n17079 ^ n17005;
  assign n17081 = ~n17006 & ~n17080;
  assign n17082 = n17081 ^ n17004;
  assign n17083 = n17082 ^ n17001;
  assign n17084 = n17002 & ~n17083;
  assign n17085 = n17084 ^ n17000;
  assign n17086 = n17085 ^ n16995;
  assign n17087 = n16998 & n17086;
  assign n17088 = n17087 ^ n16997;
  assign n17089 = n17088 ^ n16991;
  assign n17090 = ~n16994 & n17089;
  assign n17091 = n17090 ^ n16993;
  assign n17092 = n17091 ^ n16987;
  assign n17093 = ~n16990 & n17092;
  assign n17094 = n17093 ^ n16989;
  assign n17095 = n17094 ^ n16985;
  assign n17096 = n16986 & n17095;
  assign n17097 = n17096 ^ n16984;
  assign n17098 = n17097 ^ n16981;
  assign n17099 = ~n16982 & n17098;
  assign n17100 = n17099 ^ n16980;
  assign n17102 = n17101 ^ n17100;
  assign n17103 = n16267 ^ n15568;
  assign n17104 = n17103 ^ n16783;
  assign n17105 = n17104 ^ n17101;
  assign n17106 = ~n17102 & n17105;
  assign n17107 = n17106 ^ n17104;
  assign n17108 = n17107 ^ n16977;
  assign n17109 = n16978 & n17108;
  assign n17110 = n17109 ^ n16975;
  assign n17111 = n17110 ^ n16972;
  assign n17112 = ~n16973 & ~n17111;
  assign n17113 = n17112 ^ n16970;
  assign n16967 = n16724 ^ n2873;
  assign n16968 = n16967 ^ n16725;
  assign n17114 = n17113 ^ n16968;
  assign n17115 = n15668 ^ n15035;
  assign n17116 = n17115 ^ n16239;
  assign n17117 = n17116 ^ n16968;
  assign n17118 = ~n17114 & ~n17117;
  assign n17119 = n17118 ^ n17116;
  assign n17120 = n17119 ^ n16963;
  assign n17121 = n16966 & ~n17120;
  assign n17122 = n17121 ^ n16965;
  assign n16961 = n15664 ^ n15033;
  assign n16962 = n16961 ^ n16237;
  assign n17123 = n17122 ^ n16962;
  assign n16959 = n16732 ^ n1738;
  assign n16960 = n16959 ^ n16606;
  assign n17124 = n17123 ^ n16960;
  assign n17125 = n17124 ^ n14387;
  assign n17126 = n17119 ^ n16966;
  assign n17127 = n17126 ^ n14392;
  assign n17130 = n17107 ^ n16975;
  assign n17131 = n17130 ^ n16977;
  assign n17132 = n17131 ^ n14407;
  assign n17133 = n17104 ^ n17102;
  assign n17134 = n17133 ^ n14524;
  assign n17135 = n17097 ^ n16982;
  assign n17136 = n17135 ^ n14715;
  assign n17137 = n17094 ^ n16986;
  assign n17138 = n17137 ^ n14707;
  assign n17139 = n17091 ^ n16989;
  assign n17140 = n17139 ^ n16987;
  assign n17141 = n17140 ^ n14532;
  assign n17142 = n17088 ^ n16993;
  assign n17143 = n17142 ^ n16991;
  assign n17144 = n17143 ^ n14534;
  assign n17147 = n17082 ^ n17002;
  assign n17148 = n17147 ^ n14544;
  assign n17149 = n17079 ^ n17004;
  assign n17150 = n17149 ^ n17005;
  assign n17151 = n17150 ^ n14549;
  assign n17152 = n17076 ^ n17009;
  assign n17153 = n17152 ^ n17007;
  assign n17154 = n17153 ^ n14684;
  assign n17155 = n17073 ^ n17012;
  assign n17156 = n17155 ^ n16928;
  assign n17157 = n17156 ^ n14676;
  assign n17158 = n17070 ^ n17016;
  assign n17159 = n17158 ^ n14554;
  assign n17160 = n17067 ^ n17019;
  assign n17161 = n17160 ^ n14559;
  assign n17162 = n17064 ^ n17022;
  assign n17163 = n17162 ^ n14567;
  assign n17164 = n17061 ^ n17059;
  assign n17165 = n17164 ^ n14569;
  assign n17168 = n17052 ^ n17028;
  assign n17169 = n17168 ^ n14582;
  assign n17170 = n17049 ^ n17032;
  assign n17171 = n17170 ^ n14516;
  assign n17172 = n17046 ^ n17035;
  assign n17173 = n17172 ^ n17033;
  assign n17174 = n17173 ^ n14591;
  assign n17177 = n17176 ^ n14596;
  assign n17182 = n17181 ^ n17176;
  assign n17183 = ~n17177 & n17182;
  assign n17184 = n17183 ^ n14596;
  assign n17185 = n17184 ^ n17173;
  assign n17186 = n17174 & ~n17185;
  assign n17187 = n17186 ^ n14591;
  assign n17188 = n17187 ^ n17170;
  assign n17189 = ~n17171 & ~n17188;
  assign n17190 = n17189 ^ n14516;
  assign n17191 = n17190 ^ n17168;
  assign n17192 = ~n17169 & n17191;
  assign n17193 = n17192 ^ n14582;
  assign n17166 = n17055 ^ n17024;
  assign n17167 = n17166 ^ n16952;
  assign n17194 = n17193 ^ n17167;
  assign n17195 = n17167 ^ n14577;
  assign n17196 = ~n17194 & ~n17195;
  assign n17197 = n17196 ^ n14577;
  assign n17198 = n17197 ^ n17164;
  assign n17199 = ~n17165 & ~n17198;
  assign n17200 = n17199 ^ n14569;
  assign n17201 = n17200 ^ n17162;
  assign n17202 = n17163 & n17201;
  assign n17203 = n17202 ^ n14567;
  assign n17204 = n17203 ^ n17160;
  assign n17205 = n17161 & n17204;
  assign n17206 = n17205 ^ n14559;
  assign n17207 = n17206 ^ n17158;
  assign n17208 = ~n17159 & n17207;
  assign n17209 = n17208 ^ n14554;
  assign n17210 = n17209 ^ n17156;
  assign n17211 = ~n17157 & n17210;
  assign n17212 = n17211 ^ n14676;
  assign n17213 = n17212 ^ n17153;
  assign n17214 = ~n17154 & ~n17213;
  assign n17215 = n17214 ^ n14684;
  assign n17216 = n17215 ^ n17150;
  assign n17217 = n17151 & n17216;
  assign n17218 = n17217 ^ n14549;
  assign n17219 = n17218 ^ n17147;
  assign n17220 = n17148 & ~n17219;
  assign n17221 = n17220 ^ n14544;
  assign n17145 = n17085 ^ n16997;
  assign n17146 = n17145 ^ n16995;
  assign n17222 = n17221 ^ n17146;
  assign n17223 = n17146 ^ n14539;
  assign n17224 = ~n17222 & n17223;
  assign n17225 = n17224 ^ n14539;
  assign n17226 = n17225 ^ n17143;
  assign n17227 = ~n17144 & ~n17226;
  assign n17228 = n17227 ^ n14534;
  assign n17229 = n17228 ^ n17140;
  assign n17230 = n17141 & n17229;
  assign n17231 = n17230 ^ n14532;
  assign n17232 = n17231 ^ n17137;
  assign n17233 = n17138 & n17232;
  assign n17234 = n17233 ^ n14707;
  assign n17235 = n17234 ^ n17135;
  assign n17236 = ~n17136 & ~n17235;
  assign n17237 = n17236 ^ n14715;
  assign n17238 = n17237 ^ n17133;
  assign n17239 = n17134 & ~n17238;
  assign n17240 = n17239 ^ n14524;
  assign n17241 = n17240 ^ n17131;
  assign n17242 = ~n17132 & ~n17241;
  assign n17243 = n17242 ^ n14407;
  assign n17129 = n17110 ^ n16973;
  assign n17244 = n17243 ^ n17129;
  assign n17245 = n17129 ^ n14405;
  assign n17246 = n17244 & n17245;
  assign n17247 = n17246 ^ n14405;
  assign n17128 = n17116 ^ n17114;
  assign n17248 = n17247 ^ n17128;
  assign n17249 = n17128 ^ n14397;
  assign n17250 = n17248 & n17249;
  assign n17251 = n17250 ^ n14397;
  assign n17252 = n17251 ^ n17126;
  assign n17253 = ~n17127 & ~n17252;
  assign n17254 = n17253 ^ n14392;
  assign n17321 = n17254 ^ n17124;
  assign n17322 = ~n17125 & ~n17321;
  assign n17323 = n17322 ^ n14387;
  assign n17314 = n16962 ^ n16960;
  assign n17315 = n17122 ^ n16960;
  assign n17316 = ~n17314 & n17315;
  assign n17317 = n17316 ^ n16962;
  assign n17313 = n16735 ^ n16605;
  assign n17318 = n17317 ^ n17313;
  assign n17311 = n15339 ^ n15065;
  assign n17312 = n17311 ^ n16234;
  assign n17319 = n17318 ^ n17312;
  assign n17320 = n17319 ^ n14451;
  assign n17324 = n17323 ^ n17320;
  assign n17255 = n17254 ^ n17125;
  assign n17256 = n17248 ^ n14397;
  assign n17257 = n17244 ^ n14405;
  assign n17258 = n17237 ^ n17134;
  assign n17259 = n17231 ^ n14707;
  assign n17260 = n17259 ^ n17137;
  assign n17261 = n17228 ^ n17141;
  assign n17262 = n17222 ^ n14539;
  assign n17263 = n17218 ^ n14544;
  assign n17264 = n17263 ^ n17147;
  assign n17265 = n17209 ^ n14676;
  assign n17266 = n17265 ^ n17156;
  assign n17267 = n17194 ^ n14577;
  assign n17268 = n17187 ^ n17171;
  assign n17272 = ~n17270 & ~n17271;
  assign n17273 = n17184 ^ n17174;
  assign n17274 = ~n17272 & ~n17273;
  assign n17275 = n17268 & n17274;
  assign n17276 = n17190 ^ n17169;
  assign n17277 = n17275 & ~n17276;
  assign n17278 = n17267 & ~n17277;
  assign n17279 = n17197 ^ n17165;
  assign n17280 = ~n17278 & n17279;
  assign n17281 = n17200 ^ n17163;
  assign n17282 = ~n17280 & ~n17281;
  assign n17283 = n17203 ^ n17161;
  assign n17284 = ~n17282 & ~n17283;
  assign n17285 = n17206 ^ n17159;
  assign n17286 = n17284 & ~n17285;
  assign n17287 = ~n17266 & n17286;
  assign n17288 = n17212 ^ n14684;
  assign n17289 = n17288 ^ n17153;
  assign n17290 = n17287 & ~n17289;
  assign n17291 = n17215 ^ n17151;
  assign n17292 = ~n17290 & n17291;
  assign n17293 = ~n17264 & n17292;
  assign n17294 = n17262 & ~n17293;
  assign n17295 = n17225 ^ n17144;
  assign n17296 = n17294 & ~n17295;
  assign n17297 = n17261 & ~n17296;
  assign n17298 = n17260 & ~n17297;
  assign n17299 = n17234 ^ n14715;
  assign n17300 = n17299 ^ n17135;
  assign n17301 = n17298 & n17300;
  assign n17302 = ~n17258 & ~n17301;
  assign n17303 = n17240 ^ n17132;
  assign n17304 = ~n17302 & ~n17303;
  assign n17305 = ~n17257 & n17304;
  assign n17306 = n17256 & n17305;
  assign n17307 = n17251 ^ n14392;
  assign n17308 = n17307 ^ n17126;
  assign n17309 = ~n17306 & ~n17308;
  assign n17310 = ~n17255 & ~n17309;
  assign n17340 = n17324 ^ n17310;
  assign n17341 = n17340 ^ n2064;
  assign n17342 = n17309 ^ n17255;
  assign n17343 = n17342 ^ n2052;
  assign n17344 = n17308 ^ n17306;
  assign n17345 = n17344 ^ n1930;
  assign n17346 = n17305 ^ n17256;
  assign n17347 = n17346 ^ n1910;
  assign n17348 = n17304 ^ n17257;
  assign n17349 = n17348 ^ n1917;
  assign n17350 = n17303 ^ n17302;
  assign n17351 = n17350 ^ n1658;
  assign n17352 = n17301 ^ n17258;
  assign n17356 = n17355 ^ n17352;
  assign n17357 = n17300 ^ n17298;
  assign n17358 = n17357 ^ n1541;
  assign n17359 = n17297 ^ n17260;
  assign n17360 = n17359 ^ n1591;
  assign n17361 = n17296 ^ n17261;
  assign n17362 = n17361 ^ n1496;
  assign n17364 = n17293 ^ n17262;
  assign n17365 = n17364 ^ n2708;
  assign n17366 = n17292 ^ n17264;
  assign n17367 = n17366 ^ n2711;
  assign n17368 = n17291 ^ n17290;
  assign n17369 = n17368 ^ n2495;
  assign n17370 = n17289 ^ n17287;
  assign n17371 = n17370 ^ n3038;
  assign n17373 = n17285 ^ n17284;
  assign n1374 = n1268 ^ x306;
  assign n1375 = n1374 ^ x498;
  assign n1376 = n1375 ^ x242;
  assign n17374 = n17373 ^ n1376;
  assign n17375 = n17283 ^ n17282;
  assign n1456 = n1344 ^ x307;
  assign n1457 = n1456 ^ x499;
  assign n1458 = n1457 ^ x243;
  assign n17376 = n17375 ^ n1458;
  assign n17377 = n17281 ^ n17280;
  assign n1174 = n1083 ^ x308;
  assign n1175 = n1174 ^ x500;
  assign n1176 = n1175 ^ x244;
  assign n17378 = n17377 ^ n1176;
  assign n17379 = n17279 ^ n17278;
  assign n17380 = n17379 ^ n1012;
  assign n17383 = n17274 ^ n17268;
  assign n17384 = n17383 ^ n786;
  assign n17385 = n17273 ^ n17272;
  assign n17386 = n17385 ^ n773;
  assign n17388 = n17387 ^ n767;
  assign n17392 = n17391 ^ n17387;
  assign n17393 = n17388 & ~n17392;
  assign n17394 = n17393 ^ n767;
  assign n17395 = n17394 ^ n17385;
  assign n17396 = ~n17386 & n17395;
  assign n17397 = n17396 ^ n773;
  assign n17398 = n17397 ^ n17383;
  assign n17399 = ~n17384 & n17398;
  assign n17400 = n17399 ^ n786;
  assign n17382 = n17276 ^ n17275;
  assign n17401 = n17400 ^ n17382;
  assign n17402 = n17382 ^ n872;
  assign n17403 = ~n17401 & n17402;
  assign n17404 = n17403 ^ n872;
  assign n17381 = n17277 ^ n17267;
  assign n17405 = n17404 ^ n17381;
  assign n1004 = n922 ^ x310;
  assign n1005 = n1004 ^ x502;
  assign n1006 = n1005 ^ x246;
  assign n17406 = n17381 ^ n1006;
  assign n17407 = n17405 & ~n17406;
  assign n17408 = n17407 ^ n1006;
  assign n17409 = n17408 ^ n17379;
  assign n17410 = n17380 & ~n17409;
  assign n17411 = n17410 ^ n1012;
  assign n17412 = n17411 ^ n17377;
  assign n17413 = n17378 & ~n17412;
  assign n17414 = n17413 ^ n1176;
  assign n17415 = n17414 ^ n17375;
  assign n17416 = ~n17376 & n17415;
  assign n17417 = n17416 ^ n1458;
  assign n17418 = n17417 ^ n17373;
  assign n17419 = n17374 & ~n17418;
  assign n17420 = n17419 ^ n1376;
  assign n17372 = n17286 ^ n17266;
  assign n17421 = n17420 ^ n17372;
  assign n2434 = n2412 ^ x305;
  assign n2435 = n2434 ^ x497;
  assign n2436 = n2435 ^ x241;
  assign n17422 = n17372 ^ n2436;
  assign n17423 = ~n17421 & n17422;
  assign n17424 = n17423 ^ n2436;
  assign n17425 = n17424 ^ n17370;
  assign n17426 = n17371 & ~n17425;
  assign n17427 = n17426 ^ n3038;
  assign n17428 = n17427 ^ n17368;
  assign n17429 = ~n17369 & n17428;
  assign n17430 = n17429 ^ n2495;
  assign n17431 = n17430 ^ n17366;
  assign n17432 = ~n17367 & n17431;
  assign n17433 = n17432 ^ n2711;
  assign n17434 = n17433 ^ n17364;
  assign n17435 = n17365 & ~n17434;
  assign n17436 = n17435 ^ n2708;
  assign n17363 = n17295 ^ n17294;
  assign n17437 = n17436 ^ n17363;
  assign n17438 = n17363 ^ n2728;
  assign n17439 = ~n17437 & n17438;
  assign n17440 = n17439 ^ n2728;
  assign n17441 = n17440 ^ n17361;
  assign n17442 = ~n17362 & n17441;
  assign n17443 = n17442 ^ n1496;
  assign n17444 = n17443 ^ n17359;
  assign n17445 = n17360 & ~n17444;
  assign n17446 = n17445 ^ n1591;
  assign n17447 = n17446 ^ n17357;
  assign n17448 = ~n17358 & n17447;
  assign n17449 = n17448 ^ n1541;
  assign n17450 = n17449 ^ n17352;
  assign n17451 = n17356 & ~n17450;
  assign n17452 = n17451 ^ n17355;
  assign n17453 = n17452 ^ n17350;
  assign n17454 = ~n17351 & n17453;
  assign n17455 = n17454 ^ n1658;
  assign n17456 = n17455 ^ n17348;
  assign n17457 = n17349 & ~n17456;
  assign n17458 = n17457 ^ n1917;
  assign n17459 = n17458 ^ n17346;
  assign n17460 = ~n17347 & n17459;
  assign n17461 = n17460 ^ n1910;
  assign n17462 = n17461 ^ n17344;
  assign n17463 = n17345 & ~n17462;
  assign n17464 = n17463 ^ n1930;
  assign n17465 = n17464 ^ n17342;
  assign n17466 = ~n17343 & n17465;
  assign n17467 = n17466 ^ n2052;
  assign n17468 = n17467 ^ n17340;
  assign n17469 = ~n17341 & n17468;
  assign n17470 = n17469 ^ n2064;
  assign n17471 = n17470 ^ n2208;
  assign n17334 = n17323 ^ n17319;
  assign n17335 = ~n17320 & n17334;
  assign n17336 = n17335 ^ n14451;
  assign n17337 = n17336 ^ n14506;
  assign n17329 = n17313 ^ n17312;
  assign n17330 = ~n17318 & ~n17329;
  assign n17331 = n17330 ^ n17312;
  assign n17327 = n15337 ^ n14523;
  assign n17328 = n17327 ^ n16280;
  assign n17332 = n17331 ^ n17328;
  assign n17326 = n16738 ^ n16603;
  assign n17333 = n17332 ^ n17326;
  assign n17338 = n17337 ^ n17333;
  assign n17325 = n17310 & n17324;
  assign n17339 = n17338 ^ n17325;
  assign n17472 = n17471 ^ n17339;
  assign n16956 = n16317 ^ n15322;
  assign n16958 = n16957 ^ n16956;
  assign n17473 = n17472 ^ n16958;
  assign n17476 = n17467 ^ n17341;
  assign n17474 = n16310 ^ n15323;
  assign n17475 = n17474 ^ n17031;
  assign n17477 = n17476 ^ n17475;
  assign n17483 = n16039 ^ n15332;
  assign n17484 = n17483 ^ n17037;
  assign n17479 = n17458 ^ n17347;
  assign n17480 = n16041 ^ n15334;
  assign n17481 = n17480 ^ n16917;
  assign n17482 = ~n17479 & ~n17481;
  assign n17485 = n17484 ^ n17482;
  assign n17486 = n17461 ^ n17345;
  assign n17487 = n17486 ^ n17484;
  assign n17488 = ~n17485 & n17487;
  assign n17489 = n17488 ^ n17482;
  assign n17478 = n17464 ^ n17343;
  assign n17490 = n17489 ^ n17478;
  assign n17491 = n16303 ^ n15329;
  assign n17492 = n17491 ^ n17033;
  assign n17493 = n17492 ^ n17478;
  assign n17494 = n17490 & n17493;
  assign n17495 = n17494 ^ n17492;
  assign n17496 = n17495 ^ n17476;
  assign n17497 = ~n17477 & ~n17496;
  assign n17498 = n17497 ^ n17475;
  assign n17499 = n17498 ^ n17472;
  assign n17500 = ~n17473 & ~n17499;
  assign n17501 = n17500 ^ n16958;
  assign n17502 = n17501 ^ n16954;
  assign n17503 = ~n16955 & ~n17502;
  assign n17504 = n17503 ^ n16953;
  assign n17505 = n17504 ^ n16949;
  assign n17506 = ~n16950 & ~n17505;
  assign n17507 = n17506 ^ n16948;
  assign n17508 = n17507 ^ n16944;
  assign n17509 = ~n16945 & ~n17508;
  assign n17510 = n17509 ^ n16943;
  assign n17511 = n17510 ^ n16939;
  assign n17512 = ~n16940 & ~n17511;
  assign n17513 = n17512 ^ n16938;
  assign n17514 = n17513 ^ n16934;
  assign n17515 = ~n16935 & n17514;
  assign n17516 = n17515 ^ n16933;
  assign n17517 = n17516 ^ n16926;
  assign n17518 = ~n16930 & ~n17517;
  assign n17519 = n17518 ^ n16929;
  assign n17589 = n17523 ^ n17519;
  assign n17590 = n17524 & ~n17589;
  assign n17591 = n17590 ^ n17521;
  assign n17586 = n16029 ^ n15294;
  assign n17587 = n17586 ^ n17005;
  assign n17585 = n17394 ^ n17386;
  assign n17588 = n17587 ^ n17585;
  assign n17592 = n17591 ^ n17588;
  assign n17628 = n17592 ^ n15312;
  assign n17525 = n17524 ^ n17519;
  assign n17526 = n17525 ^ n15357;
  assign n17527 = n17516 ^ n16929;
  assign n17528 = n17527 ^ n16926;
  assign n17529 = n17528 ^ n15318;
  assign n17531 = n17510 ^ n16940;
  assign n17532 = n17531 ^ n15325;
  assign n17533 = n17507 ^ n16945;
  assign n17534 = n17533 ^ n15213;
  assign n17535 = n17504 ^ n16950;
  assign n17536 = n17535 ^ n15173;
  assign n17537 = n17501 ^ n16953;
  assign n17538 = n17537 ^ n16954;
  assign n17539 = n17538 ^ n15105;
  assign n17541 = n17495 ^ n17477;
  assign n17542 = n17541 ^ n14518;
  assign n17543 = n17492 ^ n17490;
  assign n17544 = n17543 ^ n14520;
  assign n17545 = n17481 ^ n17479;
  assign n17546 = ~n14522 & n17545;
  assign n17547 = n17546 ^ n14521;
  assign n17548 = n17486 ^ n17485;
  assign n17549 = n17548 ^ n17546;
  assign n17550 = ~n17547 & n17549;
  assign n17551 = n17550 ^ n14521;
  assign n17552 = n17551 ^ n17543;
  assign n17553 = ~n17544 & n17552;
  assign n17554 = n17553 ^ n14520;
  assign n17555 = n17554 ^ n17541;
  assign n17556 = n17542 & n17555;
  assign n17557 = n17556 ^ n14518;
  assign n17540 = n17498 ^ n17473;
  assign n17558 = n17557 ^ n17540;
  assign n17559 = n17540 ^ n14514;
  assign n17560 = n17558 & n17559;
  assign n17561 = n17560 ^ n14514;
  assign n17562 = n17561 ^ n17538;
  assign n17563 = ~n17539 & n17562;
  assign n17564 = n17563 ^ n15105;
  assign n17565 = n17564 ^ n17535;
  assign n17566 = n17536 & ~n17565;
  assign n17567 = n17566 ^ n15173;
  assign n17568 = n17567 ^ n17533;
  assign n17569 = ~n17534 & n17568;
  assign n17570 = n17569 ^ n15213;
  assign n17571 = n17570 ^ n17531;
  assign n17572 = ~n17532 & ~n17571;
  assign n17573 = n17572 ^ n15325;
  assign n17530 = n17513 ^ n16935;
  assign n17574 = n17573 ^ n17530;
  assign n17575 = n17530 ^ n15363;
  assign n17576 = ~n17574 & n17575;
  assign n17577 = n17576 ^ n15363;
  assign n17578 = n17577 ^ n17528;
  assign n17579 = ~n17529 & ~n17578;
  assign n17580 = n17579 ^ n15318;
  assign n17581 = n17580 ^ n17525;
  assign n17582 = ~n17526 & n17581;
  assign n17583 = n17582 ^ n15357;
  assign n17629 = n17592 ^ n17583;
  assign n17630 = ~n17628 & ~n17629;
  assign n17631 = n17630 ^ n15312;
  assign n17626 = n17397 ^ n17384;
  assign n17623 = n16373 ^ n15761;
  assign n17624 = n17623 ^ n17001;
  assign n17619 = n17591 ^ n17587;
  assign n17620 = n17591 ^ n17585;
  assign n17621 = n17619 & n17620;
  assign n17622 = n17621 ^ n17587;
  assign n17625 = n17624 ^ n17622;
  assign n17627 = n17626 ^ n17625;
  assign n17632 = n17631 ^ n17627;
  assign n17894 = n17627 ^ n15350;
  assign n17895 = ~n17632 & n17894;
  assign n17896 = n17895 ^ n15350;
  assign n17954 = n17896 ^ n15307;
  assign n17810 = n17626 ^ n17624;
  assign n17811 = n17626 ^ n17622;
  assign n17812 = n17810 & n17811;
  assign n17813 = n17812 ^ n17624;
  assign n17807 = n16995 ^ n16024;
  assign n17808 = n17807 ^ n16062;
  assign n17891 = n17813 ^ n17808;
  assign n17731 = n17401 ^ n872;
  assign n17892 = n17891 ^ n17731;
  assign n17955 = n17954 ^ n17892;
  assign n17584 = n17583 ^ n15312;
  assign n17593 = n17592 ^ n17584;
  assign n17594 = n17577 ^ n17529;
  assign n17595 = n17574 ^ n15363;
  assign n17596 = n17545 ^ n14522;
  assign n17597 = n17548 ^ n17547;
  assign n17598 = ~n17596 & n17597;
  assign n17599 = n17551 ^ n17544;
  assign n17600 = n17598 & n17599;
  assign n17601 = n17554 ^ n17542;
  assign n17602 = n17600 & ~n17601;
  assign n17603 = n17558 ^ n14514;
  assign n17604 = n17602 & n17603;
  assign n17605 = n17561 ^ n15105;
  assign n17606 = n17605 ^ n17538;
  assign n17607 = ~n17604 & ~n17606;
  assign n17608 = n17564 ^ n17536;
  assign n17609 = ~n17607 & ~n17608;
  assign n17610 = n17567 ^ n17534;
  assign n17611 = ~n17609 & ~n17610;
  assign n17612 = n17570 ^ n17532;
  assign n17613 = n17611 & ~n17612;
  assign n17614 = ~n17595 & n17613;
  assign n17615 = ~n17594 & ~n17614;
  assign n17616 = n17580 ^ n17526;
  assign n17617 = ~n17615 & ~n17616;
  assign n17618 = n17593 & ~n17617;
  assign n17633 = n17632 ^ n15350;
  assign n17956 = ~n17618 & ~n17633;
  assign n17957 = ~n17955 & n17956;
  assign n17893 = n17892 ^ n15307;
  assign n17897 = n17896 ^ n17892;
  assign n17898 = n17893 & ~n17897;
  assign n17899 = n17898 ^ n15307;
  assign n17809 = n17808 ^ n17731;
  assign n17814 = n17813 ^ n17731;
  assign n17815 = ~n17809 & n17814;
  assign n17816 = n17815 ^ n17808;
  assign n17804 = n16058 ^ n16019;
  assign n17805 = n17804 ^ n16991;
  assign n17888 = n17816 ^ n17805;
  assign n17727 = n17405 ^ n1006;
  assign n17889 = n17888 ^ n17727;
  assign n17890 = n17889 ^ n15301;
  assign n17953 = n17899 ^ n17890;
  assign n18032 = n17957 ^ n17953;
  assign n18033 = n18032 ^ n2480;
  assign n18034 = n17956 ^ n17955;
  assign n3140 = n1381 ^ x338;
  assign n3141 = n3140 ^ n1299;
  assign n3142 = n3141 ^ x274;
  assign n18035 = n18034 ^ n3142;
  assign n17635 = n17617 ^ n17593;
  assign n1120 = n1032 ^ x340;
  assign n1121 = n1120 ^ n1114;
  assign n1122 = n1121 ^ x276;
  assign n17636 = n17635 ^ n1122;
  assign n17637 = n17616 ^ n17615;
  assign n1104 = n1020 ^ x341;
  assign n1105 = n1104 ^ n992;
  assign n1106 = n1105 ^ x277;
  assign n17638 = n17637 ^ n1106;
  assign n17639 = n17614 ^ n17594;
  assign n17640 = n17639 ^ n982;
  assign n17641 = n17613 ^ n17595;
  assign n17642 = n17641 ^ n966;
  assign n17643 = n17612 ^ n17611;
  assign n17644 = n17643 ^ n960;
  assign n17646 = n17608 ^ n17607;
  assign n17650 = n17649 ^ n17646;
  assign n17651 = n17606 ^ n17604;
  assign n17652 = n17651 ^ n569;
  assign n17653 = n17603 ^ n17602;
  assign n17654 = n17653 ^ n641;
  assign n17655 = n17601 ^ n17600;
  assign n538 = n534 ^ x349;
  assign n542 = n541 ^ n538;
  assign n543 = n542 ^ x285;
  assign n17656 = n17655 ^ n543;
  assign n17657 = n2350 & n17596;
  assign n17661 = n17660 ^ n17657;
  assign n17662 = n17597 ^ n17596;
  assign n17663 = n17662 ^ n17657;
  assign n17664 = n17661 & n17663;
  assign n17665 = n17664 ^ n17660;
  assign n17666 = n17665 ^ n3278;
  assign n17667 = n17599 ^ n17598;
  assign n17668 = n17667 ^ n17665;
  assign n17669 = n17666 & ~n17668;
  assign n17670 = n17669 ^ n3278;
  assign n17671 = n17670 ^ n17655;
  assign n17672 = ~n17656 & n17671;
  assign n17673 = n17672 ^ n543;
  assign n17674 = n17673 ^ n17653;
  assign n17675 = n17654 & ~n17674;
  assign n17676 = n17675 ^ n641;
  assign n17677 = n17676 ^ n17651;
  assign n17678 = ~n17652 & n17677;
  assign n17679 = n17678 ^ n569;
  assign n17680 = n17679 ^ n17646;
  assign n17681 = n17650 & ~n17680;
  assign n17682 = n17681 ^ n17649;
  assign n17645 = n17610 ^ n17609;
  assign n17683 = n17682 ^ n17645;
  assign n17684 = n17645 ^ n735;
  assign n17685 = n17683 & ~n17684;
  assign n17686 = n17685 ^ n735;
  assign n17687 = n17686 ^ n17643;
  assign n17688 = n17644 & ~n17687;
  assign n17689 = n17688 ^ n960;
  assign n17690 = n17689 ^ n17641;
  assign n17691 = n17642 & ~n17690;
  assign n17692 = n17691 ^ n966;
  assign n17693 = n17692 ^ n17639;
  assign n17694 = n17640 & ~n17693;
  assign n17695 = n17694 ^ n982;
  assign n17696 = n17695 ^ n17637;
  assign n17697 = ~n17638 & n17696;
  assign n17698 = n17697 ^ n1106;
  assign n17699 = n17698 ^ n17635;
  assign n17700 = ~n17636 & n17699;
  assign n17701 = n17700 ^ n1122;
  assign n17634 = n17633 ^ n17618;
  assign n17702 = n17701 ^ n17634;
  assign n18036 = n17634 ^ n1292;
  assign n18037 = n17702 & ~n18036;
  assign n18038 = n18037 ^ n1292;
  assign n18039 = n18038 ^ n18034;
  assign n18040 = n18035 & ~n18039;
  assign n18041 = n18040 ^ n3142;
  assign n18042 = n18041 ^ n18032;
  assign n18043 = ~n18033 & n18042;
  assign n18044 = n18043 ^ n2480;
  assign n17958 = n17953 & n17957;
  assign n17900 = n17899 ^ n17889;
  assign n17901 = ~n17890 & ~n17900;
  assign n17902 = n17901 ^ n15301;
  assign n17806 = n17805 ^ n17727;
  assign n17817 = n17816 ^ n17727;
  assign n17818 = ~n17806 & ~n17817;
  assign n17819 = n17818 ^ n17805;
  assign n17801 = n16987 ^ n16032;
  assign n17802 = n17801 ^ n16014;
  assign n17720 = n17408 ^ n17380;
  assign n17803 = n17802 ^ n17720;
  assign n17886 = n17819 ^ n17803;
  assign n17887 = n17886 ^ n15398;
  assign n17952 = n17902 ^ n17887;
  assign n18030 = n17958 ^ n17952;
  assign n2455 = n2447 ^ x336;
  assign n2459 = n2458 ^ n2455;
  assign n2460 = n2459 ^ x272;
  assign n18031 = n18030 ^ n2460;
  assign n18474 = n18044 ^ n18031;
  assign n18472 = n16963 ^ n16765;
  assign n17763 = n17440 ^ n1496;
  assign n17764 = n17763 ^ n17361;
  assign n18473 = n18472 ^ n17764;
  assign n18475 = n18474 ^ n18473;
  assign n18303 = n18041 ^ n2480;
  assign n18304 = n18303 ^ n18032;
  assign n18301 = n16968 ^ n16598;
  assign n17768 = n17437 ^ n2728;
  assign n18302 = n18301 ^ n17768;
  assign n18305 = n18304 ^ n18302;
  assign n18194 = n16970 ^ n16401;
  assign n17772 = n17433 ^ n17365;
  assign n18195 = n18194 ^ n17772;
  assign n18192 = n18038 ^ n3142;
  assign n18193 = n18192 ^ n18034;
  assign n18196 = n18195 ^ n18193;
  assign n17705 = n17430 ^ n17367;
  assign n17704 = n16977 ^ n16008;
  assign n17706 = n17705 ^ n17704;
  assign n17703 = n17702 ^ n1292;
  assign n17707 = n17706 ^ n17703;
  assign n18175 = n17695 ^ n1106;
  assign n18176 = n18175 ^ n17637;
  assign n17710 = n17421 ^ n2436;
  assign n17711 = n17710 ^ n16019;
  assign n17712 = n17711 ^ n16985;
  assign n17709 = n17692 ^ n17640;
  assign n17713 = n17712 ^ n17709;
  assign n17715 = n17417 ^ n17374;
  assign n17716 = n17715 ^ n16987;
  assign n17717 = n17716 ^ n16024;
  assign n17714 = n17689 ^ n17642;
  assign n17718 = n17717 ^ n17714;
  assign n18156 = n17683 ^ n735;
  assign n17723 = n17679 ^ n17649;
  assign n17724 = n17723 ^ n17646;
  assign n17721 = n17720 ^ n16030;
  assign n17722 = n17721 ^ n17001;
  assign n17725 = n17724 ^ n17722;
  assign n17728 = n17727 ^ n17005;
  assign n17729 = n17728 ^ n16035;
  assign n17726 = n17676 ^ n17652;
  assign n17730 = n17729 ^ n17726;
  assign n17734 = n17673 ^ n17654;
  assign n17732 = n17731 ^ n17007;
  assign n17733 = n17732 ^ n16036;
  assign n17735 = n17734 ^ n17733;
  assign n18139 = n17670 ^ n543;
  assign n18140 = n18139 ^ n17655;
  assign n17738 = n17667 ^ n17666;
  assign n17736 = n17585 ^ n16338;
  assign n17737 = n17736 ^ n16932;
  assign n17739 = n17738 ^ n17737;
  assign n17742 = n17662 ^ n17661;
  assign n17740 = n17523 ^ n16937;
  assign n17741 = n17740 ^ n16331;
  assign n17743 = n17742 ^ n17741;
  assign n17746 = n17596 ^ n2350;
  assign n17744 = n16942 ^ n16926;
  assign n17745 = n17744 ^ n16324;
  assign n17747 = n17746 ^ n17745;
  assign n18098 = n16947 ^ n16317;
  assign n18099 = n18098 ^ n16934;
  assign n17758 = n16743 ^ n16237;
  assign n17759 = n17758 ^ n15668;
  assign n17757 = n17443 ^ n17360;
  assign n17760 = n17759 ^ n17757;
  assign n17761 = n17326 ^ n16246;
  assign n17762 = n17761 ^ n15676;
  assign n17765 = n17764 ^ n17762;
  assign n17766 = n17313 ^ n15669;
  assign n17767 = n17766 ^ n16239;
  assign n17769 = n17768 ^ n17767;
  assign n17770 = n16960 ^ n16267;
  assign n17771 = n17770 ^ n16857;
  assign n17773 = n17772 ^ n17771;
  assign n17774 = n16963 ^ n16009;
  assign n17775 = n17774 ^ n16830;
  assign n17776 = n17775 ^ n17705;
  assign n17779 = n17427 ^ n2495;
  assign n17780 = n17779 ^ n17368;
  assign n17777 = n16968 ^ n16160;
  assign n17778 = n17777 ^ n16783;
  assign n17781 = n17780 ^ n17778;
  assign n17784 = n17424 ^ n17371;
  assign n17782 = n16970 ^ n16015;
  assign n17783 = n17782 ^ n16765;
  assign n17785 = n17784 ^ n17783;
  assign n17786 = n16598 ^ n16020;
  assign n17787 = n17786 ^ n16977;
  assign n17788 = n17787 ^ n17710;
  assign n17789 = n16401 ^ n16026;
  assign n17790 = n17789 ^ n17101;
  assign n17791 = n17790 ^ n17715;
  assign n17794 = n17414 ^ n1458;
  assign n17795 = n17794 ^ n17375;
  assign n17792 = n16981 ^ n16008;
  assign n17793 = n17792 ^ n16048;
  assign n17796 = n17795 ^ n17793;
  assign n17799 = n17411 ^ n17378;
  assign n17797 = n16985 ^ n16013;
  assign n17798 = n17797 ^ n16052;
  assign n17800 = n17799 ^ n17798;
  assign n17820 = n17819 ^ n17802;
  assign n17821 = ~n17803 & n17820;
  assign n17822 = n17821 ^ n17819;
  assign n17823 = n17822 ^ n17798;
  assign n17824 = n17800 & ~n17823;
  assign n17825 = n17824 ^ n17822;
  assign n17826 = n17825 ^ n17793;
  assign n17827 = ~n17796 & ~n17826;
  assign n17828 = n17827 ^ n17825;
  assign n17829 = n17828 ^ n17715;
  assign n17830 = n17791 & ~n17829;
  assign n17831 = n17830 ^ n17790;
  assign n17832 = n17831 ^ n17787;
  assign n17833 = ~n17788 & n17832;
  assign n17834 = n17833 ^ n17710;
  assign n17835 = n17834 ^ n17784;
  assign n17836 = n17785 & ~n17835;
  assign n17837 = n17836 ^ n17783;
  assign n17838 = n17837 ^ n17780;
  assign n17839 = ~n17781 & n17838;
  assign n17840 = n17839 ^ n17778;
  assign n17841 = n17840 ^ n17775;
  assign n17842 = n17776 & n17841;
  assign n17843 = n17842 ^ n17705;
  assign n17844 = n17843 ^ n17772;
  assign n17845 = ~n17773 & n17844;
  assign n17846 = n17845 ^ n17771;
  assign n17847 = n17846 ^ n17767;
  assign n17848 = ~n17769 & ~n17847;
  assign n17849 = n17848 ^ n17768;
  assign n17850 = n17849 ^ n17762;
  assign n17851 = n17765 & n17850;
  assign n17852 = n17851 ^ n17764;
  assign n17853 = n17852 ^ n17757;
  assign n17854 = n17760 & n17853;
  assign n17855 = n17854 ^ n17759;
  assign n17754 = n16234 ^ n15667;
  assign n17755 = n17754 ^ n16772;
  assign n17753 = n17446 ^ n17358;
  assign n17756 = n17755 ^ n17753;
  assign n17860 = n17855 ^ n17756;
  assign n17861 = n17860 ^ n15034;
  assign n17862 = n17852 ^ n17760;
  assign n17863 = n17862 ^ n15035;
  assign n17864 = n17849 ^ n17765;
  assign n17865 = n17864 ^ n15043;
  assign n17866 = n17846 ^ n17769;
  assign n17867 = n17866 ^ n15036;
  assign n17868 = n17843 ^ n17771;
  assign n17869 = n17868 ^ n17772;
  assign n17870 = n17869 ^ n15568;
  assign n17871 = n17840 ^ n17776;
  assign n17872 = n17871 ^ n15553;
  assign n17873 = n17837 ^ n17778;
  assign n17874 = n17873 ^ n17780;
  assign n17875 = n17874 ^ n15437;
  assign n17876 = n17834 ^ n17783;
  assign n17877 = n17876 ^ n17784;
  assign n17878 = n17877 ^ n15342;
  assign n17880 = n17828 ^ n17791;
  assign n17881 = n17880 ^ n15417;
  assign n17882 = n17825 ^ n17796;
  assign n17883 = n17882 ^ n15343;
  assign n17884 = n17822 ^ n17800;
  assign n17885 = n17884 ^ n15296;
  assign n17903 = n17902 ^ n17886;
  assign n17904 = ~n17887 & n17903;
  assign n17905 = n17904 ^ n15398;
  assign n17906 = n17905 ^ n17884;
  assign n17907 = n17885 & ~n17906;
  assign n17908 = n17907 ^ n15296;
  assign n17909 = n17908 ^ n17882;
  assign n17910 = n17883 & n17909;
  assign n17911 = n17910 ^ n15343;
  assign n17912 = n17911 ^ n17880;
  assign n17913 = n17881 & ~n17912;
  assign n17914 = n17913 ^ n15417;
  assign n17879 = n17831 ^ n17788;
  assign n17915 = n17914 ^ n17879;
  assign n17916 = n17879 ^ n15424;
  assign n17917 = n17915 & ~n17916;
  assign n17918 = n17917 ^ n15424;
  assign n17919 = n17918 ^ n17877;
  assign n17920 = ~n17878 & ~n17919;
  assign n17921 = n17920 ^ n15342;
  assign n17922 = n17921 ^ n17874;
  assign n17923 = n17875 & ~n17922;
  assign n17924 = n17923 ^ n15437;
  assign n17925 = n17924 ^ n17871;
  assign n17926 = ~n17872 & n17925;
  assign n17927 = n17926 ^ n15553;
  assign n17928 = n17927 ^ n17869;
  assign n17929 = n17870 & n17928;
  assign n17930 = n17929 ^ n15568;
  assign n17931 = n17930 ^ n17866;
  assign n17932 = ~n17867 & ~n17931;
  assign n17933 = n17932 ^ n15036;
  assign n17934 = n17933 ^ n17864;
  assign n17935 = ~n17865 & n17934;
  assign n17936 = n17935 ^ n15043;
  assign n17937 = n17936 ^ n17862;
  assign n17938 = ~n17863 & ~n17937;
  assign n17939 = n17938 ^ n15035;
  assign n17940 = n17939 ^ n17860;
  assign n17941 = ~n17861 & n17940;
  assign n17942 = n17941 ^ n15034;
  assign n17856 = n17855 ^ n17753;
  assign n17857 = ~n17756 & n17856;
  assign n17858 = n17857 ^ n17755;
  assign n17750 = n16798 ^ n15664;
  assign n17751 = n17750 ^ n16280;
  assign n17748 = n17449 ^ n17355;
  assign n17749 = n17748 ^ n17352;
  assign n17752 = n17751 ^ n17749;
  assign n17859 = n17858 ^ n17752;
  assign n17943 = n17942 ^ n17859;
  assign n17988 = n17859 ^ n15033;
  assign n17989 = n17943 & n17988;
  assign n17990 = n17989 ^ n15033;
  assign n17991 = n17990 ^ n15065;
  assign n17985 = n17452 ^ n17351;
  assign n17982 = n17858 ^ n17749;
  assign n17983 = ~n17752 & ~n17982;
  assign n17984 = n17983 ^ n17751;
  assign n17986 = n17985 ^ n17984;
  assign n17980 = n16838 ^ n16284;
  assign n17981 = n17980 ^ n15339;
  assign n17987 = n17986 ^ n17981;
  assign n17992 = n17991 ^ n17987;
  assign n17944 = n17943 ^ n15033;
  assign n17945 = n17939 ^ n17861;
  assign n17946 = n17933 ^ n17865;
  assign n17947 = n17930 ^ n17867;
  assign n17948 = n17924 ^ n15553;
  assign n17949 = n17948 ^ n17871;
  assign n17950 = n17905 ^ n15296;
  assign n17951 = n17950 ^ n17884;
  assign n17959 = ~n17952 & n17958;
  assign n17960 = ~n17951 & ~n17959;
  assign n17961 = n17908 ^ n17883;
  assign n17962 = n17960 & ~n17961;
  assign n17963 = n17911 ^ n17881;
  assign n17964 = ~n17962 & ~n17963;
  assign n17965 = n17915 ^ n15424;
  assign n17966 = n17964 & n17965;
  assign n17967 = n17918 ^ n17878;
  assign n17968 = ~n17966 & ~n17967;
  assign n17969 = n17921 ^ n17875;
  assign n17970 = ~n17968 & n17969;
  assign n17971 = ~n17949 & n17970;
  assign n17972 = n17927 ^ n17870;
  assign n17973 = ~n17971 & ~n17972;
  assign n17974 = n17947 & ~n17973;
  assign n17975 = ~n17946 & n17974;
  assign n17976 = n17936 ^ n17863;
  assign n17977 = n17975 & ~n17976;
  assign n17978 = ~n17945 & ~n17977;
  assign n17979 = ~n17944 & ~n17978;
  assign n18008 = n17992 ^ n17979;
  assign n18009 = n18008 ^ n2169;
  assign n18010 = n17978 ^ n17944;
  assign n18011 = n18010 ^ n1955;
  assign n18012 = n17977 ^ n17945;
  assign n18013 = n18012 ^ n2176;
  assign n18015 = n17974 ^ n17946;
  assign n18016 = n18015 ^ n1703;
  assign n18017 = n17973 ^ n17947;
  assign n1725 = n1663 ^ x327;
  assign n1726 = n1725 ^ n1651;
  assign n1727 = n1726 ^ x263;
  assign n18018 = n18017 ^ n1727;
  assign n18020 = n17969 ^ n17968;
  assign n18021 = n18020 ^ n2920;
  assign n18022 = n17967 ^ n17966;
  assign n18023 = n18022 ^ n2750;
  assign n18025 = n17963 ^ n17962;
  assign n18026 = n18025 ^ n2634;
  assign n18027 = n17961 ^ n17960;
  assign n18028 = n18027 ^ n1556;
  assign n18045 = n18044 ^ n18030;
  assign n18046 = n18031 & ~n18045;
  assign n18047 = n18046 ^ n2460;
  assign n18029 = n17959 ^ n17951;
  assign n18048 = n18047 ^ n18029;
  assign n2540 = n2500 ^ x335;
  assign n2541 = n2540 ^ n2464;
  assign n2542 = n2541 ^ x271;
  assign n18049 = n18029 ^ n2542;
  assign n18050 = ~n18048 & n18049;
  assign n18051 = n18050 ^ n2542;
  assign n18052 = n18051 ^ n18027;
  assign n18053 = ~n18028 & n18052;
  assign n18054 = n18053 ^ n1556;
  assign n18055 = n18054 ^ n18025;
  assign n18056 = ~n18026 & n18055;
  assign n18057 = n18056 ^ n2634;
  assign n18024 = n17965 ^ n17964;
  assign n18058 = n18057 ^ n18024;
  assign n18059 = n18024 ^ n2906;
  assign n18060 = n18058 & ~n18059;
  assign n18061 = n18060 ^ n2906;
  assign n18062 = n18061 ^ n18022;
  assign n18063 = n18023 & ~n18062;
  assign n18064 = n18063 ^ n2750;
  assign n18065 = n18064 ^ n18020;
  assign n18066 = n18021 & ~n18065;
  assign n18067 = n18066 ^ n2920;
  assign n18019 = n17970 ^ n17949;
  assign n18068 = n18067 ^ n18019;
  assign n18069 = n18019 ^ n1637;
  assign n18070 = ~n18068 & n18069;
  assign n18071 = n18070 ^ n1637;
  assign n18072 = n18071 ^ n1646;
  assign n18073 = n17972 ^ n17971;
  assign n18074 = n18073 ^ n18071;
  assign n18075 = n18072 & ~n18074;
  assign n18076 = n18075 ^ n1646;
  assign n18077 = n18076 ^ n1727;
  assign n18078 = n18018 & ~n18077;
  assign n18079 = n18078 ^ n18017;
  assign n18080 = n18079 ^ n18015;
  assign n18081 = n18016 & ~n18080;
  assign n18082 = n18081 ^ n1703;
  assign n18014 = n17976 ^ n17975;
  assign n18083 = n18082 ^ n18014;
  assign n18084 = n18014 ^ n1811;
  assign n18085 = ~n18083 & n18084;
  assign n18086 = n18085 ^ n1811;
  assign n18087 = n18086 ^ n18012;
  assign n18088 = n18013 & ~n18087;
  assign n18089 = n18088 ^ n2176;
  assign n18090 = n18089 ^ n18010;
  assign n18091 = ~n18011 & n18090;
  assign n18092 = n18091 ^ n1955;
  assign n18093 = n18092 ^ n18008;
  assign n18094 = ~n18009 & n18093;
  assign n18095 = n18094 ^ n2169;
  assign n2199 = n2107 ^ x321;
  assign n2200 = n2199 ^ n2129;
  assign n2201 = n2200 ^ x257;
  assign n18096 = n18095 ^ n2201;
  assign n18003 = n17985 ^ n17981;
  assign n18004 = ~n17986 & n18003;
  assign n18005 = n18004 ^ n17981;
  assign n17998 = n17987 ^ n15065;
  assign n17999 = n17990 ^ n17987;
  assign n18000 = n17998 & ~n17999;
  assign n18001 = n18000 ^ n15065;
  assign n17995 = n17327 ^ n16044;
  assign n17996 = n17995 ^ n16870;
  assign n17994 = n17455 ^ n17349;
  assign n17997 = n17996 ^ n17994;
  assign n18002 = n18001 ^ n17997;
  assign n18006 = n18005 ^ n18002;
  assign n17993 = n17979 & n17992;
  assign n18007 = n18006 ^ n17993;
  assign n18097 = n18096 ^ n18007;
  assign n18100 = n18099 ^ n18097;
  assign n18102 = n16952 ^ n16310;
  assign n18103 = n18102 ^ n16939;
  assign n18101 = n18092 ^ n18009;
  assign n18104 = n18103 ^ n18101;
  assign n18107 = n16957 ^ n16303;
  assign n18108 = n18107 ^ n16944;
  assign n18105 = n18089 ^ n1955;
  assign n18106 = n18105 ^ n18010;
  assign n18109 = n18108 ^ n18106;
  assign n18114 = n17031 ^ n16949;
  assign n18115 = n18114 ^ n16039;
  assign n18110 = n17033 ^ n16954;
  assign n18111 = n18110 ^ n16041;
  assign n18112 = n18083 ^ n1811;
  assign n18113 = ~n18111 & n18112;
  assign n18116 = n18115 ^ n18113;
  assign n18117 = n18086 ^ n18013;
  assign n18118 = n18117 ^ n18115;
  assign n18119 = ~n18116 & n18118;
  assign n18120 = n18119 ^ n18113;
  assign n18121 = n18120 ^ n18106;
  assign n18122 = n18109 & n18121;
  assign n18123 = n18122 ^ n18108;
  assign n18124 = n18123 ^ n18101;
  assign n18125 = ~n18104 & ~n18124;
  assign n18126 = n18125 ^ n18103;
  assign n18127 = n18126 ^ n18097;
  assign n18128 = ~n18100 & n18127;
  assign n18129 = n18128 ^ n18099;
  assign n18130 = n18129 ^ n17746;
  assign n18131 = ~n17747 & ~n18130;
  assign n18132 = n18131 ^ n17745;
  assign n18133 = n18132 ^ n17742;
  assign n18134 = ~n17743 & ~n18133;
  assign n18135 = n18134 ^ n17741;
  assign n18136 = n18135 ^ n17737;
  assign n18137 = ~n17739 & n18136;
  assign n18138 = n18137 ^ n17738;
  assign n18141 = n18140 ^ n18138;
  assign n18142 = n17626 ^ n16345;
  assign n18143 = n18142 ^ n16928;
  assign n18144 = n18143 ^ n18140;
  assign n18145 = n18141 & n18144;
  assign n18146 = n18145 ^ n18143;
  assign n18147 = n18146 ^ n17734;
  assign n18148 = ~n17735 & n18147;
  assign n18149 = n18148 ^ n17733;
  assign n18150 = n18149 ^ n17726;
  assign n18151 = n17730 & ~n18150;
  assign n18152 = n18151 ^ n17729;
  assign n18153 = n18152 ^ n17724;
  assign n18154 = ~n17725 & n18153;
  assign n18155 = n18154 ^ n17722;
  assign n18157 = n18156 ^ n18155;
  assign n18158 = n17799 ^ n16029;
  assign n18159 = n18158 ^ n16995;
  assign n18160 = n18159 ^ n18156;
  assign n18161 = ~n18157 & ~n18160;
  assign n18162 = n18161 ^ n18159;
  assign n17719 = n17686 ^ n17644;
  assign n18163 = n18162 ^ n17719;
  assign n18164 = n17795 ^ n16991;
  assign n18165 = n18164 ^ n16373;
  assign n18166 = n18165 ^ n17719;
  assign n18167 = ~n18163 & n18166;
  assign n18168 = n18167 ^ n18165;
  assign n18169 = n18168 ^ n17714;
  assign n18170 = n17718 & ~n18169;
  assign n18171 = n18170 ^ n17717;
  assign n18172 = n18171 ^ n17712;
  assign n18173 = n17713 & ~n18172;
  assign n18174 = n18173 ^ n17709;
  assign n18177 = n18176 ^ n18174;
  assign n18178 = n16981 ^ n16014;
  assign n18179 = n18178 ^ n17784;
  assign n18180 = n18179 ^ n18176;
  assign n18181 = n18177 & n18180;
  assign n18182 = n18181 ^ n18179;
  assign n17708 = n17698 ^ n17636;
  assign n18183 = n18182 ^ n17708;
  assign n18184 = n17780 ^ n16013;
  assign n18185 = n18184 ^ n17101;
  assign n18186 = n18185 ^ n17708;
  assign n18187 = ~n18183 & n18186;
  assign n18188 = n18187 ^ n18185;
  assign n18189 = n18188 ^ n17706;
  assign n18190 = ~n17707 & n18189;
  assign n18191 = n18190 ^ n17703;
  assign n18298 = n18195 ^ n18191;
  assign n18299 = ~n18196 & ~n18298;
  assign n18300 = n18299 ^ n18193;
  assign n18469 = n18304 ^ n18300;
  assign n18470 = n18305 & n18469;
  assign n18471 = n18470 ^ n18302;
  assign n18476 = n18475 ^ n18471;
  assign n18306 = n18305 ^ n18300;
  assign n18307 = n18306 ^ n16020;
  assign n18199 = n18185 ^ n18183;
  assign n18200 = n18199 ^ n16052;
  assign n18202 = n18171 ^ n17713;
  assign n18203 = n18202 ^ n16058;
  assign n18204 = n18168 ^ n17717;
  assign n18205 = n18204 ^ n17714;
  assign n18206 = n18205 ^ n16062;
  assign n18207 = n18165 ^ n18163;
  assign n18208 = n18207 ^ n15761;
  assign n18210 = n18152 ^ n17725;
  assign n18211 = n18210 ^ n15299;
  assign n18212 = n18149 ^ n17730;
  assign n18213 = n18212 ^ n15303;
  assign n18215 = n18143 ^ n18141;
  assign n18216 = n18215 ^ n15310;
  assign n18217 = n18135 ^ n17739;
  assign n18218 = n18217 ^ n15314;
  assign n18219 = n18132 ^ n17741;
  assign n18220 = n18219 ^ n17742;
  assign n18221 = n18220 ^ n15316;
  assign n18222 = n18129 ^ n17747;
  assign n18223 = n18222 ^ n15320;
  assign n18224 = n18126 ^ n18100;
  assign n18225 = n18224 ^ n15322;
  assign n18226 = n18123 ^ n18103;
  assign n18227 = n18226 ^ n18101;
  assign n18228 = n18227 ^ n15323;
  assign n18229 = n18120 ^ n18108;
  assign n18230 = n18229 ^ n18106;
  assign n18231 = n18230 ^ n15329;
  assign n18232 = n18112 ^ n18111;
  assign n18233 = n15334 & ~n18232;
  assign n18234 = n18233 ^ n15332;
  assign n18235 = n18117 ^ n18116;
  assign n18236 = n18235 ^ n18233;
  assign n18237 = n18234 & n18236;
  assign n18238 = n18237 ^ n15332;
  assign n18239 = n18238 ^ n18230;
  assign n18240 = ~n18231 & ~n18239;
  assign n18241 = n18240 ^ n15329;
  assign n18242 = n18241 ^ n18227;
  assign n18243 = ~n18228 & n18242;
  assign n18244 = n18243 ^ n15323;
  assign n18245 = n18244 ^ n18224;
  assign n18246 = ~n18225 & ~n18245;
  assign n18247 = n18246 ^ n15322;
  assign n18248 = n18247 ^ n18222;
  assign n18249 = ~n18223 & n18248;
  assign n18250 = n18249 ^ n15320;
  assign n18251 = n18250 ^ n18220;
  assign n18252 = ~n18221 & ~n18251;
  assign n18253 = n18252 ^ n15316;
  assign n18254 = n18253 ^ n18217;
  assign n18255 = ~n18218 & ~n18254;
  assign n18256 = n18255 ^ n15314;
  assign n18257 = n18256 ^ n18215;
  assign n18258 = ~n18216 & ~n18257;
  assign n18259 = n18258 ^ n15310;
  assign n18214 = n18146 ^ n17735;
  assign n18260 = n18259 ^ n18214;
  assign n18261 = n18214 ^ n15305;
  assign n18262 = n18260 & n18261;
  assign n18263 = n18262 ^ n15305;
  assign n18264 = n18263 ^ n18212;
  assign n18265 = n18213 & n18264;
  assign n18266 = n18265 ^ n15303;
  assign n18267 = n18266 ^ n18210;
  assign n18268 = n18211 & n18267;
  assign n18269 = n18268 ^ n15299;
  assign n18209 = n18159 ^ n18157;
  assign n18270 = n18269 ^ n18209;
  assign n18271 = n18209 ^ n15294;
  assign n18272 = ~n18270 & n18271;
  assign n18273 = n18272 ^ n15294;
  assign n18274 = n18273 ^ n18207;
  assign n18275 = n18208 & ~n18274;
  assign n18276 = n18275 ^ n15761;
  assign n18277 = n18276 ^ n18205;
  assign n18278 = n18206 & ~n18277;
  assign n18279 = n18278 ^ n16062;
  assign n18280 = n18279 ^ n18202;
  assign n18281 = n18203 & ~n18280;
  assign n18282 = n18281 ^ n16058;
  assign n18201 = n18179 ^ n18177;
  assign n18283 = n18282 ^ n18201;
  assign n18284 = n18201 ^ n16032;
  assign n18285 = ~n18283 & n18284;
  assign n18286 = n18285 ^ n16032;
  assign n18287 = n18286 ^ n18199;
  assign n18288 = n18200 & n18287;
  assign n18289 = n18288 ^ n16052;
  assign n18198 = n18188 ^ n17707;
  assign n18290 = n18289 ^ n18198;
  assign n18291 = n18198 ^ n16048;
  assign n18292 = n18290 & n18291;
  assign n18293 = n18292 ^ n16048;
  assign n18197 = n18196 ^ n18191;
  assign n18294 = n18293 ^ n18197;
  assign n18295 = n18197 ^ n16026;
  assign n18296 = ~n18294 & ~n18295;
  assign n18297 = n18296 ^ n16026;
  assign n18465 = n18306 ^ n18297;
  assign n18466 = ~n18307 & n18465;
  assign n18467 = n18466 ^ n16020;
  assign n18468 = n18467 ^ n16015;
  assign n18477 = n18476 ^ n18468;
  assign n18308 = n18307 ^ n18297;
  assign n18309 = n18290 ^ n16048;
  assign n18310 = n18286 ^ n18200;
  assign n18311 = n18283 ^ n16032;
  assign n18312 = n18279 ^ n16058;
  assign n18313 = n18312 ^ n18202;
  assign n18314 = n18276 ^ n16062;
  assign n18315 = n18314 ^ n18205;
  assign n18316 = n18256 ^ n15310;
  assign n18317 = n18316 ^ n18215;
  assign n18318 = n18247 ^ n18223;
  assign n18319 = n18232 ^ n15334;
  assign n18320 = n18235 ^ n18234;
  assign n18321 = ~n18319 & ~n18320;
  assign n18322 = n18238 ^ n15329;
  assign n18323 = n18322 ^ n18230;
  assign n18324 = n18321 & ~n18323;
  assign n18325 = n18241 ^ n18228;
  assign n18326 = n18324 & n18325;
  assign n18327 = n18244 ^ n18225;
  assign n18328 = n18326 & n18327;
  assign n18329 = n18318 & ~n18328;
  assign n18330 = n18250 ^ n15316;
  assign n18331 = n18330 ^ n18220;
  assign n18332 = ~n18329 & ~n18331;
  assign n18333 = n18253 ^ n18218;
  assign n18334 = ~n18332 & ~n18333;
  assign n18335 = n18317 & n18334;
  assign n18336 = n18260 ^ n15305;
  assign n18337 = n18335 & n18336;
  assign n18338 = n18263 ^ n18213;
  assign n18339 = ~n18337 & n18338;
  assign n18340 = n18266 ^ n18211;
  assign n18341 = ~n18339 & n18340;
  assign n18342 = n18270 ^ n15294;
  assign n18343 = ~n18341 & n18342;
  assign n18344 = n18273 ^ n15761;
  assign n18345 = n18344 ^ n18207;
  assign n18346 = ~n18343 & ~n18345;
  assign n18347 = ~n18315 & n18346;
  assign n18348 = ~n18313 & n18347;
  assign n18349 = ~n18311 & n18348;
  assign n18350 = n18310 & ~n18349;
  assign n18351 = ~n18309 & n18350;
  assign n18352 = n18294 ^ n16026;
  assign n18353 = ~n18351 & n18352;
  assign n18464 = ~n18308 & n18353;
  assign n18478 = n18477 ^ n18464;
  assign n18479 = n18478 ^ n2815;
  assign n18354 = n18353 ^ n18308;
  assign n18355 = n18354 ^ n1524;
  assign n18356 = n18352 ^ n18351;
  assign n18357 = n18356 ^ n2622;
  assign n18359 = n18349 ^ n18310;
  assign n18360 = n18359 ^ n2609;
  assign n18361 = n18348 ^ n18311;
  assign n18362 = n18361 ^ n3173;
  assign n18363 = n18347 ^ n18313;
  assign n18364 = n18363 ^ n3020;
  assign n18365 = n18346 ^ n18315;
  assign n1424 = n1315 ^ x370;
  assign n1425 = n1424 ^ n1418;
  assign n1426 = n1425 ^ x306;
  assign n18366 = n18365 ^ n1426;
  assign n18367 = n18345 ^ n18343;
  assign n1260 = n1166 ^ x371;
  assign n1261 = n1260 ^ n1172;
  assign n1262 = n1261 ^ x307;
  assign n18368 = n18367 ^ n1262;
  assign n18369 = n18342 ^ n18341;
  assign n1242 = n1135 ^ x372;
  assign n1243 = n1242 ^ n1236;
  assign n1244 = n1243 ^ x308;
  assign n18370 = n18369 ^ n1244;
  assign n18371 = n18340 ^ n18339;
  assign n996 = n917 ^ x373;
  assign n1000 = n999 ^ n996;
  assign n1001 = n1000 ^ x309;
  assign n18372 = n18371 ^ n1001;
  assign n18373 = n18338 ^ n18337;
  assign n18374 = n18373 ^ n1226;
  assign n18375 = n18336 ^ n18335;
  assign n18376 = n18375 ^ n858;
  assign n18377 = n18334 ^ n18317;
  assign n18378 = n18377 ^ n760;
  assign n18380 = n18331 ^ n18329;
  assign n18381 = n18380 ^ n604;
  assign n18382 = n18328 ^ n18318;
  assign n18383 = n18382 ^ n595;
  assign n18384 = n18327 ^ n18326;
  assign n18385 = n18384 ^ n3254;
  assign n18386 = n18325 ^ n18324;
  assign n18390 = n18389 ^ n18386;
  assign n18391 = n18323 ^ n18321;
  assign n18395 = n18394 ^ n18391;
  assign n18397 = n2327 ^ x383;
  assign n18398 = n18397 ^ n13566;
  assign n18399 = n18398 ^ x319;
  assign n18396 = n687 & n18319;
  assign n18400 = n18399 ^ n18396;
  assign n18401 = n18320 ^ n18319;
  assign n18402 = n18401 ^ n18396;
  assign n18403 = n18400 & ~n18402;
  assign n18404 = n18403 ^ n18399;
  assign n18405 = n18404 ^ n18391;
  assign n18406 = ~n18395 & n18405;
  assign n18407 = n18406 ^ n18394;
  assign n18408 = n18407 ^ n18386;
  assign n18409 = n18390 & ~n18408;
  assign n18410 = n18409 ^ n18389;
  assign n18411 = n18410 ^ n18384;
  assign n18412 = n18385 & ~n18411;
  assign n18413 = n18412 ^ n3254;
  assign n18414 = n18413 ^ n18382;
  assign n18415 = n18383 & ~n18414;
  assign n18416 = n18415 ^ n595;
  assign n18417 = n18416 ^ n18380;
  assign n18418 = n18381 & ~n18417;
  assign n18419 = n18418 ^ n604;
  assign n18379 = n18333 ^ n18332;
  assign n18420 = n18419 ^ n18379;
  assign n18421 = n18379 ^ n751;
  assign n18422 = n18420 & ~n18421;
  assign n18423 = n18422 ^ n751;
  assign n18424 = n18423 ^ n18377;
  assign n18425 = ~n18378 & n18424;
  assign n18426 = n18425 ^ n760;
  assign n18427 = n18426 ^ n18375;
  assign n18428 = ~n18376 & n18427;
  assign n18429 = n18428 ^ n858;
  assign n18430 = n18429 ^ n18373;
  assign n18431 = ~n18374 & n18430;
  assign n18432 = n18431 ^ n1226;
  assign n18433 = n18432 ^ n18371;
  assign n18434 = n18372 & ~n18433;
  assign n18435 = n18434 ^ n1001;
  assign n18436 = n18435 ^ n18369;
  assign n18437 = ~n18370 & n18436;
  assign n18438 = n18437 ^ n1244;
  assign n18439 = n18438 ^ n18367;
  assign n18440 = ~n18368 & n18439;
  assign n18441 = n18440 ^ n1262;
  assign n18442 = n18441 ^ n18365;
  assign n18443 = n18366 & ~n18442;
  assign n18444 = n18443 ^ n1426;
  assign n18445 = n18444 ^ n18363;
  assign n18446 = n18364 & ~n18445;
  assign n18447 = n18446 ^ n3020;
  assign n18448 = n18447 ^ n18361;
  assign n18449 = n18362 & ~n18448;
  assign n18450 = n18449 ^ n3173;
  assign n18451 = n18450 ^ n18359;
  assign n18452 = ~n18360 & n18451;
  assign n18453 = n18452 ^ n2609;
  assign n18358 = n18350 ^ n18309;
  assign n18454 = n18453 ^ n18358;
  assign n2591 = n2559 ^ x366;
  assign n2595 = n2594 ^ n2591;
  assign n2596 = n2595 ^ x302;
  assign n18455 = n18358 ^ n2596;
  assign n18456 = n18454 & ~n18455;
  assign n18457 = n18456 ^ n2596;
  assign n18458 = n18457 ^ n18356;
  assign n18459 = n18357 & ~n18458;
  assign n18460 = n18459 ^ n2622;
  assign n18461 = n18460 ^ n18354;
  assign n18462 = n18355 & ~n18461;
  assign n18463 = n18462 ^ n1524;
  assign n18670 = n18478 ^ n18463;
  assign n18671 = ~n18479 & n18670;
  assign n18672 = n18671 ^ n2815;
  assign n18601 = ~n18464 & n18477;
  assign n18573 = n18476 ^ n16015;
  assign n18574 = n18476 ^ n18467;
  assign n18575 = ~n18573 & n18574;
  assign n18576 = n18575 ^ n16015;
  assign n18534 = n18474 ^ n18471;
  assign n18535 = ~n18475 & n18534;
  assign n18536 = n18535 ^ n18473;
  assign n18532 = n18048 ^ n2542;
  assign n18530 = n17757 ^ n16960;
  assign n18531 = n18530 ^ n16783;
  assign n18533 = n18532 ^ n18531;
  assign n18571 = n18536 ^ n18533;
  assign n18572 = n18571 ^ n16160;
  assign n18600 = n18576 ^ n18572;
  assign n18669 = n18601 ^ n18600;
  assign n18673 = n18672 ^ n18669;
  assign n18674 = n18669 ^ n1586;
  assign n18675 = n18673 & ~n18674;
  assign n18676 = n18675 ^ n1586;
  assign n18602 = ~n18600 & ~n18601;
  assign n18577 = n18576 ^ n18571;
  assign n18578 = ~n18572 & ~n18577;
  assign n18579 = n18578 ^ n16160;
  assign n18537 = n18536 ^ n18532;
  assign n18538 = n18533 & n18537;
  assign n18539 = n18538 ^ n18531;
  assign n18527 = n17753 ^ n17313;
  assign n18528 = n18527 ^ n16830;
  assign n18568 = n18539 ^ n18528;
  assign n18526 = n18051 ^ n18028;
  assign n18569 = n18568 ^ n18526;
  assign n18570 = n18569 ^ n16009;
  assign n18599 = n18579 ^ n18570;
  assign n18667 = n18602 ^ n18599;
  assign n18668 = n18667 ^ n2946;
  assign n19069 = n18676 ^ n18668;
  assign n19570 = n19069 ^ n17985;
  assign n18628 = n18076 ^ n18018;
  assign n19571 = n19570 ^ n18628;
  assign n18863 = n18304 ^ n16985;
  assign n18864 = n18863 ^ n17780;
  assign n18861 = n18429 ^ n18374;
  assign n18781 = n18426 ^ n858;
  assign n18782 = n18781 ^ n18375;
  assign n18488 = n18423 ^ n18378;
  assign n18486 = n17710 ^ n17703;
  assign n18487 = n18486 ^ n16991;
  assign n18489 = n18488 ^ n18487;
  assign n18492 = n18420 ^ n751;
  assign n18490 = n17715 ^ n16995;
  assign n18491 = n18490 ^ n17708;
  assign n18493 = n18492 ^ n18491;
  assign n18768 = n18416 ^ n18381;
  assign n18760 = n18413 ^ n595;
  assign n18761 = n18760 ^ n18382;
  assign n18495 = n17714 ^ n17007;
  assign n18496 = n18495 ^ n17720;
  assign n18494 = n18410 ^ n18385;
  assign n18497 = n18496 ^ n18494;
  assign n18502 = n18404 ^ n18394;
  assign n18503 = n18502 ^ n18391;
  assign n18500 = n18156 ^ n17731;
  assign n18501 = n18500 ^ n16932;
  assign n18504 = n18503 ^ n18501;
  assign n18741 = n18401 ^ n18400;
  assign n18507 = n18319 ^ n687;
  assign n18505 = n17726 ^ n16942;
  assign n18506 = n18505 ^ n17585;
  assign n18508 = n18507 ^ n18506;
  assign n18708 = n18140 ^ n16926;
  assign n18709 = n18708 ^ n16952;
  assign n18529 = n18528 ^ n18526;
  assign n18540 = n18539 ^ n18526;
  assign n18541 = ~n18529 & n18540;
  assign n18542 = n18541 ^ n18528;
  assign n18523 = n17749 ^ n16857;
  assign n18524 = n18523 ^ n17326;
  assign n18521 = n18054 ^ n2634;
  assign n18522 = n18521 ^ n18025;
  assign n18525 = n18524 ^ n18522;
  assign n18566 = n18542 ^ n18525;
  assign n18567 = n18566 ^ n16267;
  assign n18580 = n18579 ^ n18569;
  assign n18581 = ~n18570 & n18580;
  assign n18582 = n18581 ^ n16009;
  assign n18583 = n18582 ^ n18566;
  assign n18584 = n18567 & ~n18583;
  assign n18585 = n18584 ^ n16267;
  assign n18548 = n17985 ^ n16743;
  assign n18549 = n18548 ^ n16239;
  assign n18546 = n18058 ^ n2906;
  assign n18543 = n18542 ^ n18522;
  assign n18544 = n18525 & n18543;
  assign n18545 = n18544 ^ n18524;
  assign n18547 = n18546 ^ n18545;
  assign n18565 = n18549 ^ n18547;
  assign n18586 = n18585 ^ n18565;
  assign n18587 = n18565 ^ n15669;
  assign n18588 = n18586 & ~n18587;
  assign n18589 = n18588 ^ n15669;
  assign n18550 = n18549 ^ n18546;
  assign n18551 = ~n18547 & n18550;
  assign n18552 = n18551 ^ n18549;
  assign n18518 = n18061 ^ n2750;
  assign n18519 = n18518 ^ n18022;
  assign n18516 = n16772 ^ n16246;
  assign n18517 = n18516 ^ n17994;
  assign n18520 = n18519 ^ n18517;
  assign n18564 = n18552 ^ n18520;
  assign n18590 = n18589 ^ n18564;
  assign n18608 = n18590 ^ n15676;
  assign n18603 = n18599 & n18602;
  assign n18604 = n18582 ^ n18567;
  assign n18605 = ~n18603 & n18604;
  assign n18606 = n18586 ^ n15669;
  assign n18607 = ~n18605 & n18606;
  assign n18658 = n18608 ^ n18607;
  assign n18659 = n18658 ^ n1774;
  assign n18660 = n18606 ^ n18605;
  assign n18661 = n18660 ^ n1782;
  assign n18662 = n18604 ^ n18603;
  assign n18666 = n18665 ^ n18662;
  assign n18677 = n18676 ^ n18667;
  assign n18678 = ~n18668 & n18677;
  assign n18679 = n18678 ^ n2946;
  assign n18680 = n18679 ^ n18662;
  assign n18681 = ~n18666 & n18680;
  assign n18682 = n18681 ^ n18665;
  assign n18683 = n18682 ^ n18660;
  assign n18684 = n18661 & ~n18683;
  assign n18685 = n18684 ^ n1782;
  assign n18686 = n18685 ^ n18658;
  assign n18687 = ~n18659 & n18686;
  assign n18688 = n18687 ^ n1774;
  assign n18609 = n18607 & n18608;
  assign n18591 = n18564 ^ n15676;
  assign n18592 = ~n18590 & ~n18591;
  assign n18593 = n18592 ^ n15676;
  assign n18553 = n18552 ^ n18517;
  assign n18554 = ~n18520 & ~n18553;
  assign n18555 = n18554 ^ n18519;
  assign n18513 = n16798 ^ n16237;
  assign n18514 = n18513 ^ n17479;
  assign n18561 = n18555 ^ n18514;
  assign n18512 = n18064 ^ n18021;
  assign n18562 = n18561 ^ n18512;
  assign n18563 = n18562 ^ n15668;
  assign n18598 = n18593 ^ n18563;
  assign n18657 = n18609 ^ n18598;
  assign n18689 = n18688 ^ n18657;
  assign n18690 = n18657 ^ n1800;
  assign n18691 = n18689 & ~n18690;
  assign n18692 = n18691 ^ n1800;
  assign n18610 = n18598 & n18609;
  assign n18594 = n18593 ^ n18562;
  assign n18595 = n18563 & ~n18594;
  assign n18596 = n18595 ^ n15668;
  assign n18515 = n18514 ^ n18512;
  assign n18556 = n18555 ^ n18512;
  assign n18557 = ~n18515 & ~n18556;
  assign n18558 = n18557 ^ n18514;
  assign n18509 = n17486 ^ n16838;
  assign n18510 = n18509 ^ n16234;
  assign n18481 = n18068 ^ n1637;
  assign n18511 = n18510 ^ n18481;
  assign n18559 = n18558 ^ n18511;
  assign n18560 = n18559 ^ n15667;
  assign n18597 = n18596 ^ n18560;
  assign n18656 = n18610 ^ n18597;
  assign n18693 = n18692 ^ n18656;
  assign n18694 = n18656 ^ n1895;
  assign n18695 = ~n18693 & n18694;
  assign n18696 = n18695 ^ n1895;
  assign n18621 = n18596 ^ n18559;
  assign n18622 = n18560 & ~n18621;
  assign n18623 = n18622 ^ n15667;
  assign n18617 = n17478 ^ n16870;
  assign n18618 = n18617 ^ n16280;
  assign n18615 = n18073 ^ n18072;
  assign n18612 = n18558 ^ n18481;
  assign n18613 = n18511 & n18612;
  assign n18614 = n18613 ^ n18510;
  assign n18616 = n18615 ^ n18614;
  assign n18619 = n18618 ^ n18616;
  assign n18620 = n18619 ^ n15664;
  assign n18624 = n18623 ^ n18620;
  assign n18611 = ~n18597 & ~n18610;
  assign n18655 = n18624 ^ n18611;
  assign n18697 = n18696 ^ n18655;
  assign n18698 = n18655 ^ n2033;
  assign n18699 = ~n18697 & n18698;
  assign n18700 = n18699 ^ n2033;
  assign n18634 = n18623 ^ n18619;
  assign n18635 = n18620 & ~n18634;
  assign n18636 = n18635 ^ n15664;
  assign n18630 = n18618 ^ n18615;
  assign n18631 = ~n18616 & ~n18630;
  assign n18632 = n18631 ^ n18618;
  assign n18626 = n17476 ^ n16284;
  assign n18627 = n18626 ^ n16917;
  assign n18629 = n18628 ^ n18627;
  assign n18633 = n18632 ^ n18629;
  assign n18637 = n18636 ^ n18633;
  assign n18638 = n18637 ^ n15339;
  assign n18625 = ~n18611 & n18624;
  assign n18654 = n18638 ^ n18625;
  assign n18701 = n18700 ^ n18654;
  assign n18707 = n18701 ^ n2030;
  assign n18710 = n18709 ^ n18707;
  assign n18716 = n17742 ^ n17031;
  assign n18717 = n18716 ^ n16939;
  assign n18712 = n17746 ^ n16944;
  assign n18713 = n18712 ^ n17033;
  assign n18714 = n18689 ^ n1800;
  assign n18715 = ~n18713 & ~n18714;
  assign n18718 = n18717 ^ n18715;
  assign n18719 = n18693 ^ n1895;
  assign n18720 = n18719 ^ n18717;
  assign n18721 = n18718 & ~n18720;
  assign n18722 = n18721 ^ n18715;
  assign n18711 = n18697 ^ n2033;
  assign n18723 = n18722 ^ n18711;
  assign n18724 = n16957 ^ n16934;
  assign n18725 = n18724 ^ n17738;
  assign n18726 = n18725 ^ n18711;
  assign n18727 = ~n18723 & n18726;
  assign n18728 = n18727 ^ n18725;
  assign n18729 = n18728 ^ n18707;
  assign n18730 = n18710 & ~n18729;
  assign n18731 = n18730 ^ n18709;
  assign n18702 = n18654 ^ n2030;
  assign n18703 = ~n18701 & n18702;
  assign n18704 = n18703 ^ n2030;
  assign n18705 = n18704 ^ n2216;
  assign n18649 = n18633 ^ n15339;
  assign n18650 = n18637 & ~n18649;
  assign n18651 = n18650 ^ n15339;
  assign n18644 = n18632 ^ n18628;
  assign n18645 = ~n18629 & n18644;
  assign n18646 = n18645 ^ n18627;
  assign n18641 = n17472 ^ n17037;
  assign n18642 = n18641 ^ n16044;
  assign n18640 = n18079 ^ n18016;
  assign n18643 = n18642 ^ n18640;
  assign n18647 = n18646 ^ n18643;
  assign n18648 = n18647 ^ n15337;
  assign n18652 = n18651 ^ n18648;
  assign n18639 = n18625 & ~n18638;
  assign n18653 = n18652 ^ n18639;
  assign n18706 = n18705 ^ n18653;
  assign n18732 = n18731 ^ n18706;
  assign n18733 = n17523 ^ n16947;
  assign n18734 = n18733 ^ n17734;
  assign n18735 = n18734 ^ n18706;
  assign n18736 = n18732 & n18735;
  assign n18737 = n18736 ^ n18734;
  assign n18738 = n18737 ^ n18507;
  assign n18739 = n18508 & n18738;
  assign n18740 = n18739 ^ n18506;
  assign n18742 = n18741 ^ n18740;
  assign n18743 = n17724 ^ n16937;
  assign n18744 = n18743 ^ n17626;
  assign n18745 = n18744 ^ n18741;
  assign n18746 = ~n18742 & n18745;
  assign n18747 = n18746 ^ n18744;
  assign n18748 = n18747 ^ n18503;
  assign n18749 = n18504 & n18748;
  assign n18750 = n18749 ^ n18501;
  assign n18498 = n18407 ^ n18389;
  assign n18499 = n18498 ^ n18386;
  assign n18751 = n18750 ^ n18499;
  assign n18752 = n17727 ^ n16928;
  assign n18753 = n18752 ^ n17719;
  assign n18754 = n18753 ^ n18499;
  assign n18755 = n18751 & n18754;
  assign n18756 = n18755 ^ n18753;
  assign n18757 = n18756 ^ n18494;
  assign n18758 = n18497 & ~n18757;
  assign n18759 = n18758 ^ n18496;
  assign n18762 = n18761 ^ n18759;
  assign n18763 = n17709 ^ n17005;
  assign n18764 = n18763 ^ n17799;
  assign n18765 = n18764 ^ n18761;
  assign n18766 = ~n18762 & n18765;
  assign n18767 = n18766 ^ n18764;
  assign n18769 = n18768 ^ n18767;
  assign n18770 = n17795 ^ n17001;
  assign n18771 = n18770 ^ n18176;
  assign n18772 = n18771 ^ n18768;
  assign n18773 = ~n18769 & ~n18772;
  assign n18774 = n18773 ^ n18771;
  assign n18775 = n18774 ^ n18492;
  assign n18776 = n18493 & ~n18775;
  assign n18777 = n18776 ^ n18491;
  assign n18778 = n18777 ^ n18487;
  assign n18779 = ~n18489 & n18778;
  assign n18780 = n18779 ^ n18488;
  assign n18783 = n18782 ^ n18780;
  assign n18484 = n18193 ^ n17784;
  assign n18485 = n18484 ^ n16987;
  assign n18858 = n18782 ^ n18485;
  assign n18859 = ~n18783 & n18858;
  assign n18860 = n18859 ^ n18485;
  assign n18862 = n18861 ^ n18860;
  assign n18865 = n18864 ^ n18862;
  assign n18866 = n18865 ^ n16019;
  assign n18784 = n18783 ^ n18485;
  assign n18785 = n18784 ^ n16024;
  assign n18786 = n18777 ^ n18489;
  assign n18787 = n18786 ^ n16373;
  assign n18788 = n18774 ^ n18491;
  assign n18789 = n18788 ^ n18492;
  assign n18790 = n18789 ^ n16029;
  assign n18791 = n18771 ^ n18769;
  assign n18792 = n18791 ^ n16030;
  assign n18794 = n18756 ^ n18497;
  assign n18795 = n18794 ^ n16036;
  assign n18796 = n18753 ^ n18751;
  assign n18797 = n18796 ^ n16345;
  assign n18798 = n18747 ^ n18504;
  assign n18799 = n18798 ^ n16338;
  assign n18800 = n18744 ^ n18742;
  assign n18801 = n18800 ^ n16331;
  assign n18804 = n18734 ^ n18732;
  assign n18805 = n18804 ^ n16317;
  assign n18806 = n18728 ^ n18710;
  assign n18807 = n18806 ^ n16310;
  assign n18808 = n18725 ^ n18723;
  assign n18809 = n18808 ^ n16303;
  assign n18810 = n18714 ^ n18713;
  assign n18811 = n16041 & n18810;
  assign n18812 = n18811 ^ n16039;
  assign n18813 = n18719 ^ n18718;
  assign n18814 = n18813 ^ n18811;
  assign n18815 = n18812 & ~n18814;
  assign n18816 = n18815 ^ n16039;
  assign n18817 = n18816 ^ n18808;
  assign n18818 = n18809 & ~n18817;
  assign n18819 = n18818 ^ n16303;
  assign n18820 = n18819 ^ n18806;
  assign n18821 = n18807 & ~n18820;
  assign n18822 = n18821 ^ n16310;
  assign n18823 = n18822 ^ n18804;
  assign n18824 = ~n18805 & ~n18823;
  assign n18825 = n18824 ^ n16317;
  assign n18802 = n18737 ^ n18506;
  assign n18803 = n18802 ^ n18507;
  assign n18826 = n18825 ^ n18803;
  assign n18827 = n18803 ^ n16324;
  assign n18828 = ~n18826 & ~n18827;
  assign n18829 = n18828 ^ n16324;
  assign n18830 = n18829 ^ n18800;
  assign n18831 = ~n18801 & ~n18830;
  assign n18832 = n18831 ^ n16331;
  assign n18833 = n18832 ^ n18798;
  assign n18834 = n18799 & n18833;
  assign n18835 = n18834 ^ n16338;
  assign n18836 = n18835 ^ n18796;
  assign n18837 = n18797 & n18836;
  assign n18838 = n18837 ^ n16345;
  assign n18839 = n18838 ^ n18794;
  assign n18840 = ~n18795 & n18839;
  assign n18841 = n18840 ^ n16036;
  assign n18793 = n18764 ^ n18762;
  assign n18842 = n18841 ^ n18793;
  assign n18843 = n18793 ^ n16035;
  assign n18844 = n18842 & n18843;
  assign n18845 = n18844 ^ n16035;
  assign n18846 = n18845 ^ n18791;
  assign n18847 = ~n18792 & n18846;
  assign n18848 = n18847 ^ n16030;
  assign n18849 = n18848 ^ n18789;
  assign n18850 = ~n18790 & n18849;
  assign n18851 = n18850 ^ n16029;
  assign n18852 = n18851 ^ n18786;
  assign n18853 = n18787 & ~n18852;
  assign n18854 = n18853 ^ n16373;
  assign n18855 = n18854 ^ n18784;
  assign n18856 = n18785 & n18855;
  assign n18857 = n18856 ^ n16024;
  assign n18992 = n18865 ^ n18857;
  assign n18993 = n18866 & ~n18992;
  assign n18994 = n18993 ^ n16019;
  assign n18987 = n18864 ^ n18861;
  assign n18988 = ~n18862 & n18987;
  assign n18989 = n18988 ^ n18864;
  assign n18985 = n18432 ^ n18372;
  assign n18983 = n18474 ^ n16981;
  assign n18984 = n18983 ^ n17705;
  assign n18986 = n18985 ^ n18984;
  assign n18990 = n18989 ^ n18986;
  assign n18991 = n18990 ^ n16014;
  assign n18995 = n18994 ^ n18991;
  assign n18867 = n18866 ^ n18857;
  assign n18868 = n18854 ^ n18785;
  assign n18869 = n18851 ^ n18787;
  assign n18870 = n18845 ^ n18792;
  assign n18871 = n18842 ^ n16035;
  assign n18872 = n18838 ^ n18795;
  assign n18873 = n18835 ^ n18797;
  assign n18874 = n18810 ^ n16041;
  assign n18875 = n18813 ^ n18812;
  assign n18876 = n18874 & n18875;
  assign n18877 = n18816 ^ n18809;
  assign n18878 = n18876 & n18877;
  assign n18879 = n18819 ^ n18807;
  assign n18880 = n18878 & n18879;
  assign n18881 = n18822 ^ n18805;
  assign n18882 = n18880 & ~n18881;
  assign n18883 = n18826 ^ n16324;
  assign n18884 = ~n18882 & ~n18883;
  assign n18885 = n18829 ^ n18801;
  assign n18886 = ~n18884 & ~n18885;
  assign n18887 = n18832 ^ n18799;
  assign n18888 = ~n18886 & n18887;
  assign n18889 = ~n18873 & n18888;
  assign n18890 = ~n18872 & n18889;
  assign n18891 = ~n18871 & ~n18890;
  assign n18892 = n18870 & ~n18891;
  assign n18893 = n18848 ^ n18790;
  assign n18894 = ~n18892 & ~n18893;
  assign n18895 = ~n18869 & ~n18894;
  assign n18896 = ~n18868 & n18895;
  assign n18982 = n18867 & n18896;
  assign n18996 = n18995 ^ n18982;
  assign n2467 = n2436 ^ x400;
  assign n2471 = n2470 ^ n2467;
  assign n2472 = n2471 ^ x336;
  assign n18997 = n18996 ^ n2472;
  assign n18897 = n18896 ^ n18867;
  assign n2426 = n1376 ^ x401;
  assign n2427 = n2426 ^ n2423;
  assign n2428 = n2427 ^ x337;
  assign n18898 = n18897 ^ n2428;
  assign n18899 = n18895 ^ n18868;
  assign n2417 = n1458 ^ x402;
  assign n2418 = n2417 ^ n1279;
  assign n2419 = n2418 ^ x338;
  assign n18900 = n18899 ^ n2419;
  assign n18901 = n18894 ^ n18869;
  assign n1270 = n1176 ^ x403;
  assign n1274 = n1273 ^ n1270;
  assign n1275 = n1274 ^ x339;
  assign n18902 = n18901 ^ n1275;
  assign n18903 = n18893 ^ n18892;
  assign n18904 = n18903 ^ n1099;
  assign n18905 = n18891 ^ n18870;
  assign n1088 = n1006 ^ x405;
  assign n1089 = n1088 ^ n948;
  assign n1090 = n1089 ^ x341;
  assign n18906 = n18905 ^ n1090;
  assign n18909 = n18888 ^ n18873;
  assign n18910 = n18909 ^ n831;
  assign n18911 = n18887 ^ n18886;
  assign n18912 = n18911 ^ n822;
  assign n18913 = n18885 ^ n18884;
  assign n18914 = n18913 ^ n3270;
  assign n18915 = n18883 ^ n18882;
  assign n18919 = n18918 ^ n18915;
  assign n18922 = n16898 ^ x413;
  assign n18923 = n18922 ^ n635;
  assign n18924 = n18923 ^ x349;
  assign n18921 = n18879 ^ n18878;
  assign n18925 = n18924 ^ n18921;
  assign n18935 = n18877 ^ n18876;
  assign n18926 = n2310 & ~n18874;
  assign n18930 = n18929 ^ n18926;
  assign n18931 = n18875 ^ n18874;
  assign n18932 = n18931 ^ n18926;
  assign n18933 = n18930 & ~n18932;
  assign n18934 = n18933 ^ n18929;
  assign n18936 = n18935 ^ n18934;
  assign n525 = n524 ^ x414;
  assign n529 = n528 ^ n525;
  assign n530 = n529 ^ x350;
  assign n18937 = n18935 ^ n530;
  assign n18938 = ~n18936 & n18937;
  assign n18939 = n18938 ^ n530;
  assign n18940 = n18939 ^ n18921;
  assign n18941 = n18925 & ~n18940;
  assign n18942 = n18941 ^ n18924;
  assign n18920 = n18881 ^ n18880;
  assign n18943 = n18942 ^ n18920;
  assign n18944 = n18920 ^ n705;
  assign n18945 = n18943 & ~n18944;
  assign n18946 = n18945 ^ n705;
  assign n18947 = n18946 ^ n18915;
  assign n18948 = ~n18919 & n18947;
  assign n18949 = n18948 ^ n18918;
  assign n18950 = n18949 ^ n18913;
  assign n18951 = n18914 & ~n18950;
  assign n18952 = n18951 ^ n3270;
  assign n18953 = n18952 ^ n18911;
  assign n18954 = n18912 & ~n18953;
  assign n18955 = n18954 ^ n822;
  assign n18956 = n18955 ^ n18909;
  assign n18957 = n18910 & ~n18956;
  assign n18958 = n18957 ^ n831;
  assign n18908 = n18889 ^ n18872;
  assign n18959 = n18958 ^ n18908;
  assign n18960 = n18908 ^ n846;
  assign n18961 = ~n18959 & n18960;
  assign n18962 = n18961 ^ n846;
  assign n18907 = n18890 ^ n18871;
  assign n18963 = n18962 ^ n18907;
  assign n18964 = n18907 ^ n936;
  assign n18965 = ~n18963 & n18964;
  assign n18966 = n18965 ^ n936;
  assign n18967 = n18966 ^ n18905;
  assign n18968 = n18906 & ~n18967;
  assign n18969 = n18968 ^ n1090;
  assign n18970 = n18969 ^ n18903;
  assign n18971 = n18904 & ~n18970;
  assign n18972 = n18971 ^ n1099;
  assign n18973 = n18972 ^ n18901;
  assign n18974 = ~n18902 & n18973;
  assign n18975 = n18974 ^ n1275;
  assign n18976 = n18975 ^ n18899;
  assign n18977 = n18900 & ~n18976;
  assign n18978 = n18977 ^ n2419;
  assign n18979 = n18978 ^ n18897;
  assign n18980 = ~n18898 & n18979;
  assign n18981 = n18980 ^ n2428;
  assign n19297 = n18996 ^ n18981;
  assign n19298 = n18997 & ~n19297;
  assign n19299 = n19298 ^ n2472;
  assign n19245 = n18982 & ~n18995;
  assign n19185 = n18994 ^ n18990;
  assign n19186 = ~n18991 & n19185;
  assign n19187 = n19186 ^ n16014;
  assign n19093 = n18989 ^ n18984;
  assign n19094 = ~n18986 & ~n19093;
  assign n19095 = n19094 ^ n18985;
  assign n19090 = n18532 ^ n17772;
  assign n19091 = n19090 ^ n17101;
  assign n19089 = n18435 ^ n18370;
  assign n19092 = n19091 ^ n19089;
  assign n19183 = n19095 ^ n19092;
  assign n19184 = n19183 ^ n16013;
  assign n19244 = n19187 ^ n19184;
  assign n19296 = n19245 ^ n19244;
  assign n19300 = n19299 ^ n19296;
  assign n19301 = n19296 ^ n3050;
  assign n19302 = n19300 & ~n19301;
  assign n19303 = n19302 ^ n3050;
  assign n19246 = n19244 & ~n19245;
  assign n19188 = n19187 ^ n19183;
  assign n19189 = ~n19184 & n19188;
  assign n19190 = n19189 ^ n16013;
  assign n19242 = n19190 ^ n16008;
  assign n19100 = n17768 ^ n16977;
  assign n19101 = n19100 ^ n18526;
  assign n19096 = n19095 ^ n19089;
  assign n19097 = n19092 & n19096;
  assign n19098 = n19097 ^ n19091;
  assign n19030 = n18438 ^ n18368;
  assign n19099 = n19098 ^ n19030;
  assign n19181 = n19101 ^ n19099;
  assign n19243 = n19242 ^ n19181;
  assign n19294 = n19246 ^ n19243;
  assign n19295 = n19294 ^ n2537;
  assign n19568 = n19303 ^ n19295;
  assign n19447 = n19300 ^ n3050;
  assign n19138 = n18673 ^ n1586;
  assign n19445 = n19138 ^ n18615;
  assign n19446 = n19445 ^ n17749;
  assign n19448 = n19447 ^ n19446;
  assign n18998 = n18997 ^ n18981;
  assign n18480 = n18479 ^ n18463;
  assign n18482 = n18481 ^ n18480;
  assign n18483 = n18482 ^ n17753;
  assign n18999 = n18998 ^ n18483;
  assign n19004 = n18975 ^ n18900;
  assign n19001 = n18457 ^ n18357;
  assign n19002 = n19001 ^ n18519;
  assign n19003 = n19002 ^ n17764;
  assign n19005 = n19004 ^ n19003;
  assign n19009 = n18450 ^ n18360;
  assign n19010 = n19009 ^ n17772;
  assign n19011 = n19010 ^ n18522;
  assign n19007 = n18969 ^ n1099;
  assign n19008 = n19007 ^ n18903;
  assign n19012 = n19011 ^ n19008;
  assign n19014 = n18447 ^ n18362;
  assign n19015 = n19014 ^ n18526;
  assign n19016 = n19015 ^ n17705;
  assign n19013 = n18966 ^ n18906;
  assign n19017 = n19016 ^ n19013;
  assign n19019 = n18444 ^ n18364;
  assign n19020 = n19019 ^ n17780;
  assign n19021 = n19020 ^ n18532;
  assign n19018 = n18963 ^ n936;
  assign n19022 = n19021 ^ n19018;
  assign n19025 = n18474 ^ n17784;
  assign n19024 = n18441 ^ n18366;
  assign n19026 = n19025 ^ n19024;
  assign n19023 = n18959 ^ n846;
  assign n19027 = n19026 ^ n19023;
  assign n19031 = n19030 ^ n18304;
  assign n19032 = n19031 ^ n17710;
  assign n19028 = n18955 ^ n831;
  assign n19029 = n19028 ^ n18909;
  assign n19033 = n19032 ^ n19029;
  assign n19036 = n18985 ^ n17795;
  assign n19037 = n19036 ^ n17703;
  assign n19035 = n18949 ^ n18914;
  assign n19038 = n19037 ^ n19035;
  assign n19042 = n18782 ^ n18176;
  assign n19043 = n19042 ^ n17720;
  assign n19041 = n18943 ^ n705;
  assign n19044 = n19043 ^ n19041;
  assign n19047 = n18939 ^ n18925;
  assign n19045 = n18488 ^ n17709;
  assign n19046 = n19045 ^ n17727;
  assign n19048 = n19047 ^ n19046;
  assign n19051 = n18492 ^ n17731;
  assign n19052 = n19051 ^ n17714;
  assign n19049 = n18934 ^ n530;
  assign n19050 = n19049 ^ n18935;
  assign n19053 = n19052 ^ n19050;
  assign n19055 = n18768 ^ n17626;
  assign n19056 = n19055 ^ n17719;
  assign n19054 = n18931 ^ n18930;
  assign n19057 = n19056 ^ n19054;
  assign n19378 = n18874 ^ n2310;
  assign n19350 = n18741 ^ n18140;
  assign n19351 = n19350 ^ n16939;
  assign n19076 = n18615 ^ n17994;
  assign n19077 = n19076 ^ n17326;
  assign n19078 = n19077 ^ n19001;
  assign n19080 = n18481 ^ n17313;
  assign n19081 = n19080 ^ n17985;
  assign n19079 = n18454 ^ n2596;
  assign n19082 = n19081 ^ n19079;
  assign n19083 = n18519 ^ n16963;
  assign n19084 = n19083 ^ n17753;
  assign n19085 = n19084 ^ n19014;
  assign n19086 = n18546 ^ n17757;
  assign n19087 = n19086 ^ n16968;
  assign n19088 = n19087 ^ n19019;
  assign n19102 = n19101 ^ n19030;
  assign n19103 = ~n19099 & n19102;
  assign n19104 = n19103 ^ n19101;
  assign n19105 = n19104 ^ n19024;
  assign n19106 = n17764 ^ n16970;
  assign n19107 = n19106 ^ n18522;
  assign n19108 = n19107 ^ n19024;
  assign n19109 = n19105 & ~n19108;
  assign n19110 = n19109 ^ n19107;
  assign n19111 = n19110 ^ n19019;
  assign n19112 = n19088 & n19111;
  assign n19113 = n19112 ^ n19087;
  assign n19114 = n19113 ^ n19014;
  assign n19115 = ~n19085 & ~n19114;
  assign n19116 = n19115 ^ n19084;
  assign n19117 = n19116 ^ n19009;
  assign n19118 = n17749 ^ n16960;
  assign n19119 = n19118 ^ n18512;
  assign n19120 = n19119 ^ n19009;
  assign n19121 = ~n19117 & n19120;
  assign n19122 = n19121 ^ n19119;
  assign n19123 = n19122 ^ n19081;
  assign n19124 = n19082 & ~n19123;
  assign n19125 = n19124 ^ n19079;
  assign n19126 = n19125 ^ n19001;
  assign n19127 = ~n19078 & n19126;
  assign n19128 = n19127 ^ n19077;
  assign n19074 = n18460 ^ n1524;
  assign n19075 = n19074 ^ n18354;
  assign n19129 = n19128 ^ n19075;
  assign n19130 = n18628 ^ n16743;
  assign n19131 = n19130 ^ n17479;
  assign n19132 = n19131 ^ n19075;
  assign n19133 = n19129 & n19132;
  assign n19134 = n19133 ^ n19131;
  assign n19071 = n18640 ^ n16772;
  assign n19072 = n19071 ^ n17486;
  assign n19073 = n19072 ^ n18480;
  assign n19166 = n19134 ^ n19073;
  assign n19167 = n19166 ^ n16246;
  assign n19168 = n19131 ^ n19129;
  assign n19169 = n19168 ^ n16239;
  assign n19170 = n19125 ^ n19078;
  assign n19171 = n19170 ^ n16857;
  assign n19172 = n19122 ^ n19082;
  assign n19173 = n19172 ^ n16830;
  assign n19174 = n19119 ^ n19117;
  assign n19175 = n19174 ^ n16783;
  assign n19176 = n19113 ^ n19085;
  assign n19177 = n19176 ^ n16765;
  assign n19182 = n19181 ^ n16008;
  assign n19191 = n19190 ^ n19181;
  assign n19192 = n19182 & ~n19191;
  assign n19193 = n19192 ^ n16008;
  assign n19180 = n19107 ^ n19105;
  assign n19194 = n19193 ^ n19180;
  assign n19195 = n19180 ^ n16401;
  assign n19196 = n19194 & n19195;
  assign n19197 = n19196 ^ n16401;
  assign n19178 = n19110 ^ n19087;
  assign n19179 = n19178 ^ n19019;
  assign n19198 = n19197 ^ n19179;
  assign n19199 = n19179 ^ n16598;
  assign n19200 = n19198 & ~n19199;
  assign n19201 = n19200 ^ n16598;
  assign n19202 = n19201 ^ n19176;
  assign n19203 = ~n19177 & n19202;
  assign n19204 = n19203 ^ n16765;
  assign n19205 = n19204 ^ n19174;
  assign n19206 = n19175 & n19205;
  assign n19207 = n19206 ^ n16783;
  assign n19208 = n19207 ^ n19172;
  assign n19209 = n19173 & ~n19208;
  assign n19210 = n19209 ^ n16830;
  assign n19211 = n19210 ^ n19170;
  assign n19212 = n19171 & n19211;
  assign n19213 = n19212 ^ n16857;
  assign n19214 = n19213 ^ n19168;
  assign n19215 = n19169 & n19214;
  assign n19216 = n19215 ^ n16239;
  assign n19217 = n19216 ^ n19166;
  assign n19218 = n19167 & ~n19217;
  assign n19219 = n19218 ^ n16246;
  assign n19140 = n18112 ^ n16798;
  assign n19141 = n19140 ^ n17478;
  assign n19135 = n19134 ^ n18480;
  assign n19136 = ~n19073 & n19135;
  assign n19137 = n19136 ^ n19072;
  assign n19139 = n19138 ^ n19137;
  assign n19164 = n19141 ^ n19139;
  assign n19165 = n19164 ^ n16237;
  assign n19260 = n19219 ^ n19165;
  assign n19236 = n19210 ^ n19171;
  assign n19237 = n19204 ^ n16783;
  assign n19238 = n19237 ^ n19174;
  assign n19239 = n19201 ^ n16765;
  assign n19240 = n19239 ^ n19176;
  assign n19241 = n19198 ^ n16598;
  assign n19247 = ~n19243 & n19246;
  assign n19248 = n19194 ^ n16401;
  assign n19249 = ~n19247 & n19248;
  assign n19250 = n19241 & n19249;
  assign n19251 = ~n19240 & ~n19250;
  assign n19252 = ~n19238 & ~n19251;
  assign n19253 = n19207 ^ n19173;
  assign n19254 = n19252 & n19253;
  assign n19255 = ~n19236 & ~n19254;
  assign n19256 = n19213 ^ n19169;
  assign n19257 = ~n19255 & ~n19256;
  assign n19258 = n19216 ^ n19167;
  assign n19259 = n19257 & n19258;
  assign n19273 = n19260 ^ n19259;
  assign n19274 = n19273 ^ n1998;
  assign n19275 = n19258 ^ n19257;
  assign n19276 = n19275 ^ n1722;
  assign n19277 = n19256 ^ n19255;
  assign n19281 = n19280 ^ n19277;
  assign n19282 = n19254 ^ n19236;
  assign n19283 = n19282 ^ n1623;
  assign n19284 = n19253 ^ n19252;
  assign n19285 = n19284 ^ n1600;
  assign n19286 = n19251 ^ n19238;
  assign n19287 = n19286 ^ n1502;
  assign n19288 = n19250 ^ n19240;
  assign n19289 = n19288 ^ n2794;
  assign n19290 = n19249 ^ n19241;
  assign n19291 = n19290 ^ n2768;
  assign n19292 = n19248 ^ n19247;
  assign n19293 = n19292 ^ n2774;
  assign n19304 = n19303 ^ n19294;
  assign n19305 = ~n19295 & n19304;
  assign n19306 = n19305 ^ n2537;
  assign n19307 = n19306 ^ n19292;
  assign n19308 = n19293 & ~n19307;
  assign n19309 = n19308 ^ n2774;
  assign n19310 = n19309 ^ n19290;
  assign n19311 = ~n19291 & n19310;
  assign n19312 = n19311 ^ n2768;
  assign n19313 = n19312 ^ n19288;
  assign n19314 = n19289 & ~n19313;
  assign n19315 = n19314 ^ n2794;
  assign n19316 = n19315 ^ n19286;
  assign n19317 = ~n19287 & n19316;
  assign n19318 = n19317 ^ n1502;
  assign n19319 = n19318 ^ n19284;
  assign n19320 = ~n19285 & n19319;
  assign n19321 = n19320 ^ n1600;
  assign n19322 = n19321 ^ n1623;
  assign n19323 = n19283 & ~n19322;
  assign n19324 = n19323 ^ n19282;
  assign n19325 = n19324 ^ n19277;
  assign n19326 = ~n19281 & n19325;
  assign n19327 = n19326 ^ n19280;
  assign n19328 = n19327 ^ n19275;
  assign n19329 = ~n19276 & n19328;
  assign n19330 = n19329 ^ n1722;
  assign n19331 = n19330 ^ n1998;
  assign n19332 = ~n19274 & ~n19331;
  assign n19333 = n19332 ^ n19273;
  assign n19348 = n19333 ^ n1985;
  assign n19220 = n19219 ^ n19164;
  assign n19221 = n19165 & n19220;
  assign n19222 = n19221 ^ n16237;
  assign n19142 = n19141 ^ n19138;
  assign n19143 = n19139 & n19142;
  assign n19144 = n19143 ^ n19141;
  assign n19067 = n18117 ^ n16838;
  assign n19068 = n19067 ^ n17476;
  assign n19070 = n19069 ^ n19068;
  assign n19163 = n19144 ^ n19070;
  assign n19223 = n19222 ^ n19163;
  assign n19262 = n19223 ^ n16234;
  assign n19261 = n19259 & n19260;
  assign n19271 = n19262 ^ n19261;
  assign n19349 = n19348 ^ n19271;
  assign n19352 = n19351 ^ n19349;
  assign n19353 = n19330 ^ n19274;
  assign n19354 = n18507 ^ n16944;
  assign n19355 = n19354 ^ n17738;
  assign n19356 = ~n19353 & ~n19355;
  assign n19357 = n19356 ^ n19351;
  assign n19358 = ~n19352 & ~n19357;
  assign n19359 = n19358 ^ n19356;
  assign n19272 = n19271 ^ n1985;
  assign n19334 = n19333 ^ n19271;
  assign n19335 = n19272 & n19334;
  assign n19336 = n19335 ^ n1985;
  assign n19224 = n19163 ^ n16234;
  assign n19225 = ~n19223 & ~n19224;
  assign n19226 = n19225 ^ n16234;
  assign n19145 = n19144 ^ n19068;
  assign n19146 = ~n19070 & n19145;
  assign n19147 = n19146 ^ n19069;
  assign n19064 = n17472 ^ n16870;
  assign n19065 = n19064 ^ n18106;
  assign n19160 = n19147 ^ n19065;
  assign n19063 = n18679 ^ n18666;
  assign n19161 = n19160 ^ n19063;
  assign n19162 = n19161 ^ n16280;
  assign n19264 = n19226 ^ n19162;
  assign n19263 = ~n19261 & ~n19262;
  assign n19270 = n19264 ^ n19263;
  assign n19337 = n19336 ^ n19270;
  assign n19347 = n19337 ^ n2011;
  assign n19360 = n19359 ^ n19347;
  assign n19361 = n18503 ^ n16934;
  assign n19362 = n19361 ^ n17734;
  assign n19363 = n19362 ^ n19347;
  assign n19364 = n19360 & n19363;
  assign n19365 = n19364 ^ n19362;
  assign n19338 = n19270 ^ n2011;
  assign n19339 = n19337 & ~n19338;
  assign n19340 = n19339 ^ n2011;
  assign n19265 = ~n19263 & ~n19264;
  assign n19227 = n19226 ^ n19161;
  assign n19228 = ~n19162 & ~n19227;
  assign n19229 = n19228 ^ n16280;
  assign n19152 = n18101 ^ n16954;
  assign n19153 = n19152 ^ n16917;
  assign n19066 = n19065 ^ n19063;
  assign n19148 = n19147 ^ n19063;
  assign n19149 = n19066 & ~n19148;
  assign n19150 = n19149 ^ n19065;
  assign n19062 = n18682 ^ n18661;
  assign n19151 = n19150 ^ n19062;
  assign n19158 = n19153 ^ n19151;
  assign n19159 = n19158 ^ n16284;
  assign n19235 = n19229 ^ n19159;
  assign n19269 = n19265 ^ n19235;
  assign n19341 = n19340 ^ n19269;
  assign n19346 = n19341 ^ n2142;
  assign n19366 = n19365 ^ n19346;
  assign n19367 = n18499 ^ n16926;
  assign n19368 = n19367 ^ n17726;
  assign n19369 = n19368 ^ n19346;
  assign n19370 = ~n19366 & ~n19369;
  assign n19371 = n19370 ^ n19368;
  assign n19342 = n19269 ^ n2142;
  assign n19343 = n19341 & ~n19342;
  assign n19344 = n19343 ^ n2142;
  assign n19266 = n19235 & n19265;
  assign n19230 = n19229 ^ n19158;
  assign n19231 = ~n19159 & ~n19230;
  assign n19232 = n19231 ^ n16284;
  assign n19233 = n19232 ^ n16044;
  assign n19154 = n19153 ^ n19062;
  assign n19155 = n19151 & ~n19154;
  assign n19156 = n19155 ^ n19153;
  assign n19060 = n18685 ^ n18659;
  assign n19058 = n18097 ^ n16949;
  assign n19059 = n19058 ^ n17037;
  assign n19061 = n19060 ^ n19059;
  assign n19157 = n19156 ^ n19061;
  assign n19234 = n19233 ^ n19157;
  assign n19267 = n19266 ^ n19234;
  assign n19268 = n19267 ^ n2157;
  assign n19345 = n19344 ^ n19268;
  assign n19372 = n19371 ^ n19345;
  assign n19373 = n17724 ^ n17523;
  assign n19374 = n19373 ^ n18494;
  assign n19375 = n19374 ^ n19345;
  assign n19376 = ~n19372 & n19375;
  assign n19377 = n19376 ^ n19374;
  assign n19379 = n19378 ^ n19377;
  assign n19380 = n18761 ^ n18156;
  assign n19381 = n19380 ^ n17585;
  assign n19382 = n19381 ^ n19378;
  assign n19383 = n19379 & ~n19382;
  assign n19384 = n19383 ^ n19381;
  assign n19385 = n19384 ^ n19054;
  assign n19386 = ~n19057 & ~n19385;
  assign n19387 = n19386 ^ n19056;
  assign n19388 = n19387 ^ n19050;
  assign n19389 = ~n19053 & n19388;
  assign n19390 = n19389 ^ n19052;
  assign n19391 = n19390 ^ n19047;
  assign n19392 = n19048 & n19391;
  assign n19393 = n19392 ^ n19046;
  assign n19394 = n19393 ^ n19041;
  assign n19395 = ~n19044 & n19394;
  assign n19396 = n19395 ^ n19043;
  assign n19039 = n18946 ^ n18918;
  assign n19040 = n19039 ^ n18915;
  assign n19397 = n19396 ^ n19040;
  assign n19398 = n17799 ^ n17708;
  assign n19399 = n19398 ^ n18861;
  assign n19400 = n19399 ^ n19040;
  assign n19401 = n19397 & ~n19400;
  assign n19402 = n19401 ^ n19399;
  assign n19403 = n19402 ^ n19035;
  assign n19404 = n19038 & ~n19403;
  assign n19405 = n19404 ^ n19037;
  assign n19034 = n18952 ^ n18912;
  assign n19406 = n19405 ^ n19034;
  assign n19407 = n19089 ^ n18193;
  assign n19408 = n19407 ^ n17715;
  assign n19409 = n19408 ^ n19034;
  assign n19410 = ~n19406 & ~n19409;
  assign n19411 = n19410 ^ n19408;
  assign n19412 = n19411 ^ n19029;
  assign n19413 = n19033 & n19412;
  assign n19414 = n19413 ^ n19032;
  assign n19415 = n19414 ^ n19023;
  assign n19416 = n19027 & ~n19415;
  assign n19417 = n19416 ^ n19026;
  assign n19418 = n19417 ^ n19018;
  assign n19419 = ~n19022 & ~n19418;
  assign n19420 = n19419 ^ n19021;
  assign n19421 = n19420 ^ n19013;
  assign n19422 = n19017 & n19421;
  assign n19423 = n19422 ^ n19016;
  assign n19424 = n19423 ^ n19011;
  assign n19425 = ~n19012 & n19424;
  assign n19426 = n19425 ^ n19423;
  assign n19006 = n18972 ^ n18902;
  assign n19427 = n19426 ^ n19006;
  assign n19428 = n18546 ^ n17768;
  assign n19429 = n19428 ^ n19079;
  assign n19430 = n19429 ^ n19006;
  assign n19431 = n19427 & ~n19430;
  assign n19432 = n19431 ^ n19429;
  assign n19433 = n19432 ^ n19004;
  assign n19434 = ~n19005 & ~n19433;
  assign n19435 = n19434 ^ n19003;
  assign n19000 = n18978 ^ n18898;
  assign n19436 = n19435 ^ n19000;
  assign n19437 = n18512 ^ n17757;
  assign n19438 = n19437 ^ n19075;
  assign n19439 = n19438 ^ n19000;
  assign n19440 = ~n19436 & ~n19439;
  assign n19441 = n19440 ^ n19438;
  assign n19442 = n19441 ^ n18998;
  assign n19443 = n18999 & ~n19442;
  assign n19444 = n19443 ^ n18483;
  assign n19565 = n19447 ^ n19444;
  assign n19566 = n19448 & n19565;
  assign n19567 = n19566 ^ n19446;
  assign n19569 = n19568 ^ n19567;
  assign n19572 = n19571 ^ n19569;
  assign n19573 = n19572 ^ n17313;
  assign n19449 = n19448 ^ n19444;
  assign n19450 = n19449 ^ n16960;
  assign n19451 = n19441 ^ n18483;
  assign n19452 = n19451 ^ n18998;
  assign n19453 = n19452 ^ n16963;
  assign n19454 = n19438 ^ n19436;
  assign n19455 = n19454 ^ n16968;
  assign n19457 = n19429 ^ n19427;
  assign n19458 = n19457 ^ n16977;
  assign n19459 = n19423 ^ n19012;
  assign n19460 = n19459 ^ n17101;
  assign n19461 = n19420 ^ n19016;
  assign n19462 = n19461 ^ n19013;
  assign n19463 = n19462 ^ n16981;
  assign n19464 = n19417 ^ n19022;
  assign n19465 = n19464 ^ n16985;
  assign n19466 = n19414 ^ n19027;
  assign n19467 = n19466 ^ n16987;
  assign n19468 = n19411 ^ n19033;
  assign n19469 = n19468 ^ n16991;
  assign n19470 = n19408 ^ n19406;
  assign n19471 = n19470 ^ n16995;
  assign n19474 = n19399 ^ n19397;
  assign n19475 = n19474 ^ n17005;
  assign n19476 = n19393 ^ n19043;
  assign n19477 = n19476 ^ n19041;
  assign n19478 = n19477 ^ n17007;
  assign n19480 = n19381 ^ n19379;
  assign n19481 = n19480 ^ n16942;
  assign n19482 = n19374 ^ n19372;
  assign n19483 = n19482 ^ n16947;
  assign n19484 = n19368 ^ n19366;
  assign n19485 = n19484 ^ n16952;
  assign n19486 = n19362 ^ n19360;
  assign n19487 = n19486 ^ n16957;
  assign n19488 = n19355 ^ n19353;
  assign n19489 = n17033 & n19488;
  assign n19490 = n19489 ^ n17031;
  assign n19491 = n19356 ^ n19352;
  assign n19492 = n19491 ^ n19489;
  assign n19493 = ~n19490 & ~n19492;
  assign n19494 = n19493 ^ n17031;
  assign n19495 = n19494 ^ n19486;
  assign n19496 = n19487 & n19495;
  assign n19497 = n19496 ^ n16957;
  assign n19498 = n19497 ^ n19484;
  assign n19499 = n19485 & ~n19498;
  assign n19500 = n19499 ^ n16952;
  assign n19501 = n19500 ^ n19482;
  assign n19502 = ~n19483 & ~n19501;
  assign n19503 = n19502 ^ n16947;
  assign n19504 = n19503 ^ n19480;
  assign n19505 = ~n19481 & ~n19504;
  assign n19506 = n19505 ^ n16942;
  assign n19507 = n19506 ^ n16937;
  assign n19508 = n19384 ^ n19057;
  assign n19509 = n19508 ^ n19506;
  assign n19510 = ~n19507 & n19509;
  assign n19511 = n19510 ^ n16937;
  assign n19479 = n19387 ^ n19053;
  assign n19512 = n19511 ^ n19479;
  assign n19513 = n19479 ^ n16932;
  assign n19514 = n19512 & n19513;
  assign n19515 = n19514 ^ n16932;
  assign n19516 = n19515 ^ n16928;
  assign n19517 = n19390 ^ n19048;
  assign n19518 = n19517 ^ n19515;
  assign n19519 = ~n19516 & n19518;
  assign n19520 = n19519 ^ n16928;
  assign n19521 = n19520 ^ n19477;
  assign n19522 = ~n19478 & ~n19521;
  assign n19523 = n19522 ^ n17007;
  assign n19524 = n19523 ^ n19474;
  assign n19525 = ~n19475 & n19524;
  assign n19526 = n19525 ^ n17005;
  assign n19472 = n19402 ^ n19037;
  assign n19473 = n19472 ^ n19035;
  assign n19527 = n19526 ^ n19473;
  assign n19528 = n19473 ^ n17001;
  assign n19529 = ~n19527 & ~n19528;
  assign n19530 = n19529 ^ n17001;
  assign n19531 = n19530 ^ n19470;
  assign n19532 = ~n19471 & ~n19531;
  assign n19533 = n19532 ^ n16995;
  assign n19534 = n19533 ^ n19468;
  assign n19535 = n19469 & n19534;
  assign n19536 = n19535 ^ n16991;
  assign n19537 = n19536 ^ n19466;
  assign n19538 = ~n19467 & n19537;
  assign n19539 = n19538 ^ n16987;
  assign n19540 = n19539 ^ n19464;
  assign n19541 = n19465 & ~n19540;
  assign n19542 = n19541 ^ n16985;
  assign n19543 = n19542 ^ n19462;
  assign n19544 = ~n19463 & ~n19543;
  assign n19545 = n19544 ^ n16981;
  assign n19546 = n19545 ^ n19459;
  assign n19547 = ~n19460 & ~n19546;
  assign n19548 = n19547 ^ n17101;
  assign n19549 = n19548 ^ n19457;
  assign n19550 = ~n19458 & ~n19549;
  assign n19551 = n19550 ^ n16977;
  assign n19456 = n19432 ^ n19005;
  assign n19552 = n19551 ^ n19456;
  assign n19553 = n19456 ^ n16970;
  assign n19554 = n19552 & n19553;
  assign n19555 = n19554 ^ n16970;
  assign n19556 = n19555 ^ n19454;
  assign n19557 = ~n19455 & n19556;
  assign n19558 = n19557 ^ n16968;
  assign n19559 = n19558 ^ n19452;
  assign n19560 = n19453 & n19559;
  assign n19561 = n19560 ^ n16963;
  assign n19562 = n19561 ^ n19449;
  assign n19563 = ~n19450 & ~n19562;
  assign n19564 = n19563 ^ n16960;
  assign n19761 = n19572 ^ n19564;
  assign n19762 = n19573 & n19761;
  assign n19763 = n19762 ^ n17313;
  assign n19756 = n19571 ^ n19568;
  assign n19757 = ~n19569 & ~n19756;
  assign n19758 = n19757 ^ n19571;
  assign n19753 = n19306 ^ n2774;
  assign n19754 = n19753 ^ n19292;
  assign n19751 = n19063 ^ n18640;
  assign n19752 = n19751 ^ n17994;
  assign n19755 = n19754 ^ n19752;
  assign n19759 = n19758 ^ n19755;
  assign n19760 = n19759 ^ n17326;
  assign n19764 = n19763 ^ n19760;
  assign n19574 = n19573 ^ n19564;
  assign n19575 = n19561 ^ n19450;
  assign n19576 = n19548 ^ n16977;
  assign n19577 = n19576 ^ n19457;
  assign n19578 = n19545 ^ n19460;
  assign n19579 = n19542 ^ n19463;
  assign n19580 = n19539 ^ n19465;
  assign n19581 = n19530 ^ n16995;
  assign n19582 = n19581 ^ n19470;
  assign n19583 = n19527 ^ n17001;
  assign n19584 = n19523 ^ n19475;
  assign n19585 = n19520 ^ n19478;
  assign n19586 = n19517 ^ n19516;
  assign n19587 = n19503 ^ n19481;
  assign n19588 = n19488 ^ n17033;
  assign n19589 = n19491 ^ n19490;
  assign n19590 = n19588 & ~n19589;
  assign n19591 = n19494 ^ n16957;
  assign n19592 = n19591 ^ n19486;
  assign n19593 = n19590 & ~n19592;
  assign n19594 = n19497 ^ n19485;
  assign n19595 = n19593 & n19594;
  assign n19596 = n19500 ^ n19483;
  assign n19597 = n19595 & ~n19596;
  assign n19598 = ~n19587 & ~n19597;
  assign n19599 = n19508 ^ n16937;
  assign n19600 = n19599 ^ n19506;
  assign n19601 = ~n19598 & n19600;
  assign n19602 = n19512 ^ n16932;
  assign n19603 = ~n19601 & n19602;
  assign n19604 = ~n19586 & n19603;
  assign n19605 = ~n19585 & n19604;
  assign n19606 = ~n19584 & ~n19605;
  assign n19607 = n19583 & ~n19606;
  assign n19608 = n19582 & ~n19607;
  assign n19609 = n19533 ^ n19469;
  assign n19610 = ~n19608 & ~n19609;
  assign n19611 = n19536 ^ n19467;
  assign n19612 = n19610 & ~n19611;
  assign n19613 = n19580 & n19612;
  assign n19614 = ~n19579 & n19613;
  assign n19615 = ~n19578 & ~n19614;
  assign n19616 = n19577 & n19615;
  assign n19617 = n19552 ^ n16970;
  assign n19618 = ~n19616 & ~n19617;
  assign n19619 = n19555 ^ n16968;
  assign n19620 = n19619 ^ n19454;
  assign n19621 = n19618 & ~n19620;
  assign n19622 = n19558 ^ n19453;
  assign n19623 = ~n19621 & ~n19622;
  assign n19624 = n19575 & ~n19623;
  assign n19750 = n19574 & n19624;
  assign n19765 = n19764 ^ n19750;
  assign n19766 = n19765 ^ n1679;
  assign n19626 = n19623 ^ n19575;
  assign n19627 = n19626 ^ n2810;
  assign n19629 = n19620 ^ n19618;
  assign n19630 = n19629 ^ n2691;
  assign n19633 = n19614 ^ n19578;
  assign n2520 = n2460 ^ x431;
  assign n2521 = n2520 ^ n2517;
  assign n2522 = n2521 ^ x367;
  assign n19634 = n19633 ^ n2522;
  assign n19635 = n19613 ^ n19579;
  assign n19636 = n19635 ^ n2513;
  assign n19637 = n19612 ^ n19580;
  assign n3149 = n3142 ^ x433;
  assign n3150 = n3149 ^ n1407;
  assign n3151 = n3150 ^ x369;
  assign n19638 = n19637 ^ n3151;
  assign n19639 = n19611 ^ n19610;
  assign n19640 = n19639 ^ n1400;
  assign n19641 = n19609 ^ n19608;
  assign n1213 = n1122 ^ x435;
  assign n1214 = n1213 ^ n1207;
  assign n1215 = n1214 ^ x371;
  assign n19642 = n19641 ^ n1215;
  assign n19643 = n19607 ^ n19582;
  assign n1198 = n1106 ^ x436;
  assign n1199 = n1198 ^ n1076;
  assign n1200 = n1199 ^ x372;
  assign n19644 = n19643 ^ n1200;
  assign n19645 = n19606 ^ n19583;
  assign n1064 = n982 ^ x437;
  assign n1065 = n1064 ^ n1058;
  assign n1066 = n1065 ^ x373;
  assign n19646 = n19645 ^ n1066;
  assign n19647 = n19605 ^ n19584;
  assign n19648 = n19647 ^ n1051;
  assign n19699 = n19604 ^ n19585;
  assign n19649 = n19603 ^ n19586;
  assign n19650 = n19649 ^ n746;
  assign n19652 = n19600 ^ n19598;
  assign n19653 = n19652 ^ n587;
  assign n19654 = n19597 ^ n19587;
  assign n19655 = n19654 ^ n644;
  assign n19656 = n19596 ^ n19595;
  assign n553 = n543 ^ x444;
  assign n557 = n556 ^ n553;
  assign n558 = n557 ^ x380;
  assign n19657 = n19656 ^ n558;
  assign n19658 = n19594 ^ n19593;
  assign n19659 = n19658 ^ n3281;
  assign n19660 = n19592 ^ n19590;
  assign n19664 = n19663 ^ n19660;
  assign n2295 = n2201 ^ x416;
  assign n2296 = n2295 ^ n2225;
  assign n2297 = n2296 ^ x352;
  assign n19665 = n2297 & ~n19588;
  assign n19669 = n19668 ^ n19665;
  assign n19670 = n19589 ^ n19588;
  assign n19671 = n19670 ^ n19665;
  assign n19672 = n19669 & n19671;
  assign n19673 = n19672 ^ n19668;
  assign n19674 = n19673 ^ n19660;
  assign n19675 = ~n19664 & n19674;
  assign n19676 = n19675 ^ n19663;
  assign n19677 = n19676 ^ n19658;
  assign n19678 = n19659 & ~n19677;
  assign n19679 = n19678 ^ n3281;
  assign n19680 = n19679 ^ n19656;
  assign n19681 = ~n19657 & n19680;
  assign n19682 = n19681 ^ n558;
  assign n19683 = n19682 ^ n19654;
  assign n19684 = ~n19655 & n19683;
  assign n19685 = n19684 ^ n644;
  assign n19686 = n19685 ^ n19652;
  assign n19687 = ~n19653 & n19686;
  assign n19688 = n19687 ^ n587;
  assign n19651 = n19602 ^ n19601;
  assign n19689 = n19688 ^ n19651;
  assign n19693 = n19692 ^ n19651;
  assign n19694 = ~n19689 & n19693;
  assign n19695 = n19694 ^ n19692;
  assign n19696 = n19695 ^ n19649;
  assign n19697 = n19650 & ~n19696;
  assign n19698 = n19697 ^ n746;
  assign n19700 = n19699 ^ n19698;
  assign n19701 = n19699 ^ n1045;
  assign n19702 = ~n19700 & n19701;
  assign n19703 = n19702 ^ n1045;
  assign n19704 = n19703 ^ n19647;
  assign n19705 = n19648 & ~n19704;
  assign n19706 = n19705 ^ n1051;
  assign n19707 = n19706 ^ n19645;
  assign n19708 = n19646 & ~n19707;
  assign n19709 = n19708 ^ n1066;
  assign n19710 = n19709 ^ n19643;
  assign n19711 = ~n19644 & n19710;
  assign n19712 = n19711 ^ n1200;
  assign n19713 = n19712 ^ n19641;
  assign n19714 = ~n19642 & n19713;
  assign n19715 = n19714 ^ n1215;
  assign n19716 = n19715 ^ n19639;
  assign n19717 = n19640 & ~n19716;
  assign n19718 = n19717 ^ n1400;
  assign n19719 = n19718 ^ n19637;
  assign n19720 = ~n19638 & n19719;
  assign n19721 = n19720 ^ n3151;
  assign n19722 = n19721 ^ n19635;
  assign n19723 = n19636 & ~n19722;
  assign n19724 = n19723 ^ n2513;
  assign n19725 = n19724 ^ n19633;
  assign n19726 = n19634 & ~n19725;
  assign n19727 = n19726 ^ n2522;
  assign n19632 = n19615 ^ n19577;
  assign n19728 = n19727 ^ n19632;
  assign n2582 = n2542 ^ x430;
  assign n2583 = n2582 ^ n2529;
  assign n2584 = n2583 ^ x366;
  assign n19729 = n19632 ^ n2584;
  assign n19730 = ~n19728 & n19729;
  assign n19731 = n19730 ^ n2584;
  assign n19631 = n19617 ^ n19616;
  assign n19732 = n19731 ^ n19631;
  assign n19733 = n19631 ^ n1559;
  assign n19734 = n19732 & ~n19733;
  assign n19735 = n19734 ^ n1559;
  assign n19736 = n19735 ^ n19629;
  assign n19737 = n19630 & ~n19736;
  assign n19738 = n19737 ^ n2691;
  assign n19628 = n19622 ^ n19621;
  assign n19739 = n19738 ^ n19628;
  assign n19740 = n19628 ^ n2979;
  assign n19741 = ~n19739 & n19740;
  assign n19742 = n19741 ^ n2979;
  assign n19743 = n19742 ^ n19626;
  assign n19744 = n19627 & ~n19743;
  assign n19745 = n19744 ^ n2810;
  assign n19625 = n19624 ^ n19574;
  assign n19746 = n19745 ^ n19625;
  assign n19747 = n19625 ^ n2993;
  assign n19748 = n19746 & ~n19747;
  assign n19749 = n19748 ^ n2993;
  assign n19913 = n19765 ^ n19749;
  assign n19914 = ~n19766 & n19913;
  assign n19915 = n19914 ^ n1679;
  assign n19856 = n19763 ^ n19759;
  assign n19857 = n19760 & n19856;
  assign n19858 = n19857 ^ n17326;
  assign n19809 = n19758 ^ n19754;
  assign n19810 = ~n19755 & ~n19809;
  assign n19811 = n19810 ^ n19752;
  assign n19806 = n19062 ^ n17479;
  assign n19807 = n19806 ^ n18112;
  assign n19804 = n19309 ^ n2768;
  assign n19805 = n19804 ^ n19290;
  assign n19808 = n19807 ^ n19805;
  assign n19854 = n19811 ^ n19808;
  assign n19855 = n19854 ^ n16743;
  assign n19880 = n19858 ^ n19855;
  assign n19879 = ~n19750 & n19764;
  assign n19911 = n19880 ^ n19879;
  assign n19912 = n19911 ^ n1688;
  assign n20424 = n19915 ^ n19912;
  assign n19842 = n19324 ^ n19280;
  assign n19843 = n19842 ^ n19277;
  assign n21532 = n20424 ^ n19843;
  assign n20050 = n19138 ^ n18512;
  assign n20051 = n20050 ^ n19805;
  assign n20048 = n19718 ^ n19638;
  assign n19770 = n19754 ^ n18480;
  assign n19771 = n19770 ^ n18519;
  assign n19768 = n19715 ^ n1400;
  assign n19769 = n19768 ^ n19639;
  assign n19772 = n19771 ^ n19769;
  assign n19776 = n19447 ^ n18522;
  assign n19777 = n19776 ^ n19001;
  assign n19775 = n19709 ^ n19644;
  assign n19778 = n19777 ^ n19775;
  assign n20029 = n19706 ^ n19646;
  assign n19790 = n19676 ^ n3281;
  assign n19791 = n19790 ^ n19658;
  assign n19788 = n19029 ^ n18861;
  assign n19789 = n19788 ^ n17709;
  assign n19792 = n19791 ^ n19789;
  assign n19796 = n19035 ^ n18488;
  assign n19797 = n19796 ^ n17719;
  assign n19795 = n19670 ^ n19669;
  assign n19798 = n19797 ^ n19795;
  assign n19968 = n19588 ^ n2297;
  assign n19824 = n18106 ^ n17478;
  assign n19825 = n19824 ^ n18714;
  assign n19822 = n19315 ^ n19287;
  assign n19815 = n19312 ^ n19289;
  assign n19812 = n19811 ^ n19805;
  assign n19813 = n19808 & ~n19812;
  assign n19814 = n19813 ^ n19807;
  assign n19816 = n19815 ^ n19814;
  assign n19817 = n19060 ^ n18117;
  assign n19818 = n19817 ^ n17486;
  assign n19819 = n19818 ^ n19815;
  assign n19820 = n19816 & ~n19819;
  assign n19821 = n19820 ^ n19818;
  assign n19823 = n19822 ^ n19821;
  assign n19850 = n19825 ^ n19823;
  assign n19851 = n19850 ^ n16798;
  assign n19852 = n19818 ^ n19816;
  assign n19853 = n19852 ^ n16772;
  assign n19859 = n19858 ^ n19854;
  assign n19860 = n19855 & ~n19859;
  assign n19861 = n19860 ^ n16743;
  assign n19862 = n19861 ^ n19852;
  assign n19863 = n19853 & n19862;
  assign n19864 = n19863 ^ n16772;
  assign n19865 = n19864 ^ n19850;
  assign n19866 = ~n19851 & n19865;
  assign n19867 = n19866 ^ n16798;
  assign n19830 = n18101 ^ n17476;
  assign n19831 = n19830 ^ n18719;
  assign n19826 = n19825 ^ n19822;
  assign n19827 = ~n19823 & n19826;
  assign n19828 = n19827 ^ n19825;
  assign n19803 = n19318 ^ n19285;
  assign n19829 = n19828 ^ n19803;
  assign n19848 = n19831 ^ n19829;
  assign n19849 = n19848 ^ n16838;
  assign n19877 = n19867 ^ n19849;
  assign n19878 = n19864 ^ n19851;
  assign n19881 = ~n19879 & n19880;
  assign n19882 = n19861 ^ n19853;
  assign n19883 = n19881 & n19882;
  assign n19884 = n19878 & n19883;
  assign n19885 = ~n19877 & ~n19884;
  assign n19868 = n19867 ^ n19848;
  assign n19869 = ~n19849 & ~n19868;
  assign n19870 = n19869 ^ n16838;
  assign n19837 = n18097 ^ n17472;
  assign n19838 = n19837 ^ n18711;
  assign n19835 = n19321 ^ n19283;
  assign n19832 = n19831 ^ n19803;
  assign n19833 = ~n19829 & ~n19832;
  assign n19834 = n19833 ^ n19831;
  assign n19836 = n19835 ^ n19834;
  assign n19846 = n19838 ^ n19836;
  assign n19847 = n19846 ^ n16870;
  assign n19876 = n19870 ^ n19847;
  assign n19905 = n19885 ^ n19876;
  assign n19906 = n19905 ^ n2264;
  assign n19908 = n19883 ^ n19878;
  assign n19909 = n19908 ^ n1765;
  assign n19916 = n19915 ^ n19911;
  assign n19917 = n19912 & ~n19916;
  assign n19918 = n19917 ^ n1688;
  assign n19910 = n19882 ^ n19881;
  assign n19919 = n19918 ^ n19910;
  assign n1754 = n1727 ^ x422;
  assign n1755 = n1754 ^ n1693;
  assign n1756 = n1755 ^ x358;
  assign n19920 = n19910 ^ n1756;
  assign n19921 = n19919 & ~n19920;
  assign n19922 = n19921 ^ n1756;
  assign n19923 = n19922 ^ n19908;
  assign n19924 = ~n19909 & n19923;
  assign n19925 = n19924 ^ n1765;
  assign n19907 = n19884 ^ n19877;
  assign n19926 = n19925 ^ n19907;
  assign n19927 = n19907 ^ n1877;
  assign n19928 = ~n19926 & n19927;
  assign n19929 = n19928 ^ n1877;
  assign n19930 = n19929 ^ n19905;
  assign n19931 = ~n19906 & n19930;
  assign n19932 = n19931 ^ n2264;
  assign n19886 = ~n19876 & ~n19885;
  assign n19871 = n19870 ^ n19846;
  assign n19872 = ~n19847 & ~n19871;
  assign n19873 = n19872 ^ n16870;
  assign n19874 = n19873 ^ n16917;
  assign n19839 = n19838 ^ n19835;
  assign n19840 = ~n19836 & ~n19839;
  assign n19841 = n19840 ^ n19838;
  assign n19844 = n19843 ^ n19841;
  assign n19801 = n17746 ^ n16954;
  assign n19802 = n19801 ^ n18707;
  assign n19845 = n19844 ^ n19802;
  assign n19875 = n19874 ^ n19845;
  assign n19904 = n19886 ^ n19875;
  assign n19933 = n19932 ^ n19904;
  assign n19934 = n19904 ^ n2042;
  assign n19935 = ~n19933 & n19934;
  assign n19936 = n19935 ^ n2042;
  assign n19937 = n19936 ^ n2279;
  assign n19897 = n19845 ^ n16917;
  assign n19898 = n19873 ^ n19845;
  assign n19899 = n19897 & n19898;
  assign n19900 = n19899 ^ n16917;
  assign n19901 = n19900 ^ n17037;
  assign n19894 = n19327 ^ n1722;
  assign n19895 = n19894 ^ n19275;
  assign n19890 = n19843 ^ n19802;
  assign n19891 = ~n19844 & n19890;
  assign n19892 = n19891 ^ n19802;
  assign n19888 = n18706 ^ n17742;
  assign n19889 = n19888 ^ n16949;
  assign n19893 = n19892 ^ n19889;
  assign n19896 = n19895 ^ n19893;
  assign n19902 = n19901 ^ n19896;
  assign n19887 = ~n19875 & n19886;
  assign n19903 = n19902 ^ n19887;
  assign n19938 = n19937 ^ n19903;
  assign n19799 = n19041 ^ n18768;
  assign n19800 = n19799 ^ n17724;
  assign n19939 = n19938 ^ n19800;
  assign n19943 = n19929 ^ n19906;
  assign n19941 = n19050 ^ n18494;
  assign n19942 = n19941 ^ n17734;
  assign n19944 = n19943 ^ n19942;
  assign n19949 = n18499 ^ n18140;
  assign n19950 = n19949 ^ n19054;
  assign n19945 = n19378 ^ n17738;
  assign n19946 = n19945 ^ n18503;
  assign n19947 = n19922 ^ n19909;
  assign n19948 = n19946 & ~n19947;
  assign n19951 = n19950 ^ n19948;
  assign n19952 = n19926 ^ n1877;
  assign n19953 = n19952 ^ n19950;
  assign n19954 = ~n19951 & n19953;
  assign n19955 = n19954 ^ n19948;
  assign n19956 = n19955 ^ n19943;
  assign n19957 = ~n19944 & n19956;
  assign n19958 = n19957 ^ n19942;
  assign n19940 = n19933 ^ n2042;
  assign n19959 = n19958 ^ n19940;
  assign n19960 = n19047 ^ n18761;
  assign n19961 = n19960 ^ n17726;
  assign n19962 = n19961 ^ n19958;
  assign n19963 = ~n19959 & ~n19962;
  assign n19964 = n19963 ^ n19961;
  assign n19965 = n19964 ^ n19938;
  assign n19966 = n19939 & ~n19965;
  assign n19967 = n19966 ^ n19800;
  assign n19969 = n19968 ^ n19967;
  assign n19970 = n19040 ^ n18156;
  assign n19971 = n19970 ^ n18492;
  assign n19972 = n19971 ^ n19968;
  assign n19973 = ~n19969 & n19972;
  assign n19974 = n19973 ^ n19971;
  assign n19975 = n19974 ^ n19795;
  assign n19976 = n19798 & ~n19975;
  assign n19977 = n19976 ^ n19797;
  assign n19793 = n19673 ^ n19663;
  assign n19794 = n19793 ^ n19660;
  assign n19978 = n19977 ^ n19794;
  assign n19979 = n19034 ^ n18782;
  assign n19980 = n19979 ^ n17714;
  assign n19981 = n19980 ^ n19794;
  assign n19982 = ~n19978 & n19981;
  assign n19983 = n19982 ^ n19980;
  assign n19984 = n19983 ^ n19791;
  assign n19985 = ~n19792 & n19984;
  assign n19986 = n19985 ^ n19789;
  assign n19787 = n19679 ^ n19657;
  assign n19987 = n19986 ^ n19787;
  assign n19988 = n18985 ^ n18176;
  assign n19989 = n19988 ^ n19023;
  assign n19990 = n19989 ^ n19787;
  assign n19991 = ~n19987 & n19990;
  assign n19992 = n19991 ^ n19989;
  assign n19786 = n19682 ^ n19655;
  assign n19993 = n19992 ^ n19786;
  assign n19994 = n19089 ^ n17708;
  assign n19995 = n19994 ^ n19018;
  assign n19996 = n19995 ^ n19786;
  assign n19997 = ~n19993 & ~n19996;
  assign n19998 = n19997 ^ n19995;
  assign n19785 = n19685 ^ n19653;
  assign n19999 = n19998 ^ n19785;
  assign n20000 = n19030 ^ n17703;
  assign n20001 = n20000 ^ n19013;
  assign n20002 = n20001 ^ n19785;
  assign n20003 = n19999 & ~n20002;
  assign n20004 = n20003 ^ n20001;
  assign n19784 = n19692 ^ n19689;
  assign n20005 = n20004 ^ n19784;
  assign n20006 = n19008 ^ n18193;
  assign n20007 = n20006 ^ n19024;
  assign n20008 = n20007 ^ n19784;
  assign n20009 = ~n20005 & n20008;
  assign n20010 = n20009 ^ n20007;
  assign n19782 = n19695 ^ n746;
  assign n19783 = n19782 ^ n19649;
  assign n20011 = n20010 ^ n19783;
  assign n20012 = n19019 ^ n19006;
  assign n20013 = n20012 ^ n18304;
  assign n20014 = n20013 ^ n19783;
  assign n20015 = ~n20011 & n20014;
  assign n20016 = n20015 ^ n20013;
  assign n19780 = n19698 ^ n1045;
  assign n19781 = n19780 ^ n19699;
  assign n20017 = n20016 ^ n19781;
  assign n20018 = n19014 ^ n18474;
  assign n20019 = n20018 ^ n19004;
  assign n20020 = n20019 ^ n19781;
  assign n20021 = ~n20017 & n20020;
  assign n20022 = n20021 ^ n20019;
  assign n19779 = n19703 ^ n19648;
  assign n20023 = n20022 ^ n19779;
  assign n20024 = n19000 ^ n18532;
  assign n20025 = n20024 ^ n19009;
  assign n20026 = n20025 ^ n19779;
  assign n20027 = ~n20023 & n20026;
  assign n20028 = n20027 ^ n20025;
  assign n20030 = n20029 ^ n20028;
  assign n20031 = n18998 ^ n18526;
  assign n20032 = n20031 ^ n19079;
  assign n20033 = n20032 ^ n20029;
  assign n20034 = ~n20030 & n20033;
  assign n20035 = n20034 ^ n20032;
  assign n20036 = n20035 ^ n19775;
  assign n20037 = ~n19778 & n20036;
  assign n20038 = n20037 ^ n19777;
  assign n19773 = n19712 ^ n1215;
  assign n19774 = n19773 ^ n19641;
  assign n20039 = n20038 ^ n19774;
  assign n20040 = n19568 ^ n18546;
  assign n20041 = n20040 ^ n19075;
  assign n20042 = n20041 ^ n19774;
  assign n20043 = n20039 & ~n20042;
  assign n20044 = n20043 ^ n20041;
  assign n20045 = n20044 ^ n19769;
  assign n20046 = ~n19772 & ~n20045;
  assign n20047 = n20046 ^ n19771;
  assign n20049 = n20048 ^ n20047;
  assign n20061 = n20051 ^ n20049;
  assign n20062 = n20061 ^ n17757;
  assign n20063 = n20044 ^ n19772;
  assign n20064 = n20063 ^ n17764;
  assign n20065 = n20041 ^ n20039;
  assign n20066 = n20065 ^ n17768;
  assign n20067 = n20035 ^ n19778;
  assign n20068 = n20067 ^ n17772;
  assign n20069 = n20032 ^ n20030;
  assign n20070 = n20069 ^ n17705;
  assign n20071 = n20025 ^ n20023;
  assign n20072 = n20071 ^ n17780;
  assign n20073 = n20019 ^ n20017;
  assign n20074 = n20073 ^ n17784;
  assign n20075 = n20013 ^ n20011;
  assign n20076 = n20075 ^ n17710;
  assign n20077 = n20007 ^ n20005;
  assign n20078 = n20077 ^ n17715;
  assign n20079 = n20001 ^ n19999;
  assign n20080 = n20079 ^ n17795;
  assign n20081 = n19995 ^ n19993;
  assign n20082 = n20081 ^ n17799;
  assign n20083 = n19989 ^ n19987;
  assign n20084 = n20083 ^ n17720;
  assign n20085 = n19983 ^ n19792;
  assign n20086 = n20085 ^ n17727;
  assign n20087 = n19980 ^ n19978;
  assign n20088 = n20087 ^ n17731;
  assign n20089 = n19974 ^ n19798;
  assign n20090 = n20089 ^ n17626;
  assign n20091 = n19971 ^ n19969;
  assign n20092 = n20091 ^ n17585;
  assign n20093 = n19964 ^ n19939;
  assign n20094 = n20093 ^ n17523;
  assign n20095 = n19961 ^ n19959;
  assign n20096 = n20095 ^ n16926;
  assign n20097 = n19955 ^ n19944;
  assign n20098 = n20097 ^ n16934;
  assign n20099 = n19947 ^ n19946;
  assign n20100 = ~n16944 & ~n20099;
  assign n20101 = n20100 ^ n16939;
  assign n20102 = n19952 ^ n19951;
  assign n20103 = n20102 ^ n20100;
  assign n20104 = n20101 & n20103;
  assign n20105 = n20104 ^ n16939;
  assign n20106 = n20105 ^ n20097;
  assign n20107 = ~n20098 & n20106;
  assign n20108 = n20107 ^ n16934;
  assign n20109 = n20108 ^ n20095;
  assign n20110 = n20096 & n20109;
  assign n20111 = n20110 ^ n16926;
  assign n20112 = n20111 ^ n20093;
  assign n20113 = ~n20094 & ~n20112;
  assign n20114 = n20113 ^ n17523;
  assign n20115 = n20114 ^ n20091;
  assign n20116 = n20092 & n20115;
  assign n20117 = n20116 ^ n17585;
  assign n20118 = n20117 ^ n20089;
  assign n20119 = n20090 & ~n20118;
  assign n20120 = n20119 ^ n17626;
  assign n20121 = n20120 ^ n20087;
  assign n20122 = ~n20088 & ~n20121;
  assign n20123 = n20122 ^ n17731;
  assign n20124 = n20123 ^ n20085;
  assign n20125 = ~n20086 & ~n20124;
  assign n20126 = n20125 ^ n17727;
  assign n20127 = n20126 ^ n20083;
  assign n20128 = ~n20084 & ~n20127;
  assign n20129 = n20128 ^ n17720;
  assign n20130 = n20129 ^ n20081;
  assign n20131 = n20082 & ~n20130;
  assign n20132 = n20131 ^ n17799;
  assign n20133 = n20132 ^ n20079;
  assign n20134 = n20080 & n20133;
  assign n20135 = n20134 ^ n17795;
  assign n20136 = n20135 ^ n20077;
  assign n20137 = n20078 & n20136;
  assign n20138 = n20137 ^ n17715;
  assign n20139 = n20138 ^ n20075;
  assign n20140 = n20076 & ~n20139;
  assign n20141 = n20140 ^ n17710;
  assign n20142 = n20141 ^ n20073;
  assign n20143 = n20074 & ~n20142;
  assign n20144 = n20143 ^ n17784;
  assign n20145 = n20144 ^ n20071;
  assign n20146 = ~n20072 & ~n20145;
  assign n20147 = n20146 ^ n17780;
  assign n20148 = n20147 ^ n20069;
  assign n20149 = ~n20070 & n20148;
  assign n20150 = n20149 ^ n17705;
  assign n20151 = n20150 ^ n20067;
  assign n20152 = ~n20068 & ~n20151;
  assign n20153 = n20152 ^ n17772;
  assign n20154 = n20153 ^ n20065;
  assign n20155 = ~n20066 & n20154;
  assign n20156 = n20155 ^ n17768;
  assign n20157 = n20156 ^ n20063;
  assign n20158 = n20064 & n20157;
  assign n20159 = n20158 ^ n17764;
  assign n20160 = n20159 ^ n20061;
  assign n20161 = n20062 & n20160;
  assign n20162 = n20161 ^ n17757;
  assign n20056 = n19815 ^ n18481;
  assign n20057 = n20056 ^ n19069;
  assign n20055 = n19721 ^ n19636;
  assign n20058 = n20057 ^ n20055;
  assign n20052 = n20051 ^ n20048;
  assign n20053 = ~n20049 & ~n20052;
  assign n20054 = n20053 ^ n20051;
  assign n20059 = n20058 ^ n20054;
  assign n20060 = n20059 ^ n17753;
  assign n20176 = n20162 ^ n20060;
  assign n20177 = n20156 ^ n20064;
  assign n20178 = n20153 ^ n20066;
  assign n20179 = n20150 ^ n20068;
  assign n20180 = n20141 ^ n17784;
  assign n20181 = n20180 ^ n20073;
  assign n20182 = n20135 ^ n20078;
  assign n20183 = n20126 ^ n20084;
  assign n20184 = n20120 ^ n20088;
  assign n20185 = n20117 ^ n20090;
  assign n20186 = n20114 ^ n20092;
  assign n20187 = n20105 ^ n20098;
  assign n20188 = n20099 ^ n16944;
  assign n20189 = n20102 ^ n20101;
  assign n20190 = n20188 & ~n20189;
  assign n20191 = ~n20187 & n20190;
  assign n20192 = n20108 ^ n20096;
  assign n20193 = n20191 & n20192;
  assign n20194 = n20111 ^ n20094;
  assign n20195 = n20193 & n20194;
  assign n20196 = ~n20186 & ~n20195;
  assign n20197 = ~n20185 & ~n20196;
  assign n20198 = ~n20184 & ~n20197;
  assign n20199 = n20123 ^ n20086;
  assign n20200 = n20198 & n20199;
  assign n20201 = ~n20183 & n20200;
  assign n20202 = n20129 ^ n20082;
  assign n20203 = ~n20201 & n20202;
  assign n20204 = n20132 ^ n20080;
  assign n20205 = ~n20203 & ~n20204;
  assign n20206 = ~n20182 & ~n20205;
  assign n20207 = n20138 ^ n20076;
  assign n20208 = ~n20206 & ~n20207;
  assign n20209 = ~n20181 & n20208;
  assign n20210 = n20144 ^ n17780;
  assign n20211 = n20210 ^ n20071;
  assign n20212 = n20209 & n20211;
  assign n20213 = n20147 ^ n20070;
  assign n20214 = n20212 & ~n20213;
  assign n20215 = n20179 & ~n20214;
  assign n20216 = ~n20178 & n20215;
  assign n20217 = ~n20177 & ~n20216;
  assign n20218 = n20159 ^ n20062;
  assign n20219 = n20217 & n20218;
  assign n20220 = n20176 & ~n20219;
  assign n20171 = n19724 ^ n19634;
  assign n20169 = n19822 ^ n19063;
  assign n20170 = n20169 ^ n18615;
  assign n20172 = n20171 ^ n20170;
  assign n20166 = n20055 ^ n20054;
  assign n20167 = ~n20058 & ~n20166;
  assign n20168 = n20167 ^ n20057;
  assign n20173 = n20172 ^ n20168;
  assign n20174 = n20173 ^ n17749;
  assign n20163 = n20162 ^ n20059;
  assign n20164 = n20060 & n20163;
  assign n20165 = n20164 ^ n17753;
  assign n20175 = n20174 ^ n20165;
  assign n20236 = n20220 ^ n20175;
  assign n20237 = n20236 ^ n2880;
  assign n20239 = n20218 ^ n20217;
  assign n20240 = n20239 ^ n2679;
  assign n20242 = n20215 ^ n20178;
  assign n20243 = n20242 ^ n2657;
  assign n20244 = n20214 ^ n20179;
  assign n20245 = n20244 ^ n3185;
  assign n20246 = n20213 ^ n20212;
  assign n20247 = n20246 ^ n3029;
  assign n20248 = n20211 ^ n20209;
  assign n2409 = n1426 ^ x465;
  assign n2413 = n2412 ^ n2409;
  assign n2414 = n2413 ^ x401;
  assign n20249 = n20248 ^ n2414;
  assign n20251 = n20207 ^ n20206;
  assign n1350 = n1244 ^ x467;
  assign n1351 = n1350 ^ n1344;
  assign n1352 = n1351 ^ x403;
  assign n20252 = n20251 ^ n1352;
  assign n20253 = n20205 ^ n20182;
  assign n1080 = n1001 ^ x468;
  assign n1084 = n1083 ^ n1080;
  assign n1085 = n1084 ^ x404;
  assign n20254 = n20253 ^ n1085;
  assign n20255 = n20204 ^ n20203;
  assign n20256 = n20255 ^ n1334;
  assign n20258 = n20200 ^ n20183;
  assign n20259 = n20258 ^ n811;
  assign n20261 = n20197 ^ n20184;
  assign n20262 = n20261 ^ n631;
  assign n20263 = n20196 ^ n20185;
  assign n20264 = n20263 ^ n622;
  assign n20266 = n20194 ^ n20193;
  assign n20270 = n20269 ^ n20266;
  assign n20271 = n20192 ^ n20191;
  assign n20275 = n20274 ^ n20271;
  assign n20277 = n18399 ^ x478;
  assign n20278 = n20277 ^ n15248;
  assign n20279 = n20278 ^ x414;
  assign n20276 = n20190 ^ n20187;
  assign n20280 = n20279 ^ n20276;
  assign n20281 = n2321 & ~n20188;
  assign n20282 = n20281 ^ n690;
  assign n20283 = n20189 ^ n20188;
  assign n20284 = n20283 ^ n20281;
  assign n20285 = n20282 & n20284;
  assign n20286 = n20285 ^ n690;
  assign n20287 = n20286 ^ n20276;
  assign n20288 = ~n20280 & n20287;
  assign n20289 = n20288 ^ n20279;
  assign n20290 = n20289 ^ n20271;
  assign n20291 = n20275 & ~n20290;
  assign n20292 = n20291 ^ n20274;
  assign n20293 = n20292 ^ n20266;
  assign n20294 = n20270 & ~n20293;
  assign n20295 = n20294 ^ n20269;
  assign n20265 = n20195 ^ n20186;
  assign n20296 = n20295 ^ n20265;
  assign n20297 = n20265 ^ n3260;
  assign n20298 = n20296 & ~n20297;
  assign n20299 = n20298 ^ n3260;
  assign n20300 = n20299 ^ n20263;
  assign n20301 = n20264 & ~n20300;
  assign n20302 = n20301 ^ n622;
  assign n20303 = n20302 ^ n20261;
  assign n20304 = ~n20262 & n20303;
  assign n20305 = n20304 ^ n631;
  assign n20260 = n20199 ^ n20198;
  assign n20306 = n20305 ^ n20260;
  assign n20307 = n20260 ^ n802;
  assign n20308 = n20306 & ~n20307;
  assign n20309 = n20308 ^ n802;
  assign n20310 = n20309 ^ n20258;
  assign n20311 = n20259 & ~n20310;
  assign n20312 = n20311 ^ n811;
  assign n20257 = n20202 ^ n20201;
  assign n20313 = n20312 ^ n20257;
  assign n20314 = n20257 ^ n924;
  assign n20315 = n20313 & ~n20314;
  assign n20316 = n20315 ^ n924;
  assign n20317 = n20316 ^ n20255;
  assign n20318 = ~n20256 & n20317;
  assign n20319 = n20318 ^ n1334;
  assign n20320 = n20319 ^ n20253;
  assign n20321 = n20254 & ~n20320;
  assign n20322 = n20321 ^ n1085;
  assign n20323 = n20322 ^ n20251;
  assign n20324 = ~n20252 & n20323;
  assign n20325 = n20324 ^ n1352;
  assign n20250 = n20208 ^ n20181;
  assign n20326 = n20325 ^ n20250;
  assign n1368 = n1262 ^ x466;
  assign n1369 = n1368 ^ n1268;
  assign n1370 = n1369 ^ x402;
  assign n20327 = n20250 ^ n1370;
  assign n20328 = ~n20326 & n20327;
  assign n20329 = n20328 ^ n1370;
  assign n20330 = n20329 ^ n20248;
  assign n20331 = ~n20249 & n20330;
  assign n20332 = n20331 ^ n2414;
  assign n20333 = n20332 ^ n20246;
  assign n20334 = n20247 & ~n20333;
  assign n20335 = n20334 ^ n3029;
  assign n20336 = n20335 ^ n20244;
  assign n20337 = ~n20245 & n20336;
  assign n20338 = n20337 ^ n3185;
  assign n20339 = n20338 ^ n20242;
  assign n20340 = ~n20243 & n20339;
  assign n20341 = n20340 ^ n2657;
  assign n20241 = n20216 ^ n20177;
  assign n20342 = n20341 ^ n20241;
  assign n2662 = n2596 ^ x461;
  assign n2663 = n2662 ^ n2651;
  assign n2664 = n2663 ^ x397;
  assign n20343 = n20241 ^ n2664;
  assign n20344 = n20342 & ~n20343;
  assign n20345 = n20344 ^ n2664;
  assign n20346 = n20345 ^ n20239;
  assign n20347 = ~n20240 & n20346;
  assign n20348 = n20347 ^ n2679;
  assign n20238 = n20219 ^ n20176;
  assign n20349 = n20348 ^ n20238;
  assign n20350 = n20238 ^ n1527;
  assign n20351 = n20349 & ~n20350;
  assign n20352 = n20351 ^ n1527;
  assign n20353 = n20352 ^ n20236;
  assign n20354 = ~n20237 & n20353;
  assign n20355 = n20354 ^ n2880;
  assign n20230 = n19728 ^ n2584;
  assign n20227 = n20171 ^ n20168;
  assign n20228 = n20172 & n20227;
  assign n20229 = n20228 ^ n20170;
  assign n20231 = n20230 ^ n20229;
  assign n20225 = n19803 ^ n18628;
  assign n20226 = n20225 ^ n19062;
  assign n20232 = n20231 ^ n20226;
  assign n20233 = n20232 ^ n17985;
  assign n20222 = n20173 ^ n20165;
  assign n20223 = ~n20174 & ~n20222;
  assign n20224 = n20223 ^ n17749;
  assign n20234 = n20233 ^ n20224;
  assign n20221 = ~n20175 & ~n20220;
  assign n20235 = n20234 ^ n20221;
  assign n20356 = n20355 ^ n20235;
  assign n21002 = n20356 ^ n1595;
  assign n21533 = n21532 ^ n21002;
  assign n19767 = n19766 ^ n19749;
  assign n21496 = n19835 ^ n19767;
  assign n20995 = n20352 ^ n20237;
  assign n21497 = n21496 ^ n20995;
  assign n20635 = n19447 ^ n19009;
  assign n20636 = n20635 ^ n20048;
  assign n20399 = n20309 ^ n20259;
  assign n20397 = n19769 ^ n19014;
  assign n20398 = n20397 ^ n18998;
  assign n20400 = n20399 ^ n20398;
  assign n20624 = n20306 ^ n802;
  assign n20402 = n19775 ^ n19024;
  assign n20403 = n20402 ^ n19004;
  assign n20401 = n20302 ^ n20262;
  assign n20404 = n20403 ^ n20401;
  assign n20614 = n20299 ^ n20264;
  assign n20406 = n19089 ^ n19008;
  assign n20407 = n20406 ^ n19779;
  assign n20405 = n20296 ^ n3260;
  assign n20408 = n20407 ^ n20405;
  assign n20412 = n20289 ^ n20275;
  assign n20410 = n19783 ^ n18861;
  assign n20411 = n20410 ^ n19018;
  assign n20413 = n20412 ^ n20411;
  assign n20417 = n20283 ^ n20282;
  assign n20415 = n19785 ^ n18488;
  assign n20416 = n20415 ^ n19029;
  assign n20418 = n20417 ^ n20416;
  assign n20368 = n19060 ^ n18640;
  assign n20369 = n20368 ^ n19835;
  assign n20364 = n20230 ^ n20226;
  assign n20365 = ~n20231 & ~n20364;
  assign n20366 = n20365 ^ n20226;
  assign n20363 = n19732 ^ n1559;
  assign n20367 = n20366 ^ n20363;
  assign n20370 = n20369 ^ n20367;
  assign n20371 = n20370 ^ n17994;
  assign n20360 = n20232 ^ n20224;
  assign n20361 = n20233 & n20360;
  assign n20362 = n20361 ^ n17985;
  assign n20372 = n20371 ^ n20362;
  assign n20373 = n20221 & ~n20234;
  assign n20497 = n20372 & ~n20373;
  assign n20473 = n20370 ^ n20362;
  assign n20474 = ~n20371 & ~n20473;
  assign n20475 = n20474 ^ n17994;
  assign n20432 = n19843 ^ n18112;
  assign n20433 = n20432 ^ n18714;
  assign n20428 = n20369 ^ n20363;
  assign n20429 = ~n20367 & n20428;
  assign n20430 = n20429 ^ n20369;
  assign n20382 = n19735 ^ n19630;
  assign n20431 = n20430 ^ n20382;
  assign n20471 = n20433 ^ n20431;
  assign n20472 = n20471 ^ n17479;
  assign n20496 = n20475 ^ n20472;
  assign n20525 = n20497 ^ n20496;
  assign n20529 = n20528 ^ n20525;
  assign n20374 = n20373 ^ n20372;
  assign n20378 = n20377 ^ n20374;
  assign n20357 = n20235 ^ n1595;
  assign n20358 = ~n20356 & n20357;
  assign n20359 = n20358 ^ n1595;
  assign n20530 = n20374 ^ n20359;
  assign n20531 = ~n20378 & n20530;
  assign n20532 = n20531 ^ n20377;
  assign n20533 = n20532 ^ n20525;
  assign n20534 = ~n20529 & n20533;
  assign n20535 = n20534 ^ n20528;
  assign n20476 = n20475 ^ n20471;
  assign n20477 = n20472 & n20476;
  assign n20478 = n20477 ^ n17479;
  assign n20438 = n19895 ^ n18719;
  assign n20439 = n20438 ^ n18117;
  assign n20434 = n20433 ^ n20382;
  assign n20435 = n20431 & n20434;
  assign n20436 = n20435 ^ n20433;
  assign n20427 = n19739 ^ n2979;
  assign n20437 = n20436 ^ n20427;
  assign n20469 = n20439 ^ n20437;
  assign n20470 = n20469 ^ n17486;
  assign n20499 = n20478 ^ n20470;
  assign n20498 = ~n20496 & ~n20497;
  assign n20524 = n20499 ^ n20498;
  assign n20536 = n20535 ^ n20524;
  assign n20537 = n20524 ^ n1847;
  assign n20538 = ~n20536 & n20537;
  assign n20539 = n20538 ^ n1847;
  assign n20500 = n20498 & ~n20499;
  assign n20479 = n20478 ^ n20469;
  assign n20480 = ~n20470 & ~n20479;
  assign n20481 = n20480 ^ n17486;
  assign n20444 = n19353 ^ n18106;
  assign n20445 = n20444 ^ n18711;
  assign n20440 = n20439 ^ n20427;
  assign n20441 = ~n20437 & ~n20440;
  assign n20442 = n20441 ^ n20439;
  assign n20426 = n19742 ^ n19627;
  assign n20443 = n20442 ^ n20426;
  assign n20467 = n20445 ^ n20443;
  assign n20468 = n20467 ^ n17478;
  assign n20495 = n20481 ^ n20468;
  assign n20523 = n20500 ^ n20495;
  assign n20540 = n20539 ^ n20523;
  assign n20541 = n20523 ^ n1840;
  assign n20542 = ~n20540 & n20541;
  assign n20543 = n20542 ^ n1840;
  assign n20501 = ~n20495 & n20500;
  assign n20482 = n20481 ^ n20467;
  assign n20483 = n20468 & n20482;
  assign n20484 = n20483 ^ n17478;
  assign n20450 = n19349 ^ n18707;
  assign n20451 = n20450 ^ n18101;
  assign n20446 = n20445 ^ n20426;
  assign n20447 = n20443 & n20446;
  assign n20448 = n20447 ^ n20445;
  assign n20425 = n19746 ^ n2993;
  assign n20449 = n20448 ^ n20425;
  assign n20465 = n20451 ^ n20449;
  assign n20466 = n20465 ^ n17476;
  assign n20494 = n20484 ^ n20466;
  assign n20522 = n20501 ^ n20494;
  assign n20544 = n20543 ^ n20522;
  assign n20545 = n20522 ^ n1866;
  assign n20546 = ~n20544 & n20545;
  assign n20547 = n20546 ^ n1866;
  assign n20502 = ~n20494 & ~n20501;
  assign n20485 = n20484 ^ n20465;
  assign n20486 = n20466 & ~n20485;
  assign n20487 = n20486 ^ n17476;
  assign n20456 = n19347 ^ n18097;
  assign n20457 = n20456 ^ n18706;
  assign n20452 = n20451 ^ n20425;
  assign n20453 = n20449 & ~n20452;
  assign n20454 = n20453 ^ n20451;
  assign n20455 = n20454 ^ n19767;
  assign n20463 = n20457 ^ n20455;
  assign n20464 = n20463 ^ n17472;
  assign n20493 = n20487 ^ n20464;
  assign n20521 = n20502 ^ n20493;
  assign n20548 = n20547 ^ n20521;
  assign n20549 = n20521 ^ n1966;
  assign n20550 = ~n20548 & n20549;
  assign n20551 = n20550 ^ n1966;
  assign n20503 = n20493 & ~n20502;
  assign n20488 = n20487 ^ n20463;
  assign n20489 = n20464 & n20488;
  assign n20490 = n20489 ^ n17472;
  assign n20491 = n20490 ^ n16954;
  assign n20458 = n20457 ^ n19767;
  assign n20459 = n20455 & n20458;
  assign n20460 = n20459 ^ n20457;
  assign n20461 = n20460 ^ n20424;
  assign n20422 = n19346 ^ n18507;
  assign n20423 = n20422 ^ n17746;
  assign n20462 = n20461 ^ n20423;
  assign n20492 = n20491 ^ n20462;
  assign n20520 = n20503 ^ n20492;
  assign n20552 = n20551 ^ n20520;
  assign n20553 = n20520 ^ n2124;
  assign n20554 = n20552 & ~n20553;
  assign n20555 = n20554 ^ n2124;
  assign n20556 = n20555 ^ n2117;
  assign n20513 = n20462 ^ n16954;
  assign n20514 = n20490 ^ n20462;
  assign n20515 = ~n20513 & ~n20514;
  assign n20516 = n20515 ^ n16954;
  assign n20517 = n20516 ^ n16949;
  assign n20511 = n19919 ^ n1756;
  assign n20507 = n20424 ^ n20423;
  assign n20508 = n20461 & ~n20507;
  assign n20509 = n20508 ^ n20423;
  assign n20505 = n19345 ^ n18741;
  assign n20506 = n20505 ^ n17742;
  assign n20510 = n20509 ^ n20506;
  assign n20512 = n20511 ^ n20510;
  assign n20518 = n20517 ^ n20512;
  assign n20504 = n20492 & n20503;
  assign n20519 = n20518 ^ n20504;
  assign n20557 = n20556 ^ n20519;
  assign n20420 = n19035 ^ n18768;
  assign n20421 = n20420 ^ n19787;
  assign n20558 = n20557 ^ n20421;
  assign n20565 = n19795 ^ n18499;
  assign n20566 = n20565 ^ n19047;
  assign n20561 = n20540 ^ n1840;
  assign n20562 = n19968 ^ n19050;
  assign n20563 = n20562 ^ n18503;
  assign n20564 = n20561 & n20563;
  assign n20567 = n20566 ^ n20564;
  assign n20568 = n20544 ^ n1866;
  assign n20569 = n20568 ^ n20566;
  assign n20570 = ~n20567 & n20569;
  assign n20571 = n20570 ^ n20564;
  assign n20560 = n20548 ^ n1966;
  assign n20572 = n20571 ^ n20560;
  assign n20573 = n19041 ^ n18494;
  assign n20574 = n20573 ^ n19794;
  assign n20575 = n20574 ^ n20560;
  assign n20576 = ~n20572 & n20575;
  assign n20577 = n20576 ^ n20574;
  assign n20559 = n20552 ^ n2124;
  assign n20578 = n20577 ^ n20559;
  assign n20579 = n19791 ^ n19040;
  assign n20580 = n20579 ^ n18761;
  assign n20581 = n20580 ^ n20559;
  assign n20582 = n20578 & n20581;
  assign n20583 = n20582 ^ n20580;
  assign n20584 = n20583 ^ n20557;
  assign n20585 = n20558 & ~n20584;
  assign n20586 = n20585 ^ n20421;
  assign n20419 = n20188 ^ n2321;
  assign n20587 = n20586 ^ n20419;
  assign n20588 = n19786 ^ n18492;
  assign n20589 = n20588 ^ n19034;
  assign n20590 = n20589 ^ n20419;
  assign n20591 = ~n20587 & ~n20590;
  assign n20592 = n20591 ^ n20589;
  assign n20593 = n20592 ^ n20417;
  assign n20594 = ~n20418 & n20593;
  assign n20595 = n20594 ^ n20416;
  assign n20414 = n20286 ^ n20280;
  assign n20596 = n20595 ^ n20414;
  assign n20597 = n19784 ^ n19023;
  assign n20598 = n20597 ^ n18782;
  assign n20599 = n20598 ^ n20414;
  assign n20600 = n20596 & n20599;
  assign n20601 = n20600 ^ n20598;
  assign n20602 = n20601 ^ n20412;
  assign n20603 = ~n20413 & n20602;
  assign n20604 = n20603 ^ n20411;
  assign n20409 = n20292 ^ n20270;
  assign n20605 = n20604 ^ n20409;
  assign n20606 = n19013 ^ n18985;
  assign n20607 = n20606 ^ n19781;
  assign n20608 = n20607 ^ n20409;
  assign n20609 = n20605 & n20608;
  assign n20610 = n20609 ^ n20607;
  assign n20611 = n20610 ^ n20405;
  assign n20612 = n20408 & n20611;
  assign n20613 = n20612 ^ n20407;
  assign n20615 = n20614 ^ n20613;
  assign n20616 = n20029 ^ n19030;
  assign n20617 = n20616 ^ n19006;
  assign n20618 = n20617 ^ n20614;
  assign n20619 = n20615 & n20618;
  assign n20620 = n20619 ^ n20617;
  assign n20621 = n20620 ^ n20401;
  assign n20622 = n20404 & n20621;
  assign n20623 = n20622 ^ n20403;
  assign n20625 = n20624 ^ n20623;
  assign n20626 = n19019 ^ n19000;
  assign n20627 = n20626 ^ n19774;
  assign n20628 = n20627 ^ n20624;
  assign n20629 = ~n20625 & ~n20628;
  assign n20630 = n20629 ^ n20627;
  assign n20631 = n20630 ^ n20399;
  assign n20632 = n20400 & ~n20631;
  assign n20633 = n20632 ^ n20398;
  assign n20396 = n20313 ^ n924;
  assign n20634 = n20633 ^ n20396;
  assign n20668 = n20636 ^ n20634;
  assign n20669 = n20668 ^ n18532;
  assign n20670 = n20630 ^ n20400;
  assign n20671 = n20670 ^ n18474;
  assign n20672 = n20627 ^ n20625;
  assign n20673 = n20672 ^ n18304;
  assign n20674 = n20620 ^ n20404;
  assign n20675 = n20674 ^ n18193;
  assign n20676 = n20617 ^ n20615;
  assign n20677 = n20676 ^ n17703;
  assign n20678 = n20610 ^ n20408;
  assign n20679 = n20678 ^ n17708;
  assign n20680 = n20607 ^ n20605;
  assign n20681 = n20680 ^ n18176;
  assign n20682 = n20601 ^ n20413;
  assign n20683 = n20682 ^ n17709;
  assign n20684 = n20598 ^ n20596;
  assign n20685 = n20684 ^ n17714;
  assign n20686 = n20592 ^ n20418;
  assign n20687 = n20686 ^ n17719;
  assign n20688 = n20589 ^ n20587;
  assign n20689 = n20688 ^ n18156;
  assign n20690 = n20583 ^ n20558;
  assign n20691 = n20690 ^ n17724;
  assign n20692 = n20580 ^ n20578;
  assign n20693 = n20692 ^ n17726;
  assign n20694 = n20574 ^ n20572;
  assign n20695 = n20694 ^ n17734;
  assign n20696 = n20563 ^ n20561;
  assign n20697 = n17738 & n20696;
  assign n20698 = n20697 ^ n18140;
  assign n20699 = n20568 ^ n20567;
  assign n20700 = n20699 ^ n20697;
  assign n20701 = ~n20698 & n20700;
  assign n20702 = n20701 ^ n18140;
  assign n20703 = n20702 ^ n20694;
  assign n20704 = n20695 & n20703;
  assign n20705 = n20704 ^ n17734;
  assign n20706 = n20705 ^ n20692;
  assign n20707 = ~n20693 & ~n20706;
  assign n20708 = n20707 ^ n17726;
  assign n20709 = n20708 ^ n20690;
  assign n20710 = ~n20691 & ~n20709;
  assign n20711 = n20710 ^ n17724;
  assign n20712 = n20711 ^ n20688;
  assign n20713 = ~n20689 & ~n20712;
  assign n20714 = n20713 ^ n18156;
  assign n20715 = n20714 ^ n20686;
  assign n20716 = ~n20687 & ~n20715;
  assign n20717 = n20716 ^ n17719;
  assign n20718 = n20717 ^ n20684;
  assign n20719 = n20685 & ~n20718;
  assign n20720 = n20719 ^ n17714;
  assign n20721 = n20720 ^ n20682;
  assign n20722 = n20683 & ~n20721;
  assign n20723 = n20722 ^ n17709;
  assign n20724 = n20723 ^ n20680;
  assign n20725 = n20681 & n20724;
  assign n20726 = n20725 ^ n18176;
  assign n20727 = n20726 ^ n20678;
  assign n20728 = ~n20679 & n20727;
  assign n20729 = n20728 ^ n17708;
  assign n20730 = n20729 ^ n20676;
  assign n20731 = n20677 & ~n20730;
  assign n20732 = n20731 ^ n17703;
  assign n20733 = n20732 ^ n20674;
  assign n20734 = n20675 & n20733;
  assign n20735 = n20734 ^ n18193;
  assign n20736 = n20735 ^ n20672;
  assign n20737 = ~n20673 & ~n20736;
  assign n20738 = n20737 ^ n18304;
  assign n20739 = n20738 ^ n20670;
  assign n20740 = n20671 & n20739;
  assign n20741 = n20740 ^ n18474;
  assign n20742 = n20741 ^ n20668;
  assign n20743 = n20669 & ~n20742;
  assign n20744 = n20743 ^ n18532;
  assign n20637 = n20636 ^ n20396;
  assign n20638 = n20634 & n20637;
  assign n20639 = n20638 ^ n20636;
  assign n20393 = n19568 ^ n19079;
  assign n20394 = n20393 ^ n20055;
  assign n20392 = n20316 ^ n20256;
  assign n20395 = n20394 ^ n20392;
  assign n20666 = n20639 ^ n20395;
  assign n20667 = n20666 ^ n18526;
  assign n20804 = n20744 ^ n20667;
  assign n20773 = n20741 ^ n20669;
  assign n20774 = n20738 ^ n20671;
  assign n20775 = n20732 ^ n20675;
  assign n20776 = n20720 ^ n20683;
  assign n20777 = n20717 ^ n20685;
  assign n20778 = n20711 ^ n20689;
  assign n20779 = n20699 ^ n20698;
  assign n20780 = n20696 ^ n17738;
  assign n20781 = n20779 & n20780;
  assign n20782 = n20702 ^ n20695;
  assign n20783 = n20781 & ~n20782;
  assign n20784 = n20705 ^ n20693;
  assign n20785 = n20783 & ~n20784;
  assign n20786 = n20708 ^ n20691;
  assign n20787 = n20785 & n20786;
  assign n20788 = n20778 & ~n20787;
  assign n20789 = n20714 ^ n20687;
  assign n20790 = ~n20788 & n20789;
  assign n20791 = ~n20777 & ~n20790;
  assign n20792 = ~n20776 & n20791;
  assign n20793 = n20723 ^ n20681;
  assign n20794 = n20792 & ~n20793;
  assign n20795 = n20726 ^ n20679;
  assign n20796 = ~n20794 & n20795;
  assign n20797 = n20729 ^ n20677;
  assign n20798 = ~n20796 & n20797;
  assign n20799 = ~n20775 & ~n20798;
  assign n20800 = n20735 ^ n20673;
  assign n20801 = ~n20799 & n20800;
  assign n20802 = n20774 & n20801;
  assign n20803 = ~n20773 & n20802;
  assign n20819 = n20804 ^ n20803;
  assign n2450 = n2428 ^ x496;
  assign n2451 = n2450 ^ n2447;
  assign n2452 = n2451 ^ x432;
  assign n20820 = n20819 ^ n2452;
  assign n20821 = n20802 ^ n20773;
  assign n2441 = n2419 ^ x497;
  assign n2442 = n2441 ^ n1387;
  assign n2443 = n2442 ^ x433;
  assign n20822 = n20821 ^ n2443;
  assign n20824 = n20800 ^ n20799;
  assign n20825 = n20824 ^ n1192;
  assign n20826 = n20798 ^ n20775;
  assign n1181 = n1090 ^ x500;
  assign n1182 = n1181 ^ n1032;
  assign n1183 = n1182 ^ x436;
  assign n20827 = n20826 ^ n1183;
  assign n20828 = n20797 ^ n20796;
  assign n1023 = n936 ^ x501;
  assign n1024 = n1023 ^ n1020;
  assign n1025 = n1024 ^ x437;
  assign n20829 = n20828 ^ n1025;
  assign n20831 = n20793 ^ n20792;
  assign n20832 = n20831 ^ n897;
  assign n20834 = n20790 ^ n20777;
  assign n20835 = n20834 ^ n3301;
  assign n20836 = n20789 ^ n20788;
  assign n20840 = n20839 ^ n20836;
  assign n20843 = n18924 ^ x508;
  assign n20844 = n20843 ^ n638;
  assign n20845 = n20844 ^ x444;
  assign n20842 = n20786 ^ n20785;
  assign n20846 = n20845 ^ n20842;
  assign n20848 = n20782 ^ n20781;
  assign n20852 = n20851 ^ n20848;
  assign n20854 = n2310 ^ x511;
  assign n20855 = n20854 ^ n15939;
  assign n20856 = n20855 ^ x447;
  assign n20853 = n2251 & ~n20780;
  assign n20857 = n20856 ^ n20853;
  assign n20858 = n20780 ^ n20779;
  assign n20859 = n20858 ^ n20853;
  assign n20860 = n20857 & ~n20859;
  assign n20861 = n20860 ^ n20856;
  assign n20862 = n20861 ^ n20848;
  assign n20863 = ~n20852 & n20862;
  assign n20864 = n20863 ^ n20851;
  assign n20847 = n20784 ^ n20783;
  assign n20865 = n20864 ^ n20847;
  assign n531 = n530 ^ x509;
  assign n535 = n534 ^ n531;
  assign n536 = n535 ^ x445;
  assign n20866 = n20847 ^ n536;
  assign n20867 = n20865 & ~n20866;
  assign n20868 = n20867 ^ n536;
  assign n20869 = n20868 ^ n20842;
  assign n20870 = n20846 & ~n20869;
  assign n20871 = n20870 ^ n20845;
  assign n20841 = n20787 ^ n20778;
  assign n20872 = n20871 ^ n20841;
  assign n20873 = n20841 ^ n711;
  assign n20874 = ~n20872 & n20873;
  assign n20875 = n20874 ^ n711;
  assign n20876 = n20875 ^ n20836;
  assign n20877 = ~n20840 & n20876;
  assign n20878 = n20877 ^ n20839;
  assign n20879 = n20878 ^ n20834;
  assign n20880 = ~n20835 & n20879;
  assign n20881 = n20880 ^ n3301;
  assign n20833 = n20791 ^ n20776;
  assign n20882 = n20881 ^ n20833;
  assign n20883 = n20833 ^ n888;
  assign n20884 = ~n20882 & n20883;
  assign n20885 = n20884 ^ n888;
  assign n20886 = n20885 ^ n20831;
  assign n20887 = n20832 & ~n20886;
  assign n20888 = n20887 ^ n897;
  assign n20830 = n20795 ^ n20794;
  assign n20889 = n20888 ^ n20830;
  assign n20890 = n20830 ^ n912;
  assign n20891 = n20889 & ~n20890;
  assign n20892 = n20891 ^ n912;
  assign n20893 = n20892 ^ n20828;
  assign n20894 = n20829 & ~n20893;
  assign n20895 = n20894 ^ n1025;
  assign n20896 = n20895 ^ n20826;
  assign n20897 = n20827 & ~n20896;
  assign n20898 = n20897 ^ n1183;
  assign n20899 = n20898 ^ n20824;
  assign n20900 = n20825 & ~n20899;
  assign n20901 = n20900 ^ n1192;
  assign n20823 = n20801 ^ n20774;
  assign n20902 = n20901 ^ n20823;
  assign n1378 = n1275 ^ x498;
  assign n1382 = n1381 ^ n1378;
  assign n1383 = n1382 ^ x434;
  assign n20903 = n20823 ^ n1383;
  assign n20904 = n20902 & ~n20903;
  assign n20905 = n20904 ^ n1383;
  assign n20906 = n20905 ^ n20821;
  assign n20907 = n20822 & ~n20906;
  assign n20908 = n20907 ^ n2443;
  assign n20909 = n20908 ^ n20819;
  assign n20910 = ~n20820 & n20909;
  assign n20911 = n20910 ^ n2452;
  assign n20805 = n20803 & n20804;
  assign n20745 = n20744 ^ n20666;
  assign n20746 = ~n20667 & ~n20745;
  assign n20747 = n20746 ^ n18526;
  assign n20640 = n20639 ^ n20392;
  assign n20641 = ~n20395 & ~n20640;
  assign n20642 = n20641 ^ n20394;
  assign n20389 = n19754 ^ n19001;
  assign n20390 = n20389 ^ n20171;
  assign n20388 = n20319 ^ n20254;
  assign n20391 = n20390 ^ n20388;
  assign n20664 = n20642 ^ n20391;
  assign n20665 = n20664 ^ n18522;
  assign n20772 = n20747 ^ n20665;
  assign n20817 = n20805 ^ n20772;
  assign n2497 = n2472 ^ x495;
  assign n2501 = n2500 ^ n2497;
  assign n2502 = n2501 ^ x431;
  assign n20818 = n20817 ^ n2502;
  assign n21471 = n20911 ^ n20818;
  assign n21498 = n21497 ^ n21471;
  assign n21499 = n20425 ^ n19803;
  assign n20988 = n20349 ^ n1527;
  assign n21500 = n21499 ^ n20988;
  assign n21475 = n20908 ^ n20820;
  assign n21501 = n21500 ^ n21475;
  assign n21518 = n20905 ^ n20822;
  assign n21502 = n20427 ^ n19815;
  assign n20970 = n20342 ^ n2664;
  assign n21503 = n21502 ^ n20970;
  assign n21480 = n20902 ^ n1383;
  assign n21504 = n21503 ^ n21480;
  assign n21447 = n20363 ^ n19754;
  assign n20937 = n20335 ^ n20245;
  assign n21448 = n21447 ^ n20937;
  assign n21446 = n20895 ^ n20827;
  assign n21449 = n21448 ^ n21446;
  assign n21342 = n20892 ^ n20829;
  assign n21340 = n20230 ^ n19568;
  assign n20765 = n20332 ^ n20247;
  assign n21341 = n21340 ^ n20765;
  assign n21343 = n21342 ^ n21341;
  assign n21328 = n20889 ^ n912;
  assign n20953 = n20865 ^ n536;
  assign n20951 = n19779 ^ n19018;
  assign n20952 = n20951 ^ n20624;
  assign n20954 = n20953 ^ n20952;
  assign n20958 = n20858 ^ n20857;
  assign n20956 = n19783 ^ n19029;
  assign n20957 = n20956 ^ n20614;
  assign n20959 = n20958 ^ n20957;
  assign n20961 = n19784 ^ n19034;
  assign n20962 = n20961 ^ n20405;
  assign n20960 = n20780 ^ n2251;
  assign n20963 = n20962 ^ n20960;
  assign n21157 = n19786 ^ n19040;
  assign n21158 = n21157 ^ n20412;
  assign n21144 = n19791 ^ n19047;
  assign n21145 = n21144 ^ n20417;
  assign n21140 = n19794 ^ n19050;
  assign n21141 = n21140 ^ n20419;
  assign n20935 = n19835 ^ n19063;
  assign n20936 = n20935 ^ n20426;
  assign n20938 = n20937 ^ n20936;
  assign n20763 = n19803 ^ n19069;
  assign n20764 = n20763 ^ n20427;
  assign n20766 = n20765 ^ n20764;
  assign n20656 = n20329 ^ n20249;
  assign n20385 = n19815 ^ n18480;
  assign n20386 = n20385 ^ n20363;
  assign n20384 = n20326 ^ n1370;
  assign n20387 = n20386 ^ n20384;
  assign n20646 = n20322 ^ n20252;
  assign n20643 = n20642 ^ n20388;
  assign n20644 = n20391 & ~n20643;
  assign n20645 = n20644 ^ n20390;
  assign n20647 = n20646 ^ n20645;
  assign n20648 = n19805 ^ n19075;
  assign n20649 = n20648 ^ n20230;
  assign n20650 = n20649 ^ n20646;
  assign n20651 = n20647 & n20650;
  assign n20652 = n20651 ^ n20649;
  assign n20653 = n20652 ^ n20384;
  assign n20654 = n20387 & n20653;
  assign n20655 = n20654 ^ n20386;
  assign n20657 = n20656 ^ n20655;
  assign n20381 = n19822 ^ n19138;
  assign n20383 = n20382 ^ n20381;
  assign n20760 = n20656 ^ n20383;
  assign n20761 = n20657 & ~n20760;
  assign n20762 = n20761 ^ n20383;
  assign n20932 = n20765 ^ n20762;
  assign n20933 = n20766 & ~n20932;
  assign n20934 = n20933 ^ n20764;
  assign n20939 = n20938 ^ n20934;
  assign n20940 = n20939 ^ n18615;
  assign n20767 = n20766 ^ n20762;
  assign n20768 = n20767 ^ n18481;
  assign n20658 = n20657 ^ n20383;
  assign n20659 = n20658 ^ n18512;
  assign n20660 = n20652 ^ n20387;
  assign n20661 = n20660 ^ n18519;
  assign n20662 = n20649 ^ n20647;
  assign n20663 = n20662 ^ n18546;
  assign n20748 = n20747 ^ n20664;
  assign n20749 = ~n20665 & n20748;
  assign n20750 = n20749 ^ n18522;
  assign n20751 = n20750 ^ n20662;
  assign n20752 = ~n20663 & n20751;
  assign n20753 = n20752 ^ n18546;
  assign n20754 = n20753 ^ n20660;
  assign n20755 = ~n20661 & ~n20754;
  assign n20756 = n20755 ^ n18519;
  assign n20757 = n20756 ^ n20658;
  assign n20758 = ~n20659 & n20757;
  assign n20759 = n20758 ^ n18512;
  assign n20929 = n20767 ^ n20759;
  assign n20930 = n20768 & ~n20929;
  assign n20931 = n20930 ^ n18481;
  assign n21026 = n20939 ^ n20931;
  assign n21027 = n20940 & ~n21026;
  assign n21028 = n21027 ^ n18615;
  assign n20977 = n19843 ^ n19062;
  assign n20978 = n20977 ^ n20425;
  assign n20973 = n20937 ^ n20934;
  assign n20974 = n20938 & n20973;
  assign n20975 = n20974 ^ n20936;
  assign n20972 = n20338 ^ n20243;
  assign n20976 = n20975 ^ n20972;
  assign n21024 = n20978 ^ n20976;
  assign n21025 = n21024 ^ n18628;
  assign n21051 = n21028 ^ n21025;
  assign n20941 = n20940 ^ n20931;
  assign n20769 = n20768 ^ n20759;
  assign n20770 = n20753 ^ n20661;
  assign n20771 = n20750 ^ n20663;
  assign n20806 = n20772 & ~n20805;
  assign n20807 = n20771 & n20806;
  assign n20808 = ~n20770 & ~n20807;
  assign n20809 = n20756 ^ n20659;
  assign n20810 = n20808 & n20809;
  assign n20942 = n20769 & ~n20810;
  assign n21052 = ~n20941 & ~n20942;
  assign n21053 = ~n21051 & n21052;
  assign n21029 = n21028 ^ n21024;
  assign n21030 = n21025 & ~n21029;
  assign n21031 = n21030 ^ n18628;
  assign n20979 = n20978 ^ n20972;
  assign n20980 = ~n20976 & ~n20979;
  assign n20981 = n20980 ^ n20978;
  assign n20968 = n19895 ^ n19060;
  assign n20969 = n20968 ^ n19767;
  assign n20971 = n20970 ^ n20969;
  assign n21022 = n20981 ^ n20971;
  assign n21023 = n21022 ^ n18640;
  assign n21054 = n21031 ^ n21023;
  assign n21055 = ~n21053 & n21054;
  assign n21032 = n21031 ^ n21022;
  assign n21033 = n21023 & ~n21032;
  assign n21034 = n21033 ^ n18640;
  assign n20982 = n20981 ^ n20970;
  assign n20983 = n20971 & n20982;
  assign n20984 = n20983 ^ n20969;
  assign n20966 = n20345 ^ n20240;
  assign n20964 = n19353 ^ n18714;
  assign n20965 = n20964 ^ n20424;
  assign n20967 = n20966 ^ n20965;
  assign n21020 = n20984 ^ n20967;
  assign n21021 = n21020 ^ n18112;
  assign n21050 = n21034 ^ n21021;
  assign n21098 = n21055 ^ n21050;
  assign n21099 = n21098 ^ n1665;
  assign n21100 = n21054 ^ n21053;
  assign n21101 = n21100 ^ n1612;
  assign n20943 = n20942 ^ n20941;
  assign n20944 = n20943 ^ n2860;
  assign n20812 = n20809 ^ n20808;
  assign n20813 = n20812 ^ n2840;
  assign n20815 = n20806 ^ n20771;
  assign n20816 = n20815 ^ n3062;
  assign n20912 = n20911 ^ n20817;
  assign n20913 = ~n20818 & n20912;
  assign n20914 = n20913 ^ n2502;
  assign n20915 = n20914 ^ n20815;
  assign n20916 = n20816 & ~n20915;
  assign n20917 = n20916 ^ n3062;
  assign n20814 = n20807 ^ n20770;
  assign n20918 = n20917 ^ n20814;
  assign n20919 = n20814 ^ n2579;
  assign n20920 = n20918 & ~n20919;
  assign n20921 = n20920 ^ n2579;
  assign n20922 = n20921 ^ n20812;
  assign n20923 = ~n20813 & n20922;
  assign n20924 = n20923 ^ n2840;
  assign n20811 = n20810 ^ n20769;
  assign n20925 = n20924 ^ n20811;
  assign n20926 = n20811 ^ n2834;
  assign n20927 = n20925 & ~n20926;
  assign n20928 = n20927 ^ n2834;
  assign n21103 = n20943 ^ n20928;
  assign n21104 = ~n20944 & n21103;
  assign n21105 = n21104 ^ n2860;
  assign n21102 = n21052 ^ n21051;
  assign n21106 = n21105 ^ n21102;
  assign n21107 = n21102 ^ n1508;
  assign n21108 = ~n21106 & n21107;
  assign n21109 = n21108 ^ n1508;
  assign n21110 = n21109 ^ n21100;
  assign n21111 = ~n21101 & n21110;
  assign n21112 = n21111 ^ n1612;
  assign n21113 = n21112 ^ n21098;
  assign n21114 = ~n21099 & n21113;
  assign n21115 = n21114 ^ n1665;
  assign n21056 = ~n21050 & ~n21055;
  assign n21035 = n21034 ^ n21020;
  assign n21036 = n21021 & ~n21035;
  assign n21037 = n21036 ^ n18112;
  assign n20990 = n19349 ^ n18719;
  assign n20991 = n20990 ^ n20511;
  assign n20985 = n20984 ^ n20966;
  assign n20986 = ~n20967 & ~n20985;
  assign n20987 = n20986 ^ n20965;
  assign n20989 = n20988 ^ n20987;
  assign n21018 = n20991 ^ n20989;
  assign n21019 = n21018 ^ n18117;
  assign n21049 = n21037 ^ n21019;
  assign n21097 = n21056 ^ n21049;
  assign n21116 = n21115 ^ n21097;
  assign n21120 = n21119 ^ n21097;
  assign n21121 = n21116 & ~n21120;
  assign n21122 = n21121 ^ n21119;
  assign n21057 = n21049 & n21056;
  assign n21038 = n21037 ^ n21018;
  assign n21039 = ~n21019 & n21038;
  assign n21040 = n21039 ^ n18117;
  assign n20997 = n19347 ^ n18711;
  assign n20998 = n20997 ^ n19947;
  assign n20992 = n20991 ^ n20988;
  assign n20993 = n20989 & ~n20992;
  assign n20994 = n20993 ^ n20991;
  assign n20996 = n20995 ^ n20994;
  assign n21016 = n20998 ^ n20996;
  assign n21017 = n21016 ^ n18106;
  assign n21048 = n21040 ^ n21017;
  assign n21095 = n21057 ^ n21048;
  assign n21096 = n21095 ^ n1751;
  assign n21142 = n21122 ^ n21096;
  assign n21143 = n21141 & n21142;
  assign n21146 = n21145 ^ n21143;
  assign n21123 = n21122 ^ n21095;
  assign n21124 = n21096 & ~n21123;
  assign n21125 = n21124 ^ n1751;
  assign n21041 = n21040 ^ n21016;
  assign n21042 = n21017 & n21041;
  assign n21043 = n21042 ^ n18106;
  assign n21004 = n19346 ^ n18707;
  assign n21005 = n21004 ^ n19952;
  assign n20999 = n20998 ^ n20995;
  assign n21000 = n20996 & ~n20999;
  assign n21001 = n21000 ^ n20998;
  assign n21003 = n21002 ^ n21001;
  assign n21014 = n21005 ^ n21003;
  assign n21015 = n21014 ^ n18101;
  assign n21059 = n21043 ^ n21015;
  assign n21058 = ~n21048 & n21057;
  assign n21094 = n21059 ^ n21058;
  assign n21126 = n21125 ^ n21094;
  assign n21147 = n21126 ^ n2076;
  assign n21148 = n21147 ^ n21145;
  assign n21149 = ~n21146 & n21148;
  assign n21150 = n21149 ^ n21143;
  assign n21127 = n21094 ^ n2076;
  assign n21128 = ~n21126 & n21127;
  assign n21129 = n21128 ^ n2076;
  assign n21060 = ~n21058 & ~n21059;
  assign n21044 = n21043 ^ n21014;
  assign n21045 = n21015 & ~n21044;
  assign n21046 = n21045 ^ n18101;
  assign n21010 = n19345 ^ n18706;
  assign n21011 = n21010 ^ n19943;
  assign n21006 = n21005 ^ n21002;
  assign n21007 = ~n21003 & ~n21006;
  assign n21008 = n21007 ^ n21005;
  assign n20379 = n20378 ^ n20359;
  assign n21009 = n21008 ^ n20379;
  assign n21012 = n21011 ^ n21009;
  assign n21013 = n21012 ^ n18097;
  assign n21047 = n21046 ^ n21013;
  assign n21092 = n21060 ^ n21047;
  assign n21093 = n21092 ^ n2082;
  assign n21139 = n21129 ^ n21093;
  assign n21151 = n21150 ^ n21139;
  assign n21152 = n19787 ^ n19041;
  assign n21153 = n21152 ^ n20414;
  assign n21154 = n21153 ^ n21139;
  assign n21155 = n21151 & n21154;
  assign n21156 = n21155 ^ n21153;
  assign n21159 = n21158 ^ n21156;
  assign n21130 = n21129 ^ n21092;
  assign n21131 = ~n21093 & n21130;
  assign n21132 = n21131 ^ n2082;
  assign n21070 = n21046 ^ n21012;
  assign n21071 = ~n21013 & n21070;
  assign n21072 = n21071 ^ n18097;
  assign n21073 = n21072 ^ n17746;
  assign n21065 = n21011 ^ n20379;
  assign n21066 = ~n21009 & ~n21065;
  assign n21067 = n21066 ^ n21011;
  assign n21064 = n20532 ^ n20529;
  assign n21068 = n21067 ^ n21064;
  assign n21062 = n19378 ^ n18507;
  assign n21063 = n21062 ^ n19940;
  assign n21069 = n21068 ^ n21063;
  assign n21074 = n21073 ^ n21069;
  assign n21061 = ~n21047 & ~n21060;
  assign n21091 = n21074 ^ n21061;
  assign n21133 = n21132 ^ n21091;
  assign n21160 = n21133 ^ n2098;
  assign n21161 = n21160 ^ n21156;
  assign n21162 = ~n21159 & ~n21161;
  assign n21163 = n21162 ^ n21158;
  assign n21134 = n21091 ^ n2098;
  assign n21135 = n21133 & ~n21134;
  assign n21136 = n21135 ^ n2098;
  assign n21137 = n21136 ^ n2236;
  assign n21084 = n21069 ^ n17746;
  assign n21085 = n21072 ^ n21069;
  assign n21086 = n21084 & n21085;
  assign n21087 = n21086 ^ n17746;
  assign n21088 = n21087 ^ n17742;
  assign n21079 = n21064 ^ n21063;
  assign n21080 = n21068 & n21079;
  assign n21081 = n21080 ^ n21063;
  assign n21077 = n19054 ^ n18741;
  assign n21078 = n21077 ^ n19938;
  assign n21082 = n21081 ^ n21078;
  assign n21076 = n20536 ^ n1847;
  assign n21083 = n21082 ^ n21076;
  assign n21089 = n21088 ^ n21083;
  assign n21075 = n21061 & n21074;
  assign n21090 = n21089 ^ n21075;
  assign n21138 = n21137 ^ n21090;
  assign n21164 = n21163 ^ n21138;
  assign n21165 = n19785 ^ n19035;
  assign n21166 = n21165 ^ n20409;
  assign n21167 = n21166 ^ n21138;
  assign n21168 = ~n21164 & ~n21167;
  assign n21169 = n21168 ^ n21166;
  assign n21170 = n21169 ^ n20960;
  assign n21171 = n20963 & ~n21170;
  assign n21172 = n21171 ^ n20962;
  assign n21173 = n21172 ^ n20958;
  assign n21174 = n20959 & n21173;
  assign n21175 = n21174 ^ n20957;
  assign n20955 = n20861 ^ n20852;
  assign n21176 = n21175 ^ n20955;
  assign n21177 = n19781 ^ n19023;
  assign n21178 = n21177 ^ n20401;
  assign n21179 = n21178 ^ n20955;
  assign n21180 = n21176 & n21179;
  assign n21181 = n21180 ^ n21178;
  assign n21182 = n21181 ^ n20953;
  assign n21183 = n20954 & ~n21182;
  assign n21184 = n21183 ^ n20952;
  assign n20950 = n20868 ^ n20846;
  assign n21185 = n21184 ^ n20950;
  assign n21186 = n20029 ^ n19013;
  assign n21187 = n21186 ^ n20399;
  assign n21188 = n21187 ^ n20950;
  assign n21189 = n21185 & n21188;
  assign n21190 = n21189 ^ n21187;
  assign n20949 = n20872 ^ n711;
  assign n21191 = n21190 ^ n20949;
  assign n20947 = n19775 ^ n19008;
  assign n20948 = n20947 ^ n20396;
  assign n21248 = n20949 ^ n20948;
  assign n21249 = ~n21191 & n21248;
  assign n21250 = n21249 ^ n20948;
  assign n21247 = n20875 ^ n20840;
  assign n21251 = n21250 ^ n21247;
  assign n21245 = n19774 ^ n19006;
  assign n21246 = n21245 ^ n20392;
  assign n21283 = n21247 ^ n21246;
  assign n21284 = n21251 & n21283;
  assign n21285 = n21284 ^ n21246;
  assign n21282 = n20878 ^ n20835;
  assign n21286 = n21285 ^ n21282;
  assign n21280 = n19769 ^ n19004;
  assign n21281 = n21280 ^ n20388;
  assign n21297 = n21282 ^ n21281;
  assign n21298 = ~n21286 & ~n21297;
  assign n21299 = n21298 ^ n21281;
  assign n21296 = n20882 ^ n888;
  assign n21300 = n21299 ^ n21296;
  assign n21294 = n20048 ^ n19000;
  assign n21295 = n21294 ^ n20646;
  assign n21312 = n21296 ^ n21295;
  assign n21313 = ~n21300 & ~n21312;
  assign n21314 = n21313 ^ n21295;
  assign n21311 = n20885 ^ n20832;
  assign n21315 = n21314 ^ n21311;
  assign n21309 = n20055 ^ n18998;
  assign n21310 = n21309 ^ n20384;
  assign n21325 = n21311 ^ n21310;
  assign n21326 = n21315 & n21325;
  assign n21327 = n21326 ^ n21310;
  assign n21329 = n21328 ^ n21327;
  assign n21323 = n20171 ^ n19447;
  assign n21324 = n21323 ^ n20656;
  assign n21337 = n21328 ^ n21324;
  assign n21338 = n21329 & ~n21337;
  assign n21339 = n21338 ^ n21324;
  assign n21443 = n21342 ^ n21339;
  assign n21444 = ~n21343 & ~n21443;
  assign n21445 = n21444 ^ n21341;
  assign n21506 = n21446 ^ n21445;
  assign n21507 = n21449 & n21506;
  assign n21508 = n21507 ^ n21448;
  assign n21505 = n20898 ^ n20825;
  assign n21509 = n21508 ^ n21505;
  assign n21510 = n20382 ^ n19805;
  assign n21511 = n21510 ^ n20972;
  assign n21512 = n21511 ^ n21505;
  assign n21513 = ~n21509 & n21512;
  assign n21514 = n21513 ^ n21511;
  assign n21515 = n21514 ^ n21480;
  assign n21516 = n21504 & n21515;
  assign n21517 = n21516 ^ n21503;
  assign n21519 = n21518 ^ n21517;
  assign n21520 = n20426 ^ n19822;
  assign n21521 = n21520 ^ n20966;
  assign n21522 = n21521 ^ n21518;
  assign n21523 = n21519 & n21522;
  assign n21524 = n21523 ^ n21521;
  assign n21525 = n21524 ^ n21475;
  assign n21526 = n21501 & n21525;
  assign n21527 = n21526 ^ n21500;
  assign n21528 = n21527 ^ n21471;
  assign n21529 = ~n21498 & ~n21528;
  assign n21530 = n21529 ^ n21497;
  assign n21495 = n20914 ^ n20816;
  assign n21531 = n21530 ^ n21495;
  assign n21567 = n21533 ^ n21531;
  assign n21568 = n21567 ^ n19062;
  assign n21569 = n21527 ^ n21498;
  assign n21570 = n21569 ^ n19063;
  assign n21571 = n21524 ^ n21501;
  assign n21572 = n21571 ^ n19069;
  assign n21573 = n21521 ^ n21519;
  assign n21574 = n21573 ^ n19138;
  assign n21575 = n21514 ^ n21504;
  assign n21576 = n21575 ^ n18480;
  assign n21577 = n21511 ^ n21509;
  assign n21578 = n21577 ^ n19075;
  assign n21450 = n21449 ^ n21445;
  assign n21451 = n21450 ^ n19001;
  assign n21344 = n21343 ^ n21339;
  assign n21345 = n21344 ^ n19079;
  assign n21330 = n21329 ^ n21324;
  assign n21331 = n21330 ^ n19009;
  assign n21316 = n21315 ^ n21310;
  assign n21319 = n21316 ^ n19014;
  assign n21301 = n21300 ^ n21295;
  assign n21302 = n21301 ^ n19019;
  assign n21287 = n21286 ^ n21281;
  assign n21288 = n21287 ^ n19024;
  assign n21252 = n21251 ^ n21246;
  assign n21253 = n21252 ^ n19030;
  assign n21192 = n21191 ^ n20948;
  assign n21193 = n21192 ^ n19089;
  assign n21194 = n21187 ^ n21185;
  assign n21195 = n21194 ^ n18985;
  assign n21196 = n21181 ^ n20954;
  assign n21197 = n21196 ^ n18861;
  assign n21198 = n21178 ^ n21176;
  assign n21199 = n21198 ^ n18782;
  assign n21200 = n21172 ^ n20959;
  assign n21201 = n21200 ^ n18488;
  assign n21202 = n21169 ^ n20963;
  assign n21203 = n21202 ^ n18492;
  assign n21204 = n21166 ^ n21164;
  assign n21205 = n21204 ^ n18768;
  assign n21206 = n21160 ^ n21158;
  assign n21207 = n21206 ^ n21156;
  assign n21208 = n21207 ^ n18761;
  assign n21209 = n21153 ^ n21151;
  assign n21210 = n21209 ^ n18494;
  assign n21211 = n21142 ^ n21141;
  assign n21212 = ~n18503 & n21211;
  assign n21213 = n21212 ^ n18499;
  assign n21214 = n21147 ^ n21146;
  assign n21215 = n21214 ^ n21212;
  assign n21216 = n21213 & n21215;
  assign n21217 = n21216 ^ n18499;
  assign n21218 = n21217 ^ n21209;
  assign n21219 = n21210 & ~n21218;
  assign n21220 = n21219 ^ n18494;
  assign n21221 = n21220 ^ n21207;
  assign n21222 = n21208 & ~n21221;
  assign n21223 = n21222 ^ n18761;
  assign n21224 = n21223 ^ n21204;
  assign n21225 = ~n21205 & n21224;
  assign n21226 = n21225 ^ n18768;
  assign n21227 = n21226 ^ n21202;
  assign n21228 = n21203 & n21227;
  assign n21229 = n21228 ^ n18492;
  assign n21230 = n21229 ^ n21200;
  assign n21231 = n21201 & ~n21230;
  assign n21232 = n21231 ^ n18488;
  assign n21233 = n21232 ^ n21198;
  assign n21234 = ~n21199 & n21233;
  assign n21235 = n21234 ^ n18782;
  assign n21236 = n21235 ^ n21196;
  assign n21237 = n21197 & ~n21236;
  assign n21238 = n21237 ^ n18861;
  assign n21239 = n21238 ^ n21194;
  assign n21240 = ~n21195 & ~n21239;
  assign n21241 = n21240 ^ n18985;
  assign n21242 = n21241 ^ n21192;
  assign n21243 = ~n21193 & ~n21242;
  assign n21244 = n21243 ^ n19089;
  assign n21277 = n21252 ^ n21244;
  assign n21278 = ~n21253 & n21277;
  assign n21279 = n21278 ^ n19030;
  assign n21291 = n21287 ^ n21279;
  assign n21292 = n21288 & n21291;
  assign n21293 = n21292 ^ n19024;
  assign n21305 = n21301 ^ n21293;
  assign n21306 = ~n21302 & n21305;
  assign n21307 = n21306 ^ n19019;
  assign n21320 = n21316 ^ n21307;
  assign n21321 = ~n21319 & n21320;
  assign n21322 = n21321 ^ n19014;
  assign n21334 = n21330 ^ n21322;
  assign n21335 = n21331 & n21334;
  assign n21336 = n21335 ^ n19009;
  assign n21440 = n21344 ^ n21336;
  assign n21441 = n21345 & ~n21440;
  assign n21442 = n21441 ^ n19079;
  assign n21579 = n21450 ^ n21442;
  assign n21580 = ~n21451 & ~n21579;
  assign n21581 = n21580 ^ n19001;
  assign n21582 = n21581 ^ n21577;
  assign n21583 = n21578 & ~n21582;
  assign n21584 = n21583 ^ n19075;
  assign n21585 = n21584 ^ n21575;
  assign n21586 = ~n21576 & ~n21585;
  assign n21587 = n21586 ^ n18480;
  assign n21588 = n21587 ^ n21573;
  assign n21589 = n21574 & ~n21588;
  assign n21590 = n21589 ^ n19138;
  assign n21591 = n21590 ^ n21571;
  assign n21592 = ~n21572 & n21591;
  assign n21593 = n21592 ^ n19069;
  assign n21594 = n21593 ^ n21569;
  assign n21595 = ~n21570 & n21594;
  assign n21596 = n21595 ^ n19063;
  assign n21597 = n21596 ^ n21567;
  assign n21598 = ~n21568 & ~n21597;
  assign n21599 = n21598 ^ n19062;
  assign n21538 = n20511 ^ n19895;
  assign n21539 = n21538 ^ n20379;
  assign n21534 = n21533 ^ n21495;
  assign n21535 = ~n21531 & ~n21534;
  assign n21536 = n21535 ^ n21533;
  assign n21464 = n20918 ^ n2579;
  assign n21537 = n21536 ^ n21464;
  assign n21565 = n21539 ^ n21537;
  assign n21566 = n21565 ^ n19060;
  assign n21611 = n21599 ^ n21566;
  assign n21612 = n21593 ^ n21570;
  assign n21613 = n21581 ^ n21578;
  assign n21452 = n21451 ^ n21442;
  assign n21254 = n21253 ^ n21244;
  assign n21255 = n21241 ^ n21193;
  assign n21256 = n21238 ^ n21195;
  assign n21257 = n21235 ^ n21197;
  assign n21258 = n21232 ^ n21199;
  assign n21259 = n21229 ^ n21201;
  assign n21260 = n21223 ^ n21205;
  assign n21261 = n21217 ^ n21210;
  assign n21262 = n21211 ^ n18503;
  assign n21263 = n21214 ^ n21213;
  assign n21264 = ~n21262 & ~n21263;
  assign n21265 = n21261 & n21264;
  assign n21266 = n21220 ^ n21208;
  assign n21267 = n21265 & n21266;
  assign n21268 = ~n21260 & n21267;
  assign n21269 = n21226 ^ n21203;
  assign n21270 = ~n21268 & ~n21269;
  assign n21271 = ~n21259 & ~n21270;
  assign n21272 = ~n21258 & ~n21271;
  assign n21273 = n21257 & n21272;
  assign n21274 = ~n21256 & n21273;
  assign n21275 = ~n21255 & ~n21274;
  assign n21276 = ~n21254 & ~n21275;
  assign n21289 = n21288 ^ n21279;
  assign n21290 = ~n21276 & ~n21289;
  assign n21303 = n21302 ^ n21293;
  assign n21304 = ~n21290 & n21303;
  assign n21308 = n21307 ^ n19014;
  assign n21317 = n21316 ^ n21308;
  assign n21318 = n21304 & n21317;
  assign n21332 = n21331 ^ n21322;
  assign n21333 = n21318 & ~n21332;
  assign n21346 = n21345 ^ n21336;
  assign n21453 = n21333 & n21346;
  assign n21614 = n21452 & ~n21453;
  assign n21615 = n21613 & n21614;
  assign n21616 = n21584 ^ n21576;
  assign n21617 = ~n21615 & n21616;
  assign n21618 = n21587 ^ n21574;
  assign n21619 = n21617 & n21618;
  assign n21620 = n21590 ^ n21572;
  assign n21621 = ~n21619 & n21620;
  assign n21622 = ~n21612 & ~n21621;
  assign n21623 = n21596 ^ n21568;
  assign n21624 = n21622 & ~n21623;
  assign n21625 = n21611 & ~n21624;
  assign n21600 = n21599 ^ n21565;
  assign n21601 = n21566 & n21600;
  assign n21602 = n21601 ^ n19060;
  assign n21545 = n19947 ^ n19353;
  assign n21546 = n21545 ^ n21064;
  assign n21543 = n20921 ^ n20813;
  assign n21540 = n21539 ^ n21464;
  assign n21541 = ~n21537 & n21540;
  assign n21542 = n21541 ^ n21539;
  assign n21544 = n21543 ^ n21542;
  assign n21563 = n21546 ^ n21544;
  assign n21564 = n21563 ^ n18714;
  assign n21610 = n21602 ^ n21564;
  assign n21692 = n21625 ^ n21610;
  assign n21693 = n21692 ^ n1740;
  assign n21694 = n21624 ^ n21611;
  assign n21698 = n21697 ^ n21694;
  assign n21700 = n21621 ^ n21612;
  assign n21701 = n21700 ^ n3122;
  assign n21703 = n21618 ^ n21617;
  assign n21704 = n21703 ^ n1565;
  assign n21706 = n21614 ^ n21613;
  assign n2562 = n2522 ^ n1515;
  assign n2563 = n2562 ^ n2559;
  assign n2564 = n2563 ^ x462;
  assign n21707 = n21706 ^ n2564;
  assign n21454 = n21453 ^ n21452;
  assign n21455 = n21454 ^ n2555;
  assign n21347 = n21346 ^ n21333;
  assign n3158 = n3151 ^ n2458;
  assign n3162 = n3161 ^ n3158;
  assign n3163 = n3162 ^ x464;
  assign n21348 = n21347 ^ n3163;
  assign n21349 = n21332 ^ n21318;
  assign n21353 = n21352 ^ n21349;
  assign n21355 = n21303 ^ n21290;
  assign n1306 = n1287 ^ n1200;
  assign n1307 = n1306 ^ n1166;
  assign n1308 = n1307 ^ x467;
  assign n21356 = n21355 ^ n1308;
  assign n21357 = n21289 ^ n21276;
  assign n1154 = n1114 ^ n1066;
  assign n1155 = n1154 ^ n1135;
  assign n1156 = n1155 ^ x468;
  assign n21358 = n21357 ^ n1156;
  assign n21359 = n21275 ^ n21254;
  assign n21360 = n21359 ^ n1131;
  assign n21362 = n21273 ^ n21256;
  assign n21363 = n21362 ^ n797;
  assign n21365 = n21271 ^ n21258;
  assign n21366 = n21365 ^ n614;
  assign n21367 = n21270 ^ n21259;
  assign n21368 = n21367 ^ n650;
  assign n21370 = n21267 ^ n21260;
  assign n21371 = n21370 ^ n3284;
  assign n21372 = n21266 ^ n21265;
  assign n21376 = n21375 ^ n21372;
  assign n21377 = n21264 ^ n21261;
  assign n21381 = n21380 ^ n21377;
  assign n21382 = n2387 & n21262;
  assign n2403 = n2358 ^ n2297;
  assign n2404 = n2403 ^ n2327;
  assign n2405 = n2404 ^ x479;
  assign n21383 = n21382 ^ n2405;
  assign n21384 = n21263 ^ n21262;
  assign n21385 = n21384 ^ n21382;
  assign n21386 = n21383 & ~n21385;
  assign n21387 = n21386 ^ n2405;
  assign n21388 = n21387 ^ n21377;
  assign n21389 = n21381 & ~n21388;
  assign n21390 = n21389 ^ n21380;
  assign n21391 = n21390 ^ n21372;
  assign n21392 = n21376 & ~n21391;
  assign n21393 = n21392 ^ n21375;
  assign n21394 = n21393 ^ n21370;
  assign n21395 = ~n21371 & n21394;
  assign n21396 = n21395 ^ n3284;
  assign n21369 = n21269 ^ n21268;
  assign n21397 = n21396 ^ n21369;
  assign n571 = n567 ^ n558;
  assign n575 = n574 ^ n571;
  assign n576 = n575 ^ x475;
  assign n21398 = n21369 ^ n576;
  assign n21399 = n21397 & ~n21398;
  assign n21400 = n21399 ^ n576;
  assign n21401 = n21400 ^ n21367;
  assign n21402 = n21368 & ~n21401;
  assign n21403 = n21402 ^ n650;
  assign n21404 = n21403 ^ n21365;
  assign n21405 = ~n21366 & n21404;
  assign n21406 = n21405 ^ n614;
  assign n21364 = n21272 ^ n21257;
  assign n21407 = n21406 ^ n21364;
  assign n21411 = n21410 ^ n21364;
  assign n21412 = n21407 & ~n21411;
  assign n21413 = n21412 ^ n21410;
  assign n21414 = n21413 ^ n21362;
  assign n21415 = n21363 & ~n21414;
  assign n21416 = n21415 ^ n797;
  assign n21361 = n21274 ^ n21255;
  assign n21417 = n21416 ^ n21361;
  assign n21418 = n21361 ^ n1145;
  assign n21419 = ~n21417 & n21418;
  assign n21420 = n21419 ^ n1145;
  assign n21421 = n21420 ^ n21359;
  assign n21422 = ~n21360 & n21421;
  assign n21423 = n21422 ^ n1131;
  assign n21424 = n21423 ^ n21357;
  assign n21425 = n21358 & ~n21424;
  assign n21426 = n21425 ^ n1156;
  assign n21427 = n21426 ^ n21355;
  assign n21428 = n21356 & ~n21427;
  assign n21429 = n21428 ^ n1308;
  assign n21354 = n21317 ^ n21304;
  assign n21430 = n21429 ^ n21354;
  assign n1321 = n1315 ^ n1299;
  assign n1322 = n1321 ^ n1215;
  assign n1323 = n1322 ^ x466;
  assign n21431 = n21354 ^ n1323;
  assign n21432 = n21430 & ~n21431;
  assign n21433 = n21432 ^ n1323;
  assign n21434 = n21433 ^ n21349;
  assign n21435 = n21353 & ~n21434;
  assign n21436 = n21435 ^ n21352;
  assign n21437 = n21436 ^ n21347;
  assign n21438 = ~n21348 & n21437;
  assign n21439 = n21438 ^ n3163;
  assign n21708 = n21454 ^ n21439;
  assign n21709 = ~n21455 & n21708;
  assign n21710 = n21709 ^ n2555;
  assign n21711 = n21710 ^ n21706;
  assign n21712 = n21707 & ~n21711;
  assign n21713 = n21712 ^ n2564;
  assign n21705 = n21616 ^ n21615;
  assign n21714 = n21713 ^ n21705;
  assign n2639 = n2632 ^ n2584;
  assign n2640 = n2639 ^ n2571;
  assign n2641 = n2640 ^ x461;
  assign n21715 = n21705 ^ n2641;
  assign n21716 = ~n21714 & n21715;
  assign n21717 = n21716 ^ n2641;
  assign n21718 = n21717 ^ n21703;
  assign n21719 = ~n21704 & n21718;
  assign n21720 = n21719 ^ n1565;
  assign n21702 = n21620 ^ n21619;
  assign n21721 = n21720 ^ n21702;
  assign n21722 = n21702 ^ n2747;
  assign n21723 = n21721 & ~n21722;
  assign n21724 = n21723 ^ n2747;
  assign n21725 = n21724 ^ n21700;
  assign n21726 = ~n21701 & n21725;
  assign n21727 = n21726 ^ n3122;
  assign n21699 = n21623 ^ n21622;
  assign n21728 = n21727 ^ n21699;
  assign n21729 = n21699 ^ n2876;
  assign n21730 = ~n21728 & n21729;
  assign n21731 = n21730 ^ n2876;
  assign n21732 = n21731 ^ n21694;
  assign n21733 = ~n21698 & n21732;
  assign n21734 = n21733 ^ n21697;
  assign n21735 = n21734 ^ n21692;
  assign n21736 = n21693 & ~n21735;
  assign n21737 = n21736 ^ n1740;
  assign n21603 = n21602 ^ n21563;
  assign n21604 = n21564 & ~n21603;
  assign n21605 = n21604 ^ n18714;
  assign n21551 = n19952 ^ n19349;
  assign n21552 = n21551 ^ n21076;
  assign n21547 = n21546 ^ n21543;
  assign n21548 = ~n21544 & n21547;
  assign n21549 = n21548 ^ n21546;
  assign n21460 = n20925 ^ n2834;
  assign n21550 = n21549 ^ n21460;
  assign n21561 = n21552 ^ n21550;
  assign n21562 = n21561 ^ n18719;
  assign n21627 = n21605 ^ n21562;
  assign n21626 = n21610 & ~n21625;
  assign n21691 = n21627 ^ n21626;
  assign n21738 = n21737 ^ n21691;
  assign n21739 = n21691 ^ n1710;
  assign n21740 = ~n21738 & n21739;
  assign n21741 = n21740 ^ n1710;
  assign n21628 = n21626 & ~n21627;
  assign n21606 = n21605 ^ n21561;
  assign n21607 = ~n21562 & ~n21606;
  assign n21608 = n21607 ^ n18719;
  assign n21557 = n19943 ^ n19347;
  assign n21558 = n21557 ^ n20561;
  assign n21553 = n21552 ^ n21460;
  assign n21554 = ~n21550 & n21553;
  assign n21555 = n21554 ^ n21552;
  assign n20945 = n20944 ^ n20928;
  assign n21556 = n21555 ^ n20945;
  assign n21559 = n21558 ^ n21556;
  assign n21560 = n21559 ^ n18711;
  assign n21609 = n21608 ^ n21560;
  assign n21690 = n21628 ^ n21609;
  assign n21742 = n21741 ^ n21690;
  assign n1820 = n1808 ^ n1756;
  assign n1821 = n1820 ^ n1714;
  assign n1822 = n1821 ^ x453;
  assign n21762 = n21742 ^ n1822;
  assign n23272 = n21762 ^ n21142;
  assign n21870 = n20995 ^ n20426;
  assign n21871 = n21870 ^ n21543;
  assign n21868 = n21433 ^ n21353;
  assign n21466 = n21430 ^ n1323;
  assign n21463 = n20988 ^ n20427;
  assign n21465 = n21464 ^ n21463;
  assign n21467 = n21466 ^ n21465;
  assign n21470 = n20970 ^ n20363;
  assign n21472 = n21471 ^ n21470;
  assign n21469 = n21423 ^ n21358;
  assign n21473 = n21472 ^ n21469;
  assign n21477 = n21420 ^ n21360;
  assign n21474 = n20972 ^ n20230;
  assign n21476 = n21475 ^ n21474;
  assign n21478 = n21477 ^ n21476;
  assign n21846 = n21417 ^ n1145;
  assign n21482 = n21413 ^ n21363;
  assign n21479 = n20765 ^ n20055;
  assign n21481 = n21480 ^ n21479;
  assign n21483 = n21482 ^ n21481;
  assign n21836 = n21410 ^ n21407;
  assign n21486 = n21403 ^ n21366;
  assign n21484 = n20384 ^ n19769;
  assign n21485 = n21484 ^ n21446;
  assign n21487 = n21486 ^ n21485;
  assign n21826 = n21400 ^ n21368;
  assign n21490 = n21397 ^ n576;
  assign n21488 = n20388 ^ n19775;
  assign n21489 = n21488 ^ n21328;
  assign n21491 = n21490 ^ n21489;
  assign n21810 = n21390 ^ n21376;
  assign n21797 = n21384 ^ n21383;
  assign n21766 = n20412 ^ n19791;
  assign n21767 = n21766 ^ n20958;
  assign n21763 = n20414 ^ n19794;
  assign n21764 = n21763 ^ n20960;
  assign n21765 = n21762 & ~n21764;
  assign n21768 = n21767 ^ n21765;
  assign n21743 = n21690 ^ n1822;
  assign n21744 = ~n21742 & n21743;
  assign n21745 = n21744 ^ n1822;
  assign n21639 = n21608 ^ n21559;
  assign n21640 = n21560 & ~n21639;
  assign n21641 = n21640 ^ n18711;
  assign n21635 = n19940 ^ n19346;
  assign n21636 = n21635 ^ n20568;
  assign n21631 = n21558 ^ n20945;
  assign n21632 = ~n21556 & ~n21631;
  assign n21633 = n21632 ^ n21558;
  assign n21630 = n21106 ^ n1508;
  assign n21634 = n21633 ^ n21630;
  assign n21637 = n21636 ^ n21634;
  assign n21638 = n21637 ^ n18707;
  assign n21642 = n21641 ^ n21638;
  assign n21629 = ~n21609 & n21628;
  assign n21689 = n21642 ^ n21629;
  assign n21746 = n21745 ^ n21689;
  assign n21769 = n21746 ^ n1831;
  assign n21770 = n21769 ^ n21767;
  assign n21771 = n21768 & ~n21770;
  assign n21772 = n21771 ^ n21765;
  assign n21747 = n21689 ^ n1831;
  assign n21748 = ~n21746 & n21747;
  assign n21749 = n21748 ^ n1831;
  assign n21653 = n21641 ^ n21637;
  assign n21654 = ~n21638 & n21653;
  assign n21655 = n21654 ^ n18707;
  assign n21649 = n19938 ^ n19345;
  assign n21650 = n21649 ^ n20560;
  assign n21645 = n21636 ^ n21630;
  assign n21646 = ~n21634 & ~n21645;
  assign n21647 = n21646 ^ n21636;
  assign n21644 = n21109 ^ n21101;
  assign n21648 = n21647 ^ n21644;
  assign n21651 = n21650 ^ n21648;
  assign n21652 = n21651 ^ n18706;
  assign n21656 = n21655 ^ n21652;
  assign n21643 = ~n21629 & ~n21642;
  assign n21688 = n21656 ^ n21643;
  assign n21750 = n21749 ^ n21688;
  assign n21761 = n21750 ^ n1952;
  assign n21773 = n21772 ^ n21761;
  assign n21774 = n20409 ^ n19787;
  assign n21775 = n21774 ^ n20955;
  assign n21776 = n21775 ^ n21761;
  assign n21777 = n21773 & ~n21776;
  assign n21778 = n21777 ^ n21775;
  assign n21751 = n21688 ^ n1952;
  assign n21752 = n21750 & ~n21751;
  assign n21753 = n21752 ^ n1952;
  assign n21666 = n21655 ^ n21651;
  assign n21667 = n21652 & n21666;
  assign n21668 = n21667 ^ n18706;
  assign n21669 = n21668 ^ n18507;
  assign n21661 = n21650 ^ n21644;
  assign n21662 = ~n21648 & n21661;
  assign n21663 = n21662 ^ n21650;
  assign n21660 = n21112 ^ n21099;
  assign n21664 = n21663 ^ n21660;
  assign n21658 = n19968 ^ n19378;
  assign n21659 = n21658 ^ n20559;
  assign n21665 = n21664 ^ n21659;
  assign n21670 = n21669 ^ n21665;
  assign n21657 = ~n21643 & ~n21656;
  assign n21687 = n21670 ^ n21657;
  assign n21754 = n21753 ^ n21687;
  assign n21760 = n21754 ^ n2375;
  assign n21779 = n21778 ^ n21760;
  assign n21780 = n20405 ^ n19786;
  assign n21781 = n21780 ^ n20953;
  assign n21782 = n21781 ^ n21760;
  assign n21783 = ~n21779 & ~n21782;
  assign n21784 = n21783 ^ n21781;
  assign n21755 = n21687 ^ n2375;
  assign n21756 = ~n21754 & n21755;
  assign n21757 = n21756 ^ n2375;
  assign n2130 = n2129 ^ n2042;
  assign n2131 = n2130 ^ n2120;
  assign n2132 = n2131 ^ x449;
  assign n21758 = n21757 ^ n2132;
  assign n21680 = n21665 ^ n18507;
  assign n21681 = n21668 ^ n21665;
  assign n21682 = ~n21680 & ~n21681;
  assign n21683 = n21682 ^ n18507;
  assign n21684 = n21683 ^ n18741;
  assign n21678 = n21119 ^ n21116;
  assign n21674 = n21660 ^ n21659;
  assign n21675 = ~n21664 & n21674;
  assign n21676 = n21675 ^ n21659;
  assign n21672 = n19795 ^ n19054;
  assign n21673 = n21672 ^ n20557;
  assign n21677 = n21676 ^ n21673;
  assign n21679 = n21678 ^ n21677;
  assign n21685 = n21684 ^ n21679;
  assign n21671 = n21657 & ~n21670;
  assign n21686 = n21685 ^ n21671;
  assign n21759 = n21758 ^ n21686;
  assign n21785 = n21784 ^ n21759;
  assign n21786 = n20614 ^ n19785;
  assign n21787 = n21786 ^ n20950;
  assign n21788 = n21787 ^ n21759;
  assign n21789 = ~n21785 & n21788;
  assign n21790 = n21789 ^ n21787;
  assign n21494 = n21262 ^ n2387;
  assign n21791 = n21790 ^ n21494;
  assign n21792 = n20401 ^ n19784;
  assign n21793 = n21792 ^ n20949;
  assign n21794 = n21793 ^ n21494;
  assign n21795 = n21791 & ~n21794;
  assign n21796 = n21795 ^ n21793;
  assign n21798 = n21797 ^ n21796;
  assign n21799 = n20624 ^ n19783;
  assign n21800 = n21799 ^ n21247;
  assign n21801 = n21800 ^ n21797;
  assign n21802 = n21798 & n21801;
  assign n21803 = n21802 ^ n21800;
  assign n21493 = n21387 ^ n21381;
  assign n21804 = n21803 ^ n21493;
  assign n21805 = n20399 ^ n19781;
  assign n21806 = n21805 ^ n21282;
  assign n21807 = n21806 ^ n21493;
  assign n21808 = ~n21804 & ~n21807;
  assign n21809 = n21808 ^ n21806;
  assign n21811 = n21810 ^ n21809;
  assign n21812 = n20396 ^ n19779;
  assign n21813 = n21812 ^ n21296;
  assign n21814 = n21813 ^ n21810;
  assign n21815 = n21811 & ~n21814;
  assign n21816 = n21815 ^ n21813;
  assign n21492 = n21393 ^ n21371;
  assign n21817 = n21816 ^ n21492;
  assign n21818 = n20392 ^ n20029;
  assign n21819 = n21818 ^ n21311;
  assign n21820 = n21819 ^ n21492;
  assign n21821 = ~n21817 & n21820;
  assign n21822 = n21821 ^ n21819;
  assign n21823 = n21822 ^ n21490;
  assign n21824 = ~n21491 & ~n21823;
  assign n21825 = n21824 ^ n21489;
  assign n21827 = n21826 ^ n21825;
  assign n21828 = n20646 ^ n19774;
  assign n21829 = n21828 ^ n21342;
  assign n21830 = n21829 ^ n21826;
  assign n21831 = ~n21827 & n21830;
  assign n21832 = n21831 ^ n21829;
  assign n21833 = n21832 ^ n21486;
  assign n21834 = ~n21487 & n21833;
  assign n21835 = n21834 ^ n21485;
  assign n21837 = n21836 ^ n21835;
  assign n21838 = n20656 ^ n20048;
  assign n21839 = n21838 ^ n21505;
  assign n21840 = n21839 ^ n21836;
  assign n21841 = n21837 & ~n21840;
  assign n21842 = n21841 ^ n21839;
  assign n21843 = n21842 ^ n21482;
  assign n21844 = ~n21483 & ~n21843;
  assign n21845 = n21844 ^ n21481;
  assign n21847 = n21846 ^ n21845;
  assign n21848 = n20937 ^ n20171;
  assign n21849 = n21848 ^ n21518;
  assign n21850 = n21849 ^ n21846;
  assign n21851 = n21847 & ~n21850;
  assign n21852 = n21851 ^ n21849;
  assign n21853 = n21852 ^ n21477;
  assign n21854 = ~n21478 & ~n21853;
  assign n21855 = n21854 ^ n21476;
  assign n21856 = n21855 ^ n21469;
  assign n21857 = ~n21473 & ~n21856;
  assign n21858 = n21857 ^ n21472;
  assign n21468 = n21426 ^ n21356;
  assign n21859 = n21858 ^ n21468;
  assign n21860 = n20966 ^ n20382;
  assign n21861 = n21860 ^ n21495;
  assign n21862 = n21861 ^ n21468;
  assign n21863 = n21859 & ~n21862;
  assign n21864 = n21863 ^ n21861;
  assign n21865 = n21864 ^ n21466;
  assign n21866 = ~n21467 & ~n21865;
  assign n21867 = n21866 ^ n21465;
  assign n21869 = n21868 ^ n21867;
  assign n21900 = n21871 ^ n21869;
  assign n21901 = n21900 ^ n19822;
  assign n21902 = n21864 ^ n21467;
  assign n21903 = n21902 ^ n19815;
  assign n21904 = n21861 ^ n21859;
  assign n21905 = n21904 ^ n19805;
  assign n21906 = n21855 ^ n21473;
  assign n21907 = n21906 ^ n19754;
  assign n21908 = n21852 ^ n21478;
  assign n21909 = n21908 ^ n19568;
  assign n21910 = n21849 ^ n21847;
  assign n21911 = n21910 ^ n19447;
  assign n21912 = n21842 ^ n21483;
  assign n21913 = n21912 ^ n18998;
  assign n21914 = n21839 ^ n21837;
  assign n21915 = n21914 ^ n19000;
  assign n21916 = n21832 ^ n21487;
  assign n21917 = n21916 ^ n19004;
  assign n21918 = n21829 ^ n21827;
  assign n21919 = n21918 ^ n19006;
  assign n21920 = n21822 ^ n21491;
  assign n21921 = n21920 ^ n19008;
  assign n21922 = n21819 ^ n21817;
  assign n21923 = n21922 ^ n19013;
  assign n21924 = n21813 ^ n21811;
  assign n21925 = n21924 ^ n19018;
  assign n21926 = n21806 ^ n21804;
  assign n21927 = n21926 ^ n19023;
  assign n21928 = n21800 ^ n21798;
  assign n21929 = n21928 ^ n19029;
  assign n21930 = n21793 ^ n21791;
  assign n21931 = n21930 ^ n19034;
  assign n21932 = n21787 ^ n21785;
  assign n21933 = n21932 ^ n19035;
  assign n21934 = n21781 ^ n21779;
  assign n21935 = n21934 ^ n19040;
  assign n21936 = n21775 ^ n21773;
  assign n21937 = n21936 ^ n19041;
  assign n21938 = n21764 ^ n21762;
  assign n21939 = n19050 & ~n21938;
  assign n21940 = n21939 ^ n19047;
  assign n21941 = n21769 ^ n21768;
  assign n21942 = n21941 ^ n21939;
  assign n21943 = n21940 & ~n21942;
  assign n21944 = n21943 ^ n19047;
  assign n21945 = n21944 ^ n21936;
  assign n21946 = n21937 & n21945;
  assign n21947 = n21946 ^ n19041;
  assign n21948 = n21947 ^ n21934;
  assign n21949 = n21935 & ~n21948;
  assign n21950 = n21949 ^ n19040;
  assign n21951 = n21950 ^ n21932;
  assign n21952 = ~n21933 & ~n21951;
  assign n21953 = n21952 ^ n19035;
  assign n21954 = n21953 ^ n21930;
  assign n21955 = n21931 & ~n21954;
  assign n21956 = n21955 ^ n19034;
  assign n21957 = n21956 ^ n21928;
  assign n21958 = ~n21929 & n21957;
  assign n21959 = n21958 ^ n19029;
  assign n21960 = n21959 ^ n21926;
  assign n21961 = ~n21927 & n21960;
  assign n21962 = n21961 ^ n19023;
  assign n21963 = n21962 ^ n21924;
  assign n21964 = n21925 & ~n21963;
  assign n21965 = n21964 ^ n19018;
  assign n21966 = n21965 ^ n21922;
  assign n21967 = ~n21923 & n21966;
  assign n21968 = n21967 ^ n19013;
  assign n21969 = n21968 ^ n21920;
  assign n21970 = n21921 & ~n21969;
  assign n21971 = n21970 ^ n19008;
  assign n21972 = n21971 ^ n21918;
  assign n21973 = ~n21919 & ~n21972;
  assign n21974 = n21973 ^ n19006;
  assign n21975 = n21974 ^ n21916;
  assign n21976 = ~n21917 & ~n21975;
  assign n21977 = n21976 ^ n19004;
  assign n21978 = n21977 ^ n21914;
  assign n21979 = n21915 & n21978;
  assign n21980 = n21979 ^ n19000;
  assign n21981 = n21980 ^ n21912;
  assign n21982 = ~n21913 & ~n21981;
  assign n21983 = n21982 ^ n18998;
  assign n21984 = n21983 ^ n21910;
  assign n21985 = ~n21911 & ~n21984;
  assign n21986 = n21985 ^ n19447;
  assign n21987 = n21986 ^ n21908;
  assign n21988 = ~n21909 & n21987;
  assign n21989 = n21988 ^ n19568;
  assign n21990 = n21989 ^ n21906;
  assign n21991 = ~n21907 & ~n21990;
  assign n21992 = n21991 ^ n19754;
  assign n21993 = n21992 ^ n21904;
  assign n21994 = ~n21905 & ~n21993;
  assign n21995 = n21994 ^ n19805;
  assign n21996 = n21995 ^ n21902;
  assign n21997 = n21903 & n21996;
  assign n21998 = n21997 ^ n19815;
  assign n21999 = n21998 ^ n21900;
  assign n22000 = ~n21901 & ~n21999;
  assign n22001 = n22000 ^ n19822;
  assign n21872 = n21871 ^ n21868;
  assign n21873 = ~n21869 & n21872;
  assign n21874 = n21873 ^ n21871;
  assign n21459 = n21002 ^ n20425;
  assign n21461 = n21460 ^ n21459;
  assign n21458 = n21436 ^ n21348;
  assign n21462 = n21461 ^ n21458;
  assign n21898 = n21874 ^ n21462;
  assign n21899 = n21898 ^ n19803;
  assign n22025 = n22001 ^ n21899;
  assign n22026 = n21998 ^ n21901;
  assign n22027 = n21995 ^ n21903;
  assign n22028 = n21986 ^ n21909;
  assign n22029 = n21965 ^ n21923;
  assign n22030 = n21959 ^ n21927;
  assign n22031 = n21956 ^ n21929;
  assign n22032 = n21953 ^ n21931;
  assign n22033 = n21947 ^ n21935;
  assign n22034 = n21941 ^ n21940;
  assign n22035 = n21938 ^ n19050;
  assign n22036 = n22034 & ~n22035;
  assign n22037 = n21944 ^ n21937;
  assign n22038 = n22036 & n22037;
  assign n22039 = ~n22033 & n22038;
  assign n22040 = n21950 ^ n21933;
  assign n22041 = n22039 & n22040;
  assign n22042 = ~n22032 & ~n22041;
  assign n22043 = ~n22031 & ~n22042;
  assign n22044 = n22030 & ~n22043;
  assign n22045 = n21962 ^ n21925;
  assign n22046 = n22044 & ~n22045;
  assign n22047 = n22029 & n22046;
  assign n22048 = n21968 ^ n21921;
  assign n22049 = ~n22047 & n22048;
  assign n22050 = n21971 ^ n21919;
  assign n22051 = ~n22049 & n22050;
  assign n22052 = n21974 ^ n21917;
  assign n22053 = ~n22051 & n22052;
  assign n22054 = n21977 ^ n21915;
  assign n22055 = ~n22053 & ~n22054;
  assign n22056 = n21980 ^ n21913;
  assign n22057 = n22055 & ~n22056;
  assign n22058 = n21983 ^ n21911;
  assign n22059 = n22057 & n22058;
  assign n22060 = ~n22028 & n22059;
  assign n22061 = n21989 ^ n21907;
  assign n22062 = ~n22060 & n22061;
  assign n22063 = n21992 ^ n21905;
  assign n22064 = n22062 & ~n22063;
  assign n22065 = n22027 & ~n22064;
  assign n22066 = n22026 & n22065;
  assign n22067 = ~n22025 & ~n22066;
  assign n22002 = n22001 ^ n21898;
  assign n22003 = n21899 & ~n22002;
  assign n22004 = n22003 ^ n19803;
  assign n21875 = n21874 ^ n21458;
  assign n21876 = ~n21462 & n21875;
  assign n21877 = n21876 ^ n21461;
  assign n21456 = n21455 ^ n21439;
  assign n20380 = n20379 ^ n19767;
  assign n20946 = n20945 ^ n20380;
  assign n21457 = n21456 ^ n20946;
  assign n21896 = n21877 ^ n21457;
  assign n21897 = n21896 ^ n19835;
  assign n22068 = n22004 ^ n21897;
  assign n22069 = ~n22067 & n22068;
  assign n22005 = n22004 ^ n21896;
  assign n22006 = n21897 & n22005;
  assign n22007 = n22006 ^ n19835;
  assign n21883 = n21064 ^ n20424;
  assign n21884 = n21883 ^ n21630;
  assign n21881 = n21710 ^ n21707;
  assign n21878 = n21877 ^ n21456;
  assign n21879 = n21457 & n21878;
  assign n21880 = n21879 ^ n20946;
  assign n21882 = n21881 ^ n21880;
  assign n21894 = n21884 ^ n21882;
  assign n21895 = n21894 ^ n19843;
  assign n22070 = n22007 ^ n21895;
  assign n22071 = n22069 & n22070;
  assign n22008 = n22007 ^ n21894;
  assign n22009 = ~n21895 & ~n22008;
  assign n22010 = n22009 ^ n19843;
  assign n21890 = n21714 ^ n2641;
  assign n21888 = n21076 ^ n20511;
  assign n21889 = n21888 ^ n21644;
  assign n21891 = n21890 ^ n21889;
  assign n21885 = n21884 ^ n21881;
  assign n21886 = n21882 & ~n21885;
  assign n21887 = n21886 ^ n21884;
  assign n21892 = n21891 ^ n21887;
  assign n21893 = n21892 ^ n19895;
  assign n22024 = n22010 ^ n21893;
  assign n22093 = n22071 ^ n22024;
  assign n22094 = n22093 ^ n1607;
  assign n22096 = n22068 ^ n22067;
  assign n22097 = n22096 ^ n1529;
  assign n22099 = n22065 ^ n22026;
  assign n2719 = n2664 ^ n1490;
  assign n2720 = n2719 ^ n2708;
  assign n2721 = n2720 ^ x492;
  assign n22100 = n22099 ^ n2721;
  assign n22102 = n22063 ^ n22062;
  assign n22103 = n22102 ^ n3197;
  assign n22104 = n22061 ^ n22060;
  assign n22105 = n22104 ^ n3041;
  assign n22106 = n22059 ^ n22028;
  assign n2433 = n2432 ^ n2414;
  assign n2437 = n2436 ^ n2433;
  assign n2438 = n2437 ^ x496;
  assign n22107 = n22106 ^ n2438;
  assign n22108 = n22058 ^ n22057;
  assign n1482 = n1434 ^ n1370;
  assign n1483 = n1482 ^ n1376;
  assign n1484 = n1483 ^ x497;
  assign n22109 = n22108 ^ n1484;
  assign n22111 = n22054 ^ n22053;
  assign n1173 = n1172 ^ n1085;
  assign n1177 = n1176 ^ n1173;
  assign n1178 = n1177 ^ x499;
  assign n22112 = n22111 ^ n1178;
  assign n22113 = n22052 ^ n22051;
  assign n1446 = n1334 ^ n1236;
  assign n1447 = n1446 ^ n1012;
  assign n1448 = n1447 ^ x500;
  assign n22114 = n22113 ^ n1448;
  assign n22115 = n22050 ^ n22049;
  assign n1003 = n999 ^ n924;
  assign n1007 = n1006 ^ n1003;
  assign n1008 = n1007 ^ x501;
  assign n22116 = n22115 ^ n1008;
  assign n22120 = n22043 ^ n22030;
  assign n22121 = n22120 ^ n769;
  assign n22122 = n22042 ^ n22031;
  assign n22123 = n22122 ^ n3266;
  assign n22125 = n22040 ^ n22039;
  assign n22129 = n22128 ^ n22125;
  assign n22131 = n20279 ^ n13562;
  assign n22132 = n22131 ^ n16898;
  assign n22133 = n22132 ^ x509;
  assign n22130 = n22038 ^ n22033;
  assign n22134 = n22133 ^ n22130;
  assign n22135 = n22037 ^ n22036;
  assign n691 = n690 ^ n672;
  assign n692 = n691 ^ n524;
  assign n693 = n692 ^ x510;
  assign n22136 = n22135 ^ n693;
  assign n22137 = n2210 & n22035;
  assign n22141 = n22140 ^ n22137;
  assign n22142 = n22035 ^ n22034;
  assign n22143 = n22142 ^ n22140;
  assign n22144 = n22141 & n22143;
  assign n22145 = n22144 ^ n22137;
  assign n22146 = n22145 ^ n22135;
  assign n22147 = n22136 & ~n22146;
  assign n22148 = n22147 ^ n693;
  assign n22149 = n22148 ^ n22130;
  assign n22150 = ~n22134 & n22149;
  assign n22151 = n22150 ^ n22133;
  assign n22152 = n22151 ^ n22125;
  assign n22153 = n22129 & ~n22152;
  assign n22154 = n22153 ^ n22128;
  assign n22124 = n22041 ^ n22032;
  assign n22155 = n22154 ^ n22124;
  assign n22159 = n22158 ^ n22124;
  assign n22160 = n22155 & ~n22159;
  assign n22161 = n22160 ^ n22158;
  assign n22162 = n22161 ^ n22122;
  assign n22163 = n22123 & ~n22162;
  assign n22164 = n22163 ^ n3266;
  assign n22165 = n22164 ^ n22120;
  assign n22166 = n22121 & ~n22165;
  assign n22167 = n22166 ^ n769;
  assign n22119 = n22045 ^ n22044;
  assign n22168 = n22167 ^ n22119;
  assign n22169 = n22119 ^ n779;
  assign n22170 = ~n22168 & n22169;
  assign n22171 = n22170 ^ n779;
  assign n22118 = n22046 ^ n22029;
  assign n22172 = n22171 ^ n22118;
  assign n866 = n856 ^ n802;
  assign n867 = n866 ^ n786;
  assign n868 = n867 ^ x503;
  assign n22173 = n22118 ^ n868;
  assign n22174 = n22172 & ~n22173;
  assign n22175 = n22174 ^ n868;
  assign n22117 = n22048 ^ n22047;
  assign n22176 = n22175 ^ n22117;
  assign n22177 = n22117 ^ n877;
  assign n22178 = n22176 & ~n22177;
  assign n22179 = n22178 ^ n877;
  assign n22180 = n22179 ^ n22115;
  assign n22181 = n22116 & ~n22180;
  assign n22182 = n22181 ^ n1008;
  assign n22183 = n22182 ^ n22113;
  assign n22184 = ~n22114 & n22183;
  assign n22185 = n22184 ^ n1448;
  assign n22186 = n22185 ^ n22111;
  assign n22187 = ~n22112 & n22186;
  assign n22188 = n22187 ^ n1178;
  assign n22110 = n22056 ^ n22055;
  assign n22189 = n22188 ^ n22110;
  assign n1464 = n1418 ^ n1352;
  assign n1465 = n1464 ^ n1458;
  assign n1466 = n1465 ^ x498;
  assign n22190 = n22110 ^ n1466;
  assign n22191 = ~n22189 & n22190;
  assign n22192 = n22191 ^ n1466;
  assign n22193 = n22192 ^ n22108;
  assign n22194 = ~n22109 & n22193;
  assign n22195 = n22194 ^ n1484;
  assign n22196 = n22195 ^ n22106;
  assign n22197 = n22107 & ~n22196;
  assign n22198 = n22197 ^ n2438;
  assign n22199 = n22198 ^ n22104;
  assign n22200 = ~n22105 & n22199;
  assign n22201 = n22200 ^ n3041;
  assign n22202 = n22201 ^ n22102;
  assign n22203 = ~n22103 & n22202;
  assign n22204 = n22203 ^ n3197;
  assign n22101 = n22064 ^ n22027;
  assign n22205 = n22204 ^ n22101;
  assign n22206 = n22101 ^ n2714;
  assign n22207 = ~n22205 & n22206;
  assign n22208 = n22207 ^ n2714;
  assign n22209 = n22208 ^ n22099;
  assign n22210 = ~n22100 & n22209;
  assign n22211 = n22210 ^ n2721;
  assign n22098 = n22066 ^ n22025;
  assign n22212 = n22211 ^ n22098;
  assign n22213 = n22098 ^ n2736;
  assign n22214 = ~n22212 & n22213;
  assign n22215 = n22214 ^ n2736;
  assign n22216 = n22215 ^ n22096;
  assign n22217 = n22097 & ~n22216;
  assign n22218 = n22217 ^ n1529;
  assign n22095 = n22070 ^ n22069;
  assign n22219 = n22218 ^ n22095;
  assign n22220 = n22095 ^ n2953;
  assign n22221 = n22219 & ~n22220;
  assign n22222 = n22221 ^ n2953;
  assign n22223 = n22222 ^ n22093;
  assign n22224 = n22094 & ~n22223;
  assign n22225 = n22224 ^ n1607;
  assign n22072 = ~n22024 & ~n22071;
  assign n22018 = n20561 ^ n19947;
  assign n22019 = n22018 ^ n21660;
  assign n22017 = n21717 ^ n21704;
  assign n22020 = n22019 ^ n22017;
  assign n22014 = n21890 ^ n21887;
  assign n22015 = n21891 & n22014;
  assign n22016 = n22015 ^ n21889;
  assign n22021 = n22020 ^ n22016;
  assign n22022 = n22021 ^ n19353;
  assign n22011 = n22010 ^ n21892;
  assign n22012 = n21893 & ~n22011;
  assign n22013 = n22012 ^ n19895;
  assign n22023 = n22022 ^ n22013;
  assign n22088 = n22072 ^ n22023;
  assign n22092 = n22091 ^ n22088;
  assign n22352 = n22225 ^ n22092;
  assign n23273 = n23272 ^ n22352;
  assign n22518 = n21495 ^ n20972;
  assign n22519 = n22518 ^ n21458;
  assign n22392 = n21471 ^ n20937;
  assign n22393 = n22392 ^ n21868;
  assign n22391 = n22176 ^ n877;
  assign n22394 = n22393 ^ n22391;
  assign n22507 = n22172 ^ n868;
  assign n22397 = n22168 ^ n779;
  assign n22395 = n21518 ^ n20656;
  assign n22396 = n22395 ^ n21468;
  assign n22398 = n22397 ^ n22396;
  assign n22399 = n21480 ^ n20384;
  assign n22400 = n22399 ^ n21469;
  assign n22331 = n22164 ^ n22121;
  assign n22401 = n22400 ^ n22331;
  assign n22402 = n21446 ^ n20388;
  assign n22403 = n22402 ^ n21846;
  assign n22340 = n22158 ^ n22155;
  assign n22404 = n22403 ^ n22340;
  assign n22407 = n22148 ^ n22134;
  assign n22405 = n21328 ^ n20396;
  assign n22406 = n22405 ^ n21836;
  assign n22408 = n22407 ^ n22406;
  assign n22476 = n22145 ^ n22136;
  assign n22411 = n22142 ^ n22141;
  assign n22409 = n21296 ^ n20624;
  assign n22410 = n22409 ^ n21826;
  assign n22412 = n22411 ^ n22410;
  assign n22414 = n21490 ^ n21282;
  assign n22415 = n22414 ^ n20401;
  assign n22413 = n22035 ^ n2210;
  assign n22416 = n22415 ^ n22413;
  assign n22457 = n20949 ^ n20405;
  assign n22458 = n22457 ^ n21810;
  assign n22262 = n20953 ^ n20412;
  assign n22263 = n22262 ^ n21797;
  assign n22082 = n20568 ^ n19952;
  assign n22083 = n22082 ^ n21678;
  assign n22078 = n22017 ^ n22016;
  assign n22079 = ~n22020 & n22078;
  assign n22080 = n22079 ^ n22019;
  assign n22077 = n21721 ^ n2747;
  assign n22081 = n22080 ^ n22077;
  assign n22084 = n22083 ^ n22081;
  assign n22085 = n22084 ^ n19349;
  assign n22074 = n22021 ^ n22013;
  assign n22075 = n22022 & ~n22074;
  assign n22076 = n22075 ^ n19353;
  assign n22246 = n22084 ^ n22076;
  assign n22247 = ~n22085 & n22246;
  assign n22248 = n22247 ^ n19349;
  assign n22242 = n20560 ^ n19943;
  assign n22243 = n22242 ^ n21142;
  assign n22238 = n22083 ^ n22077;
  assign n22239 = n22081 & n22238;
  assign n22240 = n22239 ^ n22083;
  assign n22237 = n21724 ^ n21701;
  assign n22241 = n22240 ^ n22237;
  assign n22244 = n22243 ^ n22241;
  assign n22245 = n22244 ^ n19347;
  assign n22249 = n22248 ^ n22245;
  assign n22073 = n22023 & ~n22072;
  assign n22086 = n22085 ^ n22076;
  assign n22236 = n22073 & ~n22086;
  assign n22250 = n22249 ^ n22236;
  assign n22251 = n22250 ^ n1919;
  assign n22226 = n22225 ^ n22088;
  assign n22227 = n22092 & ~n22226;
  assign n22228 = n22227 ^ n22091;
  assign n22087 = n22086 ^ n22073;
  assign n22229 = n22228 ^ n22087;
  assign n22233 = n22232 ^ n22087;
  assign n22234 = ~n22229 & n22233;
  assign n22235 = n22234 ^ n22232;
  assign n22252 = n22251 ^ n22235;
  assign n22253 = n20955 ^ n20414;
  assign n22254 = n22253 ^ n21494;
  assign n22261 = ~n22252 & n22254;
  assign n22264 = n22263 ^ n22261;
  assign n22280 = n22250 ^ n22235;
  assign n22281 = ~n22251 & n22280;
  assign n22282 = n22281 ^ n1919;
  assign n22275 = n22248 ^ n22244;
  assign n22276 = n22245 & ~n22275;
  assign n22277 = n22276 ^ n19347;
  assign n22271 = n20559 ^ n19940;
  assign n22272 = n22271 ^ n21147;
  assign n22267 = n22243 ^ n22237;
  assign n22268 = ~n22241 & n22267;
  assign n22269 = n22268 ^ n22243;
  assign n22266 = n21728 ^ n2876;
  assign n22270 = n22269 ^ n22266;
  assign n22273 = n22272 ^ n22270;
  assign n22274 = n22273 ^ n19346;
  assign n22278 = n22277 ^ n22274;
  assign n22265 = n22236 & n22249;
  assign n22279 = n22278 ^ n22265;
  assign n22283 = n22282 ^ n22279;
  assign n22284 = n22283 ^ n1912;
  assign n22317 = n22284 ^ n22263;
  assign n22318 = ~n22264 & ~n22317;
  assign n22319 = n22318 ^ n22261;
  assign n22313 = n22279 ^ n1912;
  assign n22314 = n22283 & ~n22313;
  assign n22315 = n22314 ^ n1912;
  assign n22307 = n22277 ^ n22273;
  assign n22308 = ~n22274 & n22307;
  assign n22309 = n22308 ^ n19346;
  assign n22303 = n20557 ^ n19938;
  assign n22304 = n22303 ^ n21139;
  assign n22299 = n22272 ^ n22266;
  assign n22300 = n22270 & ~n22299;
  assign n22301 = n22300 ^ n22272;
  assign n22298 = n21731 ^ n21698;
  assign n22302 = n22301 ^ n22298;
  assign n22305 = n22304 ^ n22302;
  assign n22306 = n22305 ^ n19345;
  assign n22310 = n22309 ^ n22306;
  assign n22297 = ~n22265 & n22278;
  assign n22311 = n22310 ^ n22297;
  assign n22312 = n22311 ^ n1938;
  assign n22316 = n22315 ^ n22312;
  assign n22320 = n22319 ^ n22316;
  assign n22295 = n20950 ^ n20409;
  assign n22296 = n22295 ^ n21493;
  assign n22454 = n22316 ^ n22296;
  assign n22455 = n22320 & ~n22454;
  assign n22456 = n22455 ^ n22296;
  assign n22459 = n22458 ^ n22456;
  assign n22437 = n22315 ^ n22311;
  assign n22438 = ~n22312 & n22437;
  assign n22439 = n22438 ^ n1938;
  assign n22431 = ~n22297 & ~n22310;
  assign n22426 = n22309 ^ n22305;
  assign n22427 = ~n22306 & ~n22426;
  assign n22428 = n22427 ^ n19345;
  assign n22429 = n22428 ^ n19378;
  assign n22421 = n22304 ^ n22298;
  assign n22422 = ~n22302 & n22421;
  assign n22423 = n22422 ^ n22304;
  assign n22369 = n21734 ^ n21693;
  assign n22424 = n22423 ^ n22369;
  assign n22419 = n20419 ^ n19968;
  assign n22420 = n22419 ^ n21160;
  assign n22425 = n22424 ^ n22420;
  assign n22430 = n22429 ^ n22425;
  assign n22436 = n22431 ^ n22430;
  assign n22440 = n22439 ^ n22436;
  assign n22460 = n22440 ^ n2057;
  assign n22461 = n22460 ^ n22456;
  assign n22462 = ~n22459 & n22461;
  assign n22463 = n22462 ^ n22458;
  assign n22450 = n22420 ^ n22369;
  assign n22451 = n22424 & ~n22450;
  assign n22452 = n22451 ^ n22420;
  assign n22445 = n22425 ^ n19378;
  assign n22446 = n22428 ^ n22425;
  assign n22447 = ~n22445 & ~n22446;
  assign n22448 = n22447 ^ n19378;
  assign n22441 = n22436 ^ n2057;
  assign n22442 = n22440 & ~n22441;
  assign n22443 = n22442 ^ n2057;
  assign n22432 = n22430 & n22431;
  assign n22364 = n21738 ^ n1710;
  assign n22433 = n22432 ^ n22364;
  assign n22417 = n21672 ^ n20417;
  assign n22418 = n22417 ^ n21138;
  assign n22434 = n22433 ^ n22418;
  assign n22435 = n22434 ^ n2220;
  assign n22444 = n22443 ^ n22435;
  assign n22449 = n22448 ^ n22444;
  assign n22453 = n22452 ^ n22449;
  assign n22464 = n22463 ^ n22453;
  assign n22465 = n21247 ^ n20614;
  assign n22466 = n22465 ^ n21492;
  assign n22467 = n22466 ^ n22453;
  assign n22468 = ~n22464 & ~n22467;
  assign n22469 = n22468 ^ n22466;
  assign n22470 = n22469 ^ n22413;
  assign n22471 = ~n22416 & ~n22470;
  assign n22472 = n22471 ^ n22415;
  assign n22473 = n22472 ^ n22411;
  assign n22474 = n22412 & ~n22473;
  assign n22475 = n22474 ^ n22410;
  assign n22477 = n22476 ^ n22475;
  assign n22478 = n21311 ^ n20399;
  assign n22479 = n22478 ^ n21486;
  assign n22480 = n22479 ^ n22476;
  assign n22481 = n22477 & ~n22480;
  assign n22482 = n22481 ^ n22479;
  assign n22483 = n22482 ^ n22407;
  assign n22484 = n22408 & ~n22483;
  assign n22485 = n22484 ^ n22406;
  assign n22345 = n22151 ^ n22129;
  assign n22486 = n22485 ^ n22345;
  assign n22487 = n21482 ^ n21342;
  assign n22488 = n22487 ^ n20392;
  assign n22489 = n22488 ^ n22345;
  assign n22490 = n22486 & ~n22489;
  assign n22491 = n22490 ^ n22488;
  assign n22492 = n22491 ^ n22340;
  assign n22493 = ~n22404 & ~n22492;
  assign n22494 = n22493 ^ n22403;
  assign n22335 = n22161 ^ n22123;
  assign n22495 = n22494 ^ n22335;
  assign n22496 = n21505 ^ n20646;
  assign n22497 = n22496 ^ n21477;
  assign n22498 = n22497 ^ n22335;
  assign n22499 = ~n22495 & n22498;
  assign n22500 = n22499 ^ n22497;
  assign n22501 = n22500 ^ n22400;
  assign n22502 = ~n22401 & n22501;
  assign n22503 = n22502 ^ n22331;
  assign n22504 = n22503 ^ n22397;
  assign n22505 = ~n22398 & ~n22504;
  assign n22506 = n22505 ^ n22396;
  assign n22508 = n22507 ^ n22506;
  assign n22509 = n21475 ^ n20765;
  assign n22510 = n22509 ^ n21466;
  assign n22511 = n22510 ^ n22507;
  assign n22512 = ~n22508 & ~n22511;
  assign n22513 = n22512 ^ n22510;
  assign n22514 = n22513 ^ n22391;
  assign n22515 = ~n22394 & n22514;
  assign n22516 = n22515 ^ n22393;
  assign n22390 = n22179 ^ n22116;
  assign n22517 = n22516 ^ n22390;
  assign n22610 = n22519 ^ n22517;
  assign n22611 = n22610 ^ n20230;
  assign n22612 = n22513 ^ n22394;
  assign n22613 = n22612 ^ n20171;
  assign n22614 = n22510 ^ n22508;
  assign n22615 = n22614 ^ n20055;
  assign n22617 = n22497 ^ n22495;
  assign n22618 = n22617 ^ n19774;
  assign n22619 = n22491 ^ n22404;
  assign n22620 = n22619 ^ n19775;
  assign n22621 = n22488 ^ n22486;
  assign n22622 = n22621 ^ n20029;
  assign n22623 = n22482 ^ n22408;
  assign n22624 = n22623 ^ n19779;
  assign n22625 = n22479 ^ n22477;
  assign n22626 = n22625 ^ n19781;
  assign n22627 = n22472 ^ n22412;
  assign n22628 = n22627 ^ n19783;
  assign n22629 = n22469 ^ n22416;
  assign n22630 = n22629 ^ n19784;
  assign n22631 = n22466 ^ n22464;
  assign n22632 = n22631 ^ n19785;
  assign n22633 = n22460 ^ n22458;
  assign n22634 = n22633 ^ n22456;
  assign n22635 = n22634 ^ n19786;
  assign n22321 = n22320 ^ n22296;
  assign n22322 = n22321 ^ n19787;
  assign n22255 = n22254 ^ n22252;
  assign n22259 = ~n19794 & ~n22255;
  assign n22260 = n22259 ^ n19791;
  assign n22285 = n22284 ^ n22264;
  assign n22292 = n22285 ^ n22259;
  assign n22293 = n22260 & ~n22292;
  assign n22294 = n22293 ^ n19791;
  assign n22636 = n22321 ^ n22294;
  assign n22637 = n22322 & n22636;
  assign n22638 = n22637 ^ n19787;
  assign n22639 = n22638 ^ n22634;
  assign n22640 = ~n22635 & n22639;
  assign n22641 = n22640 ^ n19786;
  assign n22642 = n22641 ^ n22631;
  assign n22643 = ~n22632 & n22642;
  assign n22644 = n22643 ^ n19785;
  assign n22645 = n22644 ^ n22629;
  assign n22646 = ~n22630 & ~n22645;
  assign n22647 = n22646 ^ n19784;
  assign n22648 = n22647 ^ n22627;
  assign n22649 = ~n22628 & n22648;
  assign n22650 = n22649 ^ n19783;
  assign n22651 = n22650 ^ n22625;
  assign n22652 = n22626 & ~n22651;
  assign n22653 = n22652 ^ n19781;
  assign n22654 = n22653 ^ n22623;
  assign n22655 = ~n22624 & n22654;
  assign n22656 = n22655 ^ n19779;
  assign n22657 = n22656 ^ n22621;
  assign n22658 = n22622 & ~n22657;
  assign n22659 = n22658 ^ n20029;
  assign n22660 = n22659 ^ n22619;
  assign n22661 = ~n22620 & ~n22660;
  assign n22662 = n22661 ^ n19775;
  assign n22663 = n22662 ^ n22617;
  assign n22664 = ~n22618 & n22663;
  assign n22665 = n22664 ^ n19774;
  assign n22666 = n22665 ^ n19769;
  assign n22667 = n22500 ^ n22401;
  assign n22668 = n22667 ^ n22665;
  assign n22669 = ~n22666 & ~n22668;
  assign n22670 = n22669 ^ n19769;
  assign n22616 = n22503 ^ n22398;
  assign n22671 = n22670 ^ n22616;
  assign n22672 = n22616 ^ n20048;
  assign n22673 = n22671 & n22672;
  assign n22674 = n22673 ^ n20048;
  assign n22675 = n22674 ^ n22614;
  assign n22676 = n22615 & n22675;
  assign n22677 = n22676 ^ n20055;
  assign n22678 = n22677 ^ n22612;
  assign n22679 = ~n22613 & n22678;
  assign n22680 = n22679 ^ n20171;
  assign n22681 = n22680 ^ n22610;
  assign n22682 = n22611 & ~n22681;
  assign n22683 = n22682 ^ n20230;
  assign n22520 = n22519 ^ n22390;
  assign n22521 = ~n22517 & n22520;
  assign n22522 = n22521 ^ n22519;
  assign n22388 = n22182 ^ n22114;
  assign n22386 = n21464 ^ n20970;
  assign n22387 = n22386 ^ n21456;
  assign n22389 = n22388 ^ n22387;
  assign n22609 = n22522 ^ n22389;
  assign n22684 = n22683 ^ n22609;
  assign n22768 = n22684 ^ n20363;
  assign n22738 = n22680 ^ n22611;
  assign n22739 = n22674 ^ n22615;
  assign n22740 = n22671 ^ n20048;
  assign n22741 = n22647 ^ n22628;
  assign n22742 = n22644 ^ n22630;
  assign n22256 = n22255 ^ n19794;
  assign n22286 = n22285 ^ n22260;
  assign n22291 = n22256 & n22286;
  assign n22323 = n22322 ^ n22294;
  assign n22743 = n22291 & n22323;
  assign n22744 = n22638 ^ n22635;
  assign n22745 = n22743 & n22744;
  assign n22746 = n22641 ^ n22632;
  assign n22747 = n22745 & n22746;
  assign n22748 = ~n22742 & ~n22747;
  assign n22749 = ~n22741 & ~n22748;
  assign n22750 = n22650 ^ n22626;
  assign n22751 = ~n22749 & ~n22750;
  assign n22752 = n22653 ^ n22624;
  assign n22753 = n22751 & n22752;
  assign n22754 = n22656 ^ n22622;
  assign n22755 = n22753 & ~n22754;
  assign n22756 = n22659 ^ n22620;
  assign n22757 = ~n22755 & ~n22756;
  assign n22758 = n22662 ^ n22618;
  assign n22759 = ~n22757 & ~n22758;
  assign n22760 = n22667 ^ n19769;
  assign n22761 = n22760 ^ n22665;
  assign n22762 = ~n22759 & n22761;
  assign n22763 = ~n22740 & ~n22762;
  assign n22764 = n22739 & n22763;
  assign n22765 = n22677 ^ n22613;
  assign n22766 = n22764 & n22765;
  assign n22767 = ~n22738 & n22766;
  assign n22816 = n22768 ^ n22767;
  assign n2454 = n2452 ^ n1550;
  assign n2461 = n2460 ^ n2454;
  assign n2465 = n2464 ^ n2461;
  assign n22817 = n22816 ^ n2465;
  assign n22818 = n22766 ^ n22738;
  assign n2474 = n2470 ^ n2443;
  assign n2481 = n2480 ^ n2474;
  assign n2482 = n2481 ^ n2458;
  assign n22819 = n22818 ^ n2482;
  assign n22824 = n22756 ^ n22755;
  assign n22825 = n22824 ^ n974;
  assign n22826 = n22754 ^ n22753;
  assign n22827 = n22826 ^ n962;
  assign n22828 = n22752 ^ n22751;
  assign n22829 = n22828 ^ n3310;
  assign n22830 = n22750 ^ n22749;
  assign n22834 = n22833 ^ n22830;
  assign n22837 = n22746 ^ n22745;
  assign n537 = n536 ^ n515;
  assign n544 = n543 ^ n537;
  assign n548 = n547 ^ n544;
  assign n22838 = n22837 ^ n548;
  assign n22839 = n22744 ^ n22743;
  assign n22843 = n22842 ^ n22839;
  assign n22325 = n20856 ^ n528;
  assign n22326 = n22325 ^ n17660;
  assign n22327 = n22326 ^ n3242;
  assign n22324 = n22323 ^ n22291;
  assign n22328 = n22327 ^ n22324;
  assign n2338 = n2308 ^ n2236;
  assign n2339 = n2338 ^ n2201;
  assign n2343 = n2342 ^ n2339;
  assign n22257 = n2343 & ~n22256;
  assign n22258 = n22257 ^ n2359;
  assign n22287 = n22286 ^ n22256;
  assign n22288 = n22287 ^ n2359;
  assign n22289 = n22258 & ~n22288;
  assign n22290 = n22289 ^ n22257;
  assign n22844 = n22324 ^ n22290;
  assign n22845 = n22328 & ~n22844;
  assign n22846 = n22845 ^ n22327;
  assign n22847 = n22846 ^ n22839;
  assign n22848 = n22843 & ~n22847;
  assign n22849 = n22848 ^ n22842;
  assign n22850 = n22849 ^ n22837;
  assign n22851 = n22838 & ~n22850;
  assign n22852 = n22851 ^ n548;
  assign n22836 = n22747 ^ n22742;
  assign n22853 = n22852 ^ n22836;
  assign n22854 = n20845 ^ n14276;
  assign n22855 = n22854 ^ n641;
  assign n22856 = n22855 ^ n567;
  assign n22857 = n22856 ^ n22836;
  assign n22858 = n22853 & ~n22857;
  assign n22859 = n22858 ^ n22856;
  assign n22835 = n22748 ^ n22741;
  assign n22860 = n22859 ^ n22835;
  assign n22861 = n22835 ^ n720;
  assign n22862 = ~n22860 & n22861;
  assign n22863 = n22862 ^ n720;
  assign n22864 = n22863 ^ n22830;
  assign n22865 = ~n22834 & n22864;
  assign n22866 = n22865 ^ n22833;
  assign n22867 = n22866 ^ n22828;
  assign n22868 = ~n22829 & n22867;
  assign n22869 = n22868 ^ n3310;
  assign n22870 = n22869 ^ n22826;
  assign n22871 = n22827 & ~n22870;
  assign n22872 = n22871 ^ n962;
  assign n22873 = n22872 ^ n22824;
  assign n22874 = n22825 & ~n22873;
  assign n22875 = n22874 ^ n974;
  assign n22876 = n22875 ^ n993;
  assign n22877 = n22758 ^ n22757;
  assign n22878 = n22877 ^ n22875;
  assign n22879 = n22876 & n22878;
  assign n22880 = n22879 ^ n993;
  assign n22823 = n22761 ^ n22759;
  assign n22881 = n22880 ^ n22823;
  assign n1110 = n1094 ^ n1025;
  assign n1111 = n1110 ^ n1106;
  assign n1115 = n1114 ^ n1111;
  assign n22882 = n22880 ^ n1115;
  assign n22883 = n22881 & n22882;
  assign n22884 = n22883 ^ n1115;
  assign n22822 = n22762 ^ n22740;
  assign n22885 = n22884 ^ n22822;
  assign n1283 = n1273 ^ n1183;
  assign n1284 = n1283 ^ n1122;
  assign n1288 = n1287 ^ n1284;
  assign n22886 = n22822 ^ n1288;
  assign n22887 = n22885 & ~n22886;
  assign n22888 = n22887 ^ n1288;
  assign n22821 = n22763 ^ n22739;
  assign n22889 = n22888 ^ n22821;
  assign n22890 = n22821 ^ n1300;
  assign n22891 = n22889 & ~n22890;
  assign n22892 = n22891 ^ n1300;
  assign n22820 = n22765 ^ n22764;
  assign n22893 = n22892 ^ n22820;
  assign n3139 = n2423 ^ n1383;
  assign n3143 = n3142 ^ n3139;
  assign n3144 = n3143 ^ n2477;
  assign n22894 = n22820 ^ n3144;
  assign n22895 = n22893 & ~n22894;
  assign n22896 = n22895 ^ n3144;
  assign n22897 = n22896 ^ n22818;
  assign n22898 = n22819 & ~n22897;
  assign n22899 = n22898 ^ n2482;
  assign n22900 = n22899 ^ n22816;
  assign n22901 = n22817 & ~n22900;
  assign n22902 = n22901 ^ n2465;
  assign n22685 = n22609 ^ n20363;
  assign n22686 = ~n22684 & ~n22685;
  assign n22687 = n22686 ^ n20363;
  assign n22527 = n21543 ^ n20966;
  assign n22528 = n22527 ^ n21881;
  assign n22523 = n22522 ^ n22387;
  assign n22524 = n22389 & n22523;
  assign n22525 = n22524 ^ n22388;
  assign n22385 = n22185 ^ n22112;
  assign n22526 = n22525 ^ n22385;
  assign n22607 = n22528 ^ n22526;
  assign n22608 = n22607 ^ n20382;
  assign n22770 = n22687 ^ n22608;
  assign n22769 = ~n22767 & ~n22768;
  assign n22815 = n22770 ^ n22769;
  assign n22903 = n22902 ^ n22815;
  assign n2539 = n2535 ^ n2502;
  assign n2543 = n2542 ^ n2539;
  assign n2544 = n2543 ^ n1515;
  assign n22904 = n22902 ^ n2544;
  assign n22905 = n22903 & n22904;
  assign n22906 = n22905 ^ n2544;
  assign n22907 = n22906 ^ n3074;
  assign n22771 = n22769 & ~n22770;
  assign n22688 = n22687 ^ n22607;
  assign n22689 = n22608 & n22688;
  assign n22690 = n22689 ^ n20382;
  assign n22534 = n21460 ^ n20988;
  assign n22535 = n22534 ^ n21890;
  assign n22532 = n22189 ^ n1466;
  assign n22529 = n22528 ^ n22385;
  assign n22530 = ~n22526 & ~n22529;
  assign n22531 = n22530 ^ n22528;
  assign n22533 = n22532 ^ n22531;
  assign n22605 = n22535 ^ n22533;
  assign n22606 = n22605 ^ n20427;
  assign n22737 = n22690 ^ n22606;
  assign n22908 = n22771 ^ n22737;
  assign n22909 = n22908 ^ n3074;
  assign n22910 = n22907 & n22909;
  assign n22911 = n22910 ^ n22906;
  assign n23269 = n22911 ^ n2636;
  assign n22772 = ~n22737 & ~n22771;
  assign n22691 = n22690 ^ n22605;
  assign n22692 = n22606 & ~n22691;
  assign n22693 = n22692 ^ n20427;
  assign n22536 = n22535 ^ n22532;
  assign n22537 = ~n22533 & n22536;
  assign n22538 = n22537 ^ n22535;
  assign n22383 = n22192 ^ n22109;
  assign n22381 = n20995 ^ n20945;
  assign n22382 = n22381 ^ n22017;
  assign n22384 = n22383 ^ n22382;
  assign n22603 = n22538 ^ n22384;
  assign n22604 = n22603 ^ n20426;
  assign n22736 = n22693 ^ n22604;
  assign n22814 = n22772 ^ n22736;
  assign n23270 = n23269 ^ n22814;
  assign n23171 = n22908 ^ n22907;
  assign n23169 = n22364 ^ n21678;
  assign n22354 = n22222 ^ n22094;
  assign n23170 = n23169 ^ n22354;
  assign n23172 = n23171 ^ n23170;
  assign n23259 = n22903 ^ n2544;
  assign n23175 = n22899 ^ n22817;
  assign n23173 = n22298 ^ n21644;
  assign n22361 = n22215 ^ n22097;
  assign n23174 = n23173 ^ n22361;
  assign n23176 = n23175 ^ n23174;
  assign n23179 = n22896 ^ n22819;
  assign n23177 = n22266 ^ n21630;
  assign n22366 = n22212 ^ n2736;
  assign n23178 = n23177 ^ n22366;
  assign n23180 = n23179 ^ n23178;
  assign n23183 = n22893 ^ n3144;
  assign n23181 = n22237 ^ n20945;
  assign n22371 = n22208 ^ n22100;
  assign n23182 = n23181 ^ n22371;
  assign n23184 = n23183 ^ n23182;
  assign n23188 = n22885 ^ n1288;
  assign n23186 = n22017 ^ n21543;
  assign n22379 = n22201 ^ n22103;
  assign n23187 = n23186 ^ n22379;
  assign n23189 = n23188 ^ n23187;
  assign n23192 = n22881 ^ n1115;
  assign n23190 = n21890 ^ n21464;
  assign n22549 = n22198 ^ n22105;
  assign n23191 = n23190 ^ n22549;
  assign n23193 = n23192 ^ n23191;
  assign n23195 = n21881 ^ n21495;
  assign n22542 = n22195 ^ n22107;
  assign n23196 = n23195 ^ n22542;
  assign n23194 = n22877 ^ n22876;
  assign n23197 = n23196 ^ n23194;
  assign n23198 = n21471 ^ n21456;
  assign n23199 = n23198 ^ n22383;
  assign n23146 = n22872 ^ n22825;
  assign n23200 = n23199 ^ n23146;
  assign n23202 = n21475 ^ n21458;
  assign n23203 = n23202 ^ n22532;
  assign n23201 = n22869 ^ n22827;
  assign n23204 = n23203 ^ n23201;
  assign n23208 = n22863 ^ n22834;
  assign n23206 = n21480 ^ n21466;
  assign n23207 = n23206 ^ n22388;
  assign n23209 = n23208 ^ n23207;
  assign n23043 = n22849 ^ n22838;
  assign n23041 = n21477 ^ n21342;
  assign n23042 = n23041 ^ n22507;
  assign n23044 = n23043 ^ n23042;
  assign n22990 = n22846 ^ n22843;
  assign n22988 = n21846 ^ n21328;
  assign n22989 = n22988 ^ n22397;
  assign n22991 = n22990 ^ n22989;
  assign n22330 = n21482 ^ n21311;
  assign n22332 = n22331 ^ n22330;
  assign n22329 = n22328 ^ n22290;
  assign n22333 = n22332 ^ n22329;
  assign n22337 = n22287 ^ n22258;
  assign n22334 = n21836 ^ n21296;
  assign n22336 = n22335 ^ n22334;
  assign n22338 = n22337 ^ n22336;
  assign n22342 = n22256 ^ n2343;
  assign n22339 = n21486 ^ n21282;
  assign n22341 = n22340 ^ n22339;
  assign n22343 = n22342 ^ n22341;
  assign n22363 = n21147 ^ n20568;
  assign n22365 = n22364 ^ n22363;
  assign n22367 = n22366 ^ n22365;
  assign n22368 = n21142 ^ n20561;
  assign n22370 = n22369 ^ n22368;
  assign n22372 = n22371 ^ n22370;
  assign n22375 = n22205 ^ n2714;
  assign n22373 = n21678 ^ n21076;
  assign n22374 = n22373 ^ n22298;
  assign n22376 = n22375 ^ n22374;
  assign n22377 = n21660 ^ n21064;
  assign n22378 = n22377 ^ n22266;
  assign n22380 = n22379 ^ n22378;
  assign n22539 = n22538 ^ n22383;
  assign n22540 = n22384 & n22539;
  assign n22541 = n22540 ^ n22382;
  assign n22543 = n22542 ^ n22541;
  assign n22544 = n21630 ^ n21002;
  assign n22545 = n22544 ^ n22077;
  assign n22546 = n22545 ^ n22542;
  assign n22547 = n22543 & ~n22546;
  assign n22548 = n22547 ^ n22545;
  assign n22550 = n22549 ^ n22548;
  assign n22551 = n21644 ^ n20379;
  assign n22552 = n22551 ^ n22237;
  assign n22553 = n22552 ^ n22549;
  assign n22554 = ~n22550 & n22553;
  assign n22555 = n22554 ^ n22552;
  assign n22556 = n22555 ^ n22378;
  assign n22557 = ~n22380 & n22556;
  assign n22558 = n22557 ^ n22379;
  assign n22559 = n22558 ^ n22375;
  assign n22560 = n22376 & n22559;
  assign n22561 = n22560 ^ n22374;
  assign n22562 = n22561 ^ n22371;
  assign n22563 = ~n22372 & n22562;
  assign n22564 = n22563 ^ n22370;
  assign n22565 = n22564 ^ n22366;
  assign n22566 = n22367 & ~n22565;
  assign n22567 = n22566 ^ n22365;
  assign n22359 = n21139 ^ n20560;
  assign n22360 = n22359 ^ n21762;
  assign n22362 = n22361 ^ n22360;
  assign n22590 = n22567 ^ n22362;
  assign n22591 = n22590 ^ n19943;
  assign n22592 = n22564 ^ n22367;
  assign n22593 = n22592 ^ n19952;
  assign n22594 = n22561 ^ n22372;
  assign n22595 = n22594 ^ n19947;
  assign n22596 = n22558 ^ n22376;
  assign n22597 = n22596 ^ n20511;
  assign n22598 = n22555 ^ n22380;
  assign n22599 = n22598 ^ n20424;
  assign n22600 = n22552 ^ n22550;
  assign n22601 = n22600 ^ n19767;
  assign n22694 = n22693 ^ n22603;
  assign n22695 = n22604 & ~n22694;
  assign n22696 = n22695 ^ n20426;
  assign n22602 = n22545 ^ n22543;
  assign n22697 = n22696 ^ n22602;
  assign n22698 = n22602 ^ n20425;
  assign n22699 = ~n22697 & ~n22698;
  assign n22700 = n22699 ^ n20425;
  assign n22701 = n22700 ^ n22600;
  assign n22702 = n22601 & ~n22701;
  assign n22703 = n22702 ^ n19767;
  assign n22704 = n22703 ^ n22598;
  assign n22705 = n22599 & n22704;
  assign n22706 = n22705 ^ n20424;
  assign n22707 = n22706 ^ n22596;
  assign n22708 = n22597 & n22707;
  assign n22709 = n22708 ^ n20511;
  assign n22710 = n22709 ^ n22594;
  assign n22711 = n22595 & ~n22710;
  assign n22712 = n22711 ^ n19947;
  assign n22713 = n22712 ^ n22592;
  assign n22714 = n22593 & n22713;
  assign n22715 = n22714 ^ n19952;
  assign n22716 = n22715 ^ n22590;
  assign n22717 = n22591 & n22716;
  assign n22718 = n22717 ^ n19943;
  assign n22568 = n22567 ^ n22360;
  assign n22569 = ~n22362 & n22568;
  assign n22570 = n22569 ^ n22361;
  assign n22357 = n22219 ^ n2953;
  assign n22355 = n21160 ^ n20559;
  assign n22356 = n22355 ^ n21769;
  assign n22358 = n22357 ^ n22356;
  assign n22589 = n22570 ^ n22358;
  assign n22719 = n22718 ^ n22589;
  assign n22720 = n22589 ^ n19940;
  assign n22721 = ~n22719 & ~n22720;
  assign n22722 = n22721 ^ n19940;
  assign n22575 = n21138 ^ n20557;
  assign n22576 = n22575 ^ n21761;
  assign n22571 = n22570 ^ n22357;
  assign n22572 = ~n22358 & n22571;
  assign n22573 = n22572 ^ n22356;
  assign n22574 = n22573 ^ n22354;
  assign n22587 = n22576 ^ n22574;
  assign n22588 = n22587 ^ n19938;
  assign n22732 = n22722 ^ n22588;
  assign n22733 = n22719 ^ n19940;
  assign n22734 = n22712 ^ n22593;
  assign n22735 = n22697 ^ n20425;
  assign n22773 = ~n22736 & n22772;
  assign n22774 = ~n22735 & ~n22773;
  assign n22775 = n22700 ^ n19767;
  assign n22776 = n22775 ^ n22600;
  assign n22777 = ~n22774 & n22776;
  assign n22778 = n22703 ^ n22599;
  assign n22779 = n22777 & n22778;
  assign n22780 = n22706 ^ n20511;
  assign n22781 = n22780 ^ n22596;
  assign n22782 = ~n22779 & n22781;
  assign n22783 = n22709 ^ n22595;
  assign n22784 = ~n22782 & n22783;
  assign n22785 = n22734 & n22784;
  assign n22786 = n22715 ^ n19943;
  assign n22787 = n22786 ^ n22590;
  assign n22788 = n22785 & ~n22787;
  assign n22789 = n22733 & ~n22788;
  assign n22790 = n22732 & ~n22789;
  assign n22723 = n22722 ^ n22587;
  assign n22724 = ~n22588 & ~n22723;
  assign n22725 = n22724 ^ n19938;
  assign n22577 = n22576 ^ n22354;
  assign n22578 = ~n22574 & n22577;
  assign n22579 = n22578 ^ n22576;
  assign n22350 = n20960 ^ n20419;
  assign n22351 = n22350 ^ n21760;
  assign n22353 = n22352 ^ n22351;
  assign n22585 = n22579 ^ n22353;
  assign n22586 = n22585 ^ n19968;
  assign n22731 = n22725 ^ n22586;
  assign n22793 = n22790 ^ n22731;
  assign n22794 = n22793 ^ n2165;
  assign n22795 = n22789 ^ n22732;
  assign n22796 = n22795 ^ n2178;
  assign n22798 = n22787 ^ n22785;
  assign n22802 = n22801 ^ n22798;
  assign n22803 = n22784 ^ n22734;
  assign n1724 = n1719 ^ n1665;
  assign n1728 = n1727 ^ n1724;
  assign n1729 = n1728 ^ n1701;
  assign n22804 = n22803 ^ n1729;
  assign n22805 = n22783 ^ n22782;
  assign n22806 = n22805 ^ n1654;
  assign n22807 = n22781 ^ n22779;
  assign n1631 = n1621 ^ n1508;
  assign n1638 = n1637 ^ n1631;
  assign n1642 = n1641 ^ n1638;
  assign n22808 = n22807 ^ n1642;
  assign n22809 = n22778 ^ n22777;
  assign n22810 = n22809 ^ n2927;
  assign n22811 = n22776 ^ n22774;
  assign n22812 = n22811 ^ n2902;
  assign n22912 = n22911 ^ n22814;
  assign n22913 = n22814 ^ n2636;
  assign n22914 = ~n22912 & n22913;
  assign n22915 = n22914 ^ n2636;
  assign n22813 = n22773 ^ n22735;
  assign n22916 = n22915 ^ n22813;
  assign n22917 = n22813 ^ n2908;
  assign n22918 = ~n22916 & n22917;
  assign n22919 = n22918 ^ n2908;
  assign n22920 = n22919 ^ n22811;
  assign n22921 = n22812 & ~n22920;
  assign n22922 = n22921 ^ n2902;
  assign n22923 = n22922 ^ n22809;
  assign n22924 = ~n22810 & n22923;
  assign n22925 = n22924 ^ n2927;
  assign n22926 = n22925 ^ n1642;
  assign n22927 = ~n22808 & ~n22926;
  assign n22928 = n22927 ^ n22807;
  assign n22929 = n22928 ^ n22805;
  assign n22930 = n22806 & n22929;
  assign n22931 = n22930 ^ n1654;
  assign n22932 = n22931 ^ n22803;
  assign n22933 = ~n22804 & n22932;
  assign n22934 = n22933 ^ n1729;
  assign n22935 = n22934 ^ n22798;
  assign n22936 = n22802 & ~n22935;
  assign n22937 = n22936 ^ n22801;
  assign n22797 = n22788 ^ n22733;
  assign n22938 = n22937 ^ n22797;
  assign n22939 = n22797 ^ n1817;
  assign n22940 = n22938 & ~n22939;
  assign n22941 = n22940 ^ n1817;
  assign n22942 = n22941 ^ n2178;
  assign n22943 = n22796 & ~n22942;
  assign n22944 = n22943 ^ n22795;
  assign n22945 = n22944 ^ n22793;
  assign n22946 = n22794 & ~n22945;
  assign n22947 = n22946 ^ n2165;
  assign n22791 = ~n22731 & n22790;
  assign n22726 = n22725 ^ n22585;
  assign n22727 = ~n22586 & n22726;
  assign n22728 = n22727 ^ n19968;
  assign n22729 = n22728 ^ n19795;
  assign n22580 = n22579 ^ n22352;
  assign n22581 = n22353 & ~n22580;
  assign n22582 = n22581 ^ n22351;
  assign n22348 = n20958 ^ n20417;
  assign n22349 = n22348 ^ n21759;
  assign n22583 = n22582 ^ n22349;
  assign n22347 = n22232 ^ n22229;
  assign n22584 = n22583 ^ n22347;
  assign n22730 = n22729 ^ n22584;
  assign n22792 = n22791 ^ n22730;
  assign n22948 = n22947 ^ n22792;
  assign n2189 = n2149 ^ n2098;
  assign n2190 = n2189 ^ n2169;
  assign n2191 = n2190 ^ n2129;
  assign n22949 = n22948 ^ n2191;
  assign n22344 = n21826 ^ n21247;
  assign n22346 = n22345 ^ n22344;
  assign n22950 = n22949 ^ n22346;
  assign n22952 = n21490 ^ n20949;
  assign n22953 = n22952 ^ n22407;
  assign n22951 = n22944 ^ n22794;
  assign n22954 = n22953 ^ n22951;
  assign n22957 = n22941 ^ n22796;
  assign n22955 = n21492 ^ n20950;
  assign n22956 = n22955 ^ n22476;
  assign n22958 = n22957 ^ n22956;
  assign n22963 = n21810 ^ n20953;
  assign n22964 = n22963 ^ n22411;
  assign n22959 = n21493 ^ n20955;
  assign n22960 = n22959 ^ n22413;
  assign n22961 = n22934 ^ n22802;
  assign n22962 = ~n22960 & n22961;
  assign n22965 = n22964 ^ n22962;
  assign n22966 = n22938 ^ n1817;
  assign n22967 = n22966 ^ n22964;
  assign n22968 = n22965 & n22967;
  assign n22969 = n22968 ^ n22962;
  assign n22970 = n22969 ^ n22957;
  assign n22971 = ~n22958 & ~n22970;
  assign n22972 = n22971 ^ n22956;
  assign n22973 = n22972 ^ n22953;
  assign n22974 = n22954 & n22973;
  assign n22975 = n22974 ^ n22951;
  assign n22976 = n22975 ^ n22949;
  assign n22977 = n22950 & n22976;
  assign n22978 = n22977 ^ n22346;
  assign n22979 = n22978 ^ n22342;
  assign n22980 = n22343 & ~n22979;
  assign n22981 = n22980 ^ n22341;
  assign n22982 = n22981 ^ n22337;
  assign n22983 = ~n22338 & n22982;
  assign n22984 = n22983 ^ n22336;
  assign n22985 = n22984 ^ n22329;
  assign n22986 = n22333 & n22985;
  assign n22987 = n22986 ^ n22332;
  assign n23038 = n22990 ^ n22987;
  assign n23039 = ~n22991 & ~n23038;
  assign n23040 = n23039 ^ n22989;
  assign n23131 = n23043 ^ n23040;
  assign n23132 = n23044 & n23131;
  assign n23133 = n23132 ^ n23042;
  assign n23130 = n22856 ^ n22853;
  assign n23134 = n23133 ^ n23130;
  assign n23128 = n21469 ^ n21446;
  assign n23129 = n23128 ^ n22391;
  assign n23211 = n23130 ^ n23129;
  assign n23212 = n23134 & n23211;
  assign n23213 = n23212 ^ n23129;
  assign n23210 = n22860 ^ n720;
  assign n23214 = n23213 ^ n23210;
  assign n23215 = n21505 ^ n21468;
  assign n23216 = n23215 ^ n22390;
  assign n23217 = n23216 ^ n23210;
  assign n23218 = n23214 & n23217;
  assign n23219 = n23218 ^ n23216;
  assign n23220 = n23219 ^ n23208;
  assign n23221 = n23209 & n23220;
  assign n23222 = n23221 ^ n23207;
  assign n23205 = n22866 ^ n22829;
  assign n23223 = n23222 ^ n23205;
  assign n23224 = n21868 ^ n21518;
  assign n23225 = n23224 ^ n22385;
  assign n23226 = n23225 ^ n23205;
  assign n23227 = ~n23223 & n23226;
  assign n23228 = n23227 ^ n23225;
  assign n23229 = n23228 ^ n23201;
  assign n23230 = n23204 & n23229;
  assign n23231 = n23230 ^ n23203;
  assign n23232 = n23231 ^ n23146;
  assign n23233 = ~n23200 & ~n23232;
  assign n23234 = n23233 ^ n23199;
  assign n23235 = n23234 ^ n23194;
  assign n23236 = ~n23197 & ~n23235;
  assign n23237 = n23236 ^ n23196;
  assign n23238 = n23237 ^ n23191;
  assign n23239 = ~n23193 & ~n23238;
  assign n23240 = n23239 ^ n23192;
  assign n23241 = n23240 ^ n23188;
  assign n23242 = n23189 & ~n23241;
  assign n23243 = n23242 ^ n23187;
  assign n23185 = n22889 ^ n1300;
  assign n23244 = n23243 ^ n23185;
  assign n23245 = n22077 ^ n21460;
  assign n23246 = n23245 ^ n22375;
  assign n23247 = n23246 ^ n23185;
  assign n23248 = ~n23244 & ~n23247;
  assign n23249 = n23248 ^ n23246;
  assign n23250 = n23249 ^ n23182;
  assign n23251 = n23184 & n23250;
  assign n23252 = n23251 ^ n23183;
  assign n23253 = n23252 ^ n23179;
  assign n23254 = n23180 & n23253;
  assign n23255 = n23254 ^ n23178;
  assign n23256 = n23255 ^ n23175;
  assign n23257 = n23176 & ~n23256;
  assign n23258 = n23257 ^ n23174;
  assign n23260 = n23259 ^ n23258;
  assign n23261 = n22369 ^ n21660;
  assign n23262 = n23261 ^ n22357;
  assign n23263 = n23262 ^ n23259;
  assign n23264 = n23260 & ~n23263;
  assign n23265 = n23264 ^ n23262;
  assign n23266 = n23265 ^ n23170;
  assign n23267 = n23172 & n23266;
  assign n23268 = n23267 ^ n23171;
  assign n23271 = n23270 ^ n23268;
  assign n23296 = n23273 ^ n23271;
  assign n23297 = n23296 ^ n20561;
  assign n23298 = n23265 ^ n23172;
  assign n23299 = n23298 ^ n21076;
  assign n23300 = n23262 ^ n23260;
  assign n23301 = n23300 ^ n21064;
  assign n23302 = n23255 ^ n23174;
  assign n23303 = n23302 ^ n23175;
  assign n23304 = n23303 ^ n20379;
  assign n23305 = n23252 ^ n23180;
  assign n23306 = n23305 ^ n21002;
  assign n23307 = n23249 ^ n23184;
  assign n23308 = n23307 ^ n20995;
  assign n23309 = n23246 ^ n23244;
  assign n23310 = n23309 ^ n20988;
  assign n23312 = n23237 ^ n23193;
  assign n23313 = n23312 ^ n20970;
  assign n23314 = n23234 ^ n23196;
  assign n23315 = n23314 ^ n23194;
  assign n23316 = n23315 ^ n20972;
  assign n23317 = n23231 ^ n23200;
  assign n23318 = n23317 ^ n20937;
  assign n23319 = n23228 ^ n23204;
  assign n23320 = n23319 ^ n20765;
  assign n23321 = n23225 ^ n23223;
  assign n23322 = n23321 ^ n20656;
  assign n23323 = n23219 ^ n23207;
  assign n23324 = n23323 ^ n23208;
  assign n23325 = n23324 ^ n20384;
  assign n23326 = n23216 ^ n23214;
  assign n23327 = n23326 ^ n20646;
  assign n23045 = n23044 ^ n23040;
  assign n23136 = n23045 ^ n20392;
  assign n22992 = n22991 ^ n22987;
  assign n22993 = n22992 ^ n20396;
  assign n22995 = n22981 ^ n22336;
  assign n22996 = n22995 ^ n22337;
  assign n22997 = n22996 ^ n20624;
  assign n22998 = n22978 ^ n22343;
  assign n22999 = n22998 ^ n20401;
  assign n23000 = n22975 ^ n22346;
  assign n23001 = n23000 ^ n22949;
  assign n23002 = n23001 ^ n20614;
  assign n23003 = n22961 ^ n22960;
  assign n23004 = ~n20414 & ~n23003;
  assign n23005 = n23004 ^ n20412;
  assign n23006 = n22966 ^ n22965;
  assign n23007 = n23006 ^ n23004;
  assign n23008 = n23005 & n23007;
  assign n23009 = n23008 ^ n20412;
  assign n23010 = n23009 ^ n20409;
  assign n23011 = n22969 ^ n22956;
  assign n23012 = n23011 ^ n22957;
  assign n23013 = n23012 ^ n23009;
  assign n23014 = n23010 & n23013;
  assign n23015 = n23014 ^ n20409;
  assign n23016 = n23015 ^ n20405;
  assign n23017 = n22972 ^ n22954;
  assign n23018 = n23017 ^ n23015;
  assign n23019 = ~n23016 & n23018;
  assign n23020 = n23019 ^ n20405;
  assign n23021 = n23020 ^ n23001;
  assign n23022 = n23002 & n23021;
  assign n23023 = n23022 ^ n20614;
  assign n23024 = n23023 ^ n22998;
  assign n23025 = n22999 & n23024;
  assign n23026 = n23025 ^ n20401;
  assign n23027 = n23026 ^ n22996;
  assign n23028 = ~n22997 & n23027;
  assign n23029 = n23028 ^ n20624;
  assign n22994 = n22984 ^ n22333;
  assign n23030 = n23029 ^ n22994;
  assign n23031 = n23029 ^ n20399;
  assign n23032 = ~n23030 & ~n23031;
  assign n23033 = n23032 ^ n20399;
  assign n23034 = n23033 ^ n22992;
  assign n23035 = n22993 & n23034;
  assign n23036 = n23035 ^ n20396;
  assign n23137 = n23045 ^ n23036;
  assign n23138 = n23136 & ~n23137;
  assign n23139 = n23138 ^ n20392;
  assign n23135 = n23134 ^ n23129;
  assign n23140 = n23139 ^ n23135;
  assign n23328 = n23135 ^ n20388;
  assign n23329 = n23140 & n23328;
  assign n23330 = n23329 ^ n20388;
  assign n23331 = n23330 ^ n23326;
  assign n23332 = n23327 & n23331;
  assign n23333 = n23332 ^ n20646;
  assign n23334 = n23333 ^ n23324;
  assign n23335 = n23325 & n23334;
  assign n23336 = n23335 ^ n20384;
  assign n23337 = n23336 ^ n23321;
  assign n23338 = n23322 & n23337;
  assign n23339 = n23338 ^ n20656;
  assign n23340 = n23339 ^ n23319;
  assign n23341 = ~n23320 & ~n23340;
  assign n23342 = n23341 ^ n20765;
  assign n23343 = n23342 ^ n23317;
  assign n23344 = n23318 & n23343;
  assign n23345 = n23344 ^ n20937;
  assign n23346 = n23345 ^ n23315;
  assign n23347 = ~n23316 & n23346;
  assign n23348 = n23347 ^ n20972;
  assign n23349 = n23348 ^ n23312;
  assign n23350 = n23313 & ~n23349;
  assign n23351 = n23350 ^ n20970;
  assign n23311 = n23240 ^ n23189;
  assign n23352 = n23351 ^ n23311;
  assign n23353 = n23311 ^ n20966;
  assign n23354 = ~n23352 & n23353;
  assign n23355 = n23354 ^ n20966;
  assign n23356 = n23355 ^ n23309;
  assign n23357 = ~n23310 & n23356;
  assign n23358 = n23357 ^ n20988;
  assign n23359 = n23358 ^ n23307;
  assign n23360 = ~n23308 & n23359;
  assign n23361 = n23360 ^ n20995;
  assign n23362 = n23361 ^ n23305;
  assign n23363 = ~n23306 & ~n23362;
  assign n23364 = n23363 ^ n21002;
  assign n23365 = n23364 ^ n23303;
  assign n23366 = ~n23304 & ~n23365;
  assign n23367 = n23366 ^ n20379;
  assign n23368 = n23367 ^ n23300;
  assign n23369 = n23301 & ~n23368;
  assign n23370 = n23369 ^ n21064;
  assign n23371 = n23370 ^ n23298;
  assign n23372 = n23299 & n23371;
  assign n23373 = n23372 ^ n21076;
  assign n23374 = n23373 ^ n23296;
  assign n23375 = ~n23297 & n23374;
  assign n23376 = n23375 ^ n20561;
  assign n23274 = n23273 ^ n23270;
  assign n23275 = n23271 & n23274;
  assign n23276 = n23275 ^ n23273;
  assign n23166 = n21769 ^ n21147;
  assign n23167 = n23166 ^ n22347;
  assign n23293 = n23276 ^ n23167;
  assign n23165 = n22916 ^ n2908;
  assign n23294 = n23293 ^ n23165;
  assign n23295 = n23294 ^ n20568;
  assign n23441 = n23376 ^ n23295;
  assign n23402 = n23373 ^ n20561;
  assign n23403 = n23402 ^ n23296;
  assign n23404 = n23370 ^ n21076;
  assign n23405 = n23404 ^ n23298;
  assign n23406 = n23330 ^ n23327;
  assign n23141 = n23140 ^ n20388;
  assign n23037 = n23036 ^ n20392;
  assign n23046 = n23045 ^ n23037;
  assign n23047 = n23033 ^ n22993;
  assign n23048 = n23030 ^ n20399;
  assign n23049 = n23026 ^ n22997;
  assign n23050 = n23023 ^ n20401;
  assign n23051 = n23050 ^ n22998;
  assign n23052 = n23003 ^ n20414;
  assign n23053 = n23006 ^ n23005;
  assign n23054 = n23052 & ~n23053;
  assign n23055 = n23012 ^ n20409;
  assign n23056 = n23055 ^ n23009;
  assign n23057 = n23054 & ~n23056;
  assign n23058 = n23017 ^ n20405;
  assign n23059 = n23058 ^ n23015;
  assign n23060 = n23057 & n23059;
  assign n23061 = n23020 ^ n23002;
  assign n23062 = n23060 & ~n23061;
  assign n23063 = ~n23051 & ~n23062;
  assign n23064 = n23049 & ~n23063;
  assign n23065 = ~n23048 & ~n23064;
  assign n23066 = ~n23047 & n23065;
  assign n23142 = n23046 & n23066;
  assign n23407 = ~n23141 & ~n23142;
  assign n23408 = ~n23406 & ~n23407;
  assign n23409 = n23333 ^ n20384;
  assign n23410 = n23409 ^ n23324;
  assign n23411 = ~n23408 & ~n23410;
  assign n23412 = n23336 ^ n20656;
  assign n23413 = n23412 ^ n23321;
  assign n23414 = ~n23411 & ~n23413;
  assign n23415 = n23339 ^ n23320;
  assign n23416 = n23414 & ~n23415;
  assign n23417 = n23342 ^ n23318;
  assign n23418 = n23416 & ~n23417;
  assign n23419 = n23345 ^ n23316;
  assign n23420 = n23418 & ~n23419;
  assign n23421 = n23348 ^ n20970;
  assign n23422 = n23421 ^ n23312;
  assign n23423 = ~n23420 & ~n23422;
  assign n23424 = n23352 ^ n20966;
  assign n23425 = n23423 & ~n23424;
  assign n23426 = n23355 ^ n20988;
  assign n23427 = n23426 ^ n23309;
  assign n23428 = ~n23425 & ~n23427;
  assign n23429 = n23358 ^ n20995;
  assign n23430 = n23429 ^ n23307;
  assign n23431 = n23428 & ~n23430;
  assign n23432 = n23361 ^ n23306;
  assign n23433 = ~n23431 & n23432;
  assign n23434 = n23364 ^ n20379;
  assign n23435 = n23434 ^ n23303;
  assign n23436 = ~n23433 & n23435;
  assign n23437 = n23367 ^ n23301;
  assign n23438 = n23436 & n23437;
  assign n23439 = ~n23405 & ~n23438;
  assign n23440 = n23403 & ~n23439;
  assign n23463 = n23441 ^ n23440;
  assign n23464 = n23463 ^ n1784;
  assign n23465 = n23439 ^ n23403;
  assign n23469 = n23468 ^ n23465;
  assign n23472 = n23435 ^ n23433;
  assign n23473 = n23472 ^ n2817;
  assign n23474 = n23432 ^ n23431;
  assign n23475 = n23474 ^ n1574;
  assign n23476 = n23430 ^ n23428;
  assign n2696 = n2689 ^ n2641;
  assign n2697 = n2696 ^ n2622;
  assign n2698 = n2697 ^ n1490;
  assign n23477 = n23476 ^ n2698;
  assign n23478 = n23427 ^ n23425;
  assign n2590 = n2564 ^ n1518;
  assign n2597 = n2596 ^ n2590;
  assign n2601 = n2600 ^ n2597;
  assign n23479 = n23478 ^ n2601;
  assign n23481 = n23422 ^ n23420;
  assign n3170 = n3163 ^ n2517;
  assign n3174 = n3173 ^ n3170;
  assign n3175 = n3174 ^ n2606;
  assign n23482 = n23481 ^ n3175;
  assign n23483 = n23419 ^ n23418;
  assign n23487 = n23486 ^ n23483;
  assign n23488 = n23417 ^ n23416;
  assign n1430 = n1407 ^ n1323;
  assign n1431 = n1430 ^ n1426;
  assign n1435 = n1434 ^ n1431;
  assign n23489 = n23488 ^ n1435;
  assign n23490 = n23413 ^ n23411;
  assign n1250 = n1207 ^ n1156;
  assign n1251 = n1250 ^ n1244;
  assign n1252 = n1251 ^ n1172;
  assign n23491 = n23490 ^ n1252;
  assign n23492 = n23410 ^ n23408;
  assign n1232 = n1131 ^ n1076;
  assign n1233 = n1232 ^ n1001;
  assign n1237 = n1236 ^ n1233;
  assign n23493 = n23492 ^ n1237;
  assign n23494 = n23407 ^ n23406;
  assign n1223 = n1145 ^ n1058;
  assign n1227 = n1226 ^ n1223;
  assign n1228 = n1227 ^ n999;
  assign n23495 = n23494 ^ n1228;
  assign n23143 = n23142 ^ n23141;
  assign n23144 = n23143 ^ n863;
  assign n23067 = n23066 ^ n23046;
  assign n23071 = n23070 ^ n23067;
  assign n23072 = n23065 ^ n23047;
  assign n23073 = n23072 ^ n756;
  assign n23075 = n23063 ^ n23049;
  assign n589 = n585 ^ n576;
  assign n596 = n595 ^ n589;
  assign n600 = n599 ^ n596;
  assign n23076 = n23075 ^ n600;
  assign n23077 = n23062 ^ n23051;
  assign n23078 = n23077 ^ n3287;
  assign n23079 = n23059 ^ n23057;
  assign n23083 = n23082 ^ n23079;
  assign n2226 = n2225 ^ n2132;
  assign n2227 = n2226 ^ n2216;
  assign n2228 = n2227 ^ n518;
  assign n23085 = n2228 & ~n23052;
  assign n23089 = n23088 ^ n23085;
  assign n23090 = n23053 ^ n23052;
  assign n23091 = n23090 ^ n23088;
  assign n23092 = n23089 & n23091;
  assign n23093 = n23092 ^ n23085;
  assign n23084 = n23056 ^ n23054;
  assign n23094 = n23093 ^ n23084;
  assign n23095 = n14478 ^ n2405;
  assign n23096 = n23095 ^ n18399;
  assign n23097 = n23096 ^ n672;
  assign n23098 = n23097 ^ n23084;
  assign n23099 = n23094 & ~n23098;
  assign n23100 = n23099 ^ n23097;
  assign n23101 = n23100 ^ n23079;
  assign n23102 = n23083 & ~n23101;
  assign n23103 = n23102 ^ n23082;
  assign n23107 = n23106 ^ n23103;
  assign n23108 = n23061 ^ n23060;
  assign n23109 = n23108 ^ n23103;
  assign n23110 = n23107 & n23109;
  assign n23111 = n23110 ^ n23106;
  assign n23112 = n23111 ^ n3287;
  assign n23113 = ~n23078 & ~n23112;
  assign n23114 = n23113 ^ n23077;
  assign n23115 = n23114 ^ n23075;
  assign n23116 = ~n23076 & ~n23115;
  assign n23117 = n23116 ^ n600;
  assign n23074 = n23064 ^ n23048;
  assign n23118 = n23117 ^ n23074;
  assign n23119 = n23074 ^ n659;
  assign n23120 = n23118 & ~n23119;
  assign n23121 = n23120 ^ n659;
  assign n23122 = n23121 ^ n23072;
  assign n23123 = n23073 & ~n23122;
  assign n23124 = n23123 ^ n756;
  assign n23125 = n23124 ^ n23067;
  assign n23126 = ~n23071 & n23125;
  assign n23127 = n23126 ^ n23070;
  assign n23496 = n23143 ^ n23127;
  assign n23497 = n23144 & ~n23496;
  assign n23498 = n23497 ^ n863;
  assign n23499 = n23498 ^ n23494;
  assign n23500 = ~n23495 & n23499;
  assign n23501 = n23500 ^ n1228;
  assign n23502 = n23501 ^ n23492;
  assign n23503 = n23493 & ~n23502;
  assign n23504 = n23503 ^ n1237;
  assign n23505 = n23504 ^ n23490;
  assign n23506 = ~n23491 & n23505;
  assign n23507 = n23506 ^ n1252;
  assign n1414 = n1395 ^ n1262;
  assign n1415 = n1414 ^ n1308;
  assign n1419 = n1418 ^ n1415;
  assign n23508 = n23507 ^ n1419;
  assign n23509 = n23415 ^ n23414;
  assign n23510 = n23509 ^ n23507;
  assign n23511 = n23508 & ~n23510;
  assign n23512 = n23511 ^ n1419;
  assign n23513 = n23512 ^ n23488;
  assign n23514 = n23489 & ~n23513;
  assign n23515 = n23514 ^ n1435;
  assign n23516 = n23515 ^ n23483;
  assign n23517 = n23487 & ~n23516;
  assign n23518 = n23517 ^ n23486;
  assign n23519 = n23518 ^ n23481;
  assign n23520 = n23482 & ~n23519;
  assign n23521 = n23520 ^ n3175;
  assign n23480 = n23424 ^ n23423;
  assign n23522 = n23521 ^ n23480;
  assign n23523 = n23480 ^ n2612;
  assign n23524 = n23522 & ~n23523;
  assign n23525 = n23524 ^ n2612;
  assign n23526 = n23525 ^ n23478;
  assign n23527 = ~n23479 & n23526;
  assign n23528 = n23527 ^ n2601;
  assign n23529 = n23528 ^ n23476;
  assign n23530 = n23477 & ~n23529;
  assign n23531 = n23530 ^ n2698;
  assign n23532 = n23531 ^ n23474;
  assign n23533 = ~n23475 & n23532;
  assign n23534 = n23533 ^ n1574;
  assign n23535 = n23534 ^ n23472;
  assign n23536 = n23473 & ~n23535;
  assign n23537 = n23536 ^ n2817;
  assign n23471 = n23437 ^ n23436;
  assign n23538 = n23537 ^ n23471;
  assign n23542 = n23541 ^ n23471;
  assign n23543 = n23538 & ~n23542;
  assign n23544 = n23543 ^ n23541;
  assign n23470 = n23438 ^ n23405;
  assign n23545 = n23544 ^ n23470;
  assign n23546 = n23470 ^ n2948;
  assign n23547 = ~n23545 & n23546;
  assign n23548 = n23547 ^ n2948;
  assign n23549 = n23548 ^ n23465;
  assign n23550 = n23469 & ~n23549;
  assign n23551 = n23550 ^ n23468;
  assign n23552 = n23551 ^ n23463;
  assign n23553 = n23464 & ~n23552;
  assign n23554 = n23553 ^ n1784;
  assign n23555 = n23554 ^ n1793;
  assign n23377 = n23376 ^ n23294;
  assign n23378 = n23295 & ~n23377;
  assign n23379 = n23378 ^ n20568;
  assign n23168 = n23167 ^ n23165;
  assign n23277 = n23276 ^ n23165;
  assign n23278 = n23168 & ~n23277;
  assign n23279 = n23278 ^ n23167;
  assign n23163 = n22919 ^ n22812;
  assign n23161 = n21761 ^ n21139;
  assign n23162 = n23161 ^ n22252;
  assign n23164 = n23163 ^ n23162;
  assign n23291 = n23279 ^ n23164;
  assign n23292 = n23291 ^ n20560;
  assign n23443 = n23379 ^ n23292;
  assign n23442 = n23440 & ~n23441;
  assign n23556 = n23443 ^ n23442;
  assign n23557 = n23556 ^ n1793;
  assign n23558 = ~n23555 & ~n23557;
  assign n23559 = n23558 ^ n23556;
  assign n23380 = n23379 ^ n23291;
  assign n23381 = ~n23292 & n23380;
  assign n23382 = n23381 ^ n20560;
  assign n23280 = n23279 ^ n23163;
  assign n23281 = ~n23164 & ~n23280;
  assign n23282 = n23281 ^ n23162;
  assign n23159 = n22922 ^ n22810;
  assign n23157 = n21760 ^ n21160;
  assign n23158 = n23157 ^ n22284;
  assign n23160 = n23159 ^ n23158;
  assign n23289 = n23282 ^ n23160;
  assign n23290 = n23289 ^ n20559;
  assign n23445 = n23382 ^ n23290;
  assign n23444 = n23442 & n23443;
  assign n23461 = n23445 ^ n23444;
  assign n1886 = n1874 ^ n1822;
  assign n1887 = n1886 ^ n1800;
  assign n1891 = n1890 ^ n1887;
  assign n23462 = n23461 ^ n1891;
  assign n23591 = n23559 ^ n23462;
  assign n23588 = n22407 ^ n21810;
  assign n23589 = n23588 ^ n22337;
  assign n23584 = n23556 ^ n23555;
  assign n23585 = n22476 ^ n21493;
  assign n23586 = n23585 ^ n22342;
  assign n23587 = ~n23584 & ~n23586;
  assign n23590 = n23589 ^ n23587;
  assign n23618 = n23591 ^ n23590;
  assign n23615 = n23586 ^ n23584;
  assign n23616 = ~n20955 & n23615;
  assign n23617 = n23616 ^ n20953;
  assign n23650 = n23618 ^ n23617;
  assign n23651 = n23615 ^ n20955;
  assign n23652 = ~n23650 & ~n23651;
  assign n23592 = n23591 ^ n23589;
  assign n23593 = ~n23590 & ~n23592;
  assign n23594 = n23593 ^ n23587;
  assign n23560 = n23559 ^ n1891;
  assign n23561 = n23462 & n23560;
  assign n23562 = n23561 ^ n23461;
  assign n23446 = ~n23444 & ~n23445;
  assign n23383 = n23382 ^ n23289;
  assign n23384 = ~n23290 & ~n23383;
  assign n23385 = n23384 ^ n20559;
  assign n23287 = n22925 ^ n22808;
  assign n23283 = n23282 ^ n23159;
  assign n23284 = ~n23160 & ~n23283;
  assign n23285 = n23284 ^ n23158;
  assign n23155 = n21759 ^ n21138;
  assign n23156 = n23155 ^ n22316;
  assign n23286 = n23285 ^ n23156;
  assign n23288 = n23287 ^ n23286;
  assign n23386 = n23385 ^ n23288;
  assign n23401 = n23386 ^ n20557;
  assign n23459 = n23446 ^ n23401;
  assign n1898 = n1871 ^ n1831;
  assign n1899 = n1898 ^ n1895;
  assign n1903 = n1902 ^ n1899;
  assign n23460 = n23459 ^ n1903;
  assign n23582 = n23562 ^ n23460;
  assign n23580 = n22345 ^ n21492;
  assign n23581 = n23580 ^ n22329;
  assign n23583 = n23582 ^ n23581;
  assign n23623 = n23594 ^ n23583;
  assign n23619 = n23618 ^ n23616;
  assign n23620 = ~n23617 & ~n23619;
  assign n23621 = n23620 ^ n20953;
  assign n23622 = n23621 ^ n20950;
  assign n23649 = n23623 ^ n23622;
  assign n23702 = n23652 ^ n23649;
  assign n23692 = n2318 & n23651;
  assign n23693 = n23692 ^ n2312;
  assign n23694 = n23651 ^ n23650;
  assign n23695 = n23694 ^ n23692;
  assign n23696 = n23693 & ~n23695;
  assign n23697 = n23696 ^ n2312;
  assign n23701 = n23700 ^ n23697;
  assign n24333 = n23702 ^ n23701;
  assign n23607 = n23052 ^ n2228;
  assign n24123 = n23607 ^ n22476;
  assign n24124 = n24123 ^ n22329;
  assign n23755 = n23518 ^ n3175;
  assign n23756 = n23755 ^ n23481;
  assign n23753 = n23163 ^ n22354;
  assign n23754 = n23753 ^ n22298;
  assign n23757 = n23756 ^ n23754;
  assign n23760 = n23515 ^ n23487;
  assign n23758 = n22357 ^ n22266;
  assign n23759 = n23758 ^ n23165;
  assign n23761 = n23760 ^ n23759;
  assign n23764 = n23512 ^ n23489;
  assign n23762 = n22361 ^ n22237;
  assign n23763 = n23762 ^ n23270;
  assign n23765 = n23764 ^ n23763;
  assign n23768 = n23509 ^ n1419;
  assign n23769 = n23768 ^ n23507;
  assign n23766 = n22366 ^ n22077;
  assign n23767 = n23766 ^ n23171;
  assign n23770 = n23769 ^ n23767;
  assign n23773 = n23504 ^ n23491;
  assign n23771 = n23259 ^ n22017;
  assign n23772 = n23771 ^ n22371;
  assign n23774 = n23773 ^ n23772;
  assign n23776 = n23175 ^ n21890;
  assign n23777 = n23776 ^ n22375;
  assign n23775 = n23501 ^ n23493;
  assign n23778 = n23777 ^ n23775;
  assign n23781 = n23179 ^ n22379;
  assign n23782 = n23781 ^ n21881;
  assign n23779 = n23498 ^ n1228;
  assign n23780 = n23779 ^ n23494;
  assign n23783 = n23782 ^ n23780;
  assign n23784 = n23183 ^ n21456;
  assign n23785 = n23784 ^ n22549;
  assign n23145 = n23144 ^ n23127;
  assign n23786 = n23785 ^ n23145;
  assign n23791 = n23118 ^ n659;
  assign n23789 = n23192 ^ n21466;
  assign n23790 = n23789 ^ n22532;
  assign n23792 = n23791 ^ n23790;
  assign n23811 = n23114 ^ n23076;
  assign n23795 = n23111 ^ n23078;
  assign n23793 = n23146 ^ n21469;
  assign n23794 = n23793 ^ n22388;
  assign n23796 = n23795 ^ n23794;
  assign n23799 = n23201 ^ n22390;
  assign n23800 = n23799 ^ n21477;
  assign n23797 = n23108 ^ n23106;
  assign n23798 = n23797 ^ n23103;
  assign n23801 = n23800 ^ n23798;
  assign n23730 = n23205 ^ n22391;
  assign n23731 = n23730 ^ n21846;
  assign n23728 = n23100 ^ n23082;
  assign n23729 = n23728 ^ n23079;
  assign n23732 = n23731 ^ n23729;
  assign n23667 = n23097 ^ n23093;
  assign n23668 = n23667 ^ n23084;
  assign n23665 = n23208 ^ n21482;
  assign n23666 = n23665 ^ n22507;
  assign n23669 = n23668 ^ n23666;
  assign n23577 = n22340 ^ n21490;
  assign n23578 = n23577 ^ n22990;
  assign n23563 = n23562 ^ n23459;
  assign n23564 = n23460 & ~n23563;
  assign n23565 = n23564 ^ n1903;
  assign n2037 = n2036 ^ n1952;
  assign n2038 = n2037 ^ n2033;
  assign n2039 = n2038 ^ n2028;
  assign n23575 = n23565 ^ n2039;
  assign n23447 = n23401 & ~n23446;
  assign n23396 = n22928 ^ n22806;
  assign n23392 = n23287 ^ n23156;
  assign n23393 = n23287 ^ n23285;
  assign n23394 = ~n23392 & n23393;
  assign n23395 = n23394 ^ n23156;
  assign n23397 = n23396 ^ n23395;
  assign n23390 = n21494 ^ n20960;
  assign n23391 = n23390 ^ n22460;
  assign n23398 = n23397 ^ n23391;
  assign n23399 = n23398 ^ n20419;
  assign n23387 = n23288 ^ n20557;
  assign n23388 = ~n23386 & n23387;
  assign n23389 = n23388 ^ n20557;
  assign n23400 = n23399 ^ n23389;
  assign n23457 = n23447 ^ n23400;
  assign n23576 = n23575 ^ n23457;
  assign n23579 = n23578 ^ n23576;
  assign n23595 = n23594 ^ n23582;
  assign n23596 = ~n23583 & ~n23595;
  assign n23597 = n23596 ^ n23581;
  assign n23598 = n23597 ^ n23578;
  assign n23599 = ~n23579 & n23598;
  assign n23600 = n23599 ^ n23576;
  assign n23570 = n23389 ^ n20419;
  assign n23571 = n23398 ^ n23389;
  assign n23572 = n23570 & ~n23571;
  assign n23573 = n23572 ^ n20419;
  assign n23458 = n23457 ^ n2039;
  assign n23566 = n23565 ^ n23457;
  assign n23567 = ~n23458 & n23566;
  assign n23568 = n23567 ^ n2039;
  assign n23453 = n23396 ^ n23391;
  assign n23454 = n23397 & ~n23453;
  assign n23455 = n23454 ^ n23391;
  assign n23449 = n22931 ^ n22804;
  assign n23448 = n23400 & n23447;
  assign n23450 = n23449 ^ n23448;
  assign n23153 = n23152 ^ n22348;
  assign n23154 = n23153 ^ n21797;
  assign n23451 = n23450 ^ n23154;
  assign n23452 = n23451 ^ n22453;
  assign n23456 = n23455 ^ n23452;
  assign n23569 = n23568 ^ n23456;
  assign n23574 = n23573 ^ n23569;
  assign n23601 = n23600 ^ n23574;
  assign n23602 = n22335 ^ n21826;
  assign n23603 = n23602 ^ n23043;
  assign n23604 = n23603 ^ n23574;
  assign n23605 = ~n23601 & ~n23604;
  assign n23606 = n23605 ^ n23603;
  assign n23608 = n23607 ^ n23606;
  assign n23148 = n23130 ^ n21486;
  assign n23149 = n23148 ^ n22331;
  assign n23639 = n23607 ^ n23149;
  assign n23640 = n23608 & ~n23639;
  assign n23641 = n23640 ^ n23149;
  assign n23638 = n23090 ^ n23089;
  assign n23642 = n23641 ^ n23638;
  assign n23636 = n23210 ^ n21836;
  assign n23637 = n23636 ^ n22397;
  assign n23662 = n23638 ^ n23637;
  assign n23663 = n23642 & n23662;
  assign n23664 = n23663 ^ n23637;
  assign n23725 = n23668 ^ n23664;
  assign n23726 = ~n23669 & ~n23725;
  assign n23727 = n23726 ^ n23666;
  assign n23802 = n23731 ^ n23727;
  assign n23803 = n23732 & ~n23802;
  assign n23804 = n23803 ^ n23729;
  assign n23805 = n23804 ^ n23798;
  assign n23806 = n23801 & n23805;
  assign n23807 = n23806 ^ n23800;
  assign n23808 = n23807 ^ n23795;
  assign n23809 = n23796 & ~n23808;
  assign n23810 = n23809 ^ n23794;
  assign n23812 = n23811 ^ n23810;
  assign n23813 = n23194 ^ n22385;
  assign n23814 = n23813 ^ n21468;
  assign n23815 = n23814 ^ n23811;
  assign n23816 = n23812 & n23815;
  assign n23817 = n23816 ^ n23814;
  assign n23818 = n23817 ^ n23791;
  assign n23819 = ~n23792 & n23818;
  assign n23820 = n23819 ^ n23790;
  assign n23788 = n23121 ^ n23073;
  assign n23821 = n23820 ^ n23788;
  assign n23822 = n23188 ^ n21868;
  assign n23823 = n23822 ^ n22383;
  assign n23824 = n23823 ^ n23788;
  assign n23825 = ~n23821 & n23824;
  assign n23826 = n23825 ^ n23823;
  assign n23787 = n23124 ^ n23071;
  assign n23827 = n23826 ^ n23787;
  assign n23828 = n22542 ^ n21458;
  assign n23829 = n23828 ^ n23185;
  assign n23830 = n23829 ^ n23787;
  assign n23831 = n23827 & ~n23830;
  assign n23832 = n23831 ^ n23829;
  assign n23833 = n23832 ^ n23145;
  assign n23834 = ~n23786 & ~n23833;
  assign n23835 = n23834 ^ n23785;
  assign n23836 = n23835 ^ n23780;
  assign n23837 = n23783 & ~n23836;
  assign n23838 = n23837 ^ n23782;
  assign n23839 = n23838 ^ n23775;
  assign n23840 = n23778 & n23839;
  assign n23841 = n23840 ^ n23777;
  assign n23842 = n23841 ^ n23773;
  assign n23843 = n23774 & n23842;
  assign n23844 = n23843 ^ n23772;
  assign n23845 = n23844 ^ n23769;
  assign n23846 = n23770 & n23845;
  assign n23847 = n23846 ^ n23767;
  assign n23848 = n23847 ^ n23764;
  assign n23849 = ~n23765 & ~n23848;
  assign n23850 = n23849 ^ n23763;
  assign n23851 = n23850 ^ n23760;
  assign n23852 = ~n23761 & n23851;
  assign n23853 = n23852 ^ n23759;
  assign n23854 = n23853 ^ n23754;
  assign n23855 = ~n23757 & ~n23854;
  assign n23856 = n23855 ^ n23756;
  assign n23751 = n23522 ^ n2612;
  assign n23749 = n22369 ^ n22352;
  assign n23750 = n23749 ^ n23159;
  assign n23752 = n23751 ^ n23750;
  assign n23876 = n23856 ^ n23752;
  assign n23877 = n23876 ^ n21660;
  assign n23878 = n23853 ^ n23757;
  assign n23879 = n23878 ^ n21644;
  assign n23881 = n23847 ^ n23763;
  assign n23882 = n23881 ^ n23764;
  assign n23883 = n23882 ^ n20945;
  assign n23885 = n23841 ^ n23774;
  assign n23886 = n23885 ^ n21543;
  assign n23889 = n23832 ^ n23786;
  assign n23890 = n23889 ^ n21471;
  assign n23892 = n23823 ^ n23821;
  assign n23893 = n23892 ^ n21518;
  assign n23894 = n23817 ^ n23792;
  assign n23895 = n23894 ^ n21480;
  assign n23897 = n23807 ^ n23794;
  assign n23898 = n23897 ^ n23795;
  assign n23899 = n23898 ^ n21446;
  assign n23733 = n23732 ^ n23727;
  assign n23901 = n23733 ^ n21328;
  assign n23670 = n23669 ^ n23664;
  assign n23671 = n23670 ^ n21311;
  assign n23643 = n23642 ^ n23637;
  assign n23644 = n23643 ^ n21296;
  assign n23609 = n23608 ^ n23149;
  assign n23610 = n23609 ^ n21282;
  assign n23611 = n23603 ^ n23601;
  assign n23612 = n23611 ^ n21247;
  assign n23613 = n23597 ^ n23579;
  assign n23614 = n23613 ^ n20949;
  assign n23624 = n23623 ^ n23621;
  assign n23625 = ~n23622 & ~n23624;
  assign n23626 = n23625 ^ n20950;
  assign n23627 = n23626 ^ n23613;
  assign n23628 = n23614 & ~n23627;
  assign n23629 = n23628 ^ n20949;
  assign n23630 = n23629 ^ n23611;
  assign n23631 = ~n23612 & ~n23630;
  assign n23632 = n23631 ^ n21247;
  assign n23633 = n23632 ^ n23609;
  assign n23634 = n23610 & ~n23633;
  assign n23635 = n23634 ^ n21282;
  assign n23659 = n23643 ^ n23635;
  assign n23660 = n23644 & n23659;
  assign n23661 = n23660 ^ n21296;
  assign n23721 = n23670 ^ n23661;
  assign n23722 = n23671 & ~n23721;
  assign n23723 = n23722 ^ n21311;
  assign n23902 = n23733 ^ n23723;
  assign n23903 = ~n23901 & ~n23902;
  assign n23904 = n23903 ^ n21328;
  assign n23900 = n23804 ^ n23801;
  assign n23905 = n23904 ^ n23900;
  assign n23906 = n23900 ^ n21342;
  assign n23907 = n23905 & n23906;
  assign n23908 = n23907 ^ n21342;
  assign n23909 = n23908 ^ n23898;
  assign n23910 = ~n23899 & n23909;
  assign n23911 = n23910 ^ n21446;
  assign n23896 = n23814 ^ n23812;
  assign n23912 = n23911 ^ n23896;
  assign n23913 = n23896 ^ n21505;
  assign n23914 = n23912 & ~n23913;
  assign n23915 = n23914 ^ n21505;
  assign n23916 = n23915 ^ n23894;
  assign n23917 = n23895 & n23916;
  assign n23918 = n23917 ^ n21480;
  assign n23919 = n23918 ^ n23892;
  assign n23920 = n23893 & n23919;
  assign n23921 = n23920 ^ n21518;
  assign n23891 = n23829 ^ n23827;
  assign n23922 = n23921 ^ n23891;
  assign n23923 = n23891 ^ n21475;
  assign n23924 = n23922 & n23923;
  assign n23925 = n23924 ^ n21475;
  assign n23926 = n23925 ^ n23889;
  assign n23927 = n23890 & ~n23926;
  assign n23928 = n23927 ^ n21471;
  assign n23888 = n23835 ^ n23783;
  assign n23929 = n23928 ^ n23888;
  assign n23930 = n23888 ^ n21495;
  assign n23931 = ~n23929 & ~n23930;
  assign n23932 = n23931 ^ n21495;
  assign n23887 = n23838 ^ n23778;
  assign n23933 = n23932 ^ n23887;
  assign n23934 = n23887 ^ n21464;
  assign n23935 = n23933 & n23934;
  assign n23936 = n23935 ^ n21464;
  assign n23937 = n23936 ^ n23885;
  assign n23938 = ~n23886 & n23937;
  assign n23939 = n23938 ^ n21543;
  assign n23884 = n23844 ^ n23770;
  assign n23940 = n23939 ^ n23884;
  assign n23941 = n23884 ^ n21460;
  assign n23942 = ~n23940 & n23941;
  assign n23943 = n23942 ^ n21460;
  assign n23944 = n23943 ^ n23882;
  assign n23945 = n23883 & ~n23944;
  assign n23946 = n23945 ^ n20945;
  assign n23880 = n23850 ^ n23761;
  assign n23947 = n23946 ^ n23880;
  assign n23948 = n23880 ^ n21630;
  assign n23949 = n23947 & n23948;
  assign n23950 = n23949 ^ n21630;
  assign n23951 = n23950 ^ n23878;
  assign n23952 = ~n23879 & ~n23951;
  assign n23953 = n23952 ^ n21644;
  assign n23954 = n23953 ^ n23876;
  assign n23955 = ~n23877 & n23954;
  assign n23956 = n23955 ^ n21660;
  assign n23977 = n23956 ^ n21678;
  assign n23857 = n23856 ^ n23751;
  assign n23858 = n23752 & n23857;
  assign n23859 = n23858 ^ n23750;
  assign n23746 = n23525 ^ n2601;
  assign n23747 = n23746 ^ n23478;
  assign n23744 = n23287 ^ n22364;
  assign n23745 = n23744 ^ n22347;
  assign n23748 = n23747 ^ n23745;
  assign n23874 = n23859 ^ n23748;
  assign n23978 = n23977 ^ n23874;
  assign n23979 = n23943 ^ n23883;
  assign n23980 = n23940 ^ n21460;
  assign n23981 = n23922 ^ n21475;
  assign n23982 = n23918 ^ n23893;
  assign n23724 = n23723 ^ n21328;
  assign n23734 = n23733 ^ n23724;
  assign n23645 = n23644 ^ n23635;
  assign n23646 = n23629 ^ n21247;
  assign n23647 = n23646 ^ n23611;
  assign n23648 = n23626 ^ n23614;
  assign n23653 = n23649 & n23652;
  assign n23654 = n23648 & n23653;
  assign n23655 = ~n23647 & n23654;
  assign n23656 = n23632 ^ n23610;
  assign n23657 = ~n23655 & n23656;
  assign n23658 = ~n23645 & ~n23657;
  assign n23672 = n23671 ^ n23661;
  assign n23735 = ~n23658 & ~n23672;
  assign n23983 = n23734 & n23735;
  assign n23984 = n23905 ^ n21342;
  assign n23985 = n23983 & n23984;
  assign n23986 = n23908 ^ n21446;
  assign n23987 = n23986 ^ n23898;
  assign n23988 = ~n23985 & ~n23987;
  assign n23989 = n23912 ^ n21505;
  assign n23990 = ~n23988 & n23989;
  assign n23991 = n23915 ^ n23895;
  assign n23992 = ~n23990 & n23991;
  assign n23993 = n23982 & ~n23992;
  assign n23994 = ~n23981 & n23993;
  assign n23995 = n23925 ^ n23890;
  assign n23996 = n23994 & n23995;
  assign n23997 = n23929 ^ n21495;
  assign n23998 = n23996 & ~n23997;
  assign n23999 = n23933 ^ n21464;
  assign n24000 = ~n23998 & n23999;
  assign n24001 = n23936 ^ n23886;
  assign n24002 = n24000 & n24001;
  assign n24003 = n23980 & ~n24002;
  assign n24004 = n23979 & n24003;
  assign n24005 = n23947 ^ n21630;
  assign n24006 = ~n24004 & ~n24005;
  assign n24007 = n23950 ^ n23879;
  assign n24008 = ~n24006 & n24007;
  assign n24009 = n23953 ^ n23877;
  assign n24010 = n24008 & ~n24009;
  assign n24011 = ~n23978 & ~n24010;
  assign n23875 = n23874 ^ n21678;
  assign n23957 = n23956 ^ n23874;
  assign n23958 = n23875 & ~n23957;
  assign n23959 = n23958 ^ n21678;
  assign n23860 = n23859 ^ n23745;
  assign n23861 = n23748 & ~n23860;
  assign n23862 = n23861 ^ n23747;
  assign n23742 = n23528 ^ n23477;
  assign n23740 = n23396 ^ n22252;
  assign n23741 = n23740 ^ n21762;
  assign n23743 = n23742 ^ n23741;
  assign n23872 = n23862 ^ n23743;
  assign n23873 = n23872 ^ n21142;
  assign n24012 = n23959 ^ n23873;
  assign n24013 = ~n24011 & ~n24012;
  assign n23960 = n23959 ^ n23872;
  assign n23961 = ~n23873 & ~n23960;
  assign n23962 = n23961 ^ n21142;
  assign n23867 = n22284 ^ n21769;
  assign n23868 = n23867 ^ n23449;
  assign n23866 = n23531 ^ n23475;
  assign n23869 = n23868 ^ n23866;
  assign n23863 = n23862 ^ n23742;
  assign n23864 = n23743 & n23863;
  assign n23865 = n23864 ^ n23741;
  assign n23870 = n23869 ^ n23865;
  assign n23871 = n23870 ^ n21147;
  assign n23976 = n23962 ^ n23871;
  assign n24016 = n24013 ^ n23976;
  assign n24020 = n24019 ^ n24016;
  assign n24021 = n24012 ^ n24011;
  assign n24022 = n24021 ^ n1628;
  assign n24023 = n24010 ^ n23978;
  assign n24027 = n24026 ^ n24023;
  assign n24028 = n24007 ^ n24006;
  assign n24029 = n24028 ^ n2802;
  assign n24030 = n24005 ^ n24004;
  assign n2782 = n2721 ^ n1493;
  assign n2783 = n2782 ^ n2768;
  assign n2787 = n2786 ^ n2783;
  assign n24031 = n24030 ^ n2787;
  assign n24032 = n24003 ^ n23979;
  assign n24033 = n24032 ^ n2777;
  assign n24034 = n24002 ^ n23980;
  assign n24035 = n24034 ^ n3209;
  assign n24036 = n24001 ^ n24000;
  assign n24037 = n24036 ^ n3058;
  assign n24038 = n23999 ^ n23998;
  assign n2489 = n2488 ^ n2438;
  assign n2490 = n2489 ^ n2472;
  assign n2491 = n2490 ^ n1550;
  assign n24039 = n24038 ^ n2491;
  assign n24040 = n23997 ^ n23996;
  assign n3031 = n3026 ^ n1484;
  assign n3032 = n3031 ^ n2428;
  assign n3033 = n3032 ^ n2470;
  assign n24041 = n24040 ^ n3033;
  assign n24043 = n23993 ^ n23981;
  assign n1269 = n1268 ^ n1178;
  assign n1276 = n1275 ^ n1269;
  assign n1280 = n1279 ^ n1276;
  assign n24044 = n24043 ^ n1280;
  assign n24046 = n23991 ^ n23990;
  assign n1087 = n1083 ^ n1008;
  assign n1091 = n1090 ^ n1087;
  assign n1095 = n1094 ^ n1091;
  assign n24047 = n24046 ^ n1095;
  assign n24048 = n23989 ^ n23988;
  assign n24049 = n24048 ^ n949;
  assign n24050 = n23987 ^ n23985;
  assign n938 = n922 ^ n868;
  assign n939 = n938 ^ n846;
  assign n940 = n939 ^ n934;
  assign n24051 = n24050 ^ n940;
  assign n23736 = n23735 ^ n23734;
  assign n23737 = n23736 ^ n827;
  assign n23673 = n23672 ^ n23658;
  assign n23674 = n23673 ^ n3272;
  assign n23675 = n23657 ^ n23645;
  assign n23679 = n23678 ^ n23675;
  assign n23680 = n23656 ^ n23655;
  assign n23684 = n23683 ^ n23680;
  assign n23686 = n22133 ^ n15241;
  assign n23687 = n23686 ^ n18924;
  assign n23688 = n23687 ^ n515;
  assign n23685 = n23654 ^ n23647;
  assign n23689 = n23688 ^ n23685;
  assign n23690 = n23653 ^ n23648;
  assign n694 = n693 ^ n675;
  assign n695 = n694 ^ n530;
  assign n696 = n695 ^ n635;
  assign n23691 = n23690 ^ n696;
  assign n23703 = n23702 ^ n23697;
  assign n23704 = n23701 & ~n23703;
  assign n23705 = n23704 ^ n23700;
  assign n23706 = n23705 ^ n23690;
  assign n23707 = n23691 & ~n23706;
  assign n23708 = n23707 ^ n696;
  assign n23709 = n23708 ^ n23685;
  assign n23710 = ~n23689 & n23709;
  assign n23711 = n23710 ^ n23688;
  assign n23712 = n23711 ^ n23680;
  assign n23713 = n23684 & ~n23712;
  assign n23714 = n23713 ^ n23683;
  assign n23715 = n23714 ^ n23675;
  assign n23716 = n23679 & ~n23715;
  assign n23717 = n23716 ^ n23678;
  assign n23718 = n23717 ^ n23673;
  assign n23719 = ~n23674 & n23718;
  assign n23720 = n23719 ^ n3272;
  assign n24053 = n23736 ^ n23720;
  assign n24054 = ~n23737 & n24053;
  assign n24055 = n24054 ^ n827;
  assign n24052 = n23984 ^ n23983;
  assign n24056 = n24055 ^ n24052;
  assign n24057 = n24052 ^ n839;
  assign n24058 = n24056 & ~n24057;
  assign n24059 = n24058 ^ n839;
  assign n24060 = n24059 ^ n24050;
  assign n24061 = n24051 & ~n24060;
  assign n24062 = n24061 ^ n940;
  assign n24063 = n24062 ^ n24048;
  assign n24064 = n24049 & ~n24063;
  assign n24065 = n24064 ^ n949;
  assign n24066 = n24065 ^ n24046;
  assign n24067 = ~n24047 & n24066;
  assign n24068 = n24067 ^ n1095;
  assign n24045 = n23992 ^ n23982;
  assign n24069 = n24068 ^ n24045;
  assign n24070 = n1448 ^ n1344;
  assign n24071 = n24070 ^ n1099;
  assign n24072 = n24071 ^ n1273;
  assign n24073 = n24072 ^ n24045;
  assign n24074 = ~n24069 & n24073;
  assign n24075 = n24074 ^ n24072;
  assign n24076 = n24075 ^ n24043;
  assign n24077 = n24044 & ~n24076;
  assign n24078 = n24077 ^ n1280;
  assign n24042 = n23995 ^ n23994;
  assign n24079 = n24078 ^ n24042;
  assign n2416 = n2412 ^ n1466;
  assign n2420 = n2419 ^ n2416;
  assign n2424 = n2423 ^ n2420;
  assign n24080 = n24042 ^ n2424;
  assign n24081 = n24079 & ~n24080;
  assign n24082 = n24081 ^ n2424;
  assign n24083 = n24082 ^ n24040;
  assign n24084 = n24041 & ~n24083;
  assign n24085 = n24084 ^ n3033;
  assign n24086 = n24085 ^ n24038;
  assign n24087 = ~n24039 & n24086;
  assign n24088 = n24087 ^ n2491;
  assign n24089 = n24088 ^ n24036;
  assign n24090 = n24037 & ~n24089;
  assign n24091 = n24090 ^ n3058;
  assign n24092 = n24091 ^ n24034;
  assign n24093 = n24035 & ~n24092;
  assign n24094 = n24093 ^ n3209;
  assign n24095 = n24094 ^ n24032;
  assign n24096 = ~n24033 & n24095;
  assign n24097 = n24096 ^ n2777;
  assign n24098 = n24097 ^ n24030;
  assign n24099 = n24031 & ~n24098;
  assign n24100 = n24099 ^ n2787;
  assign n24101 = n24100 ^ n24028;
  assign n24102 = n24029 & ~n24101;
  assign n24103 = n24102 ^ n2802;
  assign n24104 = n24103 ^ n1538;
  assign n24105 = n24009 ^ n24008;
  assign n24106 = n24105 ^ n24103;
  assign n24107 = n24104 & ~n24106;
  assign n24108 = n24107 ^ n1538;
  assign n24109 = n24108 ^ n24023;
  assign n24110 = n24027 & ~n24109;
  assign n24111 = n24110 ^ n24026;
  assign n24112 = n24111 ^ n24021;
  assign n24113 = ~n24022 & n24112;
  assign n24114 = n24113 ^ n1628;
  assign n24115 = n24114 ^ n24016;
  assign n24116 = ~n24020 & n24115;
  assign n24117 = n24116 ^ n24019;
  assign n24014 = n23976 & n24013;
  assign n23971 = n23534 ^ n23473;
  assign n23969 = n22961 ^ n22316;
  assign n23970 = n23969 ^ n21761;
  assign n23972 = n23971 ^ n23970;
  assign n23966 = n23866 ^ n23865;
  assign n23967 = ~n23869 & n23966;
  assign n23968 = n23967 ^ n23868;
  assign n23973 = n23972 ^ n23968;
  assign n23974 = n23973 ^ n21139;
  assign n23963 = n23962 ^ n23870;
  assign n23964 = ~n23871 & n23963;
  assign n23965 = n23964 ^ n21147;
  assign n23975 = n23974 ^ n23965;
  assign n24015 = n24014 ^ n23975;
  assign n24118 = n24117 ^ n24015;
  assign n24122 = n24121 ^ n24118;
  assign n24125 = n24124 ^ n24122;
  assign n24186 = n24125 ^ n21493;
  assign n2285 = n2241 ^ n2191;
  assign n2286 = n2285 ^ n2279;
  assign n2287 = n2286 ^ n2225;
  assign n24255 = n24186 ^ n2287;
  assign n25538 = n24333 ^ n24255;
  assign n25539 = n25538 ^ n23668;
  assign n24305 = n24059 ^ n940;
  assign n24306 = n24305 ^ n24050;
  assign n24303 = n23764 ^ n22549;
  assign n24304 = n24303 ^ n23175;
  assign n24307 = n24306 ^ n24304;
  assign n24309 = n23773 ^ n22383;
  assign n24310 = n24309 ^ n23183;
  assign n23738 = n23737 ^ n23720;
  assign n24311 = n24310 ^ n23738;
  assign n24314 = n23717 ^ n3272;
  assign n24315 = n24314 ^ n23673;
  assign n24312 = n23775 ^ n22532;
  assign n24313 = n24312 ^ n23185;
  assign n24316 = n24315 ^ n24313;
  assign n24317 = n23188 ^ n22385;
  assign n24318 = n24317 ^ n23780;
  assign n24247 = n23714 ^ n23679;
  assign n24319 = n24318 ^ n24247;
  assign n24320 = n23145 ^ n22388;
  assign n24321 = n24320 ^ n23192;
  assign n24252 = n23711 ^ n23684;
  assign n24322 = n24321 ^ n24252;
  assign n24325 = n23708 ^ n23689;
  assign n24323 = n23787 ^ n22390;
  assign n24324 = n24323 ^ n23194;
  assign n24326 = n24325 ^ n24324;
  assign n24328 = n23788 ^ n22391;
  assign n24329 = n24328 ^ n23146;
  assign n24327 = n23705 ^ n23691;
  assign n24330 = n24329 ^ n24327;
  assign n24331 = n23791 ^ n22507;
  assign n24332 = n24331 ^ n23201;
  assign n24334 = n24333 ^ n24332;
  assign n24337 = n23694 ^ n23693;
  assign n24335 = n23811 ^ n22397;
  assign n24336 = n24335 ^ n23205;
  assign n24338 = n24337 ^ n24336;
  assign n24341 = n23651 ^ n2318;
  assign n24339 = n23208 ^ n22331;
  assign n24340 = n24339 ^ n23795;
  assign n24342 = n24341 ^ n24340;
  assign n24140 = n23541 ^ n23537;
  assign n24141 = n24140 ^ n23471;
  assign n24138 = n22966 ^ n22460;
  assign n24139 = n24138 ^ n21760;
  assign n24142 = n24141 ^ n24139;
  assign n24135 = n23970 ^ n23968;
  assign n24136 = n23972 & ~n24135;
  assign n24137 = n24136 ^ n23971;
  assign n24169 = n24141 ^ n24137;
  assign n24170 = ~n24142 & n24169;
  assign n24171 = n24170 ^ n24139;
  assign n24167 = n22453 ^ n21759;
  assign n24168 = n24167 ^ n22957;
  assign n24172 = n24171 ^ n24168;
  assign n24166 = n23545 ^ n2948;
  assign n24173 = n24172 ^ n24166;
  assign n24174 = n24173 ^ n21138;
  assign n24143 = n24142 ^ n24137;
  assign n24144 = n24143 ^ n21160;
  assign n24132 = n23973 ^ n23965;
  assign n24133 = ~n23974 & ~n24132;
  assign n24134 = n24133 ^ n21139;
  assign n24163 = n24143 ^ n24134;
  assign n24164 = n24144 & ~n24163;
  assign n24165 = n24164 ^ n21160;
  assign n24225 = n24173 ^ n24165;
  assign n24226 = n24174 & n24225;
  assign n24227 = n24226 ^ n21138;
  assign n24228 = n24227 ^ n20960;
  assign n24219 = n24168 ^ n24166;
  assign n24220 = n24171 ^ n24166;
  assign n24221 = n24219 & ~n24220;
  assign n24222 = n24221 ^ n24168;
  assign n24218 = n23548 ^ n23469;
  assign n24223 = n24222 ^ n24218;
  assign n24216 = n22413 ^ n21494;
  assign n24217 = n24216 ^ n22951;
  assign n24224 = n24223 ^ n24217;
  assign n24229 = n24228 ^ n24224;
  assign n24131 = n23975 & n24014;
  assign n24145 = n24144 ^ n24134;
  assign n24162 = ~n24131 & ~n24145;
  assign n24175 = n24174 ^ n24165;
  assign n24215 = ~n24162 & n24175;
  assign n24230 = n24229 ^ n24215;
  assign n24231 = n24230 ^ n2022;
  assign n24176 = n24175 ^ n24162;
  assign n24177 = n24176 ^ n1990;
  assign n24146 = n24145 ^ n24131;
  assign n24147 = n24146 ^ n2000;
  assign n24128 = n24121 ^ n24015;
  assign n24129 = n24118 & ~n24128;
  assign n24130 = n24129 ^ n24121;
  assign n24159 = n24146 ^ n24130;
  assign n24160 = n24147 & ~n24159;
  assign n24161 = n24160 ^ n2000;
  assign n24212 = n24176 ^ n24161;
  assign n24213 = n24177 & ~n24212;
  assign n24214 = n24213 ^ n1990;
  assign n24360 = n24230 ^ n24214;
  assign n24361 = ~n24231 & n24360;
  assign n24362 = n24361 ^ n2022;
  assign n24363 = n24362 ^ n2150;
  assign n24354 = n24224 ^ n20960;
  assign n24355 = n24227 ^ n24224;
  assign n24356 = ~n24354 & ~n24355;
  assign n24357 = n24356 ^ n20960;
  assign n24348 = n24218 ^ n24217;
  assign n24349 = ~n24223 & n24348;
  assign n24350 = n24349 ^ n24217;
  assign n24266 = n23551 ^ n1784;
  assign n24267 = n24266 ^ n23463;
  assign n24351 = n24350 ^ n24267;
  assign n24346 = n22949 ^ n21797;
  assign n24347 = n24346 ^ n22411;
  assign n24352 = n24351 ^ n24347;
  assign n24353 = n24352 ^ n20958;
  assign n24358 = n24357 ^ n24353;
  assign n24345 = n24215 & n24229;
  assign n24359 = n24358 ^ n24345;
  assign n24364 = n24363 ^ n24359;
  assign n24343 = n23210 ^ n22335;
  assign n24344 = n24343 ^ n23798;
  assign n24365 = n24364 ^ n24344;
  assign n24150 = n23638 ^ n22407;
  assign n24151 = n24150 ^ n22990;
  assign n24149 = ~n24122 & ~n24124;
  assign n24152 = n24151 ^ n24149;
  assign n24148 = n24147 ^ n24130;
  assign n24179 = n24151 ^ n24148;
  assign n24180 = n24152 & ~n24179;
  assign n24181 = n24180 ^ n24149;
  assign n24178 = n24177 ^ n24161;
  assign n24182 = n24181 ^ n24178;
  assign n24157 = n23668 ^ n23043;
  assign n24158 = n24157 ^ n22345;
  assign n24233 = n24178 ^ n24158;
  assign n24234 = ~n24182 & ~n24233;
  assign n24235 = n24234 ^ n24158;
  assign n24232 = n24231 ^ n24214;
  assign n24236 = n24235 ^ n24232;
  assign n24210 = n23729 ^ n22340;
  assign n24211 = n24210 ^ n23130;
  assign n24366 = n24232 ^ n24211;
  assign n24367 = ~n24236 & ~n24366;
  assign n24368 = n24367 ^ n24211;
  assign n24369 = n24368 ^ n24364;
  assign n24370 = ~n24365 & ~n24369;
  assign n24371 = n24370 ^ n24344;
  assign n24372 = n24371 ^ n24341;
  assign n24373 = n24342 & n24372;
  assign n24374 = n24373 ^ n24340;
  assign n24375 = n24374 ^ n24337;
  assign n24376 = ~n24338 & ~n24375;
  assign n24377 = n24376 ^ n24336;
  assign n24378 = n24377 ^ n24332;
  assign n24379 = n24334 & n24378;
  assign n24380 = n24379 ^ n24333;
  assign n24381 = n24380 ^ n24329;
  assign n24382 = ~n24330 & n24381;
  assign n24383 = n24382 ^ n24327;
  assign n24384 = n24383 ^ n24325;
  assign n24385 = ~n24326 & n24384;
  assign n24386 = n24385 ^ n24324;
  assign n24387 = n24386 ^ n24252;
  assign n24388 = n24322 & ~n24387;
  assign n24389 = n24388 ^ n24321;
  assign n24390 = n24389 ^ n24318;
  assign n24391 = ~n24319 & n24390;
  assign n24392 = n24391 ^ n24247;
  assign n24393 = n24392 ^ n24315;
  assign n24394 = n24316 & n24393;
  assign n24395 = n24394 ^ n24313;
  assign n24396 = n24395 ^ n23738;
  assign n24397 = n24311 & ~n24396;
  assign n24398 = n24397 ^ n24310;
  assign n24308 = n24056 ^ n839;
  assign n24399 = n24398 ^ n24308;
  assign n24400 = n23769 ^ n23179;
  assign n24401 = n24400 ^ n22542;
  assign n24402 = n24401 ^ n24308;
  assign n24403 = ~n24399 & ~n24402;
  assign n24404 = n24403 ^ n24401;
  assign n24405 = n24404 ^ n24306;
  assign n24406 = ~n24307 & ~n24405;
  assign n24407 = n24406 ^ n24304;
  assign n24299 = n23760 ^ n23259;
  assign n24300 = n24299 ^ n22379;
  assign n24486 = n24407 ^ n24300;
  assign n24301 = n24062 ^ n24049;
  assign n24487 = n24486 ^ n24301;
  assign n24488 = n24487 ^ n21881;
  assign n24489 = n24404 ^ n24307;
  assign n24490 = n24489 ^ n21456;
  assign n24491 = n24401 ^ n24399;
  assign n24492 = n24491 ^ n21458;
  assign n24493 = n24395 ^ n24310;
  assign n24494 = n24493 ^ n23738;
  assign n24495 = n24494 ^ n21868;
  assign n24496 = n24392 ^ n24316;
  assign n24497 = n24496 ^ n21466;
  assign n24498 = n24389 ^ n24319;
  assign n24499 = n24498 ^ n21468;
  assign n24500 = n24386 ^ n24321;
  assign n24501 = n24500 ^ n24252;
  assign n24502 = n24501 ^ n21469;
  assign n24503 = n24383 ^ n24326;
  assign n24504 = n24503 ^ n21477;
  assign n24505 = n24380 ^ n24330;
  assign n24506 = n24505 ^ n21846;
  assign n24509 = n24368 ^ n24365;
  assign n24510 = n24509 ^ n21826;
  assign n24237 = n24236 ^ n24211;
  assign n24511 = n24237 ^ n21490;
  assign n24183 = n24182 ^ n24158;
  assign n24184 = n24183 ^ n21492;
  assign n24126 = n21493 & n24125;
  assign n24127 = n24126 ^ n21810;
  assign n24153 = n24152 ^ n24148;
  assign n24154 = n24153 ^ n24126;
  assign n24155 = n24127 & ~n24154;
  assign n24156 = n24155 ^ n21810;
  assign n24206 = n24183 ^ n24156;
  assign n24207 = n24184 & n24206;
  assign n24208 = n24207 ^ n21492;
  assign n24512 = n24237 ^ n24208;
  assign n24513 = ~n24511 & n24512;
  assign n24514 = n24513 ^ n21490;
  assign n24515 = n24514 ^ n24509;
  assign n24516 = ~n24510 & ~n24515;
  assign n24517 = n24516 ^ n21826;
  assign n24508 = n24371 ^ n24342;
  assign n24518 = n24517 ^ n24508;
  assign n24519 = n24517 ^ n21486;
  assign n24520 = n24518 & ~n24519;
  assign n24521 = n24520 ^ n21486;
  assign n24522 = n24521 ^ n21836;
  assign n24523 = n24374 ^ n24336;
  assign n24524 = n24523 ^ n24337;
  assign n24525 = n24524 ^ n24521;
  assign n24526 = n24522 & ~n24525;
  assign n24527 = n24526 ^ n21836;
  assign n24507 = n24377 ^ n24334;
  assign n24528 = n24527 ^ n24507;
  assign n24529 = n24507 ^ n21482;
  assign n24530 = ~n24528 & ~n24529;
  assign n24531 = n24530 ^ n21482;
  assign n24532 = n24531 ^ n24505;
  assign n24533 = ~n24506 & n24532;
  assign n24534 = n24533 ^ n21846;
  assign n24535 = n24534 ^ n24503;
  assign n24536 = n24504 & n24535;
  assign n24537 = n24536 ^ n21477;
  assign n24538 = n24537 ^ n24501;
  assign n24539 = n24502 & n24538;
  assign n24540 = n24539 ^ n21469;
  assign n24541 = n24540 ^ n24498;
  assign n24542 = ~n24499 & n24541;
  assign n24543 = n24542 ^ n21468;
  assign n24544 = n24543 ^ n24496;
  assign n24545 = ~n24497 & ~n24544;
  assign n24546 = n24545 ^ n21466;
  assign n24547 = n24546 ^ n24494;
  assign n24548 = ~n24495 & ~n24547;
  assign n24549 = n24548 ^ n21868;
  assign n24550 = n24549 ^ n24491;
  assign n24551 = ~n24492 & ~n24550;
  assign n24552 = n24551 ^ n21458;
  assign n24553 = n24552 ^ n24489;
  assign n24554 = n24490 & ~n24553;
  assign n24555 = n24554 ^ n21456;
  assign n24556 = n24555 ^ n24487;
  assign n24557 = ~n24488 & ~n24556;
  assign n24558 = n24557 ^ n21881;
  assign n24302 = n24301 ^ n24300;
  assign n24408 = n24407 ^ n24301;
  assign n24409 = n24302 & n24408;
  assign n24410 = n24409 ^ n24300;
  assign n24296 = n24065 ^ n1095;
  assign n24297 = n24296 ^ n24046;
  assign n24294 = n23756 ^ n23171;
  assign n24295 = n24294 ^ n22375;
  assign n24298 = n24297 ^ n24295;
  assign n24485 = n24410 ^ n24298;
  assign n24559 = n24558 ^ n24485;
  assign n24643 = n24559 ^ n21890;
  assign n24612 = n24549 ^ n24492;
  assign n24613 = n24534 ^ n21477;
  assign n24614 = n24613 ^ n24503;
  assign n24615 = n24514 ^ n24510;
  assign n24209 = n24208 ^ n21490;
  assign n24238 = n24237 ^ n24209;
  assign n24185 = n24184 ^ n24156;
  assign n24187 = n24153 ^ n24127;
  assign n24188 = n24186 & n24187;
  assign n24239 = n24185 & n24188;
  assign n24616 = n24238 & n24239;
  assign n24617 = n24615 & n24616;
  assign n24618 = n24518 ^ n21486;
  assign n24619 = ~n24617 & ~n24618;
  assign n24620 = n24524 ^ n21836;
  assign n24621 = n24620 ^ n24521;
  assign n24622 = ~n24619 & ~n24621;
  assign n24623 = n24528 ^ n21482;
  assign n24624 = ~n24622 & ~n24623;
  assign n24625 = n24531 ^ n24506;
  assign n24626 = n24624 & n24625;
  assign n24627 = ~n24614 & n24626;
  assign n24628 = n24537 ^ n21469;
  assign n24629 = n24628 ^ n24501;
  assign n24630 = ~n24627 & ~n24629;
  assign n24631 = n24540 ^ n24499;
  assign n24632 = ~n24630 & n24631;
  assign n24633 = n24543 ^ n21466;
  assign n24634 = n24633 ^ n24496;
  assign n24635 = ~n24632 & ~n24634;
  assign n24636 = n24546 ^ n24495;
  assign n24637 = ~n24635 & ~n24636;
  assign n24638 = n24612 & n24637;
  assign n24639 = n24552 ^ n24490;
  assign n24640 = n24638 & n24639;
  assign n24641 = n24555 ^ n24488;
  assign n24642 = n24640 & ~n24641;
  assign n24720 = n24643 ^ n24642;
  assign n2507 = n2500 ^ n2482;
  assign n2514 = n2513 ^ n2507;
  assign n2518 = n2517 ^ n2514;
  assign n24721 = n24720 ^ n2518;
  assign n24723 = n24639 ^ n24638;
  assign n24724 = n24723 ^ n1408;
  assign n24725 = n24637 ^ n24612;
  assign n1391 = n1381 ^ n1288;
  assign n1392 = n1391 ^ n1215;
  assign n1396 = n1395 ^ n1392;
  assign n24726 = n24725 ^ n1396;
  assign n24727 = n24636 ^ n24635;
  assign n1203 = n1187 ^ n1115;
  assign n1204 = n1203 ^ n1200;
  assign n1208 = n1207 ^ n1204;
  assign n24728 = n24727 ^ n1208;
  assign n24730 = n24631 ^ n24630;
  assign n1054 = n1020 ^ n974;
  assign n1055 = n1054 ^ n1051;
  assign n1059 = n1058 ^ n1055;
  assign n24731 = n24730 ^ n1059;
  assign n24732 = n24629 ^ n24627;
  assign n24733 = n24732 ^ n1047;
  assign n24734 = n24626 ^ n24614;
  assign n24735 = n24734 ^ n3319;
  assign n24739 = n22856 ^ n15958;
  assign n24740 = n24739 ^ n644;
  assign n24741 = n24740 ^ n585;
  assign n24738 = n24621 ^ n24619;
  assign n24742 = n24741 ^ n24738;
  assign n24743 = n24618 ^ n24617;
  assign n552 = n551 ^ n548;
  assign n559 = n558 ^ n552;
  assign n563 = n562 ^ n559;
  assign n24744 = n24743 ^ n563;
  assign n24745 = n24616 ^ n24615;
  assign n24749 = n24748 ^ n24745;
  assign n24241 = n22327 ^ n534;
  assign n24242 = n24241 ^ n19663;
  assign n24243 = n24242 ^ n3245;
  assign n24240 = n24239 ^ n24238;
  assign n24244 = n24243 ^ n24240;
  assign n24191 = n15939 ^ n2343;
  assign n24192 = n24191 ^ n2297;
  assign n24193 = n24192 ^ n14474;
  assign n24190 = n2287 & ~n24186;
  assign n24194 = n24193 ^ n24190;
  assign n24195 = n24187 ^ n24186;
  assign n24196 = n24195 ^ n24190;
  assign n24197 = n24194 & ~n24196;
  assign n24198 = n24197 ^ n24193;
  assign n24189 = n24188 ^ n24185;
  assign n24199 = n24198 ^ n24189;
  assign n24203 = n24202 ^ n24198;
  assign n24204 = ~n24199 & n24203;
  assign n24205 = n24204 ^ n24202;
  assign n24750 = n24240 ^ n24205;
  assign n24751 = n24244 & ~n24750;
  assign n24752 = n24751 ^ n24243;
  assign n24753 = n24752 ^ n24745;
  assign n24754 = n24749 & ~n24753;
  assign n24755 = n24754 ^ n24748;
  assign n24756 = n24755 ^ n24743;
  assign n24757 = ~n24744 & n24756;
  assign n24758 = n24757 ^ n563;
  assign n24759 = n24758 ^ n24738;
  assign n24760 = n24742 & ~n24759;
  assign n24761 = n24760 ^ n24741;
  assign n24737 = n24623 ^ n24622;
  assign n24762 = n24761 ^ n24737;
  assign n24763 = n24737 ^ n729;
  assign n24764 = n24762 & ~n24763;
  assign n24765 = n24764 ^ n729;
  assign n24736 = n24625 ^ n24624;
  assign n24766 = n24765 ^ n24736;
  assign n24770 = n24769 ^ n24736;
  assign n24771 = n24766 & ~n24770;
  assign n24772 = n24771 ^ n24769;
  assign n24773 = n24772 ^ n24734;
  assign n24774 = n24735 & ~n24773;
  assign n24775 = n24774 ^ n3319;
  assign n24776 = n24775 ^ n24732;
  assign n24777 = n24733 & ~n24776;
  assign n24778 = n24777 ^ n1047;
  assign n24779 = n24778 ^ n24730;
  assign n24780 = n24731 & ~n24779;
  assign n24781 = n24780 ^ n1059;
  assign n24729 = n24634 ^ n24632;
  assign n24782 = n24781 ^ n24729;
  assign n1072 = n1032 ^ n993;
  assign n1073 = n1072 ^ n1066;
  assign n1077 = n1076 ^ n1073;
  assign n24783 = n24729 ^ n1077;
  assign n24784 = ~n24782 & n24783;
  assign n24785 = n24784 ^ n1077;
  assign n24786 = n24785 ^ n24727;
  assign n24787 = ~n24728 & n24786;
  assign n24788 = n24787 ^ n1208;
  assign n24789 = n24788 ^ n24725;
  assign n24790 = ~n24726 & n24789;
  assign n24791 = n24790 ^ n1396;
  assign n24792 = n24791 ^ n24723;
  assign n24793 = ~n24724 & n24792;
  assign n24794 = n24793 ^ n1408;
  assign n24722 = n24641 ^ n24640;
  assign n24795 = n24794 ^ n24722;
  assign n3148 = n3144 ^ n2447;
  assign n3152 = n3151 ^ n3148;
  assign n3153 = n3152 ^ n2510;
  assign n24796 = n24722 ^ n3153;
  assign n24797 = ~n24795 & n24796;
  assign n24798 = n24797 ^ n3153;
  assign n24799 = n24798 ^ n24720;
  assign n24800 = ~n24721 & n24799;
  assign n24801 = n24800 ^ n2518;
  assign n24560 = n24485 ^ n21890;
  assign n24561 = ~n24559 & n24560;
  assign n24562 = n24561 ^ n21890;
  assign n24411 = n24410 ^ n24297;
  assign n24412 = n24298 & n24411;
  assign n24413 = n24412 ^ n24295;
  assign n24291 = n23751 ^ n22371;
  assign n24292 = n24291 ^ n23270;
  assign n24290 = n24072 ^ n24069;
  assign n24293 = n24292 ^ n24290;
  assign n24484 = n24413 ^ n24293;
  assign n24563 = n24562 ^ n24484;
  assign n24645 = n24563 ^ n22017;
  assign n24644 = ~n24642 & n24643;
  assign n24718 = n24645 ^ n24644;
  assign n2525 = n2465 ^ n1553;
  assign n2526 = n2525 ^ n2522;
  assign n2530 = n2529 ^ n2526;
  assign n24719 = n24718 ^ n2530;
  assign n25162 = n24801 ^ n24719;
  assign n24263 = n24105 ^ n1538;
  assign n24264 = n24263 ^ n24103;
  assign n25160 = n24264 ^ n24218;
  assign n25161 = n25160 ^ n23396;
  assign n25163 = n25162 ^ n25161;
  assign n24455 = n24100 ^ n24029;
  assign n25164 = n24455 ^ n23287;
  assign n25165 = n25164 ^ n24166;
  assign n25084 = n24798 ^ n2518;
  assign n25085 = n25084 ^ n24720;
  assign n25166 = n25165 ^ n25085;
  assign n24270 = n24097 ^ n24031;
  assign n25167 = n24270 ^ n23159;
  assign n25168 = n25167 ^ n24141;
  assign n25089 = n24795 ^ n3153;
  assign n25169 = n25168 ^ n25089;
  assign n24442 = n24091 ^ n24035;
  assign n25170 = n24442 ^ n23866;
  assign n25171 = n25170 ^ n23165;
  assign n25099 = n24788 ^ n24726;
  assign n25172 = n25171 ^ n25099;
  assign n24434 = n24088 ^ n3058;
  assign n24435 = n24434 ^ n24036;
  assign n25173 = n24435 ^ n23742;
  assign n25174 = n25173 ^ n23270;
  assign n25103 = n24785 ^ n1208;
  assign n25104 = n25103 ^ n24727;
  assign n25175 = n25174 ^ n25104;
  assign n25178 = n24775 ^ n24733;
  assign n24420 = n24078 ^ n2424;
  assign n24421 = n24420 ^ n24042;
  assign n25176 = n24421 ^ n23756;
  assign n25177 = n25176 ^ n23175;
  assign n25179 = n25178 ^ n25177;
  assign n25180 = n23764 ^ n23183;
  assign n25181 = n25180 ^ n24290;
  assign n25127 = n24769 ^ n24766;
  assign n25182 = n25181 ^ n25127;
  assign n25077 = n24762 ^ n729;
  assign n25074 = n24297 ^ n23185;
  assign n25075 = n25074 ^ n23769;
  assign n25183 = n25077 ^ n25075;
  assign n24983 = n23773 ^ n23188;
  assign n24984 = n24983 ^ n24301;
  assign n24982 = n24758 ^ n24742;
  assign n24985 = n24984 ^ n24982;
  assign n24896 = n24752 ^ n24749;
  assign n24894 = n23780 ^ n23194;
  assign n24895 = n24894 ^ n24308;
  assign n24897 = n24896 ^ n24895;
  assign n24245 = n24244 ^ n24205;
  assign n23147 = n23146 ^ n23145;
  assign n23739 = n23738 ^ n23147;
  assign n24246 = n24245 ^ n23739;
  assign n24884 = n24202 ^ n24199;
  assign n24250 = n24195 ^ n24194;
  assign n24248 = n24247 ^ n23205;
  assign n24249 = n24248 ^ n23788;
  assign n24251 = n24250 ^ n24249;
  assign n24253 = n24252 ^ n23791;
  assign n24254 = n24253 ^ n23208;
  assign n24256 = n24255 ^ n24254;
  assign n24844 = n24325 ^ n23210;
  assign n24845 = n24844 ^ n23811;
  assign n24261 = n22951 ^ n22460;
  assign n24262 = n24261 ^ n23591;
  assign n24265 = n24264 ^ n24262;
  assign n24268 = n24267 ^ n22966;
  assign n24269 = n24268 ^ n22284;
  assign n24271 = n24270 ^ n24269;
  assign n24274 = n24094 ^ n24033;
  assign n24272 = n24218 ^ n22252;
  assign n24273 = n24272 ^ n22961;
  assign n24275 = n24274 ^ n24273;
  assign n24278 = n23287 ^ n22354;
  assign n24279 = n24278 ^ n23971;
  assign n24276 = n24085 ^ n2491;
  assign n24277 = n24276 ^ n24038;
  assign n24280 = n24279 ^ n24277;
  assign n24283 = n24082 ^ n24041;
  assign n24281 = n23159 ^ n22357;
  assign n24282 = n24281 ^ n23866;
  assign n24284 = n24283 ^ n24282;
  assign n24287 = n23747 ^ n23165;
  assign n24288 = n24287 ^ n22366;
  assign n24285 = n24075 ^ n1280;
  assign n24286 = n24285 ^ n24043;
  assign n24289 = n24288 ^ n24286;
  assign n24414 = n24413 ^ n24290;
  assign n24415 = n24293 & n24414;
  assign n24416 = n24415 ^ n24292;
  assign n24417 = n24416 ^ n24286;
  assign n24418 = ~n24289 & ~n24417;
  assign n24419 = n24418 ^ n24288;
  assign n24422 = n24421 ^ n24419;
  assign n24423 = n23742 ^ n23163;
  assign n24424 = n24423 ^ n22361;
  assign n24425 = n24424 ^ n24421;
  assign n24426 = ~n24422 & ~n24425;
  assign n24427 = n24426 ^ n24424;
  assign n24428 = n24427 ^ n24283;
  assign n24429 = ~n24284 & ~n24428;
  assign n24430 = n24429 ^ n24282;
  assign n24431 = n24430 ^ n24277;
  assign n24432 = n24280 & ~n24431;
  assign n24433 = n24432 ^ n24279;
  assign n24436 = n24435 ^ n24433;
  assign n24437 = n23396 ^ n22352;
  assign n24438 = n24437 ^ n24141;
  assign n24439 = n24438 ^ n24435;
  assign n24440 = n24436 & n24439;
  assign n24441 = n24440 ^ n24438;
  assign n24443 = n24442 ^ n24441;
  assign n24444 = n24166 ^ n22347;
  assign n24445 = n24444 ^ n23449;
  assign n24446 = n24445 ^ n24442;
  assign n24447 = ~n24443 & ~n24446;
  assign n24448 = n24447 ^ n24445;
  assign n24449 = n24448 ^ n24274;
  assign n24450 = n24275 & ~n24449;
  assign n24451 = n24450 ^ n24273;
  assign n24452 = n24451 ^ n24270;
  assign n24453 = n24271 & n24452;
  assign n24454 = n24453 ^ n24269;
  assign n24456 = n24455 ^ n24454;
  assign n24457 = n23584 ^ n22957;
  assign n24458 = n24457 ^ n22316;
  assign n24459 = n24458 ^ n24455;
  assign n24460 = ~n24456 & n24459;
  assign n24461 = n24460 ^ n24458;
  assign n24462 = n24461 ^ n24264;
  assign n24463 = n24265 & ~n24462;
  assign n24464 = n24463 ^ n24262;
  assign n24259 = n24108 ^ n24027;
  assign n24257 = n23582 ^ n22949;
  assign n24258 = n24257 ^ n22453;
  assign n24260 = n24259 ^ n24258;
  assign n24465 = n24464 ^ n24260;
  assign n24671 = n24465 ^ n21759;
  assign n24466 = n24461 ^ n24265;
  assign n24467 = n24466 ^ n21760;
  assign n24468 = n24458 ^ n24456;
  assign n24469 = n24468 ^ n21761;
  assign n24470 = n24451 ^ n24271;
  assign n24471 = n24470 ^ n21769;
  assign n24472 = n24448 ^ n24275;
  assign n24473 = n24472 ^ n21762;
  assign n24474 = n24445 ^ n24443;
  assign n24475 = n24474 ^ n22364;
  assign n24476 = n24438 ^ n24436;
  assign n24477 = n24476 ^ n22369;
  assign n24482 = n24416 ^ n24289;
  assign n24483 = n24482 ^ n22077;
  assign n24564 = n24484 ^ n22017;
  assign n24565 = n24563 & n24564;
  assign n24566 = n24565 ^ n22017;
  assign n24567 = n24566 ^ n24482;
  assign n24568 = n24483 & ~n24567;
  assign n24569 = n24568 ^ n22077;
  assign n24481 = n24424 ^ n24422;
  assign n24570 = n24569 ^ n24481;
  assign n24571 = n24481 ^ n22237;
  assign n24572 = n24570 & ~n24571;
  assign n24573 = n24572 ^ n22237;
  assign n24480 = n24427 ^ n24284;
  assign n24574 = n24573 ^ n24480;
  assign n24575 = n24480 ^ n22266;
  assign n24576 = ~n24574 & ~n24575;
  assign n24577 = n24576 ^ n22266;
  assign n24478 = n24430 ^ n24279;
  assign n24479 = n24478 ^ n24277;
  assign n24578 = n24577 ^ n24479;
  assign n24579 = n24479 ^ n22298;
  assign n24580 = n24578 & n24579;
  assign n24581 = n24580 ^ n22298;
  assign n24582 = n24581 ^ n24476;
  assign n24583 = ~n24477 & ~n24582;
  assign n24584 = n24583 ^ n22369;
  assign n24585 = n24584 ^ n24474;
  assign n24586 = ~n24475 & n24585;
  assign n24587 = n24586 ^ n22364;
  assign n24588 = n24587 ^ n24472;
  assign n24589 = ~n24473 & n24588;
  assign n24590 = n24589 ^ n21762;
  assign n24591 = n24590 ^ n24470;
  assign n24592 = ~n24471 & n24591;
  assign n24593 = n24592 ^ n21769;
  assign n24594 = n24593 ^ n24468;
  assign n24595 = ~n24469 & ~n24594;
  assign n24596 = n24595 ^ n21761;
  assign n24597 = n24596 ^ n24466;
  assign n24598 = n24467 & n24597;
  assign n24599 = n24598 ^ n21760;
  assign n24672 = n24599 ^ n24465;
  assign n24673 = ~n24671 & ~n24672;
  assign n24674 = n24673 ^ n21759;
  assign n24665 = n24464 ^ n24258;
  assign n24666 = n24260 & ~n24665;
  assign n24667 = n24666 ^ n24259;
  assign n24663 = n24111 ^ n1628;
  assign n24664 = n24663 ^ n24021;
  assign n24668 = n24667 ^ n24664;
  assign n24661 = n23576 ^ n22342;
  assign n24662 = n24661 ^ n22413;
  assign n24669 = n24668 ^ n24662;
  assign n24670 = n24669 ^ n21494;
  assign n24675 = n24674 ^ n24670;
  assign n24600 = n24599 ^ n21759;
  assign n24601 = n24600 ^ n24465;
  assign n24602 = n24596 ^ n24467;
  assign n24603 = n24593 ^ n21761;
  assign n24604 = n24603 ^ n24468;
  assign n24605 = n24590 ^ n21769;
  assign n24606 = n24605 ^ n24470;
  assign n24607 = n24584 ^ n24475;
  assign n24608 = n24581 ^ n24477;
  assign n24609 = n24574 ^ n22266;
  assign n24610 = n24566 ^ n22077;
  assign n24611 = n24610 ^ n24482;
  assign n24646 = n24644 & n24645;
  assign n24647 = n24611 & ~n24646;
  assign n24648 = n24570 ^ n22237;
  assign n24649 = n24647 & ~n24648;
  assign n24650 = n24609 & ~n24649;
  assign n24651 = n24578 ^ n22298;
  assign n24652 = ~n24650 & ~n24651;
  assign n24653 = ~n24608 & n24652;
  assign n24654 = ~n24607 & ~n24653;
  assign n24655 = n24587 ^ n24473;
  assign n24656 = ~n24654 & n24655;
  assign n24657 = n24606 & n24656;
  assign n24658 = n24604 & n24657;
  assign n24659 = ~n24602 & ~n24658;
  assign n24660 = n24601 & ~n24659;
  assign n24692 = n24675 ^ n24660;
  assign n24693 = n24692 ^ n2266;
  assign n24694 = n24659 ^ n24601;
  assign n24695 = n24694 ^ n1883;
  assign n24696 = n24658 ^ n24602;
  assign n24700 = n24699 ^ n24696;
  assign n24701 = n24657 ^ n24604;
  assign n1753 = n1748 ^ n1729;
  assign n1757 = n1756 ^ n1753;
  assign n1761 = n1760 ^ n1757;
  assign n24702 = n24701 ^ n1761;
  assign n24703 = n24656 ^ n24606;
  assign n24704 = n24703 ^ n1696;
  assign n24705 = n24655 ^ n24654;
  assign n1673 = n1663 ^ n1642;
  assign n1680 = n1679 ^ n1673;
  assign n1684 = n1683 ^ n1680;
  assign n24706 = n24705 ^ n1684;
  assign n24707 = n24653 ^ n24607;
  assign n24708 = n24707 ^ n3001;
  assign n24710 = n24651 ^ n24650;
  assign n24711 = n24710 ^ n2981;
  assign n24712 = n24649 ^ n24609;
  assign n24713 = n24712 ^ n2693;
  assign n24714 = n24648 ^ n24647;
  assign n24715 = n24714 ^ n3086;
  assign n24716 = n24646 ^ n24611;
  assign n2581 = n2576 ^ n2544;
  assign n2585 = n2584 ^ n2581;
  assign n2586 = n2585 ^ n1518;
  assign n24717 = n24716 ^ n2586;
  assign n24802 = n24801 ^ n24718;
  assign n24803 = n24719 & ~n24802;
  assign n24804 = n24803 ^ n2530;
  assign n24805 = n24804 ^ n24716;
  assign n24806 = n24717 & ~n24805;
  assign n24807 = n24806 ^ n2586;
  assign n24808 = n24807 ^ n24714;
  assign n24809 = n24715 & ~n24808;
  assign n24810 = n24809 ^ n3086;
  assign n24811 = n24810 ^ n24712;
  assign n24812 = ~n24713 & n24811;
  assign n24813 = n24812 ^ n2693;
  assign n24814 = n24813 ^ n24710;
  assign n24815 = ~n24711 & n24814;
  assign n24816 = n24815 ^ n2981;
  assign n24709 = n24652 ^ n24608;
  assign n24817 = n24816 ^ n24709;
  assign n24818 = n24709 ^ n2975;
  assign n24819 = ~n24817 & n24818;
  assign n24820 = n24819 ^ n2975;
  assign n24821 = n24820 ^ n24707;
  assign n24822 = n24708 & ~n24821;
  assign n24823 = n24822 ^ n3001;
  assign n24824 = n24823 ^ n24705;
  assign n24825 = n24706 & ~n24824;
  assign n24826 = n24825 ^ n1684;
  assign n24827 = n24826 ^ n24703;
  assign n24828 = ~n24704 & n24827;
  assign n24829 = n24828 ^ n1696;
  assign n24830 = n24829 ^ n1761;
  assign n24831 = ~n24702 & ~n24830;
  assign n24832 = n24831 ^ n24701;
  assign n24833 = n24832 ^ n24696;
  assign n24834 = n24700 & n24833;
  assign n24835 = n24834 ^ n24699;
  assign n24836 = n24835 ^ n24694;
  assign n24837 = n24695 & ~n24836;
  assign n24838 = n24837 ^ n1883;
  assign n24839 = n24838 ^ n24692;
  assign n24840 = n24693 & ~n24839;
  assign n24841 = n24840 ^ n2266;
  assign n2270 = n2165 ^ n2107;
  assign n2271 = n2270 ^ n2042;
  assign n2272 = n2271 ^ n681;
  assign n24842 = n24841 ^ n2272;
  assign n24686 = n24674 ^ n24669;
  assign n24687 = ~n24670 & ~n24686;
  assign n24688 = n24687 ^ n21494;
  assign n24682 = n24664 ^ n24662;
  assign n24683 = n24668 & ~n24682;
  assign n24684 = n24683 ^ n24662;
  assign n24679 = n23574 ^ n22337;
  assign n24680 = n24679 ^ n22411;
  assign n24677 = n24114 ^ n24019;
  assign n24678 = n24677 ^ n24016;
  assign n24681 = n24680 ^ n24678;
  assign n24685 = n24684 ^ n24681;
  assign n24689 = n24688 ^ n24685;
  assign n24690 = n24689 ^ n21797;
  assign n24676 = n24660 & ~n24675;
  assign n24691 = n24690 ^ n24676;
  assign n24843 = n24842 ^ n24691;
  assign n24846 = n24845 ^ n24843;
  assign n24849 = n24327 ^ n23795;
  assign n24850 = n24849 ^ n23130;
  assign n24847 = n24838 ^ n2266;
  assign n24848 = n24847 ^ n24692;
  assign n24851 = n24850 ^ n24848;
  assign n24854 = n24835 ^ n1883;
  assign n24855 = n24854 ^ n24694;
  assign n24852 = n23798 ^ n23043;
  assign n24853 = n24852 ^ n24333;
  assign n24856 = n24855 ^ n24853;
  assign n24861 = n24337 ^ n22990;
  assign n24862 = n24861 ^ n23729;
  assign n24857 = n24829 ^ n24702;
  assign n24858 = n24341 ^ n23668;
  assign n24859 = n24858 ^ n22329;
  assign n24860 = ~n24857 & ~n24859;
  assign n24863 = n24862 ^ n24860;
  assign n24864 = n24832 ^ n24699;
  assign n24865 = n24864 ^ n24696;
  assign n24866 = n24865 ^ n24862;
  assign n24867 = n24863 & n24866;
  assign n24868 = n24867 ^ n24860;
  assign n24869 = n24868 ^ n24855;
  assign n24870 = ~n24856 & ~n24869;
  assign n24871 = n24870 ^ n24853;
  assign n24872 = n24871 ^ n24848;
  assign n24873 = n24851 & n24872;
  assign n24874 = n24873 ^ n24850;
  assign n24875 = n24874 ^ n24845;
  assign n24876 = ~n24846 & n24875;
  assign n24877 = n24876 ^ n24843;
  assign n24878 = n24877 ^ n24254;
  assign n24879 = ~n24256 & ~n24878;
  assign n24880 = n24879 ^ n24255;
  assign n24881 = n24880 ^ n24250;
  assign n24882 = ~n24251 & n24881;
  assign n24883 = n24882 ^ n24249;
  assign n24885 = n24884 ^ n24883;
  assign n24886 = n24315 ^ n23201;
  assign n24887 = n24886 ^ n23787;
  assign n24888 = n24887 ^ n24884;
  assign n24889 = n24885 & n24888;
  assign n24890 = n24889 ^ n24887;
  assign n24891 = n24890 ^ n24245;
  assign n24892 = ~n24246 & ~n24891;
  assign n24893 = n24892 ^ n23739;
  assign n24950 = n24896 ^ n24893;
  assign n24951 = ~n24897 & n24950;
  assign n24952 = n24951 ^ n24895;
  assign n24948 = n24755 ^ n563;
  assign n24949 = n24948 ^ n24743;
  assign n24953 = n24952 ^ n24949;
  assign n24946 = n24306 ^ n23192;
  assign n24947 = n24946 ^ n23775;
  assign n24979 = n24949 ^ n24947;
  assign n24980 = ~n24953 & n24979;
  assign n24981 = n24980 ^ n24947;
  assign n25071 = n24982 ^ n24981;
  assign n25072 = n24985 & n25071;
  assign n25073 = n25072 ^ n24984;
  assign n25184 = n25077 ^ n25073;
  assign n25185 = ~n25183 & n25184;
  assign n25186 = n25185 ^ n25075;
  assign n25187 = n25186 ^ n25127;
  assign n25188 = n25182 & n25187;
  assign n25189 = n25188 ^ n25181;
  assign n25121 = n24772 ^ n3319;
  assign n25122 = n25121 ^ n24734;
  assign n25190 = n25189 ^ n25122;
  assign n25191 = n24286 ^ n23179;
  assign n25192 = n25191 ^ n23760;
  assign n25193 = n25192 ^ n25189;
  assign n25194 = ~n25190 & n25193;
  assign n25195 = n25194 ^ n25122;
  assign n25196 = n25195 ^ n25178;
  assign n25197 = ~n25179 & ~n25196;
  assign n25198 = n25197 ^ n25177;
  assign n25116 = n24778 ^ n24731;
  assign n25199 = n25198 ^ n25116;
  assign n25200 = n24283 ^ n23259;
  assign n25201 = n25200 ^ n23751;
  assign n25202 = n25201 ^ n25116;
  assign n25203 = n25199 & n25202;
  assign n25204 = n25203 ^ n25201;
  assign n25111 = n24782 ^ n1077;
  assign n25205 = n25204 ^ n25111;
  assign n25206 = n24277 ^ n23171;
  assign n25207 = n25206 ^ n23747;
  assign n25208 = n25207 ^ n25111;
  assign n25209 = ~n25205 & ~n25208;
  assign n25210 = n25209 ^ n25207;
  assign n25211 = n25210 ^ n25104;
  assign n25212 = ~n25175 & ~n25211;
  assign n25213 = n25212 ^ n25174;
  assign n25214 = n25213 ^ n25099;
  assign n25215 = n25172 & n25214;
  assign n25216 = n25215 ^ n25171;
  assign n25094 = n24791 ^ n24724;
  assign n25217 = n25216 ^ n25094;
  assign n25218 = n24274 ^ n23971;
  assign n25219 = n25218 ^ n23163;
  assign n25220 = n25219 ^ n25094;
  assign n25221 = ~n25217 & n25220;
  assign n25222 = n25221 ^ n25219;
  assign n25223 = n25222 ^ n25089;
  assign n25224 = n25169 & n25223;
  assign n25225 = n25224 ^ n25168;
  assign n25226 = n25225 ^ n25165;
  assign n25227 = n25166 & n25226;
  assign n25228 = n25227 ^ n25085;
  assign n25229 = n25228 ^ n25162;
  assign n25230 = ~n25163 & n25229;
  assign n25231 = n25230 ^ n25161;
  assign n25155 = n24259 ^ n23449;
  assign n25156 = n25155 ^ n24267;
  assign n25263 = n25231 ^ n25156;
  assign n25157 = n24804 ^ n2586;
  assign n25158 = n25157 ^ n24716;
  assign n25264 = n25263 ^ n25158;
  assign n25265 = n25264 ^ n22347;
  assign n25269 = n25222 ^ n25169;
  assign n25270 = n25269 ^ n22357;
  assign n25271 = n25219 ^ n25217;
  assign n25272 = n25271 ^ n22361;
  assign n25273 = n25213 ^ n25171;
  assign n25274 = n25273 ^ n25099;
  assign n25275 = n25274 ^ n22366;
  assign n25276 = n25210 ^ n25174;
  assign n25277 = n25276 ^ n25104;
  assign n25278 = n25277 ^ n22371;
  assign n25279 = n25207 ^ n25205;
  assign n25280 = n25279 ^ n22375;
  assign n25282 = n25195 ^ n25179;
  assign n25283 = n25282 ^ n22549;
  assign n25284 = n25192 ^ n25122;
  assign n25285 = n25284 ^ n25189;
  assign n25286 = n25285 ^ n22542;
  assign n25287 = n25186 ^ n25182;
  assign n25288 = n25287 ^ n22383;
  assign n25076 = n25075 ^ n25073;
  assign n25078 = n25077 ^ n25076;
  assign n25289 = n25078 ^ n22532;
  assign n24954 = n24953 ^ n24947;
  assign n24955 = n24954 ^ n22388;
  assign n24900 = n24887 ^ n24885;
  assign n24901 = n24900 ^ n22507;
  assign n24903 = n24874 ^ n24846;
  assign n24904 = n24903 ^ n22335;
  assign n24907 = n24868 ^ n24856;
  assign n24908 = n24907 ^ n22345;
  assign n24909 = n24859 ^ n24857;
  assign n24910 = n22476 & n24909;
  assign n24911 = n24910 ^ n22407;
  assign n24912 = n24865 ^ n24863;
  assign n24913 = n24912 ^ n24910;
  assign n24914 = ~n24911 & n24913;
  assign n24915 = n24914 ^ n22407;
  assign n24916 = n24915 ^ n24907;
  assign n24917 = ~n24908 & ~n24916;
  assign n24918 = n24917 ^ n22345;
  assign n24905 = n24871 ^ n24850;
  assign n24906 = n24905 ^ n24848;
  assign n24919 = n24918 ^ n24906;
  assign n24920 = n24906 ^ n22340;
  assign n24921 = n24919 & n24920;
  assign n24922 = n24921 ^ n22340;
  assign n24923 = n24922 ^ n24903;
  assign n24924 = ~n24904 & ~n24923;
  assign n24925 = n24924 ^ n22335;
  assign n24926 = n24925 ^ n22331;
  assign n24927 = n24877 ^ n24256;
  assign n24928 = n24927 ^ n24925;
  assign n24929 = n24926 & n24928;
  assign n24930 = n24929 ^ n22331;
  assign n24902 = n24880 ^ n24251;
  assign n24931 = n24930 ^ n24902;
  assign n24932 = n24902 ^ n22397;
  assign n24933 = ~n24931 & n24932;
  assign n24934 = n24933 ^ n22397;
  assign n24935 = n24934 ^ n24900;
  assign n24936 = n24901 & n24935;
  assign n24937 = n24936 ^ n22507;
  assign n24899 = n24890 ^ n24246;
  assign n24938 = n24937 ^ n24899;
  assign n24939 = n24899 ^ n22391;
  assign n24940 = ~n24938 & n24939;
  assign n24941 = n24940 ^ n22391;
  assign n24898 = n24897 ^ n24893;
  assign n24942 = n24941 ^ n24898;
  assign n24943 = n24898 ^ n22390;
  assign n24944 = n24942 & n24943;
  assign n24945 = n24944 ^ n22390;
  assign n24987 = n24954 ^ n24945;
  assign n24988 = n24955 & n24987;
  assign n24989 = n24988 ^ n22388;
  assign n24986 = n24985 ^ n24981;
  assign n24990 = n24989 ^ n24986;
  assign n25067 = n24986 ^ n22385;
  assign n25068 = ~n24990 & n25067;
  assign n25069 = n25068 ^ n22385;
  assign n25290 = n25078 ^ n25069;
  assign n25291 = ~n25289 & ~n25290;
  assign n25292 = n25291 ^ n22532;
  assign n25293 = n25292 ^ n25287;
  assign n25294 = ~n25288 & ~n25293;
  assign n25295 = n25294 ^ n22383;
  assign n25296 = n25295 ^ n25285;
  assign n25297 = ~n25286 & ~n25296;
  assign n25298 = n25297 ^ n22542;
  assign n25299 = n25298 ^ n25282;
  assign n25300 = n25283 & n25299;
  assign n25301 = n25300 ^ n22549;
  assign n25281 = n25201 ^ n25199;
  assign n25302 = n25301 ^ n25281;
  assign n25303 = n25281 ^ n22379;
  assign n25304 = ~n25302 & n25303;
  assign n25305 = n25304 ^ n22379;
  assign n25306 = n25305 ^ n25279;
  assign n25307 = ~n25280 & ~n25306;
  assign n25308 = n25307 ^ n22375;
  assign n25309 = n25308 ^ n25277;
  assign n25310 = ~n25278 & ~n25309;
  assign n25311 = n25310 ^ n22371;
  assign n25312 = n25311 ^ n25274;
  assign n25313 = n25275 & n25312;
  assign n25314 = n25313 ^ n22366;
  assign n25315 = n25314 ^ n25271;
  assign n25316 = ~n25272 & n25315;
  assign n25317 = n25316 ^ n22361;
  assign n25318 = n25317 ^ n25269;
  assign n25319 = n25270 & n25318;
  assign n25320 = n25319 ^ n22357;
  assign n25268 = n25225 ^ n25166;
  assign n25321 = n25320 ^ n25268;
  assign n25322 = n25268 ^ n22354;
  assign n25323 = n25321 & n25322;
  assign n25324 = n25323 ^ n22354;
  assign n25266 = n25228 ^ n25161;
  assign n25267 = n25266 ^ n25162;
  assign n25325 = n25324 ^ n25267;
  assign n25326 = n25267 ^ n22352;
  assign n25327 = ~n25325 & n25326;
  assign n25328 = n25327 ^ n22352;
  assign n25329 = n25328 ^ n25264;
  assign n25330 = n25265 & ~n25329;
  assign n25331 = n25330 ^ n22347;
  assign n25159 = n25158 ^ n25156;
  assign n25232 = n25231 ^ n25158;
  assign n25233 = ~n25159 & n25232;
  assign n25234 = n25233 ^ n25156;
  assign n25151 = n23584 ^ n22961;
  assign n25152 = n25151 ^ n24664;
  assign n25261 = n25234 ^ n25152;
  assign n25153 = n24807 ^ n24715;
  assign n25262 = n25261 ^ n25153;
  assign n25332 = n25331 ^ n25262;
  assign n25365 = n25332 ^ n22252;
  assign n25366 = n25328 ^ n25265;
  assign n25367 = n25321 ^ n22354;
  assign n25368 = n25317 ^ n25270;
  assign n25369 = n25311 ^ n25275;
  assign n25370 = n25308 ^ n22371;
  assign n25371 = n25370 ^ n25277;
  assign n25372 = n25302 ^ n22379;
  assign n25373 = n25295 ^ n22542;
  assign n25374 = n25373 ^ n25285;
  assign n25375 = n25292 ^ n22383;
  assign n25376 = n25375 ^ n25287;
  assign n24956 = n24955 ^ n24945;
  assign n24957 = n24934 ^ n22507;
  assign n24958 = n24957 ^ n24900;
  assign n24959 = n24927 ^ n24926;
  assign n24960 = n24922 ^ n22335;
  assign n24961 = n24960 ^ n24903;
  assign n24962 = n24919 ^ n22340;
  assign n24963 = n24915 ^ n24908;
  assign n24964 = n24909 ^ n22476;
  assign n24965 = n24912 ^ n24911;
  assign n24966 = n24964 & n24965;
  assign n24967 = n24963 & n24966;
  assign n24968 = n24962 & n24967;
  assign n24969 = n24961 & n24968;
  assign n24970 = n24959 & ~n24969;
  assign n24971 = n24931 ^ n22397;
  assign n24972 = ~n24970 & n24971;
  assign n24973 = ~n24958 & ~n24972;
  assign n24974 = n24938 ^ n22391;
  assign n24975 = n24973 & n24974;
  assign n24976 = n24942 ^ n22390;
  assign n24977 = n24975 & n24976;
  assign n24978 = n24956 & ~n24977;
  assign n24991 = n24990 ^ n22385;
  assign n25066 = ~n24978 & n24991;
  assign n25070 = n25069 ^ n22532;
  assign n25079 = n25078 ^ n25070;
  assign n25377 = ~n25066 & n25079;
  assign n25378 = n25376 & ~n25377;
  assign n25379 = ~n25374 & n25378;
  assign n25380 = n25298 ^ n22549;
  assign n25381 = n25380 ^ n25282;
  assign n25382 = n25379 & ~n25381;
  assign n25383 = n25372 & n25382;
  assign n25384 = n25305 ^ n22375;
  assign n25385 = n25384 ^ n25279;
  assign n25386 = ~n25383 & n25385;
  assign n25387 = ~n25371 & n25386;
  assign n25388 = n25369 & ~n25387;
  assign n25389 = n25314 ^ n25272;
  assign n25390 = n25388 & n25389;
  assign n25391 = n25368 & ~n25390;
  assign n25392 = n25367 & ~n25391;
  assign n25393 = n25325 ^ n22352;
  assign n25394 = n25392 & ~n25393;
  assign n25395 = n25366 & ~n25394;
  assign n25396 = ~n25365 & ~n25395;
  assign n25154 = n25153 ^ n25152;
  assign n25235 = n25234 ^ n25153;
  assign n25236 = n25154 & n25235;
  assign n25237 = n25236 ^ n25152;
  assign n25148 = n24678 ^ n23591;
  assign n25149 = n25148 ^ n22966;
  assign n25336 = n25237 ^ n25149;
  assign n25147 = n24810 ^ n24713;
  assign n25337 = n25336 ^ n25147;
  assign n25333 = n25262 ^ n22252;
  assign n25334 = n25332 & n25333;
  assign n25335 = n25334 ^ n22252;
  assign n25338 = n25337 ^ n25335;
  assign n25364 = n25338 ^ n22284;
  assign n25424 = n25396 ^ n25364;
  assign n25428 = n25427 ^ n25424;
  assign n25429 = n25395 ^ n25365;
  assign n25433 = n25432 ^ n25429;
  assign n25437 = n25389 ^ n25388;
  assign n2667 = n2601 ^ n1521;
  assign n2668 = n2667 ^ n2664;
  assign n2672 = n2671 ^ n2668;
  assign n25438 = n25437 ^ n2672;
  assign n25441 = n25385 ^ n25383;
  assign n25445 = n25444 ^ n25441;
  assign n25447 = n3161 ^ n1435;
  assign n25448 = n25447 ^ n2414;
  assign n25449 = n25448 ^ n3026;
  assign n25446 = n25382 ^ n25372;
  assign n25450 = n25449 ^ n25446;
  assign n25451 = n25381 ^ n25379;
  assign n3015 = n3014 ^ n1419;
  assign n3016 = n3015 ^ n1370;
  assign n3017 = n3016 ^ n2412;
  assign n25452 = n25451 ^ n3017;
  assign n25453 = n25378 ^ n25374;
  assign n1358 = n1315 ^ n1252;
  assign n1359 = n1358 ^ n1352;
  assign n1360 = n1359 ^ n1268;
  assign n25454 = n25453 ^ n1360;
  assign n25455 = n25377 ^ n25376;
  assign n1340 = n1166 ^ n1085;
  assign n1341 = n1340 ^ n1237;
  assign n1345 = n1344 ^ n1341;
  assign n25456 = n25455 ^ n1345;
  assign n25080 = n25079 ^ n25066;
  assign n1331 = n1228 ^ n1135;
  assign n1335 = n1334 ^ n1331;
  assign n1336 = n1335 ^ n1083;
  assign n25081 = n25080 ^ n1336;
  assign n24994 = n24976 ^ n24975;
  assign n24995 = n24994 ^ n807;
  assign n24996 = n24974 ^ n24973;
  assign n24997 = n24996 ^ n668;
  assign n24998 = n24972 ^ n24958;
  assign n616 = n612 ^ n600;
  assign n623 = n622 ^ n616;
  assign n627 = n626 ^ n623;
  assign n24999 = n24998 ^ n627;
  assign n25001 = n24969 ^ n24959;
  assign n25005 = n25004 ^ n25001;
  assign n25008 = n23097 ^ n16649;
  assign n25009 = n25008 ^ n20279;
  assign n25010 = n25009 ^ n675;
  assign n25007 = n24967 ^ n24962;
  assign n25011 = n25010 ^ n25007;
  assign n25012 = n24966 ^ n24963;
  assign n25016 = n25015 ^ n25012;
  assign n25020 = ~n24964 & n25019;
  assign n2328 = n2327 ^ n2228;
  assign n2329 = n2328 ^ n2321;
  assign n2330 = n2329 ^ n521;
  assign n25021 = n25020 ^ n2330;
  assign n25022 = n24965 ^ n24964;
  assign n25023 = n25022 ^ n2330;
  assign n25024 = n25021 & ~n25023;
  assign n25025 = n25024 ^ n25020;
  assign n25026 = n25025 ^ n25012;
  assign n25027 = n25016 & ~n25026;
  assign n25028 = n25027 ^ n25015;
  assign n25029 = n25028 ^ n25007;
  assign n25030 = n25011 & ~n25029;
  assign n25031 = n25030 ^ n25010;
  assign n25006 = n24968 ^ n24961;
  assign n25032 = n25031 ^ n25006;
  assign n25036 = n25035 ^ n25031;
  assign n25037 = ~n25032 & n25036;
  assign n25038 = n25037 ^ n25035;
  assign n25039 = n25038 ^ n25001;
  assign n25040 = n25005 & ~n25039;
  assign n25041 = n25040 ^ n25004;
  assign n25000 = n24971 ^ n24970;
  assign n25042 = n25041 ^ n25000;
  assign n25043 = n25041 ^ n3290;
  assign n25044 = n25042 & n25043;
  assign n25045 = n25044 ^ n3290;
  assign n25046 = n25045 ^ n24998;
  assign n25047 = ~n24999 & n25046;
  assign n25048 = n25047 ^ n627;
  assign n25049 = n25048 ^ n24996;
  assign n25050 = ~n24997 & n25049;
  assign n25051 = n25050 ^ n668;
  assign n25052 = n25051 ^ n24994;
  assign n25053 = ~n24995 & n25052;
  assign n25054 = n25053 ^ n807;
  assign n24993 = n24977 ^ n24956;
  assign n25055 = n25054 ^ n24993;
  assign n25059 = n25058 ^ n24993;
  assign n25060 = n25055 & ~n25059;
  assign n25061 = n25060 ^ n25058;
  assign n24992 = n24991 ^ n24978;
  assign n25062 = n25061 ^ n24992;
  assign n25063 = n24992 ^ n929;
  assign n25064 = ~n25062 & n25063;
  assign n25065 = n25064 ^ n929;
  assign n25457 = n25080 ^ n25065;
  assign n25458 = ~n25081 & n25457;
  assign n25459 = n25458 ^ n1336;
  assign n25460 = n25459 ^ n25455;
  assign n25461 = n25456 & ~n25460;
  assign n25462 = n25461 ^ n1345;
  assign n25463 = n25462 ^ n25453;
  assign n25464 = n25454 & ~n25463;
  assign n25465 = n25464 ^ n1360;
  assign n25466 = n25465 ^ n25451;
  assign n25467 = n25452 & ~n25466;
  assign n25468 = n25467 ^ n3017;
  assign n25469 = n25468 ^ n25446;
  assign n25470 = ~n25450 & n25469;
  assign n25471 = n25470 ^ n25449;
  assign n25472 = n25471 ^ n25441;
  assign n25473 = ~n25445 & n25472;
  assign n25474 = n25473 ^ n25444;
  assign n25440 = n25386 ^ n25371;
  assign n25475 = n25474 ^ n25440;
  assign n3182 = n3175 ^ n2559;
  assign n3186 = n3185 ^ n3182;
  assign n3187 = n3186 ^ n2654;
  assign n25476 = n25440 ^ n3187;
  assign n25477 = n25475 & ~n25476;
  assign n25478 = n25477 ^ n3187;
  assign n25439 = n25387 ^ n25369;
  assign n25479 = n25478 ^ n25439;
  assign n25480 = n25439 ^ n2660;
  assign n25481 = ~n25479 & n25480;
  assign n25482 = n25481 ^ n2660;
  assign n25483 = n25482 ^ n25437;
  assign n25484 = ~n25438 & n25483;
  assign n25485 = n25484 ^ n2672;
  assign n2756 = n2741 ^ n2698;
  assign n2757 = n2756 ^ n2679;
  assign n2758 = n2757 ^ n1493;
  assign n25486 = n25485 ^ n2758;
  assign n25487 = n25390 ^ n25368;
  assign n25488 = n25487 ^ n25485;
  assign n25489 = n25486 & n25488;
  assign n25490 = n25489 ^ n2758;
  assign n25436 = n25391 ^ n25367;
  assign n25491 = n25490 ^ n25436;
  assign n25492 = n25436 ^ n1583;
  assign n25493 = ~n25491 & n25492;
  assign n25494 = n25493 ^ n1583;
  assign n25435 = n25393 ^ n25392;
  assign n25495 = n25494 ^ n25435;
  assign n25496 = n25435 ^ n2883;
  assign n25497 = ~n25495 & n25496;
  assign n25498 = n25497 ^ n2883;
  assign n25434 = n25394 ^ n25366;
  assign n25499 = n25498 ^ n25434;
  assign n25503 = n25502 ^ n25434;
  assign n25504 = n25499 & ~n25503;
  assign n25505 = n25504 ^ n25502;
  assign n25506 = n25505 ^ n25429;
  assign n25507 = ~n25433 & n25506;
  assign n25508 = n25507 ^ n25432;
  assign n25509 = n25508 ^ n25424;
  assign n25510 = n25428 & ~n25509;
  assign n25511 = n25510 ^ n25427;
  assign n25536 = n25511 ^ n1849;
  assign n25397 = ~n25364 & n25396;
  assign n25339 = n25337 ^ n22284;
  assign n25340 = n25338 & ~n25339;
  assign n25341 = n25340 ^ n22284;
  assign n25150 = n25149 ^ n25147;
  assign n25238 = n25237 ^ n25147;
  assign n25239 = n25150 & n25238;
  assign n25240 = n25239 ^ n25149;
  assign n25144 = n23582 ^ n22957;
  assign n25145 = n25144 ^ n24122;
  assign n25142 = n24813 ^ n2981;
  assign n25143 = n25142 ^ n24710;
  assign n25146 = n25145 ^ n25143;
  assign n25259 = n25240 ^ n25146;
  assign n25260 = n25259 ^ n22316;
  assign n25363 = n25341 ^ n25260;
  assign n25422 = n25397 ^ n25363;
  assign n25537 = n25536 ^ n25422;
  assign n25642 = n25539 ^ n25537;
  assign n25718 = n25642 ^ n22329;
  assign n25770 = n2242 & n25718;
  assign n25774 = n25773 ^ n25770;
  assign n25423 = n25422 ^ n1849;
  assign n25512 = n25511 ^ n25422;
  assign n25513 = ~n25423 & n25512;
  assign n25514 = n25513 ^ n1849;
  assign n25398 = n25363 & n25397;
  assign n25342 = n25341 ^ n25259;
  assign n25343 = n25260 & ~n25342;
  assign n25344 = n25343 ^ n22316;
  assign n25246 = n23576 ^ n22951;
  assign n25247 = n25246 ^ n24148;
  assign n25244 = n24817 ^ n2975;
  assign n25241 = n25240 ^ n25145;
  assign n25242 = n25146 & ~n25241;
  assign n25243 = n25242 ^ n25143;
  assign n25245 = n25244 ^ n25243;
  assign n25257 = n25247 ^ n25245;
  assign n25258 = n25257 ^ n22460;
  assign n25362 = n25344 ^ n25258;
  assign n25420 = n25398 ^ n25362;
  assign n25421 = n25420 ^ n1859;
  assign n25544 = n25514 ^ n25421;
  assign n25541 = n24327 ^ n23729;
  assign n25542 = n25541 ^ n24250;
  assign n25540 = ~n25537 & n25539;
  assign n25543 = n25542 ^ n25540;
  assign n25645 = n25544 ^ n25543;
  assign n25643 = n22329 & ~n25642;
  assign n25644 = n25643 ^ n22990;
  assign n25719 = n25645 ^ n25644;
  assign n25775 = n25719 ^ n25718;
  assign n25776 = n25775 ^ n25773;
  assign n25777 = n25774 & ~n25776;
  assign n25778 = n25777 ^ n25770;
  assign n25766 = n2312 ^ n524;
  assign n25767 = n25766 ^ n20856;
  assign n25768 = n25767 ^ n3275;
  assign n25720 = ~n25718 & ~n25719;
  assign n25646 = n25645 ^ n25643;
  assign n25647 = n25644 & n25646;
  assign n25648 = n25647 ^ n22990;
  assign n25545 = n25544 ^ n25542;
  assign n25546 = n25543 & n25545;
  assign n25547 = n25546 ^ n25540;
  assign n25533 = n24884 ^ n24325;
  assign n25534 = n25533 ^ n23798;
  assign n25515 = n25514 ^ n25420;
  assign n25516 = ~n25421 & n25515;
  assign n25517 = n25516 ^ n1859;
  assign n25399 = n25362 & ~n25398;
  assign n25345 = n25344 ^ n25257;
  assign n25346 = ~n25258 & n25345;
  assign n25347 = n25346 ^ n22460;
  assign n25252 = n23574 ^ n22949;
  assign n25253 = n25252 ^ n24178;
  assign n25251 = n24820 ^ n24708;
  assign n25254 = n25253 ^ n25251;
  assign n25248 = n25247 ^ n25244;
  assign n25249 = n25245 & ~n25248;
  assign n25250 = n25249 ^ n25247;
  assign n25255 = n25254 ^ n25250;
  assign n25256 = n25255 ^ n22453;
  assign n25361 = n25347 ^ n25256;
  assign n25418 = n25399 ^ n25361;
  assign n1974 = n1946 ^ n1891;
  assign n1975 = n1974 ^ n1866;
  assign n1976 = n1975 ^ n1964;
  assign n25419 = n25418 ^ n1976;
  assign n25532 = n25517 ^ n25419;
  assign n25535 = n25534 ^ n25532;
  assign n25640 = n25547 ^ n25535;
  assign n25641 = n25640 ^ n23043;
  assign n25717 = n25648 ^ n25641;
  assign n25765 = n25720 ^ n25717;
  assign n25769 = n25768 ^ n25765;
  assign n25928 = n25778 ^ n25769;
  assign n2121 = n2120 ^ n2039;
  assign n2125 = n2124 ^ n2121;
  assign n2126 = n2125 ^ n2115;
  assign n2217 = n2216 ^ n2126;
  assign n2221 = n2220 ^ n2217;
  assign n2222 = n2221 ^ n2208;
  assign n25936 = n25718 ^ n2242;
  assign n25134 = n25025 ^ n25015;
  assign n25135 = n25134 ^ n25012;
  assign n26820 = n25936 ^ n25135;
  assign n26821 = n26820 ^ n24884;
  assign n26430 = n24865 ^ n24148;
  assign n26089 = n25508 ^ n25428;
  assign n26431 = n26430 ^ n26089;
  assign n25861 = n25158 ^ n23866;
  assign n25862 = n25861 ^ n24270;
  assign n25860 = n25462 ^ n25454;
  assign n25863 = n25862 ^ n25860;
  assign n25607 = n24274 ^ n23742;
  assign n25608 = n25607 ^ n25162;
  assign n25605 = n25459 ^ n1345;
  assign n25606 = n25605 ^ n25455;
  assign n25609 = n25608 ^ n25606;
  assign n25083 = n24442 ^ n23747;
  assign n25086 = n25085 ^ n25083;
  assign n25082 = n25081 ^ n25065;
  assign n25087 = n25086 ^ n25082;
  assign n25090 = n25089 ^ n23751;
  assign n25091 = n25090 ^ n24435;
  assign n25088 = n25062 ^ n929;
  assign n25092 = n25091 ^ n25088;
  assign n25095 = n25094 ^ n24277;
  assign n25096 = n25095 ^ n23756;
  assign n25093 = n25058 ^ n25055;
  assign n25097 = n25096 ^ n25093;
  assign n25101 = n25051 ^ n24995;
  assign n25098 = n24283 ^ n23760;
  assign n25100 = n25099 ^ n25098;
  assign n25102 = n25101 ^ n25100;
  assign n25107 = n25048 ^ n668;
  assign n25108 = n25107 ^ n24996;
  assign n25105 = n25104 ^ n24421;
  assign n25106 = n25105 ^ n23764;
  assign n25109 = n25108 ^ n25106;
  assign n25113 = n25045 ^ n24999;
  assign n25110 = n24286 ^ n23769;
  assign n25112 = n25111 ^ n25110;
  assign n25114 = n25113 ^ n25112;
  assign n25118 = n25042 ^ n3290;
  assign n25115 = n24290 ^ n23773;
  assign n25117 = n25116 ^ n25115;
  assign n25119 = n25118 ^ n25117;
  assign n25577 = n25038 ^ n25005;
  assign n25124 = n25035 ^ n25032;
  assign n25120 = n24301 ^ n23780;
  assign n25123 = n25122 ^ n25120;
  assign n25125 = n25124 ^ n25123;
  assign n25129 = n25028 ^ n25010;
  assign n25130 = n25129 ^ n25007;
  assign n25126 = n24306 ^ n23145;
  assign n25128 = n25127 ^ n25126;
  assign n25131 = n25130 ^ n25128;
  assign n25132 = n25077 ^ n24308;
  assign n25133 = n25132 ^ n23787;
  assign n25136 = n25135 ^ n25133;
  assign n25139 = n24949 ^ n23791;
  assign n25140 = n25139 ^ n24315;
  assign n25138 = n25019 ^ n24964;
  assign n25141 = n25140 ^ n25138;
  assign n25527 = n24896 ^ n24247;
  assign n25528 = n25527 ^ n23811;
  assign n25518 = n25517 ^ n25418;
  assign n25519 = n25419 & ~n25518;
  assign n25520 = n25519 ^ n1976;
  assign n25400 = n25361 & ~n25399;
  assign n25356 = n25253 ^ n25250;
  assign n25357 = n25254 & n25356;
  assign n25358 = n25357 ^ n25251;
  assign n25353 = n23607 ^ n22342;
  assign n25354 = n25353 ^ n24232;
  assign n25352 = n24823 ^ n24706;
  assign n25355 = n25354 ^ n25352;
  assign n25359 = n25358 ^ n25355;
  assign n25348 = n25347 ^ n25255;
  assign n25349 = n25256 & ~n25348;
  assign n25350 = n25349 ^ n22453;
  assign n25351 = n25350 ^ n22413;
  assign n25360 = n25359 ^ n25351;
  assign n25417 = n25400 ^ n25360;
  assign n25521 = n25520 ^ n25417;
  assign n1960 = n1943 ^ n1903;
  assign n1967 = n1966 ^ n1960;
  assign n1971 = n1970 ^ n1967;
  assign n25522 = n25417 ^ n1971;
  assign n25523 = ~n25521 & n25522;
  assign n25524 = n25523 ^ n1971;
  assign n25410 = n25359 ^ n22413;
  assign n25411 = n25359 ^ n25350;
  assign n25412 = ~n25410 & ~n25411;
  assign n25413 = n25412 ^ n22413;
  assign n25414 = n25413 ^ n22411;
  assign n25407 = n24826 ^ n24704;
  assign n25404 = n25358 ^ n25352;
  assign n25405 = ~n25355 & ~n25404;
  assign n25406 = n25405 ^ n25354;
  assign n25408 = n25407 ^ n25406;
  assign n25402 = n24364 ^ n23638;
  assign n25403 = n25402 ^ n22337;
  assign n25409 = n25408 ^ n25403;
  assign n25415 = n25414 ^ n25409;
  assign n25401 = ~n25360 & n25400;
  assign n25416 = n25415 ^ n25401;
  assign n25525 = n25524 ^ n25416;
  assign n25526 = n25525 ^ n2126;
  assign n25529 = n25528 ^ n25526;
  assign n25548 = n25547 ^ n25532;
  assign n25549 = n25535 & ~n25548;
  assign n25550 = n25549 ^ n25534;
  assign n25530 = n24245 ^ n23795;
  assign n25531 = n25530 ^ n24252;
  assign n25551 = n25550 ^ n25531;
  assign n25552 = n25521 ^ n1971;
  assign n25553 = n25552 ^ n25550;
  assign n25554 = ~n25551 & ~n25553;
  assign n25555 = n25554 ^ n25531;
  assign n25556 = n25555 ^ n25526;
  assign n25557 = ~n25529 & ~n25556;
  assign n25558 = n25557 ^ n25528;
  assign n25559 = n25558 ^ n25140;
  assign n25560 = n25141 & n25559;
  assign n25561 = n25560 ^ n25138;
  assign n25137 = n25022 ^ n25021;
  assign n25562 = n25561 ^ n25137;
  assign n25563 = n23788 ^ n23738;
  assign n25564 = n25563 ^ n24982;
  assign n25565 = n25564 ^ n25137;
  assign n25566 = n25562 & ~n25565;
  assign n25567 = n25566 ^ n25564;
  assign n25568 = n25567 ^ n25135;
  assign n25569 = ~n25136 & n25568;
  assign n25570 = n25569 ^ n25133;
  assign n25571 = n25570 ^ n25130;
  assign n25572 = ~n25131 & n25571;
  assign n25573 = n25572 ^ n25128;
  assign n25574 = n25573 ^ n25124;
  assign n25575 = ~n25125 & n25574;
  assign n25576 = n25575 ^ n25123;
  assign n25578 = n25577 ^ n25576;
  assign n25579 = n25178 ^ n23775;
  assign n25580 = n25579 ^ n24297;
  assign n25581 = n25580 ^ n25577;
  assign n25582 = n25578 & ~n25581;
  assign n25583 = n25582 ^ n25580;
  assign n25584 = n25583 ^ n25118;
  assign n25585 = n25119 & ~n25584;
  assign n25586 = n25585 ^ n25117;
  assign n25587 = n25586 ^ n25113;
  assign n25588 = ~n25114 & ~n25587;
  assign n25589 = n25588 ^ n25112;
  assign n25590 = n25589 ^ n25108;
  assign n25591 = ~n25109 & n25590;
  assign n25592 = n25591 ^ n25106;
  assign n25593 = n25592 ^ n25101;
  assign n25594 = n25102 & n25593;
  assign n25595 = n25594 ^ n25100;
  assign n25596 = n25595 ^ n25093;
  assign n25597 = ~n25097 & ~n25596;
  assign n25598 = n25597 ^ n25096;
  assign n25599 = n25598 ^ n25088;
  assign n25600 = ~n25092 & ~n25599;
  assign n25601 = n25600 ^ n25091;
  assign n25602 = n25601 ^ n25082;
  assign n25603 = ~n25087 & ~n25602;
  assign n25604 = n25603 ^ n25086;
  assign n25857 = n25606 ^ n25604;
  assign n25858 = ~n25609 & ~n25857;
  assign n25859 = n25858 ^ n25608;
  assign n25864 = n25863 ^ n25859;
  assign n25865 = n25864 ^ n23165;
  assign n25612 = n25601 ^ n25087;
  assign n25613 = n25612 ^ n23171;
  assign n25614 = n25598 ^ n25092;
  assign n25615 = n25614 ^ n23259;
  assign n25616 = n25595 ^ n25096;
  assign n25617 = n25616 ^ n25093;
  assign n25618 = n25617 ^ n23175;
  assign n25619 = n25592 ^ n25102;
  assign n25620 = n25619 ^ n23179;
  assign n25621 = n25589 ^ n25109;
  assign n25622 = n25621 ^ n23183;
  assign n25623 = n25586 ^ n25114;
  assign n25624 = n25623 ^ n23185;
  assign n25625 = n25583 ^ n25119;
  assign n25626 = n25625 ^ n23188;
  assign n25628 = n25573 ^ n25125;
  assign n25629 = n25628 ^ n23194;
  assign n25630 = n25567 ^ n25136;
  assign n25631 = n25630 ^ n23201;
  assign n25632 = n25564 ^ n25562;
  assign n25633 = n25632 ^ n23205;
  assign n25634 = n25558 ^ n25141;
  assign n25635 = n25634 ^ n23208;
  assign n25636 = n25555 ^ n25529;
  assign n25637 = n25636 ^ n23210;
  assign n25638 = n25552 ^ n25551;
  assign n25639 = n25638 ^ n23130;
  assign n25649 = n25648 ^ n25640;
  assign n25650 = n25641 & ~n25649;
  assign n25651 = n25650 ^ n23043;
  assign n25652 = n25651 ^ n25638;
  assign n25653 = n25639 & n25652;
  assign n25654 = n25653 ^ n23130;
  assign n25655 = n25654 ^ n25636;
  assign n25656 = n25637 & n25655;
  assign n25657 = n25656 ^ n23210;
  assign n25658 = n25657 ^ n25634;
  assign n25659 = ~n25635 & ~n25658;
  assign n25660 = n25659 ^ n23208;
  assign n25661 = n25660 ^ n25632;
  assign n25662 = ~n25633 & n25661;
  assign n25663 = n25662 ^ n23205;
  assign n25664 = n25663 ^ n25630;
  assign n25665 = n25631 & n25664;
  assign n25666 = n25665 ^ n23201;
  assign n25667 = n25666 ^ n23146;
  assign n25668 = n25570 ^ n25131;
  assign n25669 = n25668 ^ n25666;
  assign n25670 = n25667 & ~n25669;
  assign n25671 = n25670 ^ n23146;
  assign n25672 = n25671 ^ n25628;
  assign n25673 = ~n25629 & ~n25672;
  assign n25674 = n25673 ^ n23194;
  assign n25627 = n25580 ^ n25578;
  assign n25675 = n25674 ^ n25627;
  assign n25676 = n25627 ^ n23192;
  assign n25677 = n25675 & ~n25676;
  assign n25678 = n25677 ^ n23192;
  assign n25679 = n25678 ^ n25625;
  assign n25680 = n25626 & ~n25679;
  assign n25681 = n25680 ^ n23188;
  assign n25682 = n25681 ^ n25623;
  assign n25683 = ~n25624 & n25682;
  assign n25684 = n25683 ^ n23185;
  assign n25685 = n25684 ^ n25621;
  assign n25686 = n25622 & ~n25685;
  assign n25687 = n25686 ^ n23183;
  assign n25688 = n25687 ^ n25619;
  assign n25689 = n25620 & n25688;
  assign n25690 = n25689 ^ n23179;
  assign n25691 = n25690 ^ n25617;
  assign n25692 = n25618 & ~n25691;
  assign n25693 = n25692 ^ n23175;
  assign n25694 = n25693 ^ n25614;
  assign n25695 = n25615 & n25694;
  assign n25696 = n25695 ^ n23259;
  assign n25697 = n25696 ^ n25612;
  assign n25698 = ~n25613 & n25697;
  assign n25699 = n25698 ^ n23171;
  assign n25853 = n25699 ^ n23270;
  assign n25610 = n25609 ^ n25604;
  assign n25854 = n25699 ^ n25610;
  assign n25855 = ~n25853 & ~n25854;
  assign n25856 = n25855 ^ n23270;
  assign n25866 = n25865 ^ n25856;
  assign n25611 = n25610 ^ n23270;
  assign n25700 = n25699 ^ n25611;
  assign n25701 = n25696 ^ n25613;
  assign n25702 = n25687 ^ n23179;
  assign n25703 = n25702 ^ n25619;
  assign n25704 = n25684 ^ n25622;
  assign n25705 = n25681 ^ n25624;
  assign n25706 = n25678 ^ n23188;
  assign n25707 = n25706 ^ n25625;
  assign n25708 = n25675 ^ n23192;
  assign n25709 = n25671 ^ n25629;
  assign n25710 = n25668 ^ n25667;
  assign n25711 = n25663 ^ n25631;
  assign n25712 = n25657 ^ n23208;
  assign n25713 = n25712 ^ n25634;
  assign n25714 = n25654 ^ n25637;
  assign n25715 = n25651 ^ n23130;
  assign n25716 = n25715 ^ n25638;
  assign n25721 = n25717 & n25720;
  assign n25722 = n25716 & n25721;
  assign n25723 = ~n25714 & n25722;
  assign n25724 = n25713 & ~n25723;
  assign n25725 = n25660 ^ n23205;
  assign n25726 = n25725 ^ n25632;
  assign n25727 = ~n25724 & n25726;
  assign n25728 = n25711 & ~n25727;
  assign n25729 = ~n25710 & n25728;
  assign n25730 = n25709 & n25729;
  assign n25731 = n25708 & ~n25730;
  assign n25732 = n25707 & ~n25731;
  assign n25733 = n25705 & ~n25732;
  assign n25734 = n25704 & ~n25733;
  assign n25735 = n25703 & n25734;
  assign n25736 = n25690 ^ n25618;
  assign n25737 = n25735 & ~n25736;
  assign n25738 = n25693 ^ n25615;
  assign n25739 = n25737 & ~n25738;
  assign n25740 = n25701 & ~n25739;
  assign n25867 = n25700 & n25740;
  assign n26074 = ~n25866 & ~n25867;
  assign n26023 = n25864 ^ n25856;
  assign n26024 = n25865 & ~n26023;
  assign n26025 = n26024 ^ n23165;
  assign n25966 = n25860 ^ n25859;
  assign n25967 = ~n25863 & n25966;
  assign n25968 = n25967 ^ n25862;
  assign n25963 = n24455 ^ n23971;
  assign n25964 = n25963 ^ n25153;
  assign n25962 = n25465 ^ n25452;
  assign n25965 = n25964 ^ n25962;
  assign n26021 = n25968 ^ n25965;
  assign n26022 = n26021 ^ n23163;
  assign n26073 = n26025 ^ n26022;
  assign n26131 = n26074 ^ n26073;
  assign n26132 = n26131 ^ n3221;
  assign n25868 = n25867 ^ n25866;
  assign n25869 = n25868 ^ n3065;
  assign n25741 = n25740 ^ n25700;
  assign n2496 = n2495 ^ n2491;
  assign n2503 = n2502 ^ n2496;
  assign n2504 = n2503 ^ n1553;
  assign n25742 = n25741 ^ n2504;
  assign n25744 = n25738 ^ n25737;
  assign n2440 = n2436 ^ n2424;
  assign n2444 = n2443 ^ n2440;
  assign n2448 = n2447 ^ n2444;
  assign n25745 = n25744 ^ n2448;
  assign n25749 = n25729 ^ n25709;
  assign n25750 = n25749 ^ n893;
  assign n25751 = n25727 ^ n25711;
  assign n25755 = n25754 ^ n25751;
  assign n25758 = n25722 ^ n25714;
  assign n700 = n699 ^ n696;
  assign n701 = n700 ^ n536;
  assign n702 = n701 ^ n638;
  assign n25759 = n25758 ^ n702;
  assign n25761 = n23700 ^ n16898;
  assign n25762 = n25761 ^ n20851;
  assign n25763 = n25762 ^ n534;
  assign n25760 = n25721 ^ n25716;
  assign n25764 = n25763 ^ n25760;
  assign n25779 = n25778 ^ n25765;
  assign n25780 = n25769 & ~n25779;
  assign n25781 = n25780 ^ n25768;
  assign n25782 = n25781 ^ n25760;
  assign n25783 = n25764 & ~n25782;
  assign n25784 = n25783 ^ n25763;
  assign n25785 = n25784 ^ n25758;
  assign n25786 = ~n25759 & n25785;
  assign n25787 = n25786 ^ n702;
  assign n25757 = n25723 ^ n25713;
  assign n25788 = n25787 ^ n25757;
  assign n25789 = n23688 ^ n16883;
  assign n25790 = n25789 ^ n20845;
  assign n25791 = n25790 ^ n551;
  assign n25792 = n25791 ^ n25757;
  assign n25793 = ~n25788 & n25792;
  assign n25794 = n25793 ^ n25791;
  assign n25756 = n25726 ^ n25724;
  assign n25795 = n25794 ^ n25756;
  assign n25799 = n25798 ^ n25756;
  assign n25800 = n25795 & ~n25799;
  assign n25801 = n25800 ^ n25798;
  assign n25802 = n25801 ^ n25751;
  assign n25803 = n25755 & ~n25802;
  assign n25804 = n25803 ^ n25754;
  assign n25805 = n25804 ^ n3303;
  assign n25806 = n25728 ^ n25710;
  assign n25807 = n25806 ^ n25804;
  assign n25808 = n25805 & ~n25807;
  assign n25809 = n25808 ^ n3303;
  assign n25810 = n25809 ^ n25749;
  assign n25811 = ~n25750 & n25810;
  assign n25812 = n25811 ^ n893;
  assign n25813 = n25812 ^ n905;
  assign n25814 = n25730 ^ n25708;
  assign n25815 = n25814 ^ n25812;
  assign n25816 = n25813 & n25815;
  assign n25817 = n25816 ^ n905;
  assign n25748 = n25731 ^ n25707;
  assign n25818 = n25817 ^ n25748;
  assign n1016 = n1006 ^ n940;
  assign n1017 = n1016 ^ n912;
  assign n1021 = n1020 ^ n1017;
  assign n25819 = n25748 ^ n1021;
  assign n25820 = ~n25818 & n25819;
  assign n25821 = n25820 ^ n1021;
  assign n1028 = n1012 ^ n949;
  assign n1029 = n1028 ^ n1025;
  assign n1033 = n1032 ^ n1029;
  assign n25822 = n25821 ^ n1033;
  assign n25823 = n25732 ^ n25705;
  assign n25824 = n25823 ^ n25821;
  assign n25825 = n25822 & n25824;
  assign n25826 = n25825 ^ n1033;
  assign n1180 = n1176 ^ n1095;
  assign n1184 = n1183 ^ n1180;
  assign n1188 = n1187 ^ n1184;
  assign n25827 = n25826 ^ n1188;
  assign n25828 = n25733 ^ n25704;
  assign n25829 = n25828 ^ n25826;
  assign n25830 = n25827 & ~n25829;
  assign n25831 = n25830 ^ n1188;
  assign n25747 = n25734 ^ n25703;
  assign n25832 = n25831 ^ n25747;
  assign n25833 = n24072 ^ n1458;
  assign n25834 = n25833 ^ n1192;
  assign n25835 = n25834 ^ n1381;
  assign n25836 = n25835 ^ n25747;
  assign n25837 = n25832 & ~n25836;
  assign n25838 = n25837 ^ n25835;
  assign n25746 = n25736 ^ n25735;
  assign n25839 = n25838 ^ n25746;
  assign n1377 = n1376 ^ n1280;
  assign n1384 = n1383 ^ n1377;
  assign n1388 = n1387 ^ n1384;
  assign n25840 = n25838 ^ n1388;
  assign n25841 = ~n25839 & n25840;
  assign n25842 = n25841 ^ n1388;
  assign n25843 = n25842 ^ n25744;
  assign n25844 = n25745 & ~n25843;
  assign n25845 = n25844 ^ n2448;
  assign n25743 = n25739 ^ n25701;
  assign n25846 = n25845 ^ n25743;
  assign n3043 = n3038 ^ n3033;
  assign n3044 = n3043 ^ n2452;
  assign n3045 = n3044 ^ n2500;
  assign n25847 = n25743 ^ n3045;
  assign n25848 = n25846 & ~n25847;
  assign n25849 = n25848 ^ n3045;
  assign n25850 = n25849 ^ n25741;
  assign n25851 = n25742 & ~n25850;
  assign n25852 = n25851 ^ n2504;
  assign n26133 = n25868 ^ n25852;
  assign n26134 = ~n25869 & n26133;
  assign n26135 = n26134 ^ n3065;
  assign n26136 = n26135 ^ n26131;
  assign n26137 = ~n26132 & n26136;
  assign n26138 = n26137 ^ n3221;
  assign n26026 = n26025 ^ n26021;
  assign n26027 = ~n26022 & n26026;
  assign n26028 = n26027 ^ n23163;
  assign n25969 = n25968 ^ n25964;
  assign n25970 = n25965 & n25969;
  assign n25971 = n25970 ^ n25962;
  assign n25959 = n25147 ^ n24141;
  assign n25960 = n25959 ^ n24264;
  assign n25958 = n25468 ^ n25450;
  assign n25961 = n25960 ^ n25958;
  assign n26019 = n25971 ^ n25961;
  assign n26020 = n26019 ^ n23159;
  assign n26076 = n26028 ^ n26020;
  assign n26075 = n26073 & n26074;
  assign n26129 = n26076 ^ n26075;
  assign n26130 = n26129 ^ n2843;
  assign n26429 = n26138 ^ n26130;
  assign n26432 = n26431 ^ n26429;
  assign n26288 = n24857 ^ n24122;
  assign n26005 = n25505 ^ n25433;
  assign n26289 = n26288 ^ n26005;
  assign n26287 = n26135 ^ n26132;
  assign n26290 = n26289 ^ n26287;
  assign n25872 = n25495 ^ n2883;
  assign n25873 = n25872 ^ n24664;
  assign n25874 = n25873 ^ n25352;
  assign n25871 = n25849 ^ n25742;
  assign n25875 = n25874 ^ n25871;
  assign n25878 = n25491 ^ n1583;
  assign n25877 = n25251 ^ n24259;
  assign n25879 = n25878 ^ n25877;
  assign n25876 = n25846 ^ n3045;
  assign n25880 = n25879 ^ n25876;
  assign n25884 = n25842 ^ n2448;
  assign n25885 = n25884 ^ n25744;
  assign n25882 = n25487 ^ n25486;
  assign n25881 = n25244 ^ n24264;
  assign n25883 = n25882 ^ n25881;
  assign n25886 = n25885 ^ n25883;
  assign n26265 = n25839 ^ n1388;
  assign n25890 = n25835 ^ n25832;
  assign n25887 = n25479 ^ n2660;
  assign n25888 = n25887 ^ n24270;
  assign n25889 = n25888 ^ n25147;
  assign n25891 = n25890 ^ n25889;
  assign n25895 = n25828 ^ n25827;
  assign n25892 = n25475 ^ n3187;
  assign n25893 = n25892 ^ n24274;
  assign n25894 = n25893 ^ n25153;
  assign n25896 = n25895 ^ n25894;
  assign n25900 = n25823 ^ n25822;
  assign n25897 = n25471 ^ n25445;
  assign n25898 = n25897 ^ n25158;
  assign n25899 = n25898 ^ n24442;
  assign n25901 = n25900 ^ n25899;
  assign n26242 = n25814 ^ n905;
  assign n26243 = n26242 ^ n25812;
  assign n26235 = n25809 ^ n25750;
  assign n25905 = n25806 ^ n25805;
  assign n25903 = n25606 ^ n25094;
  assign n25904 = n25903 ^ n24421;
  assign n25906 = n25905 ^ n25904;
  assign n25909 = n25099 ^ n24286;
  assign n25910 = n25909 ^ n25082;
  assign n25907 = n25801 ^ n25754;
  assign n25908 = n25907 ^ n25751;
  assign n25911 = n25910 ^ n25908;
  assign n25913 = n25088 ^ n24290;
  assign n25914 = n25913 ^ n25104;
  assign n25912 = n25798 ^ n25795;
  assign n25915 = n25914 ^ n25912;
  assign n25917 = n25093 ^ n24297;
  assign n25918 = n25917 ^ n25111;
  assign n25916 = n25791 ^ n25788;
  assign n25919 = n25918 ^ n25916;
  assign n25924 = n25781 ^ n25764;
  assign n25922 = n25178 ^ n24306;
  assign n25923 = n25922 ^ n25108;
  assign n25925 = n25924 ^ n25923;
  assign n25926 = n25113 ^ n24308;
  assign n25927 = n25926 ^ n25122;
  assign n25929 = n25928 ^ n25927;
  assign n25932 = n25775 ^ n25774;
  assign n25930 = n25127 ^ n25118;
  assign n25931 = n25930 ^ n23738;
  assign n25933 = n25932 ^ n25931;
  assign n25934 = n25577 ^ n24315;
  assign n25935 = n25934 ^ n25077;
  assign n25937 = n25936 ^ n25935;
  assign n26172 = n25124 ^ n24247;
  assign n26173 = n26172 ^ n24982;
  assign n25942 = n24865 ^ n23576;
  assign n25943 = n25942 ^ n24232;
  assign n25944 = n25943 ^ n25872;
  assign n25945 = n25407 ^ n23591;
  assign n25946 = n25945 ^ n24148;
  assign n25947 = n25946 ^ n25882;
  assign n25950 = n25482 ^ n25438;
  assign n25948 = n25352 ^ n23584;
  assign n25949 = n25948 ^ n24122;
  assign n25951 = n25950 ^ n25949;
  assign n25952 = n25251 ^ n24678;
  assign n25953 = n25952 ^ n24267;
  assign n25954 = n25953 ^ n25887;
  assign n25955 = n25244 ^ n24664;
  assign n25956 = n25955 ^ n24218;
  assign n25957 = n25956 ^ n25892;
  assign n25972 = n25971 ^ n25958;
  assign n25973 = ~n25961 & n25972;
  assign n25974 = n25973 ^ n25960;
  assign n25975 = n25974 ^ n25897;
  assign n25976 = n25143 ^ n24166;
  assign n25977 = n25976 ^ n24259;
  assign n25978 = n25977 ^ n25897;
  assign n25979 = n25975 & n25978;
  assign n25980 = n25979 ^ n25977;
  assign n25981 = n25980 ^ n25892;
  assign n25982 = n25957 & ~n25981;
  assign n25983 = n25982 ^ n25956;
  assign n25984 = n25983 ^ n25953;
  assign n25985 = ~n25954 & ~n25984;
  assign n25986 = n25985 ^ n25887;
  assign n25987 = n25986 ^ n25949;
  assign n25988 = ~n25951 & ~n25987;
  assign n25989 = n25988 ^ n25950;
  assign n25990 = n25989 ^ n25882;
  assign n25991 = ~n25947 & ~n25990;
  assign n25992 = n25991 ^ n25946;
  assign n25993 = n25992 ^ n25878;
  assign n25994 = n24857 ^ n24178;
  assign n25995 = n25994 ^ n23582;
  assign n25996 = n25995 ^ n25878;
  assign n25997 = ~n25993 & ~n25996;
  assign n25998 = n25997 ^ n25995;
  assign n25999 = n25998 ^ n25872;
  assign n26000 = ~n25944 & n25999;
  assign n26001 = n26000 ^ n25943;
  assign n25939 = n24855 ^ n23574;
  assign n25940 = n25939 ^ n24364;
  assign n25938 = n25502 ^ n25499;
  assign n25941 = n25940 ^ n25938;
  assign n26060 = n26001 ^ n25941;
  assign n26065 = n26060 ^ n22949;
  assign n26016 = n25980 ^ n25957;
  assign n26017 = n26016 ^ n23396;
  assign n26029 = n26028 ^ n26019;
  assign n26030 = n26020 & n26029;
  assign n26031 = n26030 ^ n23159;
  assign n26018 = n25977 ^ n25975;
  assign n26032 = n26031 ^ n26018;
  assign n26033 = n26018 ^ n23287;
  assign n26034 = n26032 & ~n26033;
  assign n26035 = n26034 ^ n23287;
  assign n26036 = n26035 ^ n26016;
  assign n26037 = n26017 & ~n26036;
  assign n26038 = n26037 ^ n23396;
  assign n26015 = n25983 ^ n25954;
  assign n26039 = n26038 ^ n26015;
  assign n26040 = n26038 ^ n23449;
  assign n26041 = n26039 & n26040;
  assign n26042 = n26041 ^ n23449;
  assign n26014 = n25986 ^ n25951;
  assign n26043 = n26042 ^ n26014;
  assign n26044 = n26014 ^ n22961;
  assign n26045 = ~n26043 & ~n26044;
  assign n26046 = n26045 ^ n22961;
  assign n26013 = n25989 ^ n25947;
  assign n26047 = n26046 ^ n26013;
  assign n26048 = n26013 ^ n22966;
  assign n26049 = ~n26047 & ~n26048;
  assign n26050 = n26049 ^ n22966;
  assign n26012 = n25995 ^ n25993;
  assign n26051 = n26050 ^ n26012;
  assign n26052 = n26012 ^ n22957;
  assign n26053 = ~n26051 & ~n26052;
  assign n26054 = n26053 ^ n22957;
  assign n26011 = n25998 ^ n25944;
  assign n26055 = n26054 ^ n26011;
  assign n26056 = n26011 ^ n22951;
  assign n26057 = ~n26055 & n26056;
  assign n26058 = n26057 ^ n22951;
  assign n26066 = n26065 ^ n26058;
  assign n26067 = n26055 ^ n22951;
  assign n26068 = n26043 ^ n22961;
  assign n26069 = n26015 ^ n23449;
  assign n26070 = n26069 ^ n26038;
  assign n26071 = n26035 ^ n26017;
  assign n26072 = n26032 ^ n23287;
  assign n26077 = ~n26075 & n26076;
  assign n26078 = ~n26072 & ~n26077;
  assign n26079 = n26071 & n26078;
  assign n26080 = n26070 & ~n26079;
  assign n26081 = ~n26068 & ~n26080;
  assign n26082 = n26047 ^ n22966;
  assign n26083 = n26081 & n26082;
  assign n26084 = n26051 ^ n22957;
  assign n26085 = n26083 & ~n26084;
  assign n26086 = n26067 & ~n26085;
  assign n26087 = ~n26066 & ~n26086;
  assign n26059 = n26058 ^ n22949;
  assign n26061 = n26060 ^ n26058;
  assign n26062 = ~n26059 & n26061;
  assign n26063 = n26062 ^ n22949;
  assign n26006 = n24848 ^ n23607;
  assign n26007 = n26006 ^ n24341;
  assign n26008 = n26007 ^ n26005;
  assign n26002 = n26001 ^ n25938;
  assign n26003 = n25941 & ~n26002;
  assign n26004 = n26003 ^ n25940;
  assign n26009 = n26008 ^ n26004;
  assign n26010 = n26009 ^ n22342;
  assign n26064 = n26063 ^ n26010;
  assign n26104 = n26087 ^ n26064;
  assign n26105 = n26104 ^ n2089;
  assign n26106 = n26086 ^ n26066;
  assign n26107 = n26106 ^ n2078;
  assign n26108 = n26085 ^ n26067;
  assign n26112 = n26111 ^ n26108;
  assign n26113 = n26084 ^ n26083;
  assign n26117 = n26116 ^ n26113;
  assign n26118 = n26082 ^ n26081;
  assign n26119 = n26118 ^ n1670;
  assign n26120 = n26080 ^ n26068;
  assign n26124 = n26123 ^ n26120;
  assign n26127 = n26077 ^ n26072;
  assign n2848 = n2787 ^ n1496;
  assign n2849 = n2848 ^ n2834;
  assign n2853 = n2852 ^ n2849;
  assign n26128 = n26127 ^ n2853;
  assign n26139 = n26138 ^ n26129;
  assign n26140 = ~n26130 & n26139;
  assign n26141 = n26140 ^ n2843;
  assign n26142 = n26141 ^ n26127;
  assign n26143 = ~n26128 & n26142;
  assign n26144 = n26143 ^ n2853;
  assign n26126 = n26078 ^ n26071;
  assign n26145 = n26144 ^ n26126;
  assign n26146 = n26126 ^ n2868;
  assign n26147 = n26145 & ~n26146;
  assign n26148 = n26147 ^ n2868;
  assign n26125 = n26079 ^ n26070;
  assign n26149 = n26148 ^ n26125;
  assign n26150 = n26125 ^ n1547;
  assign n26151 = n26149 & ~n26150;
  assign n26152 = n26151 ^ n1547;
  assign n26153 = n26152 ^ n26123;
  assign n26154 = ~n26124 & ~n26153;
  assign n26155 = n26154 ^ n26120;
  assign n26156 = n26155 ^ n26118;
  assign n26157 = ~n26119 & ~n26156;
  assign n26158 = n26157 ^ n1670;
  assign n26159 = n26158 ^ n26113;
  assign n26160 = n26117 & ~n26159;
  assign n26161 = n26160 ^ n26116;
  assign n26162 = n26161 ^ n26108;
  assign n26163 = ~n26112 & n26162;
  assign n26164 = n26163 ^ n26111;
  assign n26165 = n26164 ^ n2078;
  assign n26166 = ~n26107 & ~n26165;
  assign n26167 = n26166 ^ n26106;
  assign n26168 = n26167 ^ n26104;
  assign n26169 = ~n26105 & ~n26168;
  assign n26170 = n26169 ^ n2089;
  assign n26097 = n26063 ^ n26009;
  assign n26098 = n26010 & ~n26097;
  assign n26099 = n26098 ^ n22342;
  assign n26100 = n26099 ^ n22337;
  assign n26093 = n26007 ^ n26004;
  assign n26094 = ~n26008 & n26093;
  assign n26095 = n26094 ^ n26004;
  assign n26090 = n24843 ^ n24337;
  assign n26091 = n26090 ^ n23638;
  assign n26092 = n26091 ^ n26089;
  assign n26096 = n26095 ^ n26092;
  assign n26101 = n26100 ^ n26096;
  assign n26088 = n26064 & n26087;
  assign n26102 = n26101 ^ n26088;
  assign n2103 = n2064 ^ n2022;
  assign n2104 = n2103 ^ n2098;
  assign n2108 = n2107 ^ n2104;
  assign n26103 = n26102 ^ n2108;
  assign n26171 = n26170 ^ n26103;
  assign n26174 = n26173 ^ n26171;
  assign n26177 = n26167 ^ n26105;
  assign n26175 = n25130 ^ n24252;
  assign n26176 = n26175 ^ n24949;
  assign n26178 = n26177 ^ n26176;
  assign n26183 = n25138 ^ n24333;
  assign n26184 = n26183 ^ n24884;
  assign n26185 = n26158 ^ n26116;
  assign n26186 = n26185 ^ n26113;
  assign n26187 = ~n26184 & n26186;
  assign n26181 = n25137 ^ n24245;
  assign n26182 = n26181 ^ n24327;
  assign n26188 = n26187 ^ n26182;
  assign n26189 = n26161 ^ n26111;
  assign n26190 = n26189 ^ n26108;
  assign n26191 = n26190 ^ n26187;
  assign n26192 = n26188 & n26191;
  assign n26193 = n26192 ^ n26182;
  assign n26179 = n24896 ^ n24325;
  assign n26180 = n26179 ^ n25135;
  assign n26194 = n26193 ^ n26180;
  assign n26195 = n26164 ^ n26107;
  assign n26196 = n26195 ^ n26193;
  assign n26197 = ~n26194 & n26196;
  assign n26198 = n26197 ^ n26180;
  assign n26199 = n26198 ^ n26177;
  assign n26200 = ~n26178 & n26199;
  assign n26201 = n26200 ^ n26176;
  assign n26202 = n26201 ^ n26171;
  assign n26203 = n26174 & n26202;
  assign n26204 = n26203 ^ n26173;
  assign n26205 = n26204 ^ n25936;
  assign n26206 = n25937 & ~n26205;
  assign n26207 = n26206 ^ n25935;
  assign n26208 = n26207 ^ n25932;
  assign n26209 = ~n25933 & ~n26208;
  assign n26210 = n26209 ^ n25931;
  assign n26211 = n26210 ^ n25927;
  assign n26212 = n25929 & n26211;
  assign n26213 = n26212 ^ n25928;
  assign n26214 = n26213 ^ n25924;
  assign n26215 = ~n25925 & ~n26214;
  assign n26216 = n26215 ^ n25923;
  assign n25920 = n25784 ^ n702;
  assign n25921 = n25920 ^ n25758;
  assign n26217 = n26216 ^ n25921;
  assign n26218 = n25116 ^ n25101;
  assign n26219 = n26218 ^ n24301;
  assign n26220 = n26219 ^ n25921;
  assign n26221 = ~n26217 & n26220;
  assign n26222 = n26221 ^ n26219;
  assign n26223 = n26222 ^ n25916;
  assign n26224 = n25919 & n26223;
  assign n26225 = n26224 ^ n25918;
  assign n26226 = n26225 ^ n25912;
  assign n26227 = n25915 & n26226;
  assign n26228 = n26227 ^ n25914;
  assign n26229 = n26228 ^ n25910;
  assign n26230 = n25911 & n26229;
  assign n26231 = n26230 ^ n25908;
  assign n26232 = n26231 ^ n25905;
  assign n26233 = n25906 & ~n26232;
  assign n26234 = n26233 ^ n25904;
  assign n26236 = n26235 ^ n26234;
  assign n26237 = n25860 ^ n24283;
  assign n26238 = n26237 ^ n25089;
  assign n26239 = n26238 ^ n26235;
  assign n26240 = n26236 & ~n26239;
  assign n26241 = n26240 ^ n26238;
  assign n26244 = n26243 ^ n26241;
  assign n26245 = n25962 ^ n25085;
  assign n26246 = n26245 ^ n24277;
  assign n26247 = n26246 ^ n26243;
  assign n26248 = n26244 & ~n26247;
  assign n26249 = n26248 ^ n26246;
  assign n25902 = n25818 ^ n1021;
  assign n26250 = n26249 ^ n25902;
  assign n26251 = n25162 ^ n24435;
  assign n26252 = n26251 ^ n25958;
  assign n26253 = n26252 ^ n25902;
  assign n26254 = ~n26250 & ~n26253;
  assign n26255 = n26254 ^ n26252;
  assign n26256 = n26255 ^ n25900;
  assign n26257 = n25901 & ~n26256;
  assign n26258 = n26257 ^ n25899;
  assign n26259 = n26258 ^ n25895;
  assign n26260 = n25896 & n26259;
  assign n26261 = n26260 ^ n25894;
  assign n26262 = n26261 ^ n25890;
  assign n26263 = n25891 & n26262;
  assign n26264 = n26263 ^ n25889;
  assign n26266 = n26265 ^ n26264;
  assign n26267 = n25950 ^ n25143;
  assign n26268 = n26267 ^ n24455;
  assign n26269 = n26268 ^ n26265;
  assign n26270 = n26266 & n26269;
  assign n26271 = n26270 ^ n26268;
  assign n26272 = n26271 ^ n25885;
  assign n26273 = ~n25886 & ~n26272;
  assign n26274 = n26273 ^ n25883;
  assign n26275 = n26274 ^ n25876;
  assign n26276 = ~n25880 & ~n26275;
  assign n26277 = n26276 ^ n25879;
  assign n26278 = n26277 ^ n25871;
  assign n26279 = ~n25875 & ~n26278;
  assign n26280 = n26279 ^ n25874;
  assign n25870 = n25869 ^ n25852;
  assign n26281 = n26280 ^ n25870;
  assign n26282 = n25938 ^ n24678;
  assign n26283 = n26282 ^ n25407;
  assign n26284 = n26283 ^ n25870;
  assign n26285 = ~n26281 & n26284;
  assign n26286 = n26285 ^ n26283;
  assign n26426 = n26289 ^ n26286;
  assign n26427 = n26290 & ~n26426;
  assign n26428 = n26427 ^ n26287;
  assign n26433 = n26432 ^ n26428;
  assign n26291 = n26290 ^ n26286;
  assign n26292 = n26291 ^ n23584;
  assign n26296 = n26274 ^ n25880;
  assign n26297 = n26296 ^ n24166;
  assign n26298 = n26271 ^ n25886;
  assign n26299 = n26298 ^ n24141;
  assign n26300 = n26268 ^ n26266;
  assign n26301 = n26300 ^ n23971;
  assign n26302 = n26261 ^ n25889;
  assign n26303 = n26302 ^ n25890;
  assign n26304 = n26303 ^ n23866;
  assign n26307 = n26255 ^ n25899;
  assign n26308 = n26307 ^ n25900;
  assign n26309 = n26308 ^ n23747;
  assign n26310 = n26252 ^ n26250;
  assign n26311 = n26310 ^ n23751;
  assign n26314 = n26231 ^ n25906;
  assign n26315 = n26314 ^ n23764;
  assign n26316 = n26228 ^ n25911;
  assign n26317 = n26316 ^ n23769;
  assign n26318 = n26225 ^ n25915;
  assign n26319 = n26318 ^ n23773;
  assign n26321 = n26219 ^ n26217;
  assign n26322 = n26321 ^ n23780;
  assign n26323 = n26213 ^ n25925;
  assign n26324 = n26323 ^ n23145;
  assign n26326 = n26207 ^ n25931;
  assign n26327 = n26326 ^ n25932;
  assign n26328 = n26327 ^ n23788;
  assign n26329 = n26204 ^ n25937;
  assign n26330 = n26329 ^ n23791;
  assign n26331 = n26201 ^ n26173;
  assign n26332 = n26331 ^ n26171;
  assign n26333 = n26332 ^ n23811;
  assign n26334 = n26198 ^ n26176;
  assign n26335 = n26334 ^ n26177;
  assign n26336 = n26335 ^ n23795;
  assign n26337 = n26186 ^ n26184;
  assign n26338 = ~n23668 & ~n26337;
  assign n26339 = n26338 ^ n23729;
  assign n26340 = n26190 ^ n26188;
  assign n26341 = n26340 ^ n26338;
  assign n26342 = n26339 & n26341;
  assign n26343 = n26342 ^ n23729;
  assign n26344 = n26343 ^ n23798;
  assign n26345 = n26195 ^ n26194;
  assign n26346 = n26345 ^ n26343;
  assign n26347 = ~n26344 & ~n26346;
  assign n26348 = n26347 ^ n23798;
  assign n26349 = n26348 ^ n26335;
  assign n26350 = ~n26336 & n26349;
  assign n26351 = n26350 ^ n23795;
  assign n26352 = n26351 ^ n26332;
  assign n26353 = ~n26333 & ~n26352;
  assign n26354 = n26353 ^ n23811;
  assign n26355 = n26354 ^ n26329;
  assign n26356 = ~n26330 & ~n26355;
  assign n26357 = n26356 ^ n23791;
  assign n26358 = n26357 ^ n26327;
  assign n26359 = ~n26328 & ~n26358;
  assign n26360 = n26359 ^ n23788;
  assign n26325 = n26210 ^ n25929;
  assign n26361 = n26360 ^ n26325;
  assign n26362 = n26325 ^ n23787;
  assign n26363 = n26361 & n26362;
  assign n26364 = n26363 ^ n23787;
  assign n26365 = n26364 ^ n26323;
  assign n26366 = ~n26324 & ~n26365;
  assign n26367 = n26366 ^ n23145;
  assign n26368 = n26367 ^ n26321;
  assign n26369 = n26322 & n26368;
  assign n26370 = n26369 ^ n23780;
  assign n26320 = n26222 ^ n25919;
  assign n26371 = n26370 ^ n26320;
  assign n26372 = n26320 ^ n23775;
  assign n26373 = ~n26371 & ~n26372;
  assign n26374 = n26373 ^ n23775;
  assign n26375 = n26374 ^ n26318;
  assign n26376 = ~n26319 & ~n26375;
  assign n26377 = n26376 ^ n23773;
  assign n26378 = n26377 ^ n26316;
  assign n26379 = ~n26317 & ~n26378;
  assign n26380 = n26379 ^ n23769;
  assign n26381 = n26380 ^ n26314;
  assign n26382 = n26315 & ~n26381;
  assign n26383 = n26382 ^ n23764;
  assign n26313 = n26238 ^ n26236;
  assign n26384 = n26383 ^ n26313;
  assign n26385 = n26313 ^ n23760;
  assign n26386 = n26384 & ~n26385;
  assign n26387 = n26386 ^ n23760;
  assign n26312 = n26246 ^ n26244;
  assign n26388 = n26387 ^ n26312;
  assign n26389 = n26312 ^ n23756;
  assign n26390 = n26388 & ~n26389;
  assign n26391 = n26390 ^ n23756;
  assign n26392 = n26391 ^ n26310;
  assign n26393 = n26311 & n26392;
  assign n26394 = n26393 ^ n23751;
  assign n26395 = n26394 ^ n26308;
  assign n26396 = n26309 & ~n26395;
  assign n26397 = n26396 ^ n23747;
  assign n26305 = n26258 ^ n25894;
  assign n26306 = n26305 ^ n25895;
  assign n26398 = n26397 ^ n26306;
  assign n26399 = n26306 ^ n23742;
  assign n26400 = ~n26398 & ~n26399;
  assign n26401 = n26400 ^ n23742;
  assign n26402 = n26401 ^ n26303;
  assign n26403 = ~n26304 & ~n26402;
  assign n26404 = n26403 ^ n23866;
  assign n26405 = n26404 ^ n26300;
  assign n26406 = ~n26301 & ~n26405;
  assign n26407 = n26406 ^ n23971;
  assign n26408 = n26407 ^ n26298;
  assign n26409 = n26299 & n26408;
  assign n26410 = n26409 ^ n24141;
  assign n26411 = n26410 ^ n26296;
  assign n26412 = n26297 & n26411;
  assign n26413 = n26412 ^ n24166;
  assign n26294 = n26277 ^ n25874;
  assign n26295 = n26294 ^ n25871;
  assign n26414 = n26413 ^ n26295;
  assign n26415 = n26295 ^ n24218;
  assign n26416 = n26414 & ~n26415;
  assign n26417 = n26416 ^ n24218;
  assign n26293 = n26283 ^ n26281;
  assign n26418 = n26417 ^ n26293;
  assign n26419 = n26293 ^ n24267;
  assign n26420 = n26418 & ~n26419;
  assign n26421 = n26420 ^ n24267;
  assign n26422 = n26421 ^ n26291;
  assign n26423 = n26292 & n26422;
  assign n26424 = n26423 ^ n23584;
  assign n26425 = n26424 ^ n23591;
  assign n26434 = n26433 ^ n26425;
  assign n26435 = n26421 ^ n26292;
  assign n26436 = n26414 ^ n24218;
  assign n26437 = n26410 ^ n26297;
  assign n26438 = n26401 ^ n26304;
  assign n26439 = n26388 ^ n23756;
  assign n26440 = n26380 ^ n23764;
  assign n26441 = n26440 ^ n26314;
  assign n26442 = n26377 ^ n23769;
  assign n26443 = n26442 ^ n26316;
  assign n26444 = n26374 ^ n26319;
  assign n26445 = n26371 ^ n23775;
  assign n26446 = n26361 ^ n23787;
  assign n26447 = n26357 ^ n23788;
  assign n26448 = n26447 ^ n26327;
  assign n26449 = n26351 ^ n23811;
  assign n26450 = n26449 ^ n26332;
  assign n26451 = n26348 ^ n26336;
  assign n26452 = n26337 ^ n23668;
  assign n26453 = n26340 ^ n26339;
  assign n26454 = n26452 & ~n26453;
  assign n26455 = n26345 ^ n26344;
  assign n26456 = n26454 & ~n26455;
  assign n26457 = n26451 & n26456;
  assign n26458 = n26450 & n26457;
  assign n26459 = n26354 ^ n23791;
  assign n26460 = n26459 ^ n26329;
  assign n26461 = ~n26458 & n26460;
  assign n26462 = n26448 & ~n26461;
  assign n26463 = ~n26446 & ~n26462;
  assign n26464 = n26364 ^ n26324;
  assign n26465 = n26463 & ~n26464;
  assign n26466 = n26367 ^ n26322;
  assign n26467 = n26465 & ~n26466;
  assign n26468 = n26445 & ~n26467;
  assign n26469 = n26444 & ~n26468;
  assign n26470 = n26443 & ~n26469;
  assign n26471 = ~n26441 & ~n26470;
  assign n26472 = n26384 ^ n23760;
  assign n26473 = n26471 & n26472;
  assign n26474 = n26439 & n26473;
  assign n26475 = n26391 ^ n23751;
  assign n26476 = n26475 ^ n26310;
  assign n26477 = n26474 & ~n26476;
  assign n26478 = n26394 ^ n26309;
  assign n26479 = ~n26477 & ~n26478;
  assign n26480 = n26398 ^ n23742;
  assign n26481 = n26479 & n26480;
  assign n26482 = n26438 & ~n26481;
  assign n26483 = n26404 ^ n23971;
  assign n26484 = n26483 ^ n26300;
  assign n26485 = n26482 & ~n26484;
  assign n26486 = n26407 ^ n26299;
  assign n26487 = ~n26485 & n26486;
  assign n26488 = n26437 & ~n26487;
  assign n26489 = n26436 & n26488;
  assign n26490 = n26418 ^ n24267;
  assign n26491 = ~n26489 & ~n26490;
  assign n26492 = ~n26435 & ~n26491;
  assign n26668 = n26434 & n26492;
  assign n26664 = n26141 ^ n26128;
  assign n26661 = n24855 ^ n24178;
  assign n26662 = n26661 ^ n25537;
  assign n26658 = n26431 ^ n26428;
  assign n26659 = ~n26432 & n26658;
  assign n26660 = n26659 ^ n26428;
  assign n26663 = n26662 ^ n26660;
  assign n26665 = n26664 ^ n26663;
  assign n26666 = n26665 ^ n23582;
  assign n26654 = n26433 ^ n23591;
  assign n26655 = n26433 ^ n26424;
  assign n26656 = n26654 & ~n26655;
  assign n26657 = n26656 ^ n23591;
  assign n26667 = n26666 ^ n26657;
  assign n26669 = n26668 ^ n26667;
  assign n1704 = n1703 ^ n1696;
  assign n1711 = n1710 ^ n1704;
  assign n1715 = n1714 ^ n1711;
  assign n26670 = n26669 ^ n1715;
  assign n26493 = n26492 ^ n26434;
  assign n1734 = n1727 ^ n1684;
  assign n1741 = n1740 ^ n1734;
  assign n1742 = n1741 ^ n1708;
  assign n26494 = n26493 ^ n1742;
  assign n26495 = n26490 ^ n26489;
  assign n26499 = n26498 ^ n26495;
  assign n26500 = n26488 ^ n26436;
  assign n26501 = n26500 ^ n3128;
  assign n26503 = n26486 ^ n26485;
  assign n26504 = n26503 ^ n3098;
  assign n26505 = n26484 ^ n26482;
  assign n2638 = n2634 ^ n2586;
  assign n2642 = n2641 ^ n2638;
  assign n2643 = n2642 ^ n1521;
  assign n26506 = n26505 ^ n2643;
  assign n26613 = n26478 ^ n26477;
  assign n26508 = n26476 ^ n26474;
  assign n26512 = n26511 ^ n26508;
  assign n26514 = n26472 ^ n26471;
  assign n1311 = n1292 ^ n1208;
  assign n1312 = n1311 ^ n1308;
  assign n1316 = n1315 ^ n1312;
  assign n26515 = n26514 ^ n1316;
  assign n26516 = n26470 ^ n26441;
  assign n1162 = n1122 ^ n1077;
  assign n1163 = n1162 ^ n1156;
  assign n1167 = n1166 ^ n1163;
  assign n26517 = n26516 ^ n1167;
  assign n26519 = n26468 ^ n26444;
  assign n26520 = n26519 ^ n1147;
  assign n26521 = n26467 ^ n26445;
  assign n26522 = n26521 ^ n3328;
  assign n26523 = n26466 ^ n26465;
  assign n26527 = n26526 ^ n26523;
  assign n26532 = n26462 ^ n26446;
  assign n26529 = n24741 ^ n17649;
  assign n26530 = n26529 ^ n650;
  assign n26531 = n26530 ^ n612;
  assign n26533 = n26532 ^ n26531;
  assign n26534 = n26461 ^ n26448;
  assign n570 = n569 ^ n563;
  assign n577 = n576 ^ n570;
  assign n581 = n580 ^ n577;
  assign n26535 = n26534 ^ n581;
  assign n26536 = n26460 ^ n26458;
  assign n26540 = n26539 ^ n26536;
  assign n26542 = n24243 ^ n543;
  assign n26543 = n26542 ^ n21375;
  assign n26544 = n26543 ^ n3248;
  assign n26541 = n26457 ^ n26450;
  assign n26545 = n26544 ^ n26541;
  assign n2368 = n2272 ^ n2201;
  assign n2369 = n2368 ^ n2132;
  assign n2370 = n2369 ^ n684;
  assign n26547 = n2370 & ~n26452;
  assign n2391 = n2350 ^ n2287;
  assign n2392 = n2391 ^ n2387;
  assign n2393 = n2392 ^ n2327;
  assign n26548 = n26547 ^ n2393;
  assign n26549 = n26453 ^ n26452;
  assign n26550 = n26549 ^ n2393;
  assign n26551 = n26548 & n26550;
  assign n26552 = n26551 ^ n26547;
  assign n26546 = n26455 ^ n26454;
  assign n26553 = n26552 ^ n26546;
  assign n26554 = n24193 ^ n17660;
  assign n26555 = n26554 ^ n2405;
  assign n26556 = n26555 ^ n16654;
  assign n26557 = n26556 ^ n26552;
  assign n26558 = n26553 & n26557;
  assign n26559 = n26558 ^ n26556;
  assign n26563 = n26562 ^ n26559;
  assign n26564 = n26456 ^ n26451;
  assign n26565 = n26564 ^ n26559;
  assign n26566 = n26563 & ~n26565;
  assign n26567 = n26566 ^ n26562;
  assign n26568 = n26567 ^ n26541;
  assign n26569 = n26545 & ~n26568;
  assign n26570 = n26569 ^ n26544;
  assign n26571 = n26570 ^ n26536;
  assign n26572 = n26540 & ~n26571;
  assign n26573 = n26572 ^ n26539;
  assign n26574 = n26573 ^ n26534;
  assign n26575 = ~n26535 & n26574;
  assign n26576 = n26575 ^ n581;
  assign n26577 = n26576 ^ n26532;
  assign n26578 = ~n26533 & n26577;
  assign n26579 = n26578 ^ n26531;
  assign n26528 = n26464 ^ n26463;
  assign n26580 = n26579 ^ n26528;
  assign n26581 = n26528 ^ n738;
  assign n26582 = ~n26580 & n26581;
  assign n26583 = n26582 ^ n738;
  assign n26584 = n26583 ^ n26523;
  assign n26585 = n26527 & ~n26584;
  assign n26586 = n26585 ^ n26526;
  assign n26587 = n26586 ^ n26521;
  assign n26588 = ~n26522 & n26587;
  assign n26589 = n26588 ^ n3328;
  assign n26590 = n26589 ^ n26519;
  assign n26591 = n26520 & ~n26590;
  assign n26592 = n26591 ^ n1147;
  assign n26518 = n26469 ^ n26443;
  assign n26593 = n26592 ^ n26518;
  assign n1128 = n1106 ^ n1059;
  assign n1132 = n1131 ^ n1128;
  assign n1136 = n1135 ^ n1132;
  assign n26594 = n26518 ^ n1136;
  assign n26595 = n26593 & ~n26594;
  assign n26596 = n26595 ^ n1136;
  assign n26597 = n26596 ^ n26516;
  assign n26598 = ~n26517 & n26597;
  assign n26599 = n26598 ^ n1167;
  assign n26600 = n26599 ^ n26514;
  assign n26601 = ~n26515 & n26600;
  assign n26602 = n26601 ^ n1316;
  assign n26513 = n26473 ^ n26439;
  assign n26603 = n26602 ^ n26513;
  assign n26604 = n3142 ^ n1396;
  assign n26605 = n26604 ^ n1323;
  assign n26606 = n26605 ^ n3014;
  assign n26607 = n26606 ^ n26513;
  assign n26608 = n26603 & ~n26607;
  assign n26609 = n26608 ^ n26606;
  assign n26610 = n26609 ^ n26508;
  assign n26611 = n26512 & ~n26610;
  assign n26612 = n26611 ^ n26511;
  assign n26614 = n26613 ^ n26612;
  assign n3157 = n3153 ^ n2460;
  assign n3164 = n3163 ^ n3157;
  assign n3165 = n3164 ^ n2552;
  assign n26615 = n26613 ^ n3165;
  assign n26616 = ~n26614 & n26615;
  assign n26617 = n26616 ^ n3165;
  assign n26507 = n26480 ^ n26479;
  assign n26618 = n26617 ^ n26507;
  assign n2549 = n2542 ^ n2518;
  assign n2556 = n2555 ^ n2549;
  assign n2560 = n2559 ^ n2556;
  assign n26619 = n26507 ^ n2560;
  assign n26620 = ~n26618 & n26619;
  assign n26621 = n26620 ^ n2560;
  assign n2567 = n2530 ^ n1556;
  assign n2568 = n2567 ^ n2564;
  assign n2572 = n2571 ^ n2568;
  assign n26622 = n26621 ^ n2572;
  assign n26623 = n26481 ^ n26438;
  assign n26624 = n26623 ^ n26621;
  assign n26625 = n26622 & ~n26624;
  assign n26626 = n26625 ^ n2572;
  assign n26627 = n26626 ^ n26505;
  assign n26628 = n26506 & ~n26627;
  assign n26629 = n26628 ^ n2643;
  assign n26630 = n26629 ^ n26503;
  assign n26631 = ~n26504 & n26630;
  assign n26632 = n26631 ^ n3098;
  assign n26502 = n26487 ^ n26437;
  assign n26633 = n26632 ^ n26502;
  assign n26634 = n26632 ^ n2753;
  assign n26635 = ~n26633 & n26634;
  assign n26636 = n26635 ^ n2753;
  assign n26637 = n26636 ^ n26500;
  assign n26638 = ~n26501 & n26637;
  assign n26639 = n26638 ^ n3128;
  assign n26640 = n26639 ^ n26495;
  assign n26641 = n26499 & ~n26640;
  assign n26642 = n26641 ^ n26498;
  assign n26646 = n26645 ^ n26642;
  assign n26647 = n26491 ^ n26435;
  assign n26648 = n26647 ^ n26642;
  assign n26649 = n26646 & n26648;
  assign n26650 = n26649 ^ n26645;
  assign n26651 = n26650 ^ n26493;
  assign n26652 = ~n26494 & n26651;
  assign n26653 = n26652 ^ n1742;
  assign n26671 = n26670 ^ n26653;
  assign n26956 = n26821 ^ n26671;
  assign n27047 = n26956 ^ n24333;
  assign n27144 = n2222 & ~n27047;
  assign n27148 = n27147 ^ n27144;
  assign n26801 = n26669 ^ n26653;
  assign n26802 = n26670 & ~n26801;
  assign n26803 = n26802 ^ n1715;
  assign n26788 = ~n26667 & n26668;
  assign n26769 = n26665 ^ n26657;
  assign n26770 = ~n26666 & ~n26769;
  assign n26771 = n26770 ^ n23582;
  assign n26786 = n26771 ^ n23576;
  assign n26749 = n26664 ^ n26662;
  assign n26750 = n26664 ^ n26660;
  assign n26751 = n26749 & ~n26750;
  assign n26752 = n26751 ^ n26662;
  assign n26746 = n25544 ^ n24848;
  assign n26747 = n26746 ^ n24232;
  assign n26745 = n26145 ^ n2868;
  assign n26748 = n26747 ^ n26745;
  assign n26767 = n26752 ^ n26748;
  assign n26787 = n26786 ^ n26767;
  assign n26800 = n26788 ^ n26787;
  assign n26804 = n26803 ^ n26800;
  assign n1819 = n1811 ^ n1761;
  assign n1823 = n1822 ^ n1819;
  assign n1827 = n1826 ^ n1823;
  assign n26826 = n26804 ^ n1827;
  assign n26823 = n25932 ^ n24245;
  assign n26824 = n26823 ^ n25130;
  assign n26822 = n26671 & n26821;
  assign n26825 = n26824 ^ n26822;
  assign n26959 = n26826 ^ n26825;
  assign n26957 = n24333 & n26956;
  assign n26958 = n26957 ^ n24327;
  assign n27048 = n26959 ^ n26958;
  assign n27149 = n27048 ^ n27047;
  assign n27150 = n27149 ^ n27144;
  assign n27151 = n27148 & ~n27150;
  assign n27152 = n27151 ^ n27147;
  assign n27140 = n18399 ^ n2330;
  assign n27141 = n27140 ^ n22140;
  assign n27142 = n27141 ^ n524;
  assign n27314 = n27152 ^ n27142;
  assign n26960 = n26959 ^ n26957;
  assign n26961 = n26958 & ~n26960;
  assign n26962 = n26961 ^ n24327;
  assign n26831 = n25928 ^ n24896;
  assign n26832 = n26831 ^ n25124;
  assign n26827 = n26826 ^ n26824;
  assign n26828 = n26825 & ~n26827;
  assign n26829 = n26828 ^ n26822;
  assign n26805 = n26800 ^ n1827;
  assign n26806 = ~n26804 & n26805;
  assign n26807 = n26806 ^ n1827;
  assign n26789 = ~n26787 & ~n26788;
  assign n26768 = n26767 ^ n23576;
  assign n26772 = n26771 ^ n26767;
  assign n26773 = ~n26768 & ~n26772;
  assign n26774 = n26773 ^ n23576;
  assign n26784 = n26774 ^ n23574;
  assign n26753 = n26752 ^ n26747;
  assign n26754 = ~n26748 & n26753;
  assign n26755 = n26754 ^ n26745;
  assign n26743 = n26149 ^ n1547;
  assign n26741 = n24843 ^ n24364;
  assign n26742 = n26741 ^ n25532;
  assign n26744 = n26743 ^ n26742;
  assign n26765 = n26755 ^ n26744;
  assign n26785 = n26784 ^ n26765;
  assign n26795 = n26789 ^ n26785;
  assign n26799 = n26798 ^ n26795;
  assign n26819 = n26807 ^ n26799;
  assign n26830 = n26829 ^ n26819;
  assign n26954 = n26832 ^ n26830;
  assign n26955 = n26954 ^ n24325;
  assign n27050 = n26962 ^ n26955;
  assign n27049 = n27047 & n27048;
  assign n27139 = n27050 ^ n27049;
  assign n27315 = n27314 ^ n27139;
  assign n26721 = n26556 ^ n26553;
  assign n28728 = n27315 ^ n26721;
  assign n27261 = n26626 ^ n2643;
  assign n27262 = n27261 ^ n26505;
  assign n27259 = n25537 ^ n24857;
  assign n26737 = n26152 ^ n26124;
  assign n27260 = n27259 ^ n26737;
  assign n27263 = n27262 ^ n27260;
  assign n27095 = n26623 ^ n2572;
  assign n27096 = n27095 ^ n26621;
  assign n27034 = n26618 ^ n2560;
  assign n27032 = n26005 ^ n25352;
  assign n27033 = n27032 ^ n26745;
  assign n27035 = n27034 ^ n27033;
  assign n26679 = n26609 ^ n26512;
  assign n26677 = n26429 ^ n25872;
  assign n26678 = n26677 ^ n25244;
  assign n26680 = n26679 ^ n26678;
  assign n26903 = n26606 ^ n26603;
  assign n26682 = n25882 ^ n25147;
  assign n26683 = n26682 ^ n25870;
  assign n26681 = n26599 ^ n26515;
  assign n26684 = n26683 ^ n26681;
  assign n26686 = n25950 ^ n25871;
  assign n26687 = n26686 ^ n25153;
  assign n26685 = n26596 ^ n26517;
  assign n26688 = n26687 ^ n26685;
  assign n26890 = n26593 ^ n1136;
  assign n26691 = n26589 ^ n26520;
  assign n26689 = n25892 ^ n25162;
  assign n26690 = n26689 ^ n25885;
  assign n26692 = n26691 ^ n26690;
  assign n26695 = n26586 ^ n26522;
  assign n26693 = n26265 ^ n25897;
  assign n26694 = n26693 ^ n25085;
  assign n26696 = n26695 ^ n26694;
  assign n26703 = n26576 ^ n26533;
  assign n26701 = n25900 ^ n25099;
  assign n26702 = n26701 ^ n25860;
  assign n26704 = n26703 ^ n26702;
  assign n26862 = n26573 ^ n26535;
  assign n26707 = n26243 ^ n25111;
  assign n26708 = n26707 ^ n25082;
  assign n26705 = n26570 ^ n26539;
  assign n26706 = n26705 ^ n26536;
  assign n26709 = n26708 ^ n26706;
  assign n26712 = n26567 ^ n26545;
  assign n26710 = n26235 ^ n25088;
  assign n26711 = n26710 ^ n25116;
  assign n26713 = n26712 ^ n26711;
  assign n26716 = n26564 ^ n26562;
  assign n26717 = n26716 ^ n26559;
  assign n26714 = n25905 ^ n25093;
  assign n26715 = n26714 ^ n25178;
  assign n26718 = n26717 ^ n26715;
  assign n26719 = n25122 ^ n25101;
  assign n26720 = n26719 ^ n25908;
  assign n26722 = n26721 ^ n26720;
  assign n26725 = n26549 ^ n26548;
  assign n26723 = n25912 ^ n25108;
  assign n26724 = n26723 ^ n25127;
  assign n26726 = n26725 ^ n26724;
  assign n26729 = n26452 ^ n2370;
  assign n26727 = n25916 ^ n25077;
  assign n26728 = n26727 ^ n25113;
  assign n26730 = n26729 ^ n26728;
  assign n26808 = n26807 ^ n26795;
  assign n26809 = ~n26799 & n26808;
  assign n26810 = n26809 ^ n26798;
  assign n26790 = ~n26785 & ~n26789;
  assign n26766 = n26765 ^ n23574;
  assign n26775 = n26774 ^ n26765;
  assign n26776 = ~n26766 & n26775;
  assign n26777 = n26776 ^ n23574;
  assign n26756 = n26755 ^ n26743;
  assign n26757 = ~n26744 & ~n26756;
  assign n26758 = n26757 ^ n26742;
  assign n26738 = n24341 ^ n24255;
  assign n26739 = n26738 ^ n25552;
  assign n26740 = n26739 ^ n26737;
  assign n26763 = n26758 ^ n26740;
  assign n26764 = n26763 ^ n23607;
  assign n26783 = n26777 ^ n26764;
  assign n26794 = n26790 ^ n26783;
  assign n26811 = n26810 ^ n26794;
  assign n26812 = n26794 ^ n1958;
  assign n26813 = ~n26811 & n26812;
  assign n26814 = n26813 ^ n1958;
  assign n26791 = ~n26783 & n26790;
  assign n26778 = n26777 ^ n26763;
  assign n26779 = ~n26764 & n26778;
  assign n26780 = n26779 ^ n23607;
  assign n26759 = n26758 ^ n26737;
  assign n26760 = n26740 & n26759;
  assign n26761 = n26760 ^ n26739;
  assign n26735 = n26155 ^ n26119;
  assign n26733 = n24337 ^ n24250;
  assign n26734 = n26733 ^ n25526;
  assign n26736 = n26735 ^ n26734;
  assign n26762 = n26761 ^ n26736;
  assign n26781 = n26780 ^ n26762;
  assign n26782 = n26781 ^ n23638;
  assign n26792 = n26791 ^ n26782;
  assign n26793 = n26792 ^ n2377;
  assign n26815 = n26814 ^ n26793;
  assign n26731 = n25921 ^ n24982;
  assign n26732 = n26731 ^ n25118;
  assign n26816 = n26815 ^ n26732;
  assign n26833 = n26832 ^ n26819;
  assign n26834 = n26830 & ~n26833;
  assign n26835 = n26834 ^ n26832;
  assign n26817 = n25924 ^ n24949;
  assign n26818 = n26817 ^ n25577;
  assign n26836 = n26835 ^ n26818;
  assign n26837 = n26811 ^ n1958;
  assign n26838 = n26837 ^ n26835;
  assign n26839 = ~n26836 & ~n26838;
  assign n26840 = n26839 ^ n26818;
  assign n26841 = n26840 ^ n26815;
  assign n26842 = ~n26816 & ~n26841;
  assign n26843 = n26842 ^ n26732;
  assign n26844 = n26843 ^ n26729;
  assign n26845 = ~n26730 & n26844;
  assign n26846 = n26845 ^ n26728;
  assign n26847 = n26846 ^ n26725;
  assign n26848 = n26726 & n26847;
  assign n26849 = n26848 ^ n26724;
  assign n26850 = n26849 ^ n26721;
  assign n26851 = n26722 & ~n26850;
  assign n26852 = n26851 ^ n26720;
  assign n26853 = n26852 ^ n26717;
  assign n26854 = ~n26718 & n26853;
  assign n26855 = n26854 ^ n26715;
  assign n26856 = n26855 ^ n26712;
  assign n26857 = ~n26713 & n26856;
  assign n26858 = n26857 ^ n26711;
  assign n26859 = n26858 ^ n26706;
  assign n26860 = n26709 & n26859;
  assign n26861 = n26860 ^ n26708;
  assign n26863 = n26862 ^ n26861;
  assign n26864 = n25902 ^ n25606;
  assign n26865 = n26864 ^ n25104;
  assign n26866 = n26865 ^ n26862;
  assign n26867 = n26863 & n26866;
  assign n26868 = n26867 ^ n26865;
  assign n26869 = n26868 ^ n26703;
  assign n26870 = ~n26704 & ~n26869;
  assign n26871 = n26870 ^ n26702;
  assign n26699 = n26579 ^ n738;
  assign n26700 = n26699 ^ n26528;
  assign n26872 = n26871 ^ n26700;
  assign n26873 = n25962 ^ n25895;
  assign n26874 = n26873 ^ n25094;
  assign n26875 = n26874 ^ n26700;
  assign n26876 = ~n26872 & ~n26875;
  assign n26877 = n26876 ^ n26874;
  assign n26697 = n26583 ^ n26526;
  assign n26698 = n26697 ^ n26523;
  assign n26878 = n26877 ^ n26698;
  assign n26879 = n25958 ^ n25890;
  assign n26880 = n26879 ^ n25089;
  assign n26881 = n26880 ^ n26698;
  assign n26882 = n26878 & n26881;
  assign n26883 = n26882 ^ n26880;
  assign n26884 = n26883 ^ n26695;
  assign n26885 = ~n26696 & n26884;
  assign n26886 = n26885 ^ n26694;
  assign n26887 = n26886 ^ n26690;
  assign n26888 = ~n26692 & n26887;
  assign n26889 = n26888 ^ n26691;
  assign n26891 = n26890 ^ n26889;
  assign n26892 = n25887 ^ n25876;
  assign n26893 = n26892 ^ n25158;
  assign n26894 = n26893 ^ n26890;
  assign n26895 = n26891 & n26894;
  assign n26896 = n26895 ^ n26893;
  assign n26897 = n26896 ^ n26685;
  assign n26898 = n26688 & ~n26897;
  assign n26899 = n26898 ^ n26687;
  assign n26900 = n26899 ^ n26681;
  assign n26901 = n26684 & ~n26900;
  assign n26902 = n26901 ^ n26683;
  assign n26904 = n26903 ^ n26902;
  assign n26905 = n26287 ^ n25878;
  assign n26906 = n26905 ^ n25143;
  assign n26907 = n26906 ^ n26903;
  assign n26908 = ~n26904 & ~n26907;
  assign n26909 = n26908 ^ n26906;
  assign n26910 = n26909 ^ n26678;
  assign n26911 = ~n26680 & n26910;
  assign n26912 = n26911 ^ n26679;
  assign n26675 = n26612 ^ n3165;
  assign n26676 = n26675 ^ n26613;
  assign n26913 = n26912 ^ n26676;
  assign n26673 = n26664 ^ n25251;
  assign n26674 = n26673 ^ n25938;
  assign n27029 = n26676 ^ n26674;
  assign n27030 = ~n26913 & n27029;
  assign n27031 = n27030 ^ n26674;
  assign n27092 = n27034 ^ n27031;
  assign n27093 = n27035 & ~n27092;
  assign n27094 = n27093 ^ n27033;
  assign n27097 = n27096 ^ n27094;
  assign n27090 = n26089 ^ n25407;
  assign n27091 = n27090 ^ n26743;
  assign n27256 = n27096 ^ n27091;
  assign n27257 = ~n27097 & n27256;
  assign n27258 = n27257 ^ n27091;
  assign n27264 = n27263 ^ n27258;
  assign n27265 = n27264 ^ n24122;
  assign n27098 = n27097 ^ n27091;
  assign n27099 = n27098 ^ n24678;
  assign n27036 = n27035 ^ n27031;
  assign n27037 = n27036 ^ n24664;
  assign n26914 = n26913 ^ n26674;
  assign n26915 = n26914 ^ n24259;
  assign n26916 = n26909 ^ n26680;
  assign n26917 = n26916 ^ n24264;
  assign n26918 = n26906 ^ n26904;
  assign n26919 = n26918 ^ n24455;
  assign n26920 = n26899 ^ n26684;
  assign n26921 = n26920 ^ n24270;
  assign n26922 = n26896 ^ n26688;
  assign n26923 = n26922 ^ n24274;
  assign n26924 = n26893 ^ n26891;
  assign n26925 = n26924 ^ n24442;
  assign n26926 = n26886 ^ n26692;
  assign n26927 = n26926 ^ n24435;
  assign n26928 = n26883 ^ n26696;
  assign n26929 = n26928 ^ n24277;
  assign n26931 = n26874 ^ n26872;
  assign n26932 = n26931 ^ n24421;
  assign n26933 = n26868 ^ n26702;
  assign n26934 = n26933 ^ n26703;
  assign n26935 = n26934 ^ n24286;
  assign n26936 = n26865 ^ n26863;
  assign n26937 = n26936 ^ n24290;
  assign n26941 = n26852 ^ n26715;
  assign n26942 = n26941 ^ n26717;
  assign n26943 = n26942 ^ n24306;
  assign n26944 = n26849 ^ n26722;
  assign n26945 = n26944 ^ n24308;
  assign n26946 = n26846 ^ n26726;
  assign n26947 = n26946 ^ n23738;
  assign n26948 = n26843 ^ n26730;
  assign n26949 = n26948 ^ n24315;
  assign n26950 = n26840 ^ n26816;
  assign n26951 = n26950 ^ n24247;
  assign n26952 = n26837 ^ n26836;
  assign n26953 = n26952 ^ n24252;
  assign n26963 = n26962 ^ n26954;
  assign n26964 = n26955 & n26963;
  assign n26965 = n26964 ^ n24325;
  assign n26966 = n26965 ^ n26952;
  assign n26967 = ~n26953 & ~n26966;
  assign n26968 = n26967 ^ n24252;
  assign n26969 = n26968 ^ n26950;
  assign n26970 = n26951 & ~n26969;
  assign n26971 = n26970 ^ n24247;
  assign n26972 = n26971 ^ n26948;
  assign n26973 = n26949 & n26972;
  assign n26974 = n26973 ^ n24315;
  assign n26975 = n26974 ^ n26946;
  assign n26976 = ~n26947 & n26975;
  assign n26977 = n26976 ^ n23738;
  assign n26978 = n26977 ^ n26944;
  assign n26979 = n26945 & ~n26978;
  assign n26980 = n26979 ^ n24308;
  assign n26981 = n26980 ^ n26942;
  assign n26982 = n26943 & n26981;
  assign n26983 = n26982 ^ n24306;
  assign n26940 = n26855 ^ n26713;
  assign n26984 = n26983 ^ n26940;
  assign n26985 = n26940 ^ n24301;
  assign n26986 = ~n26984 & n26985;
  assign n26987 = n26986 ^ n24301;
  assign n26938 = n26858 ^ n26708;
  assign n26939 = n26938 ^ n26706;
  assign n26988 = n26987 ^ n26939;
  assign n26989 = n26939 ^ n24297;
  assign n26990 = n26988 & n26989;
  assign n26991 = n26990 ^ n24297;
  assign n26992 = n26991 ^ n26936;
  assign n26993 = n26937 & n26992;
  assign n26994 = n26993 ^ n24290;
  assign n26995 = n26994 ^ n26934;
  assign n26996 = n26935 & ~n26995;
  assign n26997 = n26996 ^ n24286;
  assign n26998 = n26997 ^ n26931;
  assign n26999 = n26932 & n26998;
  assign n27000 = n26999 ^ n24421;
  assign n26930 = n26880 ^ n26878;
  assign n27001 = n27000 ^ n26930;
  assign n27002 = n26930 ^ n24283;
  assign n27003 = ~n27001 & ~n27002;
  assign n27004 = n27003 ^ n24283;
  assign n27005 = n27004 ^ n26928;
  assign n27006 = n26929 & n27005;
  assign n27007 = n27006 ^ n24277;
  assign n27008 = n27007 ^ n26926;
  assign n27009 = ~n26927 & ~n27008;
  assign n27010 = n27009 ^ n24435;
  assign n27011 = n27010 ^ n26924;
  assign n27012 = n26925 & ~n27011;
  assign n27013 = n27012 ^ n24442;
  assign n27014 = n27013 ^ n26922;
  assign n27015 = n26923 & n27014;
  assign n27016 = n27015 ^ n24274;
  assign n27017 = n27016 ^ n26920;
  assign n27018 = ~n26921 & ~n27017;
  assign n27019 = n27018 ^ n24270;
  assign n27020 = n27019 ^ n26918;
  assign n27021 = n26919 & ~n27020;
  assign n27022 = n27021 ^ n24455;
  assign n27023 = n27022 ^ n26916;
  assign n27024 = ~n26917 & n27023;
  assign n27025 = n27024 ^ n24264;
  assign n27026 = n27025 ^ n26914;
  assign n27027 = n26915 & ~n27026;
  assign n27028 = n27027 ^ n24259;
  assign n27087 = n27036 ^ n27028;
  assign n27088 = ~n27037 & ~n27087;
  assign n27089 = n27088 ^ n24664;
  assign n27253 = n27098 ^ n27089;
  assign n27254 = ~n27099 & n27253;
  assign n27255 = n27254 ^ n24678;
  assign n27371 = n27264 ^ n27255;
  assign n27372 = n27265 & ~n27371;
  assign n27373 = n27372 ^ n24122;
  assign n27341 = n27260 ^ n27258;
  assign n27342 = ~n27263 & n27341;
  assign n27343 = n27342 ^ n27262;
  assign n27336 = n26735 ^ n25544;
  assign n27337 = n27336 ^ n24865;
  assign n27368 = n27343 ^ n27337;
  assign n27338 = n26629 ^ n3098;
  assign n27339 = n27338 ^ n26503;
  assign n27369 = n27368 ^ n27339;
  assign n27370 = n27369 ^ n24148;
  assign n27392 = n27373 ^ n27370;
  assign n27266 = n27265 ^ n27255;
  assign n27038 = n27037 ^ n27028;
  assign n27039 = n27025 ^ n26915;
  assign n27040 = n27022 ^ n26917;
  assign n27041 = n27010 ^ n26925;
  assign n27042 = n27007 ^ n26927;
  assign n27043 = n27004 ^ n26929;
  assign n27044 = n26997 ^ n26932;
  assign n27045 = n26984 ^ n24301;
  assign n27046 = n26968 ^ n26951;
  assign n27051 = n27049 & n27050;
  assign n27052 = n26965 ^ n26953;
  assign n27053 = n27051 & n27052;
  assign n27054 = n27046 & n27053;
  assign n27055 = n26971 ^ n24315;
  assign n27056 = n27055 ^ n26948;
  assign n27057 = ~n27054 & ~n27056;
  assign n27058 = n26974 ^ n26947;
  assign n27059 = ~n27057 & n27058;
  assign n27060 = n26977 ^ n26945;
  assign n27061 = ~n27059 & n27060;
  assign n27062 = n26980 ^ n26943;
  assign n27063 = n27061 & n27062;
  assign n27064 = ~n27045 & n27063;
  assign n27065 = n26988 ^ n24297;
  assign n27066 = ~n27064 & n27065;
  assign n27067 = n26991 ^ n24290;
  assign n27068 = n27067 ^ n26936;
  assign n27069 = ~n27066 & n27068;
  assign n27070 = n26994 ^ n26935;
  assign n27071 = ~n27069 & n27070;
  assign n27072 = ~n27044 & ~n27071;
  assign n27073 = n27001 ^ n24283;
  assign n27074 = n27072 & ~n27073;
  assign n27075 = ~n27043 & n27074;
  assign n27076 = ~n27042 & n27075;
  assign n27077 = n27041 & ~n27076;
  assign n27078 = n27013 ^ n26923;
  assign n27079 = n27077 & n27078;
  assign n27080 = n27016 ^ n26921;
  assign n27081 = ~n27079 & ~n27080;
  assign n27082 = n27019 ^ n26919;
  assign n27083 = n27081 & ~n27082;
  assign n27084 = ~n27040 & ~n27083;
  assign n27085 = ~n27039 & ~n27084;
  assign n27086 = n27038 & n27085;
  assign n27100 = n27099 ^ n27089;
  assign n27267 = ~n27086 & n27100;
  assign n27391 = n27266 & ~n27267;
  assign n27418 = n27392 ^ n27391;
  assign n27422 = n27421 ^ n27418;
  assign n27268 = n27267 ^ n27266;
  assign n27101 = n27100 ^ n27086;
  assign n27102 = n27101 ^ n2955;
  assign n27106 = n27082 ^ n27081;
  assign n27107 = n27106 ^ n2717;
  assign n27108 = n27078 ^ n27077;
  assign n27112 = n27111 ^ n27108;
  assign n27114 = n25449 ^ n3173;
  assign n27115 = n27114 ^ n2438;
  assign n27116 = n27115 ^ n3038;
  assign n27113 = n27076 ^ n27041;
  assign n27117 = n27116 ^ n27113;
  assign n27118 = n27075 ^ n27042;
  assign n3021 = n3020 ^ n3017;
  assign n3022 = n3021 ^ n1484;
  assign n3023 = n3022 ^ n2436;
  assign n27119 = n27118 ^ n3023;
  assign n27121 = n27073 ^ n27072;
  assign n1454 = n1345 ^ n1262;
  assign n1455 = n1454 ^ n1178;
  assign n1459 = n1458 ^ n1455;
  assign n27122 = n27121 ^ n1459;
  assign n27123 = n27071 ^ n27044;
  assign n1445 = n1336 ^ n1244;
  assign n1449 = n1448 ^ n1445;
  assign n1450 = n1449 ^ n1176;
  assign n27124 = n27123 ^ n1450;
  assign n27125 = n27070 ^ n27069;
  assign n1002 = n1001 ^ n929;
  assign n1009 = n1008 ^ n1002;
  assign n1013 = n1012 ^ n1009;
  assign n27126 = n27125 ^ n1013;
  assign n27128 = n25058 ^ n1226;
  assign n27129 = n27128 ^ n877;
  assign n27130 = n27129 ^ n1006;
  assign n27127 = n27068 ^ n27066;
  assign n27131 = n27130 ^ n27127;
  assign n27132 = n27065 ^ n27064;
  assign n865 = n858 ^ n807;
  assign n869 = n868 ^ n865;
  assign n873 = n872 ^ n869;
  assign n27133 = n27132 ^ n873;
  assign n27156 = n25015 ^ n18394;
  assign n27157 = n27156 ^ n693;
  assign n27158 = n27157 ^ n16898;
  assign n27143 = n27142 ^ n27139;
  assign n27153 = n27152 ^ n27139;
  assign n27154 = n27143 & ~n27153;
  assign n27155 = n27154 ^ n27142;
  assign n27159 = n27158 ^ n27155;
  assign n27160 = n27052 ^ n27051;
  assign n27161 = n27160 ^ n27155;
  assign n27162 = n27159 & ~n27161;
  assign n27163 = n27162 ^ n27158;
  assign n27138 = n27053 ^ n27046;
  assign n27164 = n27163 ^ n27138;
  assign n27165 = n25010 ^ n18389;
  assign n27166 = n27165 ^ n22133;
  assign n27167 = n27166 ^ n699;
  assign n27168 = n27167 ^ n27138;
  assign n27169 = ~n27164 & n27168;
  assign n27170 = n27169 ^ n27167;
  assign n27137 = n27056 ^ n27054;
  assign n27171 = n27170 ^ n27137;
  assign n27175 = n27174 ^ n27137;
  assign n27176 = n27171 & ~n27175;
  assign n27177 = n27176 ^ n27174;
  assign n27136 = n27058 ^ n27057;
  assign n27178 = n27177 ^ n27136;
  assign n27182 = n27181 ^ n27136;
  assign n27183 = n27178 & ~n27182;
  assign n27184 = n27183 ^ n27181;
  assign n27185 = n27184 ^ n3293;
  assign n27186 = n27060 ^ n27059;
  assign n27187 = n27186 ^ n27184;
  assign n27188 = n27185 & ~n27187;
  assign n27189 = n27188 ^ n3293;
  assign n27135 = n27062 ^ n27061;
  assign n27190 = n27189 ^ n27135;
  assign n763 = n751 ^ n627;
  assign n770 = n769 ^ n763;
  assign n774 = n773 ^ n770;
  assign n27191 = n27189 ^ n774;
  assign n27192 = n27190 & n27191;
  assign n27193 = n27192 ^ n774;
  assign n27134 = n27063 ^ n27045;
  assign n27194 = n27193 ^ n27134;
  assign n27195 = n27134 ^ n787;
  assign n27196 = ~n27194 & n27195;
  assign n27197 = n27196 ^ n787;
  assign n27198 = n27197 ^ n27132;
  assign n27199 = ~n27133 & n27198;
  assign n27200 = n27199 ^ n873;
  assign n27201 = n27200 ^ n27127;
  assign n27202 = n27131 & ~n27201;
  assign n27203 = n27202 ^ n27130;
  assign n27204 = n27203 ^ n27125;
  assign n27205 = ~n27126 & n27204;
  assign n27206 = n27205 ^ n1013;
  assign n27207 = n27206 ^ n27123;
  assign n27208 = ~n27124 & n27207;
  assign n27209 = n27208 ^ n1450;
  assign n27210 = n27209 ^ n27121;
  assign n27211 = n27122 & ~n27210;
  assign n27212 = n27211 ^ n1459;
  assign n27120 = n27074 ^ n27043;
  assign n27213 = n27212 ^ n27120;
  assign n1472 = n1426 ^ n1360;
  assign n1473 = n1472 ^ n1466;
  assign n1474 = n1473 ^ n1376;
  assign n27214 = n27212 ^ n1474;
  assign n27215 = ~n27213 & n27214;
  assign n27216 = n27215 ^ n1474;
  assign n27217 = n27216 ^ n27118;
  assign n27218 = n27119 & ~n27217;
  assign n27219 = n27218 ^ n3023;
  assign n27220 = n27219 ^ n27113;
  assign n27221 = ~n27117 & n27220;
  assign n27222 = n27221 ^ n27116;
  assign n27223 = n27222 ^ n27108;
  assign n27224 = n27112 & ~n27223;
  assign n27225 = n27224 ^ n27111;
  assign n3194 = n3187 ^ n2596;
  assign n3198 = n3197 ^ n3194;
  assign n3199 = n3198 ^ n2711;
  assign n27226 = n27225 ^ n3199;
  assign n27227 = n27080 ^ n27079;
  assign n27228 = n27227 ^ n27225;
  assign n27229 = n27226 & n27228;
  assign n27230 = n27229 ^ n3199;
  assign n27231 = n27230 ^ n27106;
  assign n27232 = n27107 & ~n27231;
  assign n27233 = n27232 ^ n2717;
  assign n27105 = n27083 ^ n27040;
  assign n27234 = n27233 ^ n27105;
  assign n2724 = n2672 ^ n1524;
  assign n2725 = n2724 ^ n2721;
  assign n2729 = n2728 ^ n2725;
  assign n27235 = n27105 ^ n2729;
  assign n27236 = ~n27234 & n27235;
  assign n27237 = n27236 ^ n2729;
  assign n27104 = n27084 ^ n27039;
  assign n27238 = n27237 ^ n27104;
  assign n2822 = n2815 ^ n2758;
  assign n2823 = n2822 ^ n2736;
  assign n2824 = n2823 ^ n1496;
  assign n27239 = n27237 ^ n2824;
  assign n27240 = n27238 & n27239;
  assign n27241 = n27240 ^ n2824;
  assign n27103 = n27085 ^ n27038;
  assign n27242 = n27241 ^ n27103;
  assign n27243 = n27241 ^ n1592;
  assign n27244 = n27242 & n27243;
  assign n27245 = n27244 ^ n1592;
  assign n27246 = n27245 ^ n27101;
  assign n27247 = ~n27102 & n27246;
  assign n27248 = n27247 ^ n2955;
  assign n27423 = n27268 ^ n27248;
  assign n27424 = n27268 ^ n27251;
  assign n27425 = ~n27423 & n27424;
  assign n27426 = n27425 ^ n27251;
  assign n27427 = n27426 ^ n27418;
  assign n27428 = n27422 & ~n27427;
  assign n27429 = n27428 ^ n27421;
  assign n27393 = n27391 & ~n27392;
  assign n27374 = n27373 ^ n27369;
  assign n27375 = ~n27370 & ~n27374;
  assign n27376 = n27375 ^ n24148;
  assign n27340 = n27339 ^ n27337;
  assign n27344 = n27343 ^ n27339;
  assign n27345 = ~n27340 & n27344;
  assign n27346 = n27345 ^ n27337;
  assign n27333 = n25532 ^ n24855;
  assign n27334 = n27333 ^ n26186;
  assign n27365 = n27346 ^ n27334;
  assign n27332 = n26633 ^ n2753;
  assign n27366 = n27365 ^ n27332;
  assign n27367 = n27366 ^ n24178;
  assign n27390 = n27376 ^ n27367;
  assign n27417 = n27393 ^ n27390;
  assign n27430 = n27429 ^ n27417;
  assign n27469 = n27433 ^ n27430;
  assign n27465 = n25928 ^ n25135;
  assign n27466 = n26729 ^ n25928;
  assign n27467 = n27465 & n27466;
  assign n27468 = n27467 ^ n25135;
  assign n27583 = n27469 ^ n27468;
  assign n27765 = n27583 ^ n24884;
  assign n2197 = n2157 ^ n2108;
  assign n2198 = n2197 ^ n2191;
  assign n2202 = n2201 ^ n2198;
  assign n28246 = n27765 ^ n2202;
  assign n28729 = n28246 ^ n27315;
  assign n28730 = ~n28728 & ~n28729;
  assign n28731 = n28730 ^ n26721;
  assign n27283 = n26265 ^ n25962;
  assign n27284 = n26685 ^ n26265;
  assign n27285 = n27283 & n27284;
  assign n27286 = n27285 ^ n25962;
  assign n27282 = n27190 ^ n774;
  assign n27287 = n27286 ^ n27282;
  assign n27290 = n25890 ^ n25860;
  assign n27291 = n26890 ^ n25890;
  assign n27292 = ~n27290 & ~n27291;
  assign n27293 = n27292 ^ n25860;
  assign n27288 = n27186 ^ n3293;
  assign n27289 = n27288 ^ n27184;
  assign n27294 = n27293 ^ n27289;
  assign n27296 = n25895 ^ n25606;
  assign n27297 = n26691 ^ n25895;
  assign n27298 = n27296 & ~n27297;
  assign n27299 = n27298 ^ n25606;
  assign n27295 = n27181 ^ n27178;
  assign n27300 = n27299 ^ n27295;
  assign n27302 = n25900 ^ n25082;
  assign n27303 = n26695 ^ n25900;
  assign n27304 = n27302 & ~n27303;
  assign n27305 = n27304 ^ n25082;
  assign n27301 = n27174 ^ n27171;
  assign n27306 = n27305 ^ n27301;
  assign n27310 = n26235 ^ n25101;
  assign n27311 = n26703 ^ n26235;
  assign n27312 = n27310 & ~n27311;
  assign n27313 = n27312 ^ n25101;
  assign n27316 = n27315 ^ n27313;
  assign n27318 = n25905 ^ n25108;
  assign n27319 = n26862 ^ n25905;
  assign n27320 = ~n27318 & n27319;
  assign n27321 = n27320 ^ n25108;
  assign n27317 = n27149 ^ n27148;
  assign n27322 = n27321 ^ n27317;
  assign n27453 = n25912 ^ n25118;
  assign n27454 = n26712 ^ n25912;
  assign n27455 = n27453 & n27454;
  assign n27456 = n27455 ^ n25118;
  assign n27358 = n26647 ^ n26645;
  assign n27359 = n27358 ^ n26642;
  assign n27356 = n26177 ^ n24255;
  assign n27357 = n27356 ^ n25138;
  assign n27360 = n27359 ^ n27357;
  assign n27326 = n26639 ^ n26499;
  assign n27324 = n25526 ^ n24843;
  assign n27325 = n27324 ^ n26195;
  assign n27327 = n27326 ^ n27325;
  assign n27330 = n26636 ^ n26501;
  assign n27328 = n26190 ^ n24848;
  assign n27329 = n27328 ^ n25552;
  assign n27331 = n27330 ^ n27329;
  assign n27335 = n27334 ^ n27332;
  assign n27347 = n27346 ^ n27332;
  assign n27348 = n27335 & ~n27347;
  assign n27349 = n27348 ^ n27334;
  assign n27350 = n27349 ^ n27330;
  assign n27351 = n27331 & n27350;
  assign n27352 = n27351 ^ n27329;
  assign n27353 = n27352 ^ n27325;
  assign n27354 = n27327 & n27353;
  assign n27355 = n27354 ^ n27326;
  assign n27449 = n27359 ^ n27355;
  assign n27450 = ~n27360 & n27449;
  assign n27451 = n27450 ^ n27357;
  assign n27377 = n27376 ^ n27366;
  assign n27378 = n27367 & ~n27377;
  assign n27379 = n27378 ^ n24178;
  assign n27395 = n27379 ^ n24232;
  assign n27362 = n27349 ^ n27329;
  assign n27363 = n27362 ^ n27330;
  assign n27396 = n27395 ^ n27363;
  assign n27394 = ~n27390 & n27393;
  assign n27415 = n27396 ^ n27394;
  assign n27416 = n27415 ^ n1921;
  assign n27434 = n27433 ^ n27429;
  assign n27435 = ~n27430 & n27434;
  assign n27436 = n27435 ^ n27433;
  assign n27437 = n27436 ^ n27415;
  assign n27438 = n27416 & ~n27437;
  assign n27439 = n27438 ^ n1921;
  assign n27384 = n27352 ^ n27327;
  assign n27398 = n27384 ^ n24364;
  assign n27364 = n27363 ^ n24232;
  assign n27380 = n27379 ^ n27363;
  assign n27381 = ~n27364 & ~n27380;
  assign n27382 = n27381 ^ n24232;
  assign n27399 = n27398 ^ n27382;
  assign n27397 = ~n27394 & ~n27396;
  assign n27414 = n27399 ^ n27397;
  assign n27440 = n27439 ^ n27414;
  assign n27441 = n27439 ^ n1931;
  assign n27442 = n27440 & n27441;
  assign n27443 = n27442 ^ n1931;
  assign n27400 = ~n27397 & ~n27399;
  assign n27383 = n27382 ^ n24364;
  assign n27385 = n27384 ^ n27382;
  assign n27386 = ~n27383 & ~n27385;
  assign n27387 = n27386 ^ n24364;
  assign n27388 = n27387 ^ n24341;
  assign n27361 = n27360 ^ n27355;
  assign n27389 = n27388 ^ n27361;
  assign n27413 = n27400 ^ n27389;
  assign n27444 = n27443 ^ n27413;
  assign n2048 = n2033 ^ n1976;
  assign n2049 = n2048 ^ n1938;
  assign n2053 = n2052 ^ n2049;
  assign n27445 = n27413 ^ n2053;
  assign n27446 = n27444 & ~n27445;
  assign n27447 = n27446 ^ n2053;
  assign n27408 = n27361 ^ n24341;
  assign n27409 = n27387 ^ n27361;
  assign n27410 = ~n27408 & n27409;
  assign n27411 = n27410 ^ n24341;
  assign n27406 = n26650 ^ n26494;
  assign n27401 = n27389 & n27400;
  assign n27402 = n27401 ^ n26171;
  assign n2060 = n2030 ^ n1971;
  assign n2061 = n2060 ^ n2057;
  assign n2065 = n2064 ^ n2061;
  assign n27403 = n27402 ^ n2065;
  assign n27404 = n27403 ^ n26733;
  assign n27405 = n27404 ^ n25137;
  assign n27407 = n27406 ^ n27405;
  assign n27412 = n27411 ^ n27407;
  assign n27448 = n27447 ^ n27412;
  assign n27452 = n27451 ^ n27448;
  assign n27457 = n27456 ^ n27452;
  assign n27459 = n25916 ^ n25577;
  assign n27460 = n26717 ^ n25916;
  assign n27461 = n27459 & ~n27460;
  assign n27462 = n27461 ^ n25577;
  assign n27458 = n27444 ^ n2053;
  assign n27463 = n27462 ^ n27458;
  assign n27471 = n25924 ^ n25130;
  assign n27472 = n26725 ^ n25924;
  assign n27473 = n27471 & n27472;
  assign n27474 = n27473 ^ n25130;
  assign n27470 = n27468 & n27469;
  assign n27475 = n27474 ^ n27470;
  assign n27476 = n27436 ^ n27416;
  assign n27477 = n27476 ^ n27474;
  assign n27478 = n27475 & ~n27477;
  assign n27479 = n27478 ^ n27470;
  assign n27464 = n27440 ^ n1931;
  assign n27480 = n27479 ^ n27464;
  assign n27481 = n25921 ^ n25124;
  assign n27482 = n26721 ^ n25921;
  assign n27483 = ~n27481 & ~n27482;
  assign n27484 = n27483 ^ n25124;
  assign n27485 = n27484 ^ n27464;
  assign n27486 = n27480 & ~n27485;
  assign n27487 = n27486 ^ n27484;
  assign n27488 = n27487 ^ n27458;
  assign n27489 = ~n27463 & n27488;
  assign n27490 = n27489 ^ n27462;
  assign n27491 = n27490 ^ n27456;
  assign n27492 = ~n27457 & n27491;
  assign n27493 = n27492 ^ n27452;
  assign n27323 = n27047 ^ n2222;
  assign n27494 = n27493 ^ n27323;
  assign n27495 = n25908 ^ n25113;
  assign n27496 = n26706 ^ n25908;
  assign n27497 = ~n27495 & ~n27496;
  assign n27498 = n27497 ^ n25113;
  assign n27499 = n27498 ^ n27323;
  assign n27500 = n27494 & n27499;
  assign n27501 = n27500 ^ n27498;
  assign n27502 = n27501 ^ n27321;
  assign n27503 = ~n27322 & ~n27502;
  assign n27504 = n27503 ^ n27317;
  assign n27505 = n27504 ^ n27313;
  assign n27506 = ~n27316 & n27505;
  assign n27507 = n27506 ^ n27315;
  assign n27309 = n27160 ^ n27159;
  assign n27508 = n27507 ^ n27309;
  assign n27509 = n26243 ^ n25093;
  assign n27510 = n26700 ^ n26243;
  assign n27511 = n27509 & n27510;
  assign n27512 = n27511 ^ n25093;
  assign n27513 = n27512 ^ n27507;
  assign n27514 = n27508 & n27513;
  assign n27515 = n27514 ^ n27309;
  assign n27307 = n27167 ^ n27163;
  assign n27308 = n27307 ^ n27138;
  assign n27516 = n27515 ^ n27308;
  assign n27517 = n25902 ^ n25088;
  assign n27518 = n26698 ^ n25902;
  assign n27519 = n27517 & ~n27518;
  assign n27520 = n27519 ^ n25088;
  assign n27521 = n27520 ^ n27308;
  assign n27522 = ~n27516 & n27521;
  assign n27523 = n27522 ^ n27520;
  assign n27524 = n27523 ^ n27305;
  assign n27525 = n27306 & n27524;
  assign n27526 = n27525 ^ n27301;
  assign n27527 = n27526 ^ n27295;
  assign n27528 = ~n27300 & ~n27527;
  assign n27529 = n27528 ^ n27299;
  assign n27530 = n27529 ^ n27289;
  assign n27531 = n27294 & ~n27530;
  assign n27532 = n27531 ^ n27293;
  assign n27533 = n27532 ^ n27282;
  assign n27534 = ~n27287 & n27533;
  assign n27535 = n27534 ^ n27286;
  assign n27277 = n25958 ^ n25885;
  assign n27278 = n26681 ^ n25885;
  assign n27279 = ~n27277 & n27278;
  assign n27280 = n27279 ^ n25958;
  assign n27276 = n27194 ^ n787;
  assign n27281 = n27280 ^ n27276;
  assign n27564 = n27535 ^ n27281;
  assign n27565 = n27564 ^ n25089;
  assign n27566 = n27532 ^ n27287;
  assign n27567 = n27566 ^ n25094;
  assign n27568 = n27526 ^ n27300;
  assign n27569 = n27568 ^ n25104;
  assign n27570 = n27520 ^ n27516;
  assign n27571 = n27570 ^ n25116;
  assign n27573 = n27501 ^ n27322;
  assign n27574 = n27573 ^ n25127;
  assign n27575 = n27498 ^ n27494;
  assign n27576 = n27575 ^ n25077;
  assign n27577 = n27490 ^ n27457;
  assign n27578 = n27577 ^ n24982;
  assign n27579 = n27487 ^ n27462;
  assign n27580 = n27579 ^ n27458;
  assign n27581 = n27580 ^ n24949;
  assign n27584 = n24884 & n27583;
  assign n27585 = n27584 ^ n24245;
  assign n27586 = n27476 ^ n27475;
  assign n27587 = n27586 ^ n27584;
  assign n27588 = n27585 & ~n27587;
  assign n27589 = n27588 ^ n24245;
  assign n27582 = n27484 ^ n27480;
  assign n27590 = n27589 ^ n27582;
  assign n27591 = n27582 ^ n24896;
  assign n27592 = n27590 & ~n27591;
  assign n27593 = n27592 ^ n24896;
  assign n27594 = n27593 ^ n27580;
  assign n27595 = n27581 & n27594;
  assign n27596 = n27595 ^ n24949;
  assign n27597 = n27596 ^ n27577;
  assign n27598 = ~n27578 & ~n27597;
  assign n27599 = n27598 ^ n24982;
  assign n27600 = n27599 ^ n27575;
  assign n27601 = ~n27576 & ~n27600;
  assign n27602 = n27601 ^ n25077;
  assign n27603 = n27602 ^ n27573;
  assign n27604 = ~n27574 & n27603;
  assign n27605 = n27604 ^ n25127;
  assign n27572 = n27504 ^ n27316;
  assign n27606 = n27605 ^ n27572;
  assign n27607 = n27572 ^ n25122;
  assign n27608 = ~n27606 & ~n27607;
  assign n27609 = n27608 ^ n25122;
  assign n27610 = n27609 ^ n25178;
  assign n27611 = n27512 ^ n27309;
  assign n27612 = n27611 ^ n27507;
  assign n27613 = n27612 ^ n27609;
  assign n27614 = n27610 & n27613;
  assign n27615 = n27614 ^ n25178;
  assign n27616 = n27615 ^ n27570;
  assign n27617 = n27571 & ~n27616;
  assign n27618 = n27617 ^ n25116;
  assign n27619 = n27618 ^ n25111;
  assign n27620 = n27523 ^ n27306;
  assign n27621 = n27620 ^ n27618;
  assign n27622 = n27619 & ~n27621;
  assign n27623 = n27622 ^ n25111;
  assign n27624 = n27623 ^ n27568;
  assign n27625 = ~n27569 & ~n27624;
  assign n27626 = n27625 ^ n25104;
  assign n27627 = n27626 ^ n25099;
  assign n27628 = n27529 ^ n27294;
  assign n27629 = n27628 ^ n27626;
  assign n27630 = n27627 & n27629;
  assign n27631 = n27630 ^ n25099;
  assign n27632 = n27631 ^ n27566;
  assign n27633 = n27567 & ~n27632;
  assign n27634 = n27633 ^ n25094;
  assign n27635 = n27634 ^ n27564;
  assign n27636 = ~n27565 & ~n27635;
  assign n27637 = n27636 ^ n25089;
  assign n27540 = n25897 ^ n25876;
  assign n27541 = n26903 ^ n25876;
  assign n27542 = n27540 & ~n27541;
  assign n27543 = n27542 ^ n25897;
  assign n27536 = n27535 ^ n27276;
  assign n27537 = ~n27281 & ~n27536;
  assign n27538 = n27537 ^ n27280;
  assign n27275 = n27197 ^ n27133;
  assign n27539 = n27538 ^ n27275;
  assign n27563 = n27543 ^ n27539;
  assign n27638 = n27637 ^ n27563;
  assign n27639 = n27563 ^ n25085;
  assign n27640 = n27638 & n27639;
  assign n27641 = n27640 ^ n25085;
  assign n27677 = n27641 ^ n25162;
  assign n27548 = n25892 ^ n25871;
  assign n27549 = n26679 ^ n25871;
  assign n27550 = ~n27548 & ~n27549;
  assign n27551 = n27550 ^ n25892;
  assign n27544 = n27543 ^ n27275;
  assign n27545 = ~n27539 & n27544;
  assign n27546 = n27545 ^ n27543;
  assign n27274 = n27200 ^ n27131;
  assign n27547 = n27546 ^ n27274;
  assign n27561 = n27551 ^ n27547;
  assign n27678 = n27677 ^ n27561;
  assign n27647 = n27620 ^ n25111;
  assign n27648 = n27647 ^ n27618;
  assign n27649 = n27602 ^ n27574;
  assign n27650 = n27599 ^ n27576;
  assign n27651 = n27590 ^ n24896;
  assign n27652 = n27593 ^ n27581;
  assign n27653 = n27651 & ~n27652;
  assign n27654 = n27596 ^ n24982;
  assign n27655 = n27654 ^ n27577;
  assign n27656 = n27653 & ~n27655;
  assign n27657 = ~n27650 & ~n27656;
  assign n27658 = ~n27649 & ~n27657;
  assign n27659 = n27606 ^ n25122;
  assign n27660 = n27658 & ~n27659;
  assign n27661 = n27612 ^ n27610;
  assign n27662 = ~n27660 & ~n27661;
  assign n27663 = n27615 ^ n27571;
  assign n27664 = n27662 & n27663;
  assign n27665 = ~n27648 & ~n27664;
  assign n27666 = n27623 ^ n27569;
  assign n27667 = n27665 & n27666;
  assign n27668 = n27628 ^ n25099;
  assign n27669 = n27668 ^ n27626;
  assign n27670 = n27667 & ~n27669;
  assign n27671 = n27631 ^ n27567;
  assign n27672 = n27670 & n27671;
  assign n27673 = n27634 ^ n27565;
  assign n27674 = ~n27672 & n27673;
  assign n27675 = n27638 ^ n25085;
  assign n27676 = ~n27674 & ~n27675;
  assign n27719 = n27678 ^ n27676;
  assign n3138 = n2428 ^ n1388;
  assign n3145 = n3144 ^ n3138;
  assign n3146 = n3145 ^ n2480;
  assign n27720 = n27719 ^ n3146;
  assign n27722 = n25835 ^ n2419;
  assign n27723 = n27722 ^ n1300;
  assign n27724 = n27723 ^ n3142;
  assign n27721 = n27675 ^ n27674;
  assign n27725 = n27724 ^ n27721;
  assign n27727 = n27671 ^ n27670;
  assign n1118 = n1099 ^ n1033;
  assign n1119 = n1118 ^ n1115;
  assign n1123 = n1122 ^ n1119;
  assign n27728 = n27727 ^ n1123;
  assign n27729 = n27669 ^ n27667;
  assign n1102 = n1090 ^ n1021;
  assign n1103 = n1102 ^ n993;
  assign n1107 = n1106 ^ n1103;
  assign n27730 = n27729 ^ n1107;
  assign n27732 = n27664 ^ n27648;
  assign n27733 = n27732 ^ n967;
  assign n27734 = n27661 ^ n27660;
  assign n27738 = n27737 ^ n27734;
  assign n27739 = n27659 ^ n27658;
  assign n27743 = n27742 ^ n27739;
  assign n27745 = n25791 ^ n18918;
  assign n27746 = n27745 ^ n22856;
  assign n27747 = n27746 ^ n569;
  assign n27744 = n27657 ^ n27649;
  assign n27748 = n27747 ^ n27744;
  assign n27749 = n27656 ^ n27650;
  assign n706 = n705 ^ n702;
  assign n707 = n706 ^ n548;
  assign n708 = n707 ^ n641;
  assign n27750 = n27749 ^ n708;
  assign n27754 = n27655 ^ n27653;
  assign n27751 = n25763 ^ n18924;
  assign n27752 = n27751 ^ n22842;
  assign n27753 = n27752 ^ n543;
  assign n27755 = n27754 ^ n27753;
  assign n27757 = n25768 ^ n530;
  assign n27758 = n27757 ^ n22327;
  assign n27759 = n27758 ^ n3278;
  assign n27756 = n27652 ^ n27651;
  assign n27760 = n27759 ^ n27756;
  assign n27764 = n27763 ^ n27651;
  assign n27766 = n2202 & n27765;
  assign n2346 = n2310 ^ n2242;
  assign n2347 = n2346 ^ n2343;
  assign n2351 = n2350 ^ n2347;
  assign n27767 = n27766 ^ n2351;
  assign n27768 = n27586 ^ n27585;
  assign n27769 = n27768 ^ n27766;
  assign n27770 = n27767 & ~n27769;
  assign n27771 = n27770 ^ n2351;
  assign n27772 = n27771 ^ n27763;
  assign n27773 = n27764 & ~n27772;
  assign n27774 = n27773 ^ n27651;
  assign n27775 = n27774 ^ n27756;
  assign n27776 = n27760 & ~n27775;
  assign n27777 = n27776 ^ n27759;
  assign n27778 = n27777 ^ n27754;
  assign n27779 = n27755 & ~n27778;
  assign n27780 = n27779 ^ n27753;
  assign n27781 = n27780 ^ n27749;
  assign n27782 = n27750 & ~n27781;
  assign n27783 = n27782 ^ n708;
  assign n27784 = n27783 ^ n27744;
  assign n27785 = ~n27748 & n27784;
  assign n27786 = n27785 ^ n27747;
  assign n27787 = n27786 ^ n27739;
  assign n27788 = n27743 & ~n27787;
  assign n27789 = n27788 ^ n27742;
  assign n27790 = n27789 ^ n27734;
  assign n27791 = n27738 & ~n27790;
  assign n27792 = n27791 ^ n27737;
  assign n27793 = n27792 ^ n3312;
  assign n27794 = n27663 ^ n27662;
  assign n27795 = n27794 ^ n27792;
  assign n27796 = n27793 & ~n27795;
  assign n27797 = n27796 ^ n3312;
  assign n27798 = n27797 ^ n27732;
  assign n27799 = ~n27733 & n27798;
  assign n27800 = n27799 ^ n967;
  assign n27731 = n27666 ^ n27665;
  assign n27801 = n27800 ^ n27731;
  assign n27802 = n27800 ^ n983;
  assign n27803 = n27801 & n27802;
  assign n27804 = n27803 ^ n983;
  assign n27805 = n27804 ^ n27729;
  assign n27806 = n27730 & ~n27805;
  assign n27807 = n27806 ^ n1107;
  assign n27808 = n27807 ^ n27727;
  assign n27809 = ~n27728 & n27808;
  assign n27810 = n27809 ^ n1123;
  assign n27726 = n27673 ^ n27672;
  assign n27811 = n27810 ^ n27726;
  assign n1282 = n1275 ^ n1188;
  assign n1289 = n1288 ^ n1282;
  assign n1293 = n1292 ^ n1289;
  assign n27812 = n27726 ^ n1293;
  assign n27813 = n27811 & ~n27812;
  assign n27814 = n27813 ^ n1293;
  assign n27815 = n27814 ^ n27721;
  assign n27816 = ~n27725 & n27815;
  assign n27817 = n27816 ^ n27724;
  assign n27818 = n27817 ^ n27719;
  assign n27819 = ~n27720 & n27818;
  assign n27820 = n27819 ^ n3146;
  assign n2473 = n2472 ^ n2448;
  assign n2483 = n2482 ^ n2473;
  assign n2484 = n2483 ^ n2460;
  assign n27871 = n27820 ^ n2484;
  assign n27679 = n27676 & n27678;
  assign n27562 = n27561 ^ n25162;
  assign n27642 = n27641 ^ n27561;
  assign n27643 = n27562 & n27642;
  assign n27644 = n27643 ^ n25162;
  assign n27556 = n25887 ^ n25870;
  assign n27557 = n26676 ^ n25870;
  assign n27558 = ~n27556 & n27557;
  assign n27559 = n27558 ^ n25887;
  assign n27552 = n27551 ^ n27274;
  assign n27553 = n27547 & ~n27552;
  assign n27554 = n27553 ^ n27551;
  assign n27273 = n27203 ^ n27126;
  assign n27555 = n27554 ^ n27273;
  assign n27560 = n27559 ^ n27555;
  assign n27645 = n27644 ^ n27560;
  assign n27646 = n27645 ^ n25158;
  assign n27717 = n27679 ^ n27646;
  assign n27872 = n27871 ^ n27717;
  assign n27866 = n27326 ^ n26743;
  assign n27867 = n27238 ^ n2824;
  assign n27868 = n27867 ^ n27326;
  assign n27869 = ~n27866 & n27868;
  assign n27870 = n27869 ^ n26743;
  assign n27873 = n27872 ^ n27870;
  assign n27879 = n27817 ^ n27720;
  assign n27874 = n27330 ^ n26745;
  assign n27875 = n27234 ^ n2729;
  assign n27876 = n27875 ^ n27330;
  assign n27877 = n27874 & n27876;
  assign n27878 = n27877 ^ n26745;
  assign n27880 = n27879 ^ n27878;
  assign n28308 = n27814 ^ n27725;
  assign n27886 = n27811 ^ n1293;
  assign n27881 = n27339 ^ n26429;
  assign n27882 = n27227 ^ n27226;
  assign n27883 = n27882 ^ n27339;
  assign n27884 = n27881 & ~n27883;
  assign n27885 = n27884 ^ n26429;
  assign n27887 = n27886 ^ n27885;
  assign n27893 = n27807 ^ n27728;
  assign n27888 = n27262 ^ n26287;
  assign n27889 = n27222 ^ n27112;
  assign n27890 = n27889 ^ n27262;
  assign n27891 = ~n27888 & ~n27890;
  assign n27892 = n27891 ^ n26287;
  assign n27894 = n27893 ^ n27892;
  assign n27901 = n27804 ^ n1107;
  assign n27902 = n27901 ^ n27729;
  assign n27895 = n27096 ^ n25870;
  assign n27896 = n27219 ^ n27116;
  assign n27897 = n27896 ^ n27113;
  assign n27898 = n27897 ^ n27096;
  assign n27899 = ~n27895 & n27898;
  assign n27900 = n27899 ^ n25870;
  assign n27903 = n27902 ^ n27900;
  assign n28290 = n27801 ^ n983;
  assign n27908 = n27797 ^ n967;
  assign n27909 = n27908 ^ n27732;
  assign n27904 = n26676 ^ n25876;
  assign n27837 = n27213 ^ n1474;
  assign n27905 = n27837 ^ n26676;
  assign n27906 = ~n27904 & ~n27905;
  assign n27907 = n27906 ^ n25876;
  assign n27910 = n27909 ^ n27907;
  assign n27915 = n27794 ^ n27793;
  assign n27911 = n26679 ^ n25885;
  assign n27697 = n27209 ^ n27122;
  assign n27912 = n27697 ^ n26679;
  assign n27913 = n27911 & ~n27912;
  assign n27914 = n27913 ^ n25885;
  assign n27916 = n27915 ^ n27914;
  assign n27918 = n26903 ^ n26265;
  assign n27681 = n27206 ^ n27124;
  assign n27919 = n27681 ^ n26903;
  assign n27920 = ~n27918 & ~n27919;
  assign n27921 = n27920 ^ n26265;
  assign n27917 = n27789 ^ n27738;
  assign n27922 = n27921 ^ n27917;
  assign n27924 = n26681 ^ n25890;
  assign n27925 = n27273 ^ n26681;
  assign n27926 = n27924 & ~n27925;
  assign n27927 = n27926 ^ n25890;
  assign n27923 = n27786 ^ n27743;
  assign n27928 = n27927 ^ n27923;
  assign n27931 = n26685 ^ n25895;
  assign n27932 = n27274 ^ n26685;
  assign n27933 = ~n27931 & n27932;
  assign n27934 = n27933 ^ n25895;
  assign n27929 = n27783 ^ n27747;
  assign n27930 = n27929 ^ n27744;
  assign n27935 = n27934 ^ n27930;
  assign n27937 = n26890 ^ n25900;
  assign n27938 = n27275 ^ n26890;
  assign n27939 = n27937 & ~n27938;
  assign n27940 = n27939 ^ n25900;
  assign n27936 = n27780 ^ n27750;
  assign n27941 = n27940 ^ n27936;
  assign n27946 = n27777 ^ n27755;
  assign n27942 = n26691 ^ n25902;
  assign n27943 = n27276 ^ n26691;
  assign n27944 = n27942 & ~n27943;
  assign n27945 = n27944 ^ n25902;
  assign n27947 = n27946 ^ n27945;
  assign n27950 = n26698 ^ n26235;
  assign n27951 = n27289 ^ n26698;
  assign n27952 = ~n27950 & ~n27951;
  assign n27953 = n27952 ^ n26235;
  assign n27949 = n27771 ^ n27764;
  assign n27954 = n27953 ^ n27949;
  assign n27956 = n26700 ^ n25905;
  assign n27957 = n27295 ^ n26700;
  assign n27958 = n27956 & n27957;
  assign n27959 = n27958 ^ n25905;
  assign n27955 = n27768 ^ n27767;
  assign n27960 = n27959 ^ n27955;
  assign n27975 = n26195 ^ n25532;
  assign n27976 = n26671 ^ n26195;
  assign n27977 = ~n27975 & n27976;
  assign n27978 = n27977 ^ n25532;
  assign n27979 = n27978 ^ n27867;
  assign n27980 = n26190 ^ n25544;
  assign n27981 = n27406 ^ n26190;
  assign n27982 = n27980 & ~n27981;
  assign n27983 = n27982 ^ n25544;
  assign n27984 = n27983 ^ n27875;
  assign n27986 = n26735 ^ n26089;
  assign n27987 = n27326 ^ n26735;
  assign n27988 = n27986 & ~n27987;
  assign n27989 = n27988 ^ n26089;
  assign n27990 = n27989 ^ n27882;
  assign n27991 = n26737 ^ n26005;
  assign n27992 = n27330 ^ n26737;
  assign n27993 = n27991 & ~n27992;
  assign n27994 = n27993 ^ n26005;
  assign n27995 = n27994 ^ n27889;
  assign n27996 = n26743 ^ n25938;
  assign n27997 = n27332 ^ n26743;
  assign n27998 = n27996 & n27997;
  assign n27999 = n27998 ^ n25938;
  assign n28000 = n27999 ^ n27897;
  assign n28003 = n26745 ^ n25872;
  assign n28004 = n27339 ^ n26745;
  assign n28005 = ~n28003 & ~n28004;
  assign n28006 = n28005 ^ n25872;
  assign n28001 = n27216 ^ n3023;
  assign n28002 = n28001 ^ n27118;
  assign n28007 = n28006 ^ n28002;
  assign n27838 = n26664 ^ n25878;
  assign n27839 = n27262 ^ n26664;
  assign n27840 = ~n27838 & n27839;
  assign n27841 = n27840 ^ n25878;
  assign n27842 = n27841 ^ n27837;
  assign n27698 = n26429 ^ n25882;
  assign n27699 = n27096 ^ n26429;
  assign n27700 = n27698 & n27699;
  assign n27701 = n27700 ^ n25882;
  assign n27702 = n27701 ^ n27697;
  assign n27682 = n26287 ^ n25950;
  assign n27683 = n27034 ^ n26287;
  assign n27684 = n27682 & n27683;
  assign n27685 = n27684 ^ n25950;
  assign n27703 = n27685 ^ n27681;
  assign n27686 = n27559 ^ n27273;
  assign n27687 = ~n27555 & ~n27686;
  assign n27688 = n27687 ^ n27559;
  assign n27704 = n27688 ^ n27681;
  assign n27705 = n27703 & n27704;
  assign n27706 = n27705 ^ n27685;
  assign n27834 = n27706 ^ n27697;
  assign n27835 = ~n27702 & n27834;
  assign n27836 = n27835 ^ n27701;
  assign n28008 = n27837 ^ n27836;
  assign n28009 = n27842 & n28008;
  assign n28010 = n28009 ^ n27841;
  assign n28011 = n28010 ^ n28002;
  assign n28012 = n28007 & ~n28011;
  assign n28013 = n28012 ^ n28006;
  assign n28014 = n28013 ^ n27999;
  assign n28015 = n28000 & n28014;
  assign n28016 = n28015 ^ n27897;
  assign n28017 = n28016 ^ n27889;
  assign n28018 = ~n27995 & n28017;
  assign n28019 = n28018 ^ n27994;
  assign n28020 = n28019 ^ n27882;
  assign n28021 = ~n27990 & ~n28020;
  assign n28022 = n28021 ^ n27989;
  assign n27985 = n27230 ^ n27107;
  assign n28023 = n28022 ^ n27985;
  assign n28024 = n26186 ^ n25537;
  assign n28025 = n27359 ^ n26186;
  assign n28026 = ~n28024 & n28025;
  assign n28027 = n28026 ^ n25537;
  assign n28028 = n28027 ^ n27985;
  assign n28029 = ~n28023 & ~n28028;
  assign n28030 = n28029 ^ n28027;
  assign n28031 = n28030 ^ n27875;
  assign n28032 = ~n27984 & n28031;
  assign n28033 = n28032 ^ n27983;
  assign n28034 = n28033 ^ n27867;
  assign n28035 = ~n27979 & ~n28034;
  assign n28036 = n28035 ^ n27978;
  assign n27970 = n26177 ^ n25552;
  assign n27971 = n26826 ^ n26177;
  assign n27972 = n27970 & ~n27971;
  assign n27973 = n27972 ^ n25552;
  assign n28041 = n28036 ^ n27973;
  assign n27859 = n27242 ^ n1592;
  assign n28042 = n28041 ^ n27859;
  assign n28043 = n28042 ^ n24848;
  assign n28044 = n28033 ^ n27978;
  assign n28045 = n28044 ^ n27867;
  assign n28046 = n28045 ^ n24855;
  assign n28047 = n28030 ^ n27984;
  assign n28048 = n28047 ^ n24865;
  assign n28049 = n28027 ^ n28023;
  assign n28050 = n28049 ^ n24857;
  assign n28072 = n28019 ^ n27989;
  assign n28073 = n28072 ^ n27882;
  assign n28051 = n28016 ^ n27994;
  assign n28052 = n28051 ^ n27889;
  assign n28053 = n28052 ^ n25352;
  assign n28054 = n28013 ^ n28000;
  assign n28055 = n28054 ^ n25251;
  assign n28056 = n28010 ^ n28006;
  assign n28057 = n28056 ^ n28002;
  assign n28058 = n28057 ^ n25244;
  assign n27843 = n27842 ^ n27836;
  assign n28059 = n27843 ^ n25143;
  assign n27691 = n27560 ^ n25158;
  assign n27692 = ~n27645 & n27691;
  assign n27693 = n27692 ^ n25158;
  assign n27689 = n27688 ^ n27685;
  assign n27690 = n27689 ^ n27681;
  assign n27694 = n27693 ^ n27690;
  assign n27708 = n27690 ^ n25153;
  assign n27709 = ~n27694 & n27708;
  assign n27710 = n27709 ^ n25153;
  assign n27707 = n27706 ^ n27702;
  assign n27711 = n27710 ^ n27707;
  assign n27830 = n27707 ^ n25147;
  assign n27831 = ~n27711 & ~n27830;
  assign n27832 = n27831 ^ n25147;
  assign n28060 = n27843 ^ n27832;
  assign n28061 = n28059 & ~n28060;
  assign n28062 = n28061 ^ n25143;
  assign n28063 = n28062 ^ n28057;
  assign n28064 = n28058 & n28063;
  assign n28065 = n28064 ^ n25244;
  assign n28066 = n28065 ^ n28054;
  assign n28067 = n28055 & ~n28066;
  assign n28068 = n28067 ^ n25251;
  assign n28069 = n28068 ^ n28052;
  assign n28070 = n28053 & ~n28069;
  assign n28071 = n28070 ^ n25352;
  assign n28074 = n28073 ^ n28071;
  assign n28075 = n28073 ^ n25407;
  assign n28076 = ~n28074 & ~n28075;
  assign n28077 = n28076 ^ n25407;
  assign n28078 = n28077 ^ n28049;
  assign n28079 = n28050 & ~n28078;
  assign n28080 = n28079 ^ n24857;
  assign n28081 = n28080 ^ n28047;
  assign n28082 = ~n28048 & n28081;
  assign n28083 = n28082 ^ n24865;
  assign n28084 = n28083 ^ n28045;
  assign n28085 = n28046 & n28084;
  assign n28086 = n28085 ^ n24855;
  assign n28087 = n28086 ^ n28042;
  assign n28088 = ~n28043 & n28087;
  assign n28089 = n28088 ^ n24848;
  assign n27974 = n27973 ^ n27859;
  assign n28037 = n28036 ^ n27859;
  assign n28038 = ~n27974 & n28037;
  assign n28039 = n28038 ^ n27973;
  assign n27965 = n26171 ^ n25526;
  assign n27966 = n26819 ^ n26171;
  assign n27967 = ~n27965 & n27966;
  assign n27968 = n27967 ^ n25526;
  assign n27851 = n27245 ^ n2955;
  assign n27852 = n27851 ^ n27101;
  assign n27969 = n27968 ^ n27852;
  assign n28040 = n28039 ^ n27969;
  assign n28090 = n28089 ^ n28040;
  assign n28122 = n28040 ^ n24843;
  assign n28123 = ~n28090 & n28122;
  assign n28124 = n28123 ^ n24843;
  assign n28115 = n25936 ^ n25138;
  assign n28116 = n26837 ^ n25936;
  assign n28117 = ~n28115 & ~n28116;
  assign n28118 = n28117 ^ n25138;
  assign n27252 = n27251 ^ n27248;
  assign n27269 = n27268 ^ n27252;
  assign n28119 = n28118 ^ n27269;
  assign n28112 = n28039 ^ n27852;
  assign n28113 = n27969 & n28112;
  assign n28114 = n28113 ^ n27968;
  assign n28120 = n28119 ^ n28114;
  assign n28121 = n28120 ^ n24255;
  assign n28125 = n28124 ^ n28121;
  assign n28091 = n28090 ^ n24843;
  assign n28092 = n28086 ^ n24848;
  assign n28093 = n28092 ^ n28042;
  assign n28094 = n28083 ^ n28046;
  assign n28095 = n28077 ^ n28050;
  assign n28096 = n28074 ^ n25407;
  assign n28097 = n28068 ^ n25352;
  assign n28098 = n28097 ^ n28052;
  assign n28099 = n28065 ^ n28055;
  assign n28100 = n28062 ^ n28058;
  assign n27833 = n27832 ^ n25143;
  assign n27844 = n27843 ^ n27833;
  assign n27680 = ~n27646 & n27679;
  assign n27695 = n27694 ^ n25153;
  assign n27696 = ~n27680 & n27695;
  assign n27712 = n27711 ^ n25147;
  assign n27845 = ~n27696 & n27712;
  assign n28101 = n27844 & n27845;
  assign n28102 = ~n28100 & ~n28101;
  assign n28103 = n28099 & n28102;
  assign n28104 = n28098 & n28103;
  assign n28105 = n28096 & ~n28104;
  assign n28106 = n28095 & n28105;
  assign n28107 = n28080 ^ n28048;
  assign n28108 = n28106 & ~n28107;
  assign n28109 = n28094 & n28108;
  assign n28110 = ~n28093 & ~n28109;
  assign n28111 = n28091 & n28110;
  assign n28145 = n28125 ^ n28111;
  assign n28146 = n28145 ^ n2180;
  assign n28147 = n28110 ^ n28091;
  assign n28151 = n28150 ^ n28147;
  assign n28152 = n28109 ^ n28093;
  assign n28156 = n28155 ^ n28152;
  assign n28159 = n26123 ^ n19280;
  assign n28160 = n28159 ^ n1654;
  assign n28161 = n28160 ^ n1727;
  assign n28158 = n28107 ^ n28106;
  assign n28162 = n28161 ^ n28158;
  assign n28163 = n28105 ^ n28095;
  assign n1630 = n1623 ^ n1547;
  assign n1643 = n1642 ^ n1630;
  assign n1647 = n1646 ^ n1643;
  assign n28164 = n28163 ^ n1647;
  assign n28165 = n28104 ^ n28096;
  assign n28166 = n28165 ^ n2937;
  assign n28167 = n28103 ^ n28098;
  assign n2916 = n2853 ^ n1502;
  assign n2917 = n2916 ^ n2902;
  assign n2921 = n2920 ^ n2917;
  assign n28168 = n28167 ^ n2921;
  assign n28169 = n28102 ^ n28099;
  assign n28170 = n28169 ^ n2911;
  assign n28171 = n28101 ^ n28100;
  assign n28172 = n28171 ^ n3233;
  assign n27846 = n27845 ^ n27844;
  assign n27847 = n27846 ^ n3077;
  assign n27713 = n27712 ^ n27696;
  assign n2538 = n2537 ^ n2504;
  assign n2545 = n2544 ^ n2538;
  assign n2546 = n2545 ^ n1556;
  assign n27714 = n27713 ^ n2546;
  assign n27715 = n27695 ^ n27680;
  assign n3051 = n3050 ^ n3045;
  assign n3052 = n3051 ^ n2465;
  assign n3053 = n3052 ^ n2542;
  assign n27716 = n27715 ^ n3053;
  assign n27718 = n27717 ^ n2484;
  assign n27821 = n27820 ^ n27717;
  assign n27822 = n27718 & ~n27821;
  assign n27823 = n27822 ^ n2484;
  assign n27824 = n27823 ^ n27715;
  assign n27825 = ~n27716 & n27824;
  assign n27826 = n27825 ^ n3053;
  assign n27827 = n27826 ^ n27713;
  assign n27828 = n27714 & ~n27827;
  assign n27829 = n27828 ^ n2546;
  assign n28173 = n27846 ^ n27829;
  assign n28174 = ~n27847 & n28173;
  assign n28175 = n28174 ^ n3077;
  assign n28176 = n28175 ^ n28171;
  assign n28177 = n28172 & ~n28176;
  assign n28178 = n28177 ^ n3233;
  assign n28179 = n28178 ^ n2911;
  assign n28180 = n28170 & ~n28179;
  assign n28181 = n28180 ^ n28169;
  assign n28182 = n28181 ^ n28167;
  assign n28183 = n28168 & ~n28182;
  assign n28184 = n28183 ^ n2921;
  assign n28185 = n28184 ^ n28165;
  assign n28186 = n28166 & ~n28185;
  assign n28187 = n28186 ^ n2937;
  assign n28188 = n28187 ^ n28163;
  assign n28189 = ~n28164 & n28188;
  assign n28190 = n28189 ^ n1647;
  assign n28191 = n28190 ^ n28158;
  assign n28192 = n28162 & ~n28191;
  assign n28193 = n28192 ^ n28161;
  assign n28157 = n28108 ^ n28094;
  assign n28194 = n28193 ^ n28157;
  assign n1723 = n1722 ^ n1670;
  assign n1730 = n1729 ^ n1723;
  assign n1731 = n1730 ^ n1703;
  assign n28195 = n28157 ^ n1731;
  assign n28196 = n28194 & ~n28195;
  assign n28197 = n28196 ^ n1731;
  assign n28198 = n28197 ^ n28155;
  assign n28199 = n28156 & ~n28198;
  assign n28200 = n28199 ^ n28152;
  assign n28201 = n28200 ^ n28147;
  assign n28202 = n28151 & ~n28201;
  assign n28203 = n28202 ^ n28150;
  assign n28204 = n28203 ^ n28145;
  assign n28205 = ~n28146 & n28204;
  assign n28206 = n28205 ^ n2180;
  assign n28139 = n28124 ^ n28120;
  assign n28140 = ~n28121 & ~n28139;
  assign n28141 = n28140 ^ n24255;
  assign n28133 = n28114 ^ n27269;
  assign n28134 = ~n28119 & n28133;
  assign n28135 = n28134 ^ n28118;
  assign n28129 = n25932 ^ n25137;
  assign n28130 = n26815 ^ n25932;
  assign n28131 = n28129 & n28130;
  assign n28132 = n28131 ^ n25137;
  assign n28136 = n28135 ^ n28132;
  assign n28127 = n27426 ^ n27421;
  assign n28128 = n28127 ^ n27418;
  assign n28137 = n28136 ^ n28128;
  assign n28138 = n28137 ^ n24250;
  assign n28142 = n28141 ^ n28138;
  assign n28126 = n28111 & ~n28125;
  assign n28143 = n28142 ^ n28126;
  assign n2162 = n2142 ^ n2089;
  assign n2166 = n2165 ^ n2162;
  assign n2170 = n2169 ^ n2166;
  assign n28144 = n28143 ^ n2170;
  assign n28207 = n28206 ^ n28144;
  assign n27961 = n26862 ^ n25912;
  assign n27962 = n27308 ^ n26862;
  assign n27963 = n27961 & n27962;
  assign n27964 = n27963 ^ n25912;
  assign n28208 = n28207 ^ n27964;
  assign n28213 = n28203 ^ n28146;
  assign n28209 = n26706 ^ n25916;
  assign n28210 = n27309 ^ n26706;
  assign n28211 = n28209 & ~n28210;
  assign n28212 = n28211 ^ n25916;
  assign n28214 = n28213 ^ n28212;
  assign n28219 = n28200 ^ n28150;
  assign n28220 = n28219 ^ n28147;
  assign n28215 = n26712 ^ n25921;
  assign n28216 = n27315 ^ n26712;
  assign n28217 = ~n28215 & ~n28216;
  assign n28218 = n28217 ^ n25921;
  assign n28221 = n28220 ^ n28218;
  assign n28226 = n28194 ^ n1731;
  assign n28227 = n26721 ^ n25928;
  assign n28228 = n27323 ^ n26721;
  assign n28229 = ~n28227 & ~n28228;
  assign n28230 = n28229 ^ n25928;
  assign n28231 = ~n28226 & n28230;
  assign n28222 = n26717 ^ n25924;
  assign n28223 = n27317 ^ n26717;
  assign n28224 = n28222 & ~n28223;
  assign n28225 = n28224 ^ n25924;
  assign n28232 = n28231 ^ n28225;
  assign n28233 = n28197 ^ n28156;
  assign n28234 = n28233 ^ n28231;
  assign n28235 = n28232 & ~n28234;
  assign n28236 = n28235 ^ n28225;
  assign n28237 = n28236 ^ n28220;
  assign n28238 = ~n28221 & ~n28237;
  assign n28239 = n28238 ^ n28218;
  assign n28240 = n28239 ^ n28213;
  assign n28241 = ~n28214 & ~n28240;
  assign n28242 = n28241 ^ n28212;
  assign n28243 = n28242 ^ n28207;
  assign n28244 = n28208 & n28243;
  assign n28245 = n28244 ^ n27964;
  assign n28247 = n28246 ^ n28245;
  assign n28248 = n26703 ^ n25908;
  assign n28249 = n27301 ^ n26703;
  assign n28250 = ~n28248 & ~n28249;
  assign n28251 = n28250 ^ n25908;
  assign n28252 = n28251 ^ n28245;
  assign n28253 = ~n28247 & n28252;
  assign n28254 = n28253 ^ n28246;
  assign n28255 = n28254 ^ n27955;
  assign n28256 = n27960 & ~n28255;
  assign n28257 = n28256 ^ n27959;
  assign n28258 = n28257 ^ n27949;
  assign n28259 = ~n27954 & ~n28258;
  assign n28260 = n28259 ^ n27953;
  assign n27948 = n27774 ^ n27760;
  assign n28261 = n28260 ^ n27948;
  assign n28262 = n26695 ^ n26243;
  assign n28263 = n27282 ^ n26695;
  assign n28264 = n28262 & ~n28263;
  assign n28265 = n28264 ^ n26243;
  assign n28266 = n28265 ^ n28260;
  assign n28267 = ~n28261 & ~n28266;
  assign n28268 = n28267 ^ n27948;
  assign n28269 = n28268 ^ n27946;
  assign n28270 = n27947 & ~n28269;
  assign n28271 = n28270 ^ n27945;
  assign n28272 = n28271 ^ n27940;
  assign n28273 = ~n27941 & n28272;
  assign n28274 = n28273 ^ n27936;
  assign n28275 = n28274 ^ n27934;
  assign n28276 = ~n27935 & ~n28275;
  assign n28277 = n28276 ^ n27930;
  assign n28278 = n28277 ^ n27927;
  assign n28279 = ~n27928 & ~n28278;
  assign n28280 = n28279 ^ n27923;
  assign n28281 = n28280 ^ n27921;
  assign n28282 = n27922 & ~n28281;
  assign n28283 = n28282 ^ n27917;
  assign n28284 = n28283 ^ n27915;
  assign n28285 = n27916 & ~n28284;
  assign n28286 = n28285 ^ n27914;
  assign n28287 = n28286 ^ n27909;
  assign n28288 = n27910 & n28287;
  assign n28289 = n28288 ^ n27907;
  assign n28291 = n28290 ^ n28289;
  assign n28292 = n27034 ^ n25871;
  assign n28293 = n28002 ^ n27034;
  assign n28294 = n28292 & ~n28293;
  assign n28295 = n28294 ^ n25871;
  assign n28296 = n28295 ^ n28290;
  assign n28297 = ~n28291 & ~n28296;
  assign n28298 = n28297 ^ n28295;
  assign n28299 = n28298 ^ n27902;
  assign n28300 = ~n27903 & ~n28299;
  assign n28301 = n28300 ^ n27900;
  assign n28302 = n28301 ^ n27892;
  assign n28303 = n27894 & ~n28302;
  assign n28304 = n28303 ^ n27893;
  assign n28305 = n28304 ^ n27886;
  assign n28306 = n27887 & ~n28305;
  assign n28307 = n28306 ^ n27885;
  assign n28309 = n28308 ^ n28307;
  assign n28310 = n27332 ^ n26664;
  assign n28311 = n27985 ^ n27332;
  assign n28312 = ~n28310 & ~n28311;
  assign n28313 = n28312 ^ n26664;
  assign n28314 = n28313 ^ n28308;
  assign n28315 = ~n28309 & n28314;
  assign n28316 = n28315 ^ n28313;
  assign n28317 = n28316 ^ n27879;
  assign n28318 = n27880 & ~n28317;
  assign n28319 = n28318 ^ n27878;
  assign n28320 = n28319 ^ n27872;
  assign n28321 = ~n27873 & n28320;
  assign n28322 = n28321 ^ n27870;
  assign n27858 = n27359 ^ n26737;
  assign n27860 = n27859 ^ n27359;
  assign n27861 = n27858 & ~n27860;
  assign n27862 = n27861 ^ n26737;
  assign n28342 = n28322 ^ n27862;
  assign n27863 = n27823 ^ n3053;
  assign n27864 = n27863 ^ n27715;
  assign n28343 = n28342 ^ n27864;
  assign n28344 = n28343 ^ n26005;
  assign n28345 = n28319 ^ n27870;
  assign n28346 = n28345 ^ n27872;
  assign n28347 = n28346 ^ n25938;
  assign n28348 = n28316 ^ n27878;
  assign n28349 = n28348 ^ n27879;
  assign n28350 = n28349 ^ n25872;
  assign n28351 = n28313 ^ n28309;
  assign n28352 = n28351 ^ n25878;
  assign n28353 = n28304 ^ n27885;
  assign n28354 = n28353 ^ n27886;
  assign n28355 = n28354 ^ n25882;
  assign n28356 = n28301 ^ n27894;
  assign n28357 = n28356 ^ n25950;
  assign n28358 = n28298 ^ n27903;
  assign n28359 = n28358 ^ n25887;
  assign n28360 = n28295 ^ n28291;
  assign n28361 = n28360 ^ n25892;
  assign n28364 = n28283 ^ n27916;
  assign n28365 = n28364 ^ n25958;
  assign n28432 = n28280 ^ n27922;
  assign n28366 = n28277 ^ n27928;
  assign n28367 = n28366 ^ n25860;
  assign n28368 = n28274 ^ n27935;
  assign n28369 = n28368 ^ n25606;
  assign n28370 = n28271 ^ n27941;
  assign n28371 = n28370 ^ n25082;
  assign n28372 = n28268 ^ n27947;
  assign n28373 = n28372 ^ n25088;
  assign n28374 = n28265 ^ n27948;
  assign n28375 = n28374 ^ n28260;
  assign n28376 = n28375 ^ n25093;
  assign n28377 = n28257 ^ n27953;
  assign n28378 = n28377 ^ n27949;
  assign n28379 = n28378 ^ n25101;
  assign n28382 = n28242 ^ n28208;
  assign n28383 = n28382 ^ n25118;
  assign n28384 = n28239 ^ n28214;
  assign n28385 = n28384 ^ n25577;
  assign n28386 = n28230 ^ n28226;
  assign n28387 = n25135 & ~n28386;
  assign n28388 = n28387 ^ n25130;
  assign n28389 = n28233 ^ n28232;
  assign n28390 = n28389 ^ n28387;
  assign n28391 = n28388 & ~n28390;
  assign n28392 = n28391 ^ n25130;
  assign n28393 = n28392 ^ n25124;
  assign n28394 = n28236 ^ n28221;
  assign n28395 = n28394 ^ n28392;
  assign n28396 = n28393 & n28395;
  assign n28397 = n28396 ^ n25124;
  assign n28398 = n28397 ^ n28384;
  assign n28399 = n28385 & ~n28398;
  assign n28400 = n28399 ^ n25577;
  assign n28401 = n28400 ^ n28382;
  assign n28402 = ~n28383 & ~n28401;
  assign n28403 = n28402 ^ n25118;
  assign n28380 = n28251 ^ n28246;
  assign n28381 = n28380 ^ n28245;
  assign n28404 = n28403 ^ n28381;
  assign n28405 = n28381 ^ n25113;
  assign n28406 = ~n28404 & n28405;
  assign n28407 = n28406 ^ n25113;
  assign n28408 = n28407 ^ n25108;
  assign n28409 = n28254 ^ n27959;
  assign n28410 = n28409 ^ n27955;
  assign n28411 = n28410 ^ n28407;
  assign n28412 = n28408 & n28411;
  assign n28413 = n28412 ^ n25108;
  assign n28414 = n28413 ^ n28378;
  assign n28415 = n28379 & ~n28414;
  assign n28416 = n28415 ^ n25101;
  assign n28417 = n28416 ^ n28375;
  assign n28418 = ~n28376 & n28417;
  assign n28419 = n28418 ^ n25093;
  assign n28420 = n28419 ^ n28372;
  assign n28421 = n28373 & n28420;
  assign n28422 = n28421 ^ n25088;
  assign n28423 = n28422 ^ n28370;
  assign n28424 = n28371 & n28423;
  assign n28425 = n28424 ^ n25082;
  assign n28426 = n28425 ^ n28368;
  assign n28427 = ~n28369 & ~n28426;
  assign n28428 = n28427 ^ n25606;
  assign n28429 = n28428 ^ n28366;
  assign n28430 = n28367 & ~n28429;
  assign n28431 = n28430 ^ n25860;
  assign n28433 = n28432 ^ n28431;
  assign n28434 = n28431 ^ n25962;
  assign n28435 = ~n28433 & n28434;
  assign n28436 = n28435 ^ n25962;
  assign n28437 = n28436 ^ n28364;
  assign n28438 = ~n28365 & ~n28437;
  assign n28439 = n28438 ^ n25958;
  assign n28362 = n28286 ^ n27907;
  assign n28363 = n28362 ^ n27909;
  assign n28440 = n28439 ^ n28363;
  assign n28441 = n28363 ^ n25897;
  assign n28442 = n28440 & ~n28441;
  assign n28443 = n28442 ^ n25897;
  assign n28444 = n28443 ^ n28360;
  assign n28445 = ~n28361 & n28444;
  assign n28446 = n28445 ^ n25892;
  assign n28447 = n28446 ^ n28358;
  assign n28448 = ~n28359 & ~n28447;
  assign n28449 = n28448 ^ n25887;
  assign n28450 = n28449 ^ n28356;
  assign n28451 = n28357 & n28450;
  assign n28452 = n28451 ^ n25950;
  assign n28453 = n28452 ^ n28354;
  assign n28454 = n28355 & ~n28453;
  assign n28455 = n28454 ^ n25882;
  assign n28456 = n28455 ^ n28351;
  assign n28457 = ~n28352 & ~n28456;
  assign n28458 = n28457 ^ n25878;
  assign n28459 = n28458 ^ n28349;
  assign n28460 = ~n28350 & n28459;
  assign n28461 = n28460 ^ n25872;
  assign n28462 = n28461 ^ n28346;
  assign n28463 = ~n28347 & ~n28462;
  assign n28464 = n28463 ^ n25938;
  assign n28465 = n28464 ^ n28343;
  assign n28466 = n28344 & ~n28465;
  assign n28467 = n28466 ^ n26005;
  assign n27865 = n27864 ^ n27862;
  assign n28323 = n28322 ^ n27864;
  assign n28324 = n27865 & ~n28323;
  assign n28325 = n28324 ^ n27862;
  assign n27856 = n27826 ^ n27714;
  assign n27850 = n27406 ^ n26735;
  assign n27853 = n27852 ^ n27406;
  assign n27854 = ~n27850 & ~n27853;
  assign n27855 = n27854 ^ n26735;
  assign n27857 = n27856 ^ n27855;
  assign n28341 = n28325 ^ n27857;
  assign n28468 = n28467 ^ n28341;
  assign n28495 = n28468 ^ n26089;
  assign n28496 = n28464 ^ n28344;
  assign n28497 = n28458 ^ n25872;
  assign n28498 = n28497 ^ n28349;
  assign n28499 = n28455 ^ n25878;
  assign n28500 = n28499 ^ n28351;
  assign n28501 = n28452 ^ n25882;
  assign n28502 = n28501 ^ n28354;
  assign n28503 = n28428 ^ n28367;
  assign n28504 = n28422 ^ n28371;
  assign n28505 = n28410 ^ n25108;
  assign n28506 = n28505 ^ n28407;
  assign n28507 = n28404 ^ n25113;
  assign n28508 = n28400 ^ n28383;
  assign n28509 = n28394 ^ n28393;
  assign n28510 = n28397 ^ n28385;
  assign n28511 = n28509 & ~n28510;
  assign n28512 = n28508 & n28511;
  assign n28513 = ~n28507 & ~n28512;
  assign n28514 = ~n28506 & ~n28513;
  assign n28515 = n28413 ^ n28379;
  assign n28516 = n28514 & n28515;
  assign n28517 = n28416 ^ n28376;
  assign n28518 = ~n28516 & n28517;
  assign n28519 = n28419 ^ n28373;
  assign n28520 = n28518 & ~n28519;
  assign n28521 = ~n28504 & ~n28520;
  assign n28522 = n28425 ^ n28369;
  assign n28523 = n28521 & ~n28522;
  assign n28524 = ~n28503 & n28523;
  assign n28525 = n28432 ^ n25962;
  assign n28526 = n28525 ^ n28431;
  assign n28527 = n28524 & ~n28526;
  assign n28528 = n28436 ^ n25958;
  assign n28529 = n28528 ^ n28364;
  assign n28530 = ~n28527 & ~n28529;
  assign n28531 = n28440 ^ n25897;
  assign n28532 = ~n28530 & ~n28531;
  assign n28533 = n28443 ^ n25892;
  assign n28534 = n28533 ^ n28360;
  assign n28535 = n28532 & ~n28534;
  assign n28536 = n28446 ^ n28359;
  assign n28537 = n28535 & ~n28536;
  assign n28538 = n28449 ^ n25950;
  assign n28539 = n28538 ^ n28356;
  assign n28540 = ~n28537 & n28539;
  assign n28541 = n28502 & ~n28540;
  assign n28542 = ~n28500 & n28541;
  assign n28543 = ~n28498 & ~n28542;
  assign n28544 = n28461 ^ n28347;
  assign n28545 = n28543 & ~n28544;
  assign n28546 = ~n28496 & n28545;
  assign n28547 = ~n28495 & ~n28546;
  assign n28326 = n28325 ^ n27856;
  assign n28327 = ~n27857 & ~n28326;
  assign n28328 = n28327 ^ n28325;
  assign n27848 = n27847 ^ n27829;
  assign n26672 = n26671 ^ n26186;
  assign n27270 = n27269 ^ n26671;
  assign n27271 = n26672 & ~n27270;
  assign n27272 = n27271 ^ n26186;
  assign n27849 = n27848 ^ n27272;
  assign n28473 = n28328 ^ n27849;
  assign n28548 = n28473 ^ n25537;
  assign n28469 = n28341 ^ n26089;
  assign n28470 = ~n28468 & ~n28469;
  assign n28471 = n28470 ^ n26089;
  assign n28549 = n28548 ^ n28471;
  assign n28550 = n28547 & n28549;
  assign n28472 = n28471 ^ n25537;
  assign n28474 = n28473 ^ n28471;
  assign n28475 = ~n28472 & ~n28474;
  assign n28476 = n28475 ^ n25537;
  assign n28493 = n28476 ^ n25544;
  assign n28337 = n28175 ^ n3233;
  assign n28338 = n28337 ^ n28171;
  assign n28332 = n26826 ^ n26190;
  assign n28333 = n28128 ^ n26826;
  assign n28334 = ~n28332 & ~n28333;
  assign n28335 = n28334 ^ n26190;
  assign n28329 = n28328 ^ n27848;
  assign n28330 = ~n27849 & ~n28329;
  assign n28331 = n28330 ^ n27272;
  assign n28336 = n28335 ^ n28331;
  assign n28339 = n28338 ^ n28336;
  assign n28494 = n28493 ^ n28339;
  assign n28553 = n28550 ^ n28494;
  assign n28557 = n28556 ^ n28553;
  assign n28558 = n28549 ^ n28547;
  assign n28562 = n28561 ^ n28558;
  assign n28563 = n28546 ^ n28495;
  assign n28567 = n28566 ^ n28563;
  assign n28568 = n28545 ^ n28496;
  assign n28569 = n28568 ^ n2819;
  assign n28570 = n28544 ^ n28543;
  assign n28571 = n28570 ^ n3110;
  assign n28572 = n28542 ^ n28498;
  assign n2695 = n2691 ^ n2643;
  assign n2699 = n2698 ^ n2695;
  assign n2700 = n2699 ^ n1524;
  assign n28573 = n28572 ^ n2700;
  assign n28574 = n28541 ^ n28500;
  assign n2618 = n2572 ^ n1559;
  assign n2619 = n2618 ^ n2601;
  assign n2623 = n2622 ^ n2619;
  assign n28575 = n28574 ^ n2623;
  assign n28576 = n28540 ^ n28502;
  assign n2603 = n2584 ^ n2560;
  assign n2613 = n2612 ^ n2603;
  assign n2614 = n2613 ^ n2596;
  assign n28577 = n28576 ^ n2614;
  assign n28578 = n28539 ^ n28537;
  assign n3169 = n3165 ^ n2522;
  assign n3176 = n3175 ^ n3169;
  assign n3177 = n3176 ^ n2609;
  assign n28579 = n28578 ^ n3177;
  assign n28580 = n28536 ^ n28535;
  assign n28584 = n28583 ^ n28580;
  assign n28586 = n26606 ^ n3151;
  assign n28587 = n28586 ^ n1435;
  assign n28588 = n28587 ^ n3020;
  assign n28585 = n28534 ^ n28532;
  assign n28589 = n28588 ^ n28585;
  assign n28590 = n28531 ^ n28530;
  assign n1422 = n1400 ^ n1316;
  assign n1423 = n1422 ^ n1419;
  assign n1427 = n1426 ^ n1423;
  assign n28591 = n28590 ^ n1427;
  assign n28592 = n28529 ^ n28527;
  assign n1258 = n1215 ^ n1167;
  assign n1259 = n1258 ^ n1252;
  assign n1263 = n1262 ^ n1259;
  assign n28593 = n28592 ^ n1263;
  assign n28594 = n28526 ^ n28524;
  assign n1240 = n1200 ^ n1136;
  assign n1241 = n1240 ^ n1237;
  assign n1245 = n1244 ^ n1241;
  assign n28595 = n28594 ^ n1245;
  assign n28596 = n28523 ^ n28503;
  assign n1222 = n1147 ^ n1066;
  assign n1229 = n1228 ^ n1222;
  assign n1230 = n1229 ^ n1001;
  assign n28597 = n28596 ^ n1230;
  assign n28600 = n28519 ^ n28518;
  assign n28601 = n28600 ^ n761;
  assign n28605 = n28517 ^ n28516;
  assign n28602 = n26531 ^ n19692;
  assign n28603 = n28602 ^ n659;
  assign n28604 = n28603 ^ n751;
  assign n28606 = n28605 ^ n28604;
  assign n28608 = n28513 ^ n28506;
  assign n28612 = n28611 ^ n28608;
  assign n28614 = n26544 ^ n558;
  assign n28615 = n28614 ^ n23106;
  assign n28616 = n28615 ^ n3254;
  assign n28613 = n28512 ^ n28507;
  assign n28617 = n28616 ^ n28613;
  assign n28619 = n26556 ^ n19663;
  assign n28620 = n28619 ^ n23097;
  assign n28621 = n28620 ^ n18394;
  assign n28618 = n28510 ^ n28509;
  assign n28622 = n28621 ^ n28618;
  assign n28629 = n28386 ^ n25135;
  assign n28630 = n28628 & ~n28629;
  assign n28623 = n2370 ^ n2297;
  assign n28624 = n28623 ^ n2228;
  assign n28625 = n28624 ^ n687;
  assign n28631 = n28630 ^ n28625;
  assign n28632 = n28389 ^ n28388;
  assign n28633 = n28632 ^ n28625;
  assign n28634 = n28631 & ~n28633;
  assign n28635 = n28634 ^ n28630;
  assign n28636 = n28635 ^ n28509;
  assign n28637 = n19668 ^ n2393;
  assign n28638 = n28637 ^ n23088;
  assign n28639 = n28638 ^ n18399;
  assign n28640 = n28639 ^ n28635;
  assign n28641 = ~n28636 & n28640;
  assign n28642 = n28641 ^ n28639;
  assign n28643 = n28642 ^ n28618;
  assign n28644 = n28622 & ~n28643;
  assign n28645 = n28644 ^ n28621;
  assign n28649 = n28648 ^ n28645;
  assign n28650 = n28511 ^ n28508;
  assign n28651 = n28650 ^ n28648;
  assign n28652 = n28649 & n28651;
  assign n28653 = n28652 ^ n28645;
  assign n28654 = n28653 ^ n28613;
  assign n28655 = n28617 & ~n28654;
  assign n28656 = n28655 ^ n28616;
  assign n28657 = n28656 ^ n28608;
  assign n28658 = ~n28612 & n28657;
  assign n28659 = n28658 ^ n28611;
  assign n28607 = n28515 ^ n28514;
  assign n28660 = n28659 ^ n28607;
  assign n588 = n587 ^ n581;
  assign n601 = n600 ^ n588;
  assign n605 = n604 ^ n601;
  assign n28661 = n28607 ^ n605;
  assign n28662 = n28660 & ~n28661;
  assign n28663 = n28662 ^ n605;
  assign n28664 = n28663 ^ n28604;
  assign n28665 = ~n28606 & ~n28664;
  assign n28666 = n28665 ^ n28605;
  assign n28667 = n28666 ^ n28600;
  assign n28668 = ~n28601 & ~n28667;
  assign n28669 = n28668 ^ n761;
  assign n28599 = n28520 ^ n28504;
  assign n28670 = n28669 ^ n28599;
  assign n28674 = n28673 ^ n28599;
  assign n28675 = n28670 & ~n28674;
  assign n28676 = n28675 ^ n28673;
  assign n28598 = n28522 ^ n28521;
  assign n28677 = n28676 ^ n28598;
  assign n28678 = n28598 ^ n3337;
  assign n28679 = ~n28677 & n28678;
  assign n28680 = n28679 ^ n3337;
  assign n28681 = n28680 ^ n28596;
  assign n28682 = n28597 & ~n28681;
  assign n28683 = n28682 ^ n1230;
  assign n28684 = n28683 ^ n28594;
  assign n28685 = n28595 & ~n28684;
  assign n28686 = n28685 ^ n1245;
  assign n28687 = n28686 ^ n28592;
  assign n28688 = n28593 & ~n28687;
  assign n28689 = n28688 ^ n1263;
  assign n28690 = n28689 ^ n28590;
  assign n28691 = ~n28591 & n28690;
  assign n28692 = n28691 ^ n1427;
  assign n28693 = n28692 ^ n28585;
  assign n28694 = n28589 & ~n28693;
  assign n28695 = n28694 ^ n28588;
  assign n28696 = n28695 ^ n28580;
  assign n28697 = n28584 & ~n28696;
  assign n28698 = n28697 ^ n28583;
  assign n28699 = n28698 ^ n28578;
  assign n28700 = ~n28579 & n28699;
  assign n28701 = n28700 ^ n3177;
  assign n28702 = n28701 ^ n28576;
  assign n28703 = n28577 & ~n28702;
  assign n28704 = n28703 ^ n2614;
  assign n28705 = n28704 ^ n28574;
  assign n28706 = n28575 & ~n28705;
  assign n28707 = n28706 ^ n2623;
  assign n28708 = n28707 ^ n28572;
  assign n28709 = n28573 & ~n28708;
  assign n28710 = n28709 ^ n2700;
  assign n28711 = n28710 ^ n28570;
  assign n28712 = ~n28571 & n28711;
  assign n28713 = n28712 ^ n3110;
  assign n28714 = n28713 ^ n28568;
  assign n28715 = ~n28569 & n28714;
  assign n28716 = n28715 ^ n2819;
  assign n28717 = n28716 ^ n28563;
  assign n28718 = ~n28567 & n28717;
  assign n28719 = n28718 ^ n28566;
  assign n28720 = n28719 ^ n28558;
  assign n28721 = ~n28562 & n28720;
  assign n28722 = n28721 ^ n28561;
  assign n28723 = n28722 ^ n28553;
  assign n28724 = ~n28557 & n28723;
  assign n28725 = n28724 ^ n28556;
  assign n28551 = n28494 & n28550;
  assign n28485 = n26819 ^ n26195;
  assign n28486 = n27469 ^ n26819;
  assign n28487 = n28485 & n28486;
  assign n28488 = n28487 ^ n26195;
  assign n28484 = n28178 ^ n28170;
  assign n28489 = n28488 ^ n28484;
  assign n28480 = n28338 ^ n28335;
  assign n28481 = n28338 ^ n28331;
  assign n28482 = ~n28480 & ~n28481;
  assign n28483 = n28482 ^ n28335;
  assign n28490 = n28489 ^ n28483;
  assign n28491 = n28490 ^ n25532;
  assign n28340 = n28339 ^ n25544;
  assign n28477 = n28476 ^ n28339;
  assign n28478 = n28340 & ~n28477;
  assign n28479 = n28478 ^ n25544;
  assign n28492 = n28491 ^ n28479;
  assign n28552 = n28551 ^ n28492;
  assign n28726 = n28725 ^ n28552;
  assign n1775 = n1756 ^ n1742;
  assign n1785 = n1784 ^ n1775;
  assign n1786 = n1785 ^ n1774;
  assign n28727 = n28726 ^ n1786;
  assign n28732 = n28731 ^ n28727;
  assign n28765 = n25928 & n28732;
  assign n28766 = n28765 ^ n25924;
  assign n28759 = n27309 ^ n26717;
  assign n28760 = n27955 ^ n27309;
  assign n28761 = n28759 & ~n28760;
  assign n28762 = n28761 ^ n26717;
  assign n28758 = ~n28727 & ~n28731;
  assign n28763 = n28762 ^ n28758;
  assign n28750 = n28181 ^ n28168;
  assign n28746 = n26837 ^ n26177;
  assign n28747 = n27476 ^ n26837;
  assign n28748 = n28746 & ~n28747;
  assign n28749 = n28748 ^ n26177;
  assign n28751 = n28750 ^ n28749;
  assign n28743 = n28484 ^ n28483;
  assign n28744 = ~n28489 & n28743;
  assign n28745 = n28744 ^ n28488;
  assign n28752 = n28751 ^ n28745;
  assign n28753 = n28752 ^ n25552;
  assign n28740 = n28490 ^ n28479;
  assign n28741 = n28491 & n28740;
  assign n28742 = n28741 ^ n25532;
  assign n28754 = n28753 ^ n28742;
  assign n28739 = n28492 & n28551;
  assign n28755 = n28754 ^ n28739;
  assign n1796 = n1765 ^ n1715;
  assign n1797 = n1796 ^ n1793;
  assign n1801 = n1800 ^ n1797;
  assign n28756 = n28755 ^ n1801;
  assign n28736 = n28552 ^ n1786;
  assign n28737 = n28726 & ~n28736;
  assign n28738 = n28737 ^ n1786;
  assign n28757 = n28756 ^ n28738;
  assign n28764 = n28763 ^ n28757;
  assign n28802 = n28765 ^ n28764;
  assign n28803 = n28766 & ~n28802;
  assign n28804 = n28803 ^ n25924;
  assign n28790 = n26815 ^ n26171;
  assign n28791 = n27464 ^ n26815;
  assign n28792 = ~n28790 & ~n28791;
  assign n28793 = n28792 ^ n26171;
  assign n28789 = n28184 ^ n28166;
  assign n28794 = n28793 ^ n28789;
  assign n28786 = n28750 ^ n28745;
  assign n28787 = n28751 & n28786;
  assign n28788 = n28787 ^ n28749;
  assign n28795 = n28794 ^ n28788;
  assign n28782 = n28752 ^ n28742;
  assign n28783 = ~n28753 & n28782;
  assign n28784 = n28783 ^ n25552;
  assign n28785 = n28784 ^ n25526;
  assign n28796 = n28795 ^ n28785;
  assign n28781 = ~n28739 & ~n28754;
  assign n28797 = n28796 ^ n28781;
  assign n1885 = n1877 ^ n1827;
  assign n1892 = n1891 ^ n1885;
  assign n1896 = n1895 ^ n1892;
  assign n28798 = n28797 ^ n1896;
  assign n28778 = n28755 ^ n28738;
  assign n28779 = n28756 & ~n28778;
  assign n28780 = n28779 ^ n1801;
  assign n28799 = n28798 ^ n28780;
  assign n28774 = n27308 ^ n26712;
  assign n28775 = n27949 ^ n27308;
  assign n28776 = n28774 & ~n28775;
  assign n28777 = n28776 ^ n26712;
  assign n28800 = n28799 ^ n28777;
  assign n28771 = n28762 ^ n28757;
  assign n28772 = n28763 & ~n28771;
  assign n28773 = n28772 ^ n28758;
  assign n28801 = n28800 ^ n28773;
  assign n28805 = n28804 ^ n28801;
  assign n28806 = n28805 ^ n25921;
  assign n28810 = n28809 ^ n28806;
  assign n2153 = n2117 ^ n2065;
  assign n2154 = n2153 ^ n2150;
  assign n2158 = n2157 ^ n2154;
  assign n28733 = n28732 ^ n25928;
  assign n28734 = n2158 & n28733;
  assign n2322 = n2321 ^ n2222;
  assign n2323 = n2322 ^ n2318;
  assign n2324 = n2323 ^ n2310;
  assign n28735 = n28734 ^ n2324;
  assign n28767 = n28766 ^ n28764;
  assign n28768 = n28767 ^ n2324;
  assign n28769 = n28735 & ~n28768;
  assign n28770 = n28769 ^ n28734;
  assign n28811 = n28810 ^ n28770;
  assign n30524 = n28625 ^ n2405;
  assign n30525 = n30524 ^ n2330;
  assign n30526 = n30525 ^ n690;
  assign n29137 = n27889 ^ n27034;
  assign n29138 = n27889 ^ n27879;
  assign n29139 = n29137 & n29138;
  assign n29140 = n29139 ^ n27034;
  assign n29136 = n28677 ^ n3337;
  assign n29141 = n29140 ^ n29136;
  assign n29143 = n27897 ^ n26676;
  assign n29144 = n28308 ^ n27897;
  assign n29145 = ~n29143 & ~n29144;
  assign n29146 = n29145 ^ n26676;
  assign n29142 = n28673 ^ n28670;
  assign n29147 = n29146 ^ n29142;
  assign n29149 = n28002 ^ n26679;
  assign n29150 = n28002 ^ n27886;
  assign n29151 = n29149 & n29150;
  assign n29152 = n29151 ^ n26679;
  assign n29148 = n28666 ^ n28601;
  assign n29153 = n29152 ^ n29148;
  assign n29155 = n27837 ^ n26903;
  assign n29156 = n27893 ^ n27837;
  assign n29157 = ~n29155 & n29156;
  assign n29158 = n29157 ^ n26903;
  assign n29154 = n28663 ^ n28606;
  assign n29159 = n29158 ^ n29154;
  assign n29086 = n28659 ^ n605;
  assign n29087 = n29086 ^ n28607;
  assign n29081 = n27697 ^ n26681;
  assign n29082 = n27902 ^ n27697;
  assign n29083 = ~n29081 & ~n29082;
  assign n29084 = n29083 ^ n26681;
  assign n29160 = n29087 ^ n29084;
  assign n28987 = n27681 ^ n26685;
  assign n28988 = n28290 ^ n27681;
  assign n28989 = n28987 & ~n28988;
  assign n28990 = n28989 ^ n26685;
  assign n28986 = n28656 ^ n28612;
  assign n28991 = n28990 ^ n28986;
  assign n28822 = n27274 ^ n26691;
  assign n28823 = n27915 ^ n27274;
  assign n28824 = n28822 & ~n28823;
  assign n28825 = n28824 ^ n26691;
  assign n28821 = n28650 ^ n28649;
  assign n28826 = n28825 ^ n28821;
  assign n28831 = n28642 ^ n28621;
  assign n28832 = n28831 ^ n28618;
  assign n28827 = n27275 ^ n26695;
  assign n28828 = n27917 ^ n27275;
  assign n28829 = n28827 & n28828;
  assign n28830 = n28829 ^ n26695;
  assign n28833 = n28832 ^ n28830;
  assign n28921 = n28639 ^ n28636;
  assign n28838 = n28632 ^ n28631;
  assign n28834 = n27282 ^ n26700;
  assign n28835 = n27930 ^ n27282;
  assign n28836 = ~n28834 & ~n28835;
  assign n28837 = n28836 ^ n26700;
  assign n28839 = n28838 ^ n28837;
  assign n28844 = n28629 ^ n28628;
  assign n28840 = n27289 ^ n26703;
  assign n28841 = n27936 ^ n27289;
  assign n28842 = ~n28840 & ~n28841;
  assign n28843 = n28842 ^ n26703;
  assign n28845 = n28844 ^ n28843;
  assign n28895 = n27295 ^ n26862;
  assign n28896 = n27946 ^ n27295;
  assign n28897 = n28895 & n28896;
  assign n28898 = n28897 ^ n26862;
  assign n28883 = n26798 ^ n2264;
  assign n28884 = n28883 ^ n1903;
  assign n28885 = n28884 ^ n2033;
  assign n28862 = n28781 & ~n28796;
  assign n28855 = n28789 ^ n28788;
  assign n28856 = n28794 & ~n28855;
  assign n28857 = n28856 ^ n28793;
  assign n28851 = n26729 ^ n25936;
  assign n28852 = n27458 ^ n26729;
  assign n28853 = ~n28851 & ~n28852;
  assign n28854 = n28853 ^ n25936;
  assign n28858 = n28857 ^ n28854;
  assign n28850 = n28187 ^ n28164;
  assign n28859 = n28858 ^ n28850;
  assign n28860 = n28859 ^ n25138;
  assign n28846 = n28795 ^ n25526;
  assign n28847 = n28795 ^ n28784;
  assign n28848 = ~n28846 & ~n28847;
  assign n28849 = n28848 ^ n25526;
  assign n28861 = n28860 ^ n28849;
  assign n28882 = n28862 ^ n28861;
  assign n28886 = n28885 ^ n28882;
  assign n28887 = n28797 ^ n28780;
  assign n28888 = ~n28798 & n28887;
  assign n28889 = n28888 ^ n1896;
  assign n28890 = n28889 ^ n28882;
  assign n28891 = ~n28886 & n28890;
  assign n28892 = n28891 ^ n28885;
  assign n2043 = n2042 ^ n1958;
  assign n2044 = n2043 ^ n2039;
  assign n2045 = n2044 ^ n2030;
  assign n28893 = n28892 ^ n2045;
  assign n28875 = n28849 ^ n25138;
  assign n28876 = n28859 ^ n28849;
  assign n28877 = n28875 & ~n28876;
  assign n28878 = n28877 ^ n25138;
  assign n28870 = n26725 ^ n25932;
  assign n28871 = n27452 ^ n26725;
  assign n28872 = ~n28870 & n28871;
  assign n28873 = n28872 ^ n25932;
  assign n28865 = n28854 ^ n28850;
  assign n28866 = n28857 ^ n28850;
  assign n28867 = ~n28865 & n28866;
  assign n28868 = n28867 ^ n28854;
  assign n28864 = n28190 ^ n28162;
  assign n28869 = n28868 ^ n28864;
  assign n28874 = n28873 ^ n28869;
  assign n28879 = n28878 ^ n28874;
  assign n28880 = n28879 ^ n25137;
  assign n28863 = ~n28861 & n28862;
  assign n28881 = n28880 ^ n28863;
  assign n28894 = n28893 ^ n28881;
  assign n28899 = n28898 ^ n28894;
  assign n28901 = n27301 ^ n26706;
  assign n28902 = n27948 ^ n27301;
  assign n28903 = ~n28901 & n28902;
  assign n28904 = n28903 ^ n26706;
  assign n28900 = n28889 ^ n28886;
  assign n28905 = n28904 ^ n28900;
  assign n28906 = n28799 ^ n28773;
  assign n28907 = ~n28800 & n28906;
  assign n28908 = n28907 ^ n28777;
  assign n28909 = n28908 ^ n28900;
  assign n28910 = ~n28905 & n28909;
  assign n28911 = n28910 ^ n28904;
  assign n28912 = n28911 ^ n28894;
  assign n28913 = ~n28899 & ~n28912;
  assign n28914 = n28913 ^ n28898;
  assign n28915 = n28914 ^ n28844;
  assign n28916 = n28845 & ~n28915;
  assign n28917 = n28916 ^ n28843;
  assign n28918 = n28917 ^ n28838;
  assign n28919 = n28839 & n28918;
  assign n28920 = n28919 ^ n28837;
  assign n28922 = n28921 ^ n28920;
  assign n28923 = n27276 ^ n26698;
  assign n28924 = n27923 ^ n27276;
  assign n28925 = n28923 & ~n28924;
  assign n28926 = n28925 ^ n26698;
  assign n28927 = n28926 ^ n28921;
  assign n28928 = ~n28922 & n28927;
  assign n28929 = n28928 ^ n28926;
  assign n28930 = n28929 ^ n28832;
  assign n28931 = ~n28833 & ~n28930;
  assign n28932 = n28931 ^ n28830;
  assign n28933 = n28932 ^ n28825;
  assign n28934 = ~n28826 & n28933;
  assign n28935 = n28934 ^ n28821;
  assign n28819 = n28653 ^ n28617;
  assign n28982 = n28935 ^ n28819;
  assign n28815 = n27273 ^ n26890;
  assign n28816 = n27909 ^ n27273;
  assign n28817 = n28815 & ~n28816;
  assign n28818 = n28817 ^ n26890;
  assign n28983 = n28935 ^ n28818;
  assign n28984 = ~n28982 & ~n28983;
  assign n28985 = n28984 ^ n28819;
  assign n29078 = n28986 ^ n28985;
  assign n29079 = n28991 & n29078;
  assign n29080 = n29079 ^ n28990;
  assign n29161 = n29087 ^ n29080;
  assign n29162 = n29160 & ~n29161;
  assign n29163 = n29162 ^ n29084;
  assign n29164 = n29163 ^ n29154;
  assign n29165 = n29159 & ~n29164;
  assign n29166 = n29165 ^ n29158;
  assign n29167 = n29166 ^ n29148;
  assign n29168 = n29153 & n29167;
  assign n29169 = n29168 ^ n29152;
  assign n29170 = n29169 ^ n29142;
  assign n29171 = ~n29147 & n29170;
  assign n29172 = n29171 ^ n29146;
  assign n29173 = n29172 ^ n29140;
  assign n29174 = n29141 & ~n29173;
  assign n29175 = n29174 ^ n29136;
  assign n29132 = n27882 ^ n27096;
  assign n29133 = n27882 ^ n27872;
  assign n29134 = ~n29132 & n29133;
  assign n29135 = n29134 ^ n27096;
  assign n29176 = n29175 ^ n29135;
  assign n29177 = n28680 ^ n1230;
  assign n29178 = n29177 ^ n28596;
  assign n29179 = n29178 ^ n29175;
  assign n29180 = ~n29176 & n29179;
  assign n29181 = n29180 ^ n29178;
  assign n29127 = n27985 ^ n27262;
  assign n29128 = n27985 ^ n27864;
  assign n29129 = n29127 & n29128;
  assign n29130 = n29129 ^ n27262;
  assign n29101 = n28683 ^ n28595;
  assign n29131 = n29130 ^ n29101;
  assign n29239 = n29181 ^ n29131;
  assign n29240 = n29239 ^ n26287;
  assign n29241 = n29178 ^ n29135;
  assign n29242 = n29241 ^ n29175;
  assign n29243 = n29242 ^ n25870;
  assign n29244 = n29172 ^ n29141;
  assign n29245 = n29244 ^ n25871;
  assign n29246 = n29169 ^ n29147;
  assign n29247 = n29246 ^ n25876;
  assign n29250 = n29163 ^ n29158;
  assign n29251 = n29250 ^ n29154;
  assign n29252 = n29251 ^ n26265;
  assign n29085 = n29084 ^ n29080;
  assign n29088 = n29087 ^ n29085;
  assign n29089 = n29088 ^ n25890;
  assign n28992 = n28991 ^ n28985;
  assign n28993 = n28992 ^ n25895;
  assign n28820 = n28819 ^ n28818;
  assign n28936 = n28935 ^ n28820;
  assign n28937 = n28936 ^ n25900;
  assign n28938 = n28929 ^ n28830;
  assign n28939 = n28938 ^ n28832;
  assign n28940 = n28939 ^ n26243;
  assign n28943 = n28914 ^ n28845;
  assign n28944 = n28943 ^ n25908;
  assign n28945 = n28911 ^ n28898;
  assign n28946 = n28945 ^ n28894;
  assign n28947 = n28946 ^ n25912;
  assign n28948 = n28908 ^ n28904;
  assign n28949 = n28948 ^ n28900;
  assign n28950 = n28949 ^ n25916;
  assign n28951 = n28801 ^ n25921;
  assign n28952 = n28805 & n28951;
  assign n28953 = n28952 ^ n25921;
  assign n28954 = n28953 ^ n28949;
  assign n28955 = ~n28950 & ~n28954;
  assign n28956 = n28955 ^ n25916;
  assign n28957 = n28956 ^ n28946;
  assign n28958 = n28947 & n28957;
  assign n28959 = n28958 ^ n25912;
  assign n28960 = n28959 ^ n28943;
  assign n28961 = ~n28944 & ~n28960;
  assign n28962 = n28961 ^ n25908;
  assign n28942 = n28917 ^ n28839;
  assign n28963 = n28962 ^ n28942;
  assign n28964 = n28942 ^ n25905;
  assign n28965 = n28963 & ~n28964;
  assign n28966 = n28965 ^ n25905;
  assign n28941 = n28926 ^ n28922;
  assign n28967 = n28966 ^ n28941;
  assign n28968 = n28941 ^ n26235;
  assign n28969 = ~n28967 & ~n28968;
  assign n28970 = n28969 ^ n26235;
  assign n28971 = n28970 ^ n28939;
  assign n28972 = n28940 & ~n28971;
  assign n28973 = n28972 ^ n26243;
  assign n28974 = n28973 ^ n25902;
  assign n28975 = n28932 ^ n28826;
  assign n28976 = n28975 ^ n28973;
  assign n28977 = ~n28974 & n28976;
  assign n28978 = n28977 ^ n25902;
  assign n28979 = n28978 ^ n28936;
  assign n28980 = ~n28937 & ~n28979;
  assign n28981 = n28980 ^ n25900;
  assign n29075 = n28992 ^ n28981;
  assign n29076 = n28993 & n29075;
  assign n29077 = n29076 ^ n25895;
  assign n29253 = n29088 ^ n29077;
  assign n29254 = n29089 & n29253;
  assign n29255 = n29254 ^ n25890;
  assign n29256 = n29255 ^ n29251;
  assign n29257 = ~n29252 & ~n29256;
  assign n29258 = n29257 ^ n26265;
  assign n29248 = n29166 ^ n29152;
  assign n29249 = n29248 ^ n29148;
  assign n29259 = n29258 ^ n29249;
  assign n29260 = n29249 ^ n25885;
  assign n29261 = n29259 & ~n29260;
  assign n29262 = n29261 ^ n25885;
  assign n29263 = n29262 ^ n29246;
  assign n29264 = n29247 & n29263;
  assign n29265 = n29264 ^ n25876;
  assign n29266 = n29265 ^ n29244;
  assign n29267 = n29245 & n29266;
  assign n29268 = n29267 ^ n25871;
  assign n29269 = n29268 ^ n29242;
  assign n29270 = ~n29243 & ~n29269;
  assign n29271 = n29270 ^ n25870;
  assign n29272 = n29271 ^ n29239;
  assign n29273 = ~n29240 & n29272;
  assign n29274 = n29273 ^ n26287;
  assign n29186 = n27875 ^ n27339;
  assign n29187 = n27875 ^ n27856;
  assign n29188 = ~n29186 & ~n29187;
  assign n29189 = n29188 ^ n27339;
  assign n28812 = n28686 ^ n1263;
  assign n28813 = n28812 ^ n28592;
  assign n29236 = n29189 ^ n28813;
  assign n29182 = n29181 ^ n29101;
  assign n29183 = n29131 & ~n29182;
  assign n29184 = n29183 ^ n29130;
  assign n29237 = n29236 ^ n29184;
  assign n29238 = n29237 ^ n26429;
  assign n29330 = n29274 ^ n29238;
  assign n29331 = n29265 ^ n29245;
  assign n29332 = n29262 ^ n29247;
  assign n29333 = n29259 ^ n25885;
  assign n29090 = n29089 ^ n29077;
  assign n28994 = n28993 ^ n28981;
  assign n28995 = n28975 ^ n25902;
  assign n28996 = n28995 ^ n28973;
  assign n28997 = n28970 ^ n28940;
  assign n28998 = n28953 ^ n28950;
  assign n28999 = ~n28806 & ~n28998;
  assign n29000 = n28956 ^ n28947;
  assign n29001 = n28999 & ~n29000;
  assign n29002 = n28959 ^ n28944;
  assign n29003 = ~n29001 & n29002;
  assign n29004 = n28963 ^ n25905;
  assign n29005 = ~n29003 & n29004;
  assign n29006 = n28967 ^ n26235;
  assign n29007 = n29005 & n29006;
  assign n29008 = ~n28997 & ~n29007;
  assign n29009 = ~n28996 & n29008;
  assign n29010 = n28978 ^ n28937;
  assign n29011 = ~n29009 & n29010;
  assign n29091 = n28994 & n29011;
  assign n29334 = ~n29090 & n29091;
  assign n29335 = n29255 ^ n29252;
  assign n29336 = n29334 & ~n29335;
  assign n29337 = ~n29333 & ~n29336;
  assign n29338 = ~n29332 & ~n29337;
  assign n29339 = n29331 & n29338;
  assign n29340 = n29268 ^ n29243;
  assign n29341 = n29339 & n29340;
  assign n29342 = n29271 ^ n29240;
  assign n29343 = ~n29341 & n29342;
  assign n29344 = n29330 & ~n29343;
  assign n29275 = n29274 ^ n29237;
  assign n29276 = n29238 & ~n29275;
  assign n29277 = n29276 ^ n26429;
  assign n29194 = n27867 ^ n27332;
  assign n29195 = n27867 ^ n27848;
  assign n29196 = ~n29194 & ~n29195;
  assign n29197 = n29196 ^ n27332;
  assign n29185 = n29184 ^ n28813;
  assign n29190 = n29189 ^ n29184;
  assign n29191 = n29185 & n29190;
  assign n29192 = n29191 ^ n28813;
  assign n29126 = n28689 ^ n28591;
  assign n29193 = n29192 ^ n29126;
  assign n29234 = n29197 ^ n29193;
  assign n29235 = n29234 ^ n26664;
  assign n29329 = n29277 ^ n29235;
  assign n29400 = n29344 ^ n29329;
  assign n3206 = n3199 ^ n2664;
  assign n3210 = n3209 ^ n3206;
  assign n3211 = n3210 ^ n2774;
  assign n29401 = n29400 ^ n3211;
  assign n29402 = n29343 ^ n29330;
  assign n29406 = n29405 ^ n29402;
  assign n29408 = n27116 ^ n3185;
  assign n29409 = n29408 ^ n2491;
  assign n29410 = n29409 ^ n3050;
  assign n29407 = n29342 ^ n29341;
  assign n29411 = n29410 ^ n29407;
  assign n29412 = n29340 ^ n29339;
  assign n3030 = n3029 ^ n3023;
  assign n3034 = n3033 ^ n3030;
  assign n3035 = n3034 ^ n2472;
  assign n29413 = n29412 ^ n3035;
  assign n29414 = n29338 ^ n29331;
  assign n2415 = n2414 ^ n1474;
  assign n2425 = n2424 ^ n2415;
  assign n2429 = n2428 ^ n2425;
  assign n29415 = n29414 ^ n2429;
  assign n29419 = n29337 ^ n29332;
  assign n29416 = n1459 ^ n1370;
  assign n29417 = n29416 ^ n1280;
  assign n29418 = n29417 ^ n2419;
  assign n29420 = n29419 ^ n29418;
  assign n29422 = n1450 ^ n1352;
  assign n29423 = n29422 ^ n24072;
  assign n29424 = n29423 ^ n1275;
  assign n29421 = n29336 ^ n29333;
  assign n29425 = n29424 ^ n29421;
  assign n29426 = n29335 ^ n29334;
  assign n1086 = n1085 ^ n1013;
  assign n1096 = n1095 ^ n1086;
  assign n1100 = n1099 ^ n1096;
  assign n29427 = n29426 ^ n1100;
  assign n29093 = n27130 ^ n1334;
  assign n29094 = n29093 ^ n949;
  assign n29095 = n29094 ^ n1090;
  assign n29092 = n29091 ^ n29090;
  assign n29096 = n29095 ^ n29092;
  assign n29012 = n29011 ^ n28994;
  assign n937 = n936 ^ n873;
  assign n941 = n940 ^ n937;
  assign n942 = n941 ^ n924;
  assign n29013 = n29012 ^ n942;
  assign n29016 = n29007 ^ n28997;
  assign n29017 = n29016 ^ n3296;
  assign n29018 = n29006 ^ n29005;
  assign n29022 = n29021 ^ n29018;
  assign n29023 = n29004 ^ n29003;
  assign n29027 = n29026 ^ n29023;
  assign n29029 = n27167 ^ n20269;
  assign n29030 = n29029 ^ n23688;
  assign n29031 = n29030 ^ n705;
  assign n29028 = n29002 ^ n29001;
  assign n29032 = n29031 ^ n29028;
  assign n29037 = n27142 ^ n20279;
  assign n29038 = n29037 ^ n23700;
  assign n29039 = n29038 ^ n530;
  assign n29036 = n28998 ^ n28806;
  assign n29040 = n29039 ^ n29036;
  assign n29041 = n28806 ^ n28770;
  assign n29042 = ~n28810 & n29041;
  assign n29043 = n29042 ^ n28809;
  assign n29044 = n29043 ^ n29036;
  assign n29045 = ~n29040 & n29044;
  assign n29046 = n29045 ^ n29039;
  assign n29033 = n27158 ^ n20274;
  assign n29034 = n29033 ^ n696;
  assign n29035 = n29034 ^ n18924;
  assign n29047 = n29046 ^ n29035;
  assign n29048 = n29000 ^ n28999;
  assign n29049 = n29048 ^ n29046;
  assign n29050 = n29047 & ~n29049;
  assign n29051 = n29050 ^ n29035;
  assign n29052 = n29051 ^ n29028;
  assign n29053 = ~n29032 & n29052;
  assign n29054 = n29053 ^ n29031;
  assign n29055 = n29054 ^ n29023;
  assign n29056 = n29027 & ~n29055;
  assign n29057 = n29056 ^ n29026;
  assign n29058 = n29057 ^ n29018;
  assign n29059 = ~n29022 & n29058;
  assign n29060 = n29059 ^ n29021;
  assign n29061 = n29060 ^ n3296;
  assign n29062 = n29017 & ~n29061;
  assign n29063 = n29062 ^ n29016;
  assign n29015 = n29008 ^ n28996;
  assign n29064 = n29063 ^ n29015;
  assign n815 = n802 ^ n774;
  assign n828 = n827 ^ n815;
  assign n832 = n831 ^ n828;
  assign n29065 = n29063 ^ n832;
  assign n29066 = n29064 & n29065;
  assign n29067 = n29066 ^ n832;
  assign n29014 = n29010 ^ n29009;
  assign n29068 = n29067 ^ n29014;
  assign n29069 = n29014 ^ n847;
  assign n29070 = ~n29068 & n29069;
  assign n29071 = n29070 ^ n847;
  assign n29072 = n29071 ^ n29012;
  assign n29073 = ~n29013 & n29072;
  assign n29074 = n29073 ^ n942;
  assign n29428 = n29092 ^ n29074;
  assign n29429 = n29096 & ~n29428;
  assign n29430 = n29429 ^ n29095;
  assign n29431 = n29430 ^ n29426;
  assign n29432 = n29427 & ~n29431;
  assign n29433 = n29432 ^ n1100;
  assign n29434 = n29433 ^ n29421;
  assign n29435 = n29425 & ~n29434;
  assign n29436 = n29435 ^ n29424;
  assign n29437 = n29436 ^ n29419;
  assign n29438 = ~n29420 & n29437;
  assign n29439 = n29438 ^ n29418;
  assign n29440 = n29439 ^ n29414;
  assign n29441 = ~n29415 & n29440;
  assign n29442 = n29441 ^ n2429;
  assign n29443 = n29442 ^ n29412;
  assign n29444 = ~n29413 & n29443;
  assign n29445 = n29444 ^ n3035;
  assign n29446 = n29445 ^ n29407;
  assign n29447 = ~n29411 & n29446;
  assign n29448 = n29447 ^ n29410;
  assign n29449 = n29448 ^ n29405;
  assign n29450 = n29406 & ~n29449;
  assign n29451 = n29450 ^ n29402;
  assign n29452 = n29451 ^ n3211;
  assign n29453 = ~n29401 & ~n29452;
  assign n29454 = n29453 ^ n29400;
  assign n29345 = n29329 & n29344;
  assign n29278 = n29277 ^ n29234;
  assign n29279 = n29235 & ~n29278;
  assign n29280 = n29279 ^ n26664;
  assign n29198 = n29197 ^ n29126;
  assign n29199 = n29193 & ~n29198;
  assign n29200 = n29199 ^ n29197;
  assign n29123 = n28692 ^ n28588;
  assign n29124 = n29123 ^ n28585;
  assign n29119 = n27859 ^ n27330;
  assign n29120 = n28338 ^ n27859;
  assign n29121 = n29119 & n29120;
  assign n29122 = n29121 ^ n27330;
  assign n29125 = n29124 ^ n29122;
  assign n29232 = n29200 ^ n29125;
  assign n29233 = n29232 ^ n26745;
  assign n29328 = n29280 ^ n29233;
  assign n29398 = n29345 ^ n29328;
  assign n29399 = n29398 ^ n2780;
  assign n29735 = n29454 ^ n29399;
  assign n29731 = n28233 ^ n27476;
  assign n29576 = n28722 ^ n28556;
  assign n29577 = n29576 ^ n28553;
  assign n29732 = n29577 ^ n28233;
  assign n29733 = n29731 & n29732;
  assign n29734 = n29733 ^ n27476;
  assign n29736 = n29735 ^ n29734;
  assign n29741 = n29451 ^ n29401;
  assign n29737 = n28226 ^ n27469;
  assign n29531 = n28719 ^ n28561;
  assign n29532 = n29531 ^ n28558;
  assign n29738 = n29532 ^ n28226;
  assign n29739 = ~n29737 & ~n29738;
  assign n29740 = n29739 ^ n27469;
  assign n29742 = n29741 ^ n29740;
  assign n29746 = n28850 ^ n27269;
  assign n29360 = n28713 ^ n28569;
  assign n29747 = n29360 ^ n28850;
  assign n29748 = ~n29746 & ~n29747;
  assign n29749 = n29748 ^ n27269;
  assign n29744 = n29445 ^ n29410;
  assign n29745 = n29744 ^ n29407;
  assign n29750 = n29749 ^ n29745;
  assign n29884 = n29442 ^ n29413;
  assign n29875 = n29439 ^ n29415;
  assign n29756 = n29433 ^ n29425;
  assign n29752 = n28338 ^ n27875;
  assign n29111 = n28701 ^ n28577;
  assign n29753 = n29111 ^ n28338;
  assign n29754 = n29752 & ~n29753;
  assign n29755 = n29754 ^ n27875;
  assign n29757 = n29756 ^ n29755;
  assign n29762 = n29430 ^ n29427;
  assign n29758 = n27985 ^ n27848;
  assign n29207 = n28698 ^ n28579;
  assign n29759 = n29207 ^ n27848;
  assign n29760 = ~n29758 & ~n29759;
  assign n29761 = n29760 ^ n27985;
  assign n29763 = n29762 ^ n29761;
  assign n29768 = n27889 ^ n27864;
  assign n29769 = n29124 ^ n27864;
  assign n29770 = ~n29768 & n29769;
  assign n29771 = n29770 ^ n27889;
  assign n29103 = n29071 ^ n29013;
  assign n29772 = n29771 ^ n29103;
  assign n29773 = n27897 ^ n27872;
  assign n29774 = n29126 ^ n27872;
  assign n29775 = ~n29773 & n29774;
  assign n29776 = n29775 ^ n27897;
  assign n29683 = n29068 ^ n847;
  assign n29777 = n29776 ^ n29683;
  assign n29778 = n28002 ^ n27879;
  assign n29779 = n28813 ^ n27879;
  assign n29780 = ~n29778 & n29779;
  assign n29781 = n29780 ^ n28002;
  assign n29690 = n29064 ^ n832;
  assign n29782 = n29781 ^ n29690;
  assign n29787 = n29060 ^ n29017;
  assign n29783 = n28308 ^ n27837;
  assign n29784 = n29101 ^ n28308;
  assign n29785 = ~n29783 & n29784;
  assign n29786 = n29785 ^ n27837;
  assign n29788 = n29787 ^ n29786;
  assign n29789 = n27886 ^ n27697;
  assign n29790 = n29178 ^ n27886;
  assign n29791 = ~n29789 & n29790;
  assign n29792 = n29791 ^ n27697;
  assign n29698 = n29057 ^ n29021;
  assign n29699 = n29698 ^ n29018;
  assign n29793 = n29792 ^ n29699;
  assign n29795 = n27893 ^ n27681;
  assign n29796 = n29136 ^ n27893;
  assign n29797 = n29795 & n29796;
  assign n29798 = n29797 ^ n27681;
  assign n29794 = n29054 ^ n29027;
  assign n29799 = n29798 ^ n29794;
  assign n29804 = n29051 ^ n29032;
  assign n29800 = n27902 ^ n27273;
  assign n29801 = n29142 ^ n27902;
  assign n29802 = ~n29800 & n29801;
  assign n29803 = n29802 ^ n27273;
  assign n29805 = n29804 ^ n29803;
  assign n29810 = n29048 ^ n29047;
  assign n29806 = n28290 ^ n27274;
  assign n29807 = n29148 ^ n28290;
  assign n29808 = ~n29806 & n29807;
  assign n29809 = n29808 ^ n27274;
  assign n29811 = n29810 ^ n29809;
  assign n29816 = n29043 ^ n29039;
  assign n29817 = n29816 ^ n29036;
  assign n29812 = n27909 ^ n27275;
  assign n29813 = n29154 ^ n27909;
  assign n29814 = n29812 & ~n29813;
  assign n29815 = n29814 ^ n27275;
  assign n29818 = n29817 ^ n29815;
  assign n29613 = n27923 ^ n27289;
  assign n29614 = n28819 ^ n27923;
  assign n29615 = n29613 & ~n29614;
  assign n29616 = n29615 ^ n27289;
  assign n29612 = n28733 ^ n2158;
  assign n29617 = n29616 ^ n29612;
  assign n29545 = n27936 ^ n27301;
  assign n29546 = n28832 ^ n27936;
  assign n29547 = ~n29545 & ~n29546;
  assign n29548 = n29547 ^ n27301;
  assign n29307 = n28707 ^ n28573;
  assign n29302 = n27476 ^ n26826;
  assign n29303 = n28864 ^ n27476;
  assign n29304 = n29302 & ~n29303;
  assign n29305 = n29304 ^ n26826;
  assign n29319 = n29307 ^ n29305;
  assign n29224 = n28704 ^ n28575;
  assign n29219 = n27469 ^ n26671;
  assign n29220 = n28850 ^ n27469;
  assign n29221 = n29219 & n29220;
  assign n29222 = n29221 ^ n26671;
  assign n29298 = n29224 ^ n29222;
  assign n29107 = n28128 ^ n27406;
  assign n29108 = n28789 ^ n28128;
  assign n29109 = ~n29107 & ~n29108;
  assign n29110 = n29109 ^ n27406;
  assign n29112 = n29111 ^ n29110;
  assign n29114 = n27852 ^ n27326;
  assign n29115 = n28484 ^ n27852;
  assign n29116 = ~n29114 & n29115;
  assign n29117 = n29116 ^ n27326;
  assign n29113 = n28695 ^ n28584;
  assign n29118 = n29117 ^ n29113;
  assign n29201 = n29200 ^ n29122;
  assign n29202 = ~n29125 & n29201;
  assign n29203 = n29202 ^ n29124;
  assign n29204 = n29203 ^ n29113;
  assign n29205 = n29118 & ~n29204;
  assign n29206 = n29205 ^ n29117;
  assign n29208 = n29207 ^ n29206;
  assign n29209 = n27359 ^ n27269;
  assign n29210 = n28750 ^ n27269;
  assign n29211 = ~n29209 & ~n29210;
  assign n29212 = n29211 ^ n27359;
  assign n29213 = n29212 ^ n29207;
  assign n29214 = n29208 & n29213;
  assign n29215 = n29214 ^ n29212;
  assign n29216 = n29215 ^ n29110;
  assign n29217 = ~n29112 & ~n29216;
  assign n29218 = n29217 ^ n29111;
  assign n29299 = n29224 ^ n29218;
  assign n29300 = n29298 & ~n29299;
  assign n29301 = n29300 ^ n29222;
  assign n29320 = n29307 ^ n29301;
  assign n29321 = n29319 & ~n29320;
  assign n29322 = n29321 ^ n29305;
  assign n29315 = n27464 ^ n26819;
  assign n29316 = n28226 ^ n27464;
  assign n29317 = n29315 & ~n29316;
  assign n29318 = n29317 ^ n26819;
  assign n29323 = n29322 ^ n29318;
  assign n29314 = n28710 ^ n28571;
  assign n29324 = n29323 ^ n29314;
  assign n29306 = n29305 ^ n29301;
  assign n29308 = n29307 ^ n29306;
  assign n29226 = n29215 ^ n29112;
  assign n29227 = n29226 ^ n26735;
  assign n29228 = n29212 ^ n29208;
  assign n29229 = n29228 ^ n26737;
  assign n29281 = n29280 ^ n29232;
  assign n29282 = n29233 & ~n29281;
  assign n29283 = n29282 ^ n26745;
  assign n29230 = n29203 ^ n29117;
  assign n29231 = n29230 ^ n29113;
  assign n29284 = n29283 ^ n29231;
  assign n29285 = n29231 ^ n26743;
  assign n29286 = n29284 & ~n29285;
  assign n29287 = n29286 ^ n26743;
  assign n29288 = n29287 ^ n29228;
  assign n29289 = ~n29229 & n29288;
  assign n29290 = n29289 ^ n26737;
  assign n29291 = n29290 ^ n29226;
  assign n29292 = n29227 & n29291;
  assign n29293 = n29292 ^ n26735;
  assign n29223 = n29222 ^ n29218;
  assign n29225 = n29224 ^ n29223;
  assign n29294 = n29293 ^ n29225;
  assign n29295 = n29225 ^ n26186;
  assign n29296 = ~n29294 & n29295;
  assign n29297 = n29296 ^ n26186;
  assign n29309 = n29308 ^ n29297;
  assign n29310 = n29308 ^ n26190;
  assign n29311 = ~n29309 & ~n29310;
  assign n29312 = n29311 ^ n26190;
  assign n29313 = n29312 ^ n26195;
  assign n29325 = n29324 ^ n29313;
  assign n29326 = n29294 ^ n26186;
  assign n29327 = n29284 ^ n26743;
  assign n29346 = ~n29328 & ~n29345;
  assign n29347 = n29327 & n29346;
  assign n29348 = n29287 ^ n29229;
  assign n29349 = n29347 & n29348;
  assign n29350 = n29290 ^ n29227;
  assign n29351 = ~n29349 & n29350;
  assign n29352 = ~n29326 & n29351;
  assign n29353 = n29309 ^ n26190;
  assign n29354 = n29352 & n29353;
  assign n29355 = ~n29325 & n29354;
  assign n29368 = n29324 ^ n26195;
  assign n29369 = n29324 ^ n29312;
  assign n29370 = ~n29368 & n29369;
  assign n29371 = n29370 ^ n26195;
  assign n29362 = n27458 ^ n26837;
  assign n29363 = n28233 ^ n27458;
  assign n29364 = ~n29362 & n29363;
  assign n29365 = n29364 ^ n26837;
  assign n29356 = n29318 ^ n29314;
  assign n29357 = n29322 ^ n29314;
  assign n29358 = n29356 & n29357;
  assign n29359 = n29358 ^ n29318;
  assign n29361 = n29360 ^ n29359;
  assign n29366 = n29365 ^ n29361;
  assign n29367 = n29366 ^ n26177;
  assign n29372 = n29371 ^ n29367;
  assign n29495 = ~n29355 & ~n29372;
  assign n29490 = n29371 ^ n29366;
  assign n29491 = n29367 & n29490;
  assign n29492 = n29491 ^ n26177;
  assign n29485 = n27452 ^ n26815;
  assign n29486 = n28220 ^ n27452;
  assign n29487 = ~n29485 & ~n29486;
  assign n29488 = n29487 ^ n26815;
  assign n29481 = n29365 ^ n29360;
  assign n29482 = ~n29361 & ~n29481;
  assign n29483 = n29482 ^ n29365;
  assign n29480 = n28716 ^ n28567;
  assign n29484 = n29483 ^ n29480;
  assign n29489 = n29488 ^ n29484;
  assign n29493 = n29492 ^ n29489;
  assign n29494 = n29493 ^ n26171;
  assign n29496 = n29495 ^ n29494;
  assign n29497 = n29496 ^ n2002;
  assign n29373 = n29372 ^ n29355;
  assign n29377 = n29376 ^ n29373;
  assign n29378 = n29354 ^ n29325;
  assign n29382 = n29381 ^ n29378;
  assign n29383 = n29353 ^ n29352;
  assign n29387 = n29386 ^ n29383;
  assign n29388 = n29351 ^ n29326;
  assign n29392 = n29391 ^ n29388;
  assign n29393 = n29350 ^ n29349;
  assign n29394 = n29393 ^ n1601;
  assign n29395 = n29348 ^ n29347;
  assign n2888 = n2880 ^ n2824;
  assign n2889 = n2888 ^ n2802;
  assign n2890 = n2889 ^ n1502;
  assign n29396 = n29395 ^ n2890;
  assign n29455 = n29454 ^ n29398;
  assign n29456 = n29399 & n29455;
  assign n29457 = n29456 ^ n2780;
  assign n29397 = n29346 ^ n29327;
  assign n29458 = n29457 ^ n29397;
  assign n2790 = n2729 ^ n1527;
  assign n2791 = n2790 ^ n2787;
  assign n2795 = n2794 ^ n2791;
  assign n29459 = n29397 ^ n2795;
  assign n29460 = ~n29458 & n29459;
  assign n29461 = n29460 ^ n2795;
  assign n29462 = n29461 ^ n29395;
  assign n29463 = n29396 & ~n29462;
  assign n29464 = n29463 ^ n2890;
  assign n29465 = n29464 ^ n29393;
  assign n29466 = n29394 & ~n29465;
  assign n29467 = n29466 ^ n1601;
  assign n29468 = n29467 ^ n29388;
  assign n29469 = n29392 & ~n29468;
  assign n29470 = n29469 ^ n29391;
  assign n29471 = n29470 ^ n29383;
  assign n29472 = ~n29387 & n29471;
  assign n29473 = n29472 ^ n29386;
  assign n29474 = n29473 ^ n29378;
  assign n29475 = n29382 & ~n29474;
  assign n29476 = n29475 ^ n29381;
  assign n29477 = n29476 ^ n29373;
  assign n29478 = n29377 & ~n29477;
  assign n29479 = n29478 ^ n29376;
  assign n29540 = n29496 ^ n29479;
  assign n29541 = n29497 & ~n29540;
  assign n29542 = n29541 ^ n2002;
  assign n29535 = n29489 ^ n26171;
  assign n29536 = ~n29493 & n29535;
  assign n29537 = n29536 ^ n26171;
  assign n29527 = n29488 ^ n29480;
  assign n29528 = n29484 & n29527;
  assign n29529 = n29528 ^ n29488;
  assign n29523 = n27323 ^ n26729;
  assign n29524 = n28213 ^ n27323;
  assign n29525 = n29523 & ~n29524;
  assign n29526 = n29525 ^ n26729;
  assign n29530 = n29529 ^ n29526;
  assign n29533 = n29532 ^ n29530;
  assign n29534 = n29533 ^ n25936;
  assign n29538 = n29537 ^ n29534;
  assign n29522 = n29494 & n29495;
  assign n29539 = n29538 ^ n29522;
  assign n29543 = n29542 ^ n29539;
  assign n29544 = n29543 ^ n2012;
  assign n29549 = n29548 ^ n29544;
  assign n29499 = n27946 ^ n27308;
  assign n29500 = n28921 ^ n27946;
  assign n29501 = n29499 & ~n29500;
  assign n29502 = n29501 ^ n27308;
  assign n29498 = n29497 ^ n29479;
  assign n29503 = n29502 ^ n29498;
  assign n29505 = n27948 ^ n27309;
  assign n29506 = n28838 ^ n27948;
  assign n29507 = n29505 & ~n29506;
  assign n29508 = n29507 ^ n27309;
  assign n29504 = n29476 ^ n29377;
  assign n29509 = n29508 ^ n29504;
  assign n29510 = n29473 ^ n29382;
  assign n29511 = n27949 ^ n27315;
  assign n29512 = n28844 ^ n27949;
  assign n29513 = n29511 & n29512;
  assign n29514 = n29513 ^ n27315;
  assign n29515 = n29510 & n29514;
  assign n29516 = n29515 ^ n29504;
  assign n29517 = ~n29509 & n29516;
  assign n29518 = n29517 ^ n29515;
  assign n29519 = n29518 ^ n29502;
  assign n29520 = n29503 & ~n29519;
  assign n29521 = n29520 ^ n29498;
  assign n29596 = n29544 ^ n29521;
  assign n29597 = n29549 & n29596;
  assign n29598 = n29597 ^ n29548;
  assign n29591 = n29539 ^ n2012;
  assign n29592 = n29543 & ~n29591;
  assign n29593 = n29592 ^ n2012;
  assign n2138 = n2124 ^ n2053;
  assign n2139 = n2138 ^ n2022;
  assign n2143 = n2142 ^ n2139;
  assign n29594 = n29593 ^ n2143;
  assign n29589 = n29522 & ~n29538;
  assign n29584 = n29537 ^ n29533;
  assign n29585 = ~n29534 & n29584;
  assign n29586 = n29585 ^ n25936;
  assign n29587 = n29586 ^ n25932;
  assign n29579 = n27317 ^ n26725;
  assign n29580 = n28207 ^ n27317;
  assign n29581 = ~n29579 & n29580;
  assign n29582 = n29581 ^ n26725;
  assign n29572 = n29532 ^ n29526;
  assign n29573 = n29532 ^ n29529;
  assign n29574 = n29572 & ~n29573;
  assign n29575 = n29574 ^ n29526;
  assign n29578 = n29577 ^ n29575;
  assign n29583 = n29582 ^ n29578;
  assign n29588 = n29587 ^ n29583;
  assign n29590 = n29589 ^ n29588;
  assign n29595 = n29594 ^ n29590;
  assign n29599 = n29598 ^ n29595;
  assign n29568 = n27930 ^ n27295;
  assign n29569 = n28821 ^ n27930;
  assign n29570 = n29568 & ~n29569;
  assign n29571 = n29570 ^ n27295;
  assign n29609 = n29595 ^ n29571;
  assign n29610 = n29599 & ~n29609;
  assign n29611 = n29610 ^ n29571;
  assign n29633 = n29616 ^ n29611;
  assign n29634 = n29617 & n29633;
  assign n29635 = n29634 ^ n29612;
  assign n29632 = n28767 ^ n28735;
  assign n29636 = n29635 ^ n29632;
  assign n29628 = n27917 ^ n27282;
  assign n29629 = n28986 ^ n27917;
  assign n29630 = ~n29628 & n29629;
  assign n29631 = n29630 ^ n27282;
  assign n29819 = n29632 ^ n29631;
  assign n29820 = ~n29636 & ~n29819;
  assign n29821 = n29820 ^ n29631;
  assign n29822 = n29821 ^ n28811;
  assign n29823 = n27915 ^ n27276;
  assign n29824 = n29087 ^ n27915;
  assign n29825 = n29823 & n29824;
  assign n29826 = n29825 ^ n27276;
  assign n29827 = n29826 ^ n28811;
  assign n29828 = ~n29822 & ~n29827;
  assign n29829 = n29828 ^ n29826;
  assign n29830 = n29829 ^ n29817;
  assign n29831 = n29818 & n29830;
  assign n29832 = n29831 ^ n29815;
  assign n29833 = n29832 ^ n29809;
  assign n29834 = n29811 & n29833;
  assign n29835 = n29834 ^ n29810;
  assign n29836 = n29835 ^ n29803;
  assign n29837 = n29805 & n29836;
  assign n29838 = n29837 ^ n29804;
  assign n29839 = n29838 ^ n29794;
  assign n29840 = ~n29799 & n29839;
  assign n29841 = n29840 ^ n29798;
  assign n29842 = n29841 ^ n29792;
  assign n29843 = ~n29793 & n29842;
  assign n29844 = n29843 ^ n29699;
  assign n29845 = n29844 ^ n29787;
  assign n29846 = n29788 & n29845;
  assign n29847 = n29846 ^ n29786;
  assign n29848 = n29847 ^ n29690;
  assign n29849 = ~n29782 & n29848;
  assign n29850 = n29849 ^ n29781;
  assign n29851 = n29850 ^ n29776;
  assign n29852 = ~n29777 & n29851;
  assign n29853 = n29852 ^ n29683;
  assign n29854 = n29853 ^ n29103;
  assign n29855 = ~n29772 & n29854;
  assign n29856 = n29855 ^ n29771;
  assign n29764 = n27882 ^ n27856;
  assign n29765 = n29113 ^ n27856;
  assign n29766 = ~n29764 & ~n29765;
  assign n29767 = n29766 ^ n27882;
  assign n29857 = n29856 ^ n29767;
  assign n29097 = n29096 ^ n29074;
  assign n29858 = n29856 ^ n29097;
  assign n29859 = ~n29857 & ~n29858;
  assign n29860 = n29859 ^ n29767;
  assign n29861 = n29860 ^ n29761;
  assign n29862 = n29763 & n29861;
  assign n29863 = n29862 ^ n29762;
  assign n29864 = n29863 ^ n29756;
  assign n29865 = n29757 & ~n29864;
  assign n29866 = n29865 ^ n29755;
  assign n29751 = n29436 ^ n29420;
  assign n29867 = n29866 ^ n29751;
  assign n29868 = n28484 ^ n27867;
  assign n29869 = n29224 ^ n28484;
  assign n29870 = ~n29868 & ~n29869;
  assign n29871 = n29870 ^ n27867;
  assign n29872 = n29871 ^ n29751;
  assign n29873 = n29867 & n29872;
  assign n29874 = n29873 ^ n29871;
  assign n29876 = n29875 ^ n29874;
  assign n29877 = n28750 ^ n27859;
  assign n29878 = n29307 ^ n28750;
  assign n29879 = ~n29877 & ~n29878;
  assign n29880 = n29879 ^ n27859;
  assign n29881 = n29880 ^ n29874;
  assign n29882 = n29876 & ~n29881;
  assign n29883 = n29882 ^ n29875;
  assign n29885 = n29884 ^ n29883;
  assign n29886 = n28789 ^ n27852;
  assign n29887 = n29314 ^ n28789;
  assign n29888 = ~n29886 & n29887;
  assign n29889 = n29888 ^ n27852;
  assign n29890 = n29889 ^ n29883;
  assign n29891 = n29885 & ~n29890;
  assign n29892 = n29891 ^ n29884;
  assign n29893 = n29892 ^ n29745;
  assign n29894 = ~n29750 & ~n29893;
  assign n29895 = n29894 ^ n29749;
  assign n29743 = n29448 ^ n29406;
  assign n29896 = n29895 ^ n29743;
  assign n29897 = n28864 ^ n28128;
  assign n29898 = n29480 ^ n28864;
  assign n29899 = n29897 & n29898;
  assign n29900 = n29899 ^ n28128;
  assign n29901 = n29900 ^ n29743;
  assign n29902 = ~n29896 & n29901;
  assign n29903 = n29902 ^ n29900;
  assign n29904 = n29903 ^ n29741;
  assign n29905 = ~n29742 & n29904;
  assign n29906 = n29905 ^ n29740;
  assign n29907 = n29906 ^ n29735;
  assign n29908 = ~n29736 & n29907;
  assign n29909 = n29908 ^ n29734;
  assign n29725 = n28220 ^ n27464;
  assign n29726 = n28727 ^ n28220;
  assign n29727 = ~n29725 & n29726;
  assign n29728 = n29727 ^ n27464;
  assign n29938 = n29909 ^ n29728;
  assign n29729 = n29458 ^ n2795;
  assign n29939 = n29938 ^ n29729;
  assign n29940 = n29939 ^ n26819;
  assign n29941 = n29906 ^ n29736;
  assign n29942 = n29941 ^ n26826;
  assign n29943 = n29903 ^ n29740;
  assign n29944 = n29943 ^ n29741;
  assign n29945 = n29944 ^ n26671;
  assign n29946 = n29900 ^ n29896;
  assign n29947 = n29946 ^ n27406;
  assign n29950 = n29889 ^ n29884;
  assign n29951 = n29950 ^ n29883;
  assign n29952 = n29951 ^ n27326;
  assign n29953 = n29880 ^ n29875;
  assign n29954 = n29953 ^ n29874;
  assign n29955 = n29954 ^ n27330;
  assign n29956 = n29871 ^ n29867;
  assign n29957 = n29956 ^ n27332;
  assign n29958 = n29863 ^ n29757;
  assign n29959 = n29958 ^ n27339;
  assign n29960 = n29860 ^ n29763;
  assign n29961 = n29960 ^ n27262;
  assign n29964 = n29853 ^ n29771;
  assign n29965 = n29964 ^ n29103;
  assign n29966 = n29965 ^ n27034;
  assign n29968 = n29847 ^ n29781;
  assign n29969 = n29968 ^ n29690;
  assign n29970 = n29969 ^ n26679;
  assign n29971 = n29844 ^ n29788;
  assign n29972 = n29971 ^ n26903;
  assign n29974 = n29838 ^ n29799;
  assign n29975 = n29974 ^ n26685;
  assign n29977 = n29829 ^ n29818;
  assign n29978 = n29977 ^ n26695;
  assign n29979 = n29826 ^ n29822;
  assign n29980 = n29979 ^ n26698;
  assign n29637 = n29636 ^ n29631;
  assign n29638 = n29637 ^ n26700;
  assign n29600 = n29599 ^ n29571;
  assign n29601 = n29600 ^ n26862;
  assign n29550 = n29549 ^ n29521;
  assign n29551 = n29550 ^ n26706;
  assign n29552 = n29518 ^ n29503;
  assign n29553 = n29552 ^ n26712;
  assign n29554 = n29514 ^ n29510;
  assign n29555 = ~n26721 & n29554;
  assign n29556 = n29555 ^ n26717;
  assign n29557 = n29515 ^ n29508;
  assign n29558 = n29557 ^ n29504;
  assign n29559 = n29558 ^ n29555;
  assign n29560 = n29556 & ~n29559;
  assign n29561 = n29560 ^ n26717;
  assign n29562 = n29561 ^ n29552;
  assign n29563 = n29553 & ~n29562;
  assign n29564 = n29563 ^ n26712;
  assign n29565 = n29564 ^ n29550;
  assign n29566 = n29551 & ~n29565;
  assign n29567 = n29566 ^ n26706;
  assign n29619 = n29600 ^ n29567;
  assign n29620 = ~n29601 & ~n29619;
  assign n29621 = n29620 ^ n26862;
  assign n29622 = n29621 ^ n26703;
  assign n29618 = n29617 ^ n29611;
  assign n29625 = n29621 ^ n29618;
  assign n29626 = n29622 & ~n29625;
  assign n29627 = n29626 ^ n26703;
  assign n29981 = n29637 ^ n29627;
  assign n29982 = ~n29638 & ~n29981;
  assign n29983 = n29982 ^ n26700;
  assign n29984 = n29983 ^ n29979;
  assign n29985 = n29980 & ~n29984;
  assign n29986 = n29985 ^ n26698;
  assign n29987 = n29986 ^ n29977;
  assign n29988 = ~n29978 & ~n29987;
  assign n29989 = n29988 ^ n26695;
  assign n29990 = n29989 ^ n26691;
  assign n29991 = n29832 ^ n29811;
  assign n29992 = n29991 ^ n29989;
  assign n29993 = ~n29990 & ~n29992;
  assign n29994 = n29993 ^ n26691;
  assign n29976 = n29835 ^ n29805;
  assign n29995 = n29994 ^ n29976;
  assign n29996 = n29976 ^ n26890;
  assign n29997 = ~n29995 & ~n29996;
  assign n29998 = n29997 ^ n26890;
  assign n29999 = n29998 ^ n29974;
  assign n30000 = ~n29975 & n29999;
  assign n30001 = n30000 ^ n26685;
  assign n29973 = n29841 ^ n29793;
  assign n30002 = n30001 ^ n29973;
  assign n30003 = n29973 ^ n26681;
  assign n30004 = n30002 & ~n30003;
  assign n30005 = n30004 ^ n26681;
  assign n30006 = n30005 ^ n29971;
  assign n30007 = n29972 & ~n30006;
  assign n30008 = n30007 ^ n26903;
  assign n30009 = n30008 ^ n29969;
  assign n30010 = ~n29970 & ~n30009;
  assign n30011 = n30010 ^ n26679;
  assign n29967 = n29850 ^ n29777;
  assign n30012 = n30011 ^ n29967;
  assign n30013 = n29967 ^ n26676;
  assign n30014 = n30012 & ~n30013;
  assign n30015 = n30014 ^ n26676;
  assign n30016 = n30015 ^ n29965;
  assign n30017 = ~n29966 & n30016;
  assign n30018 = n30017 ^ n27034;
  assign n29962 = n29767 ^ n29097;
  assign n29963 = n29962 ^ n29856;
  assign n30019 = n30018 ^ n29963;
  assign n30020 = n30018 ^ n27096;
  assign n30021 = n30019 & n30020;
  assign n30022 = n30021 ^ n27096;
  assign n30023 = n30022 ^ n29960;
  assign n30024 = ~n29961 & n30023;
  assign n30025 = n30024 ^ n27262;
  assign n30026 = n30025 ^ n29958;
  assign n30027 = ~n29959 & ~n30026;
  assign n30028 = n30027 ^ n27339;
  assign n30029 = n30028 ^ n29956;
  assign n30030 = n29957 & n30029;
  assign n30031 = n30030 ^ n27332;
  assign n30032 = n30031 ^ n29954;
  assign n30033 = n29955 & n30032;
  assign n30034 = n30033 ^ n27330;
  assign n30035 = n30034 ^ n29951;
  assign n30036 = ~n29952 & ~n30035;
  assign n30037 = n30036 ^ n27326;
  assign n29948 = n29892 ^ n29749;
  assign n29949 = n29948 ^ n29745;
  assign n30038 = n30037 ^ n29949;
  assign n30039 = n29949 ^ n27359;
  assign n30040 = ~n30038 & ~n30039;
  assign n30041 = n30040 ^ n27359;
  assign n30042 = n30041 ^ n29946;
  assign n30043 = ~n29947 & n30042;
  assign n30044 = n30043 ^ n27406;
  assign n30045 = n30044 ^ n29944;
  assign n30046 = ~n29945 & ~n30045;
  assign n30047 = n30046 ^ n26671;
  assign n30048 = n30047 ^ n29941;
  assign n30049 = ~n29942 & n30048;
  assign n30050 = n30049 ^ n26826;
  assign n30051 = n30050 ^ n29939;
  assign n30052 = n29940 & n30051;
  assign n30053 = n30052 ^ n26819;
  assign n29730 = n29729 ^ n29728;
  assign n29910 = n29909 ^ n29729;
  assign n29911 = ~n29730 & ~n29910;
  assign n29912 = n29911 ^ n29728;
  assign n29720 = n28213 ^ n27458;
  assign n29721 = n28757 ^ n28213;
  assign n29722 = n29720 & n29721;
  assign n29723 = n29722 ^ n27458;
  assign n29935 = n29912 ^ n29723;
  assign n29718 = n29461 ^ n2890;
  assign n29719 = n29718 ^ n29395;
  assign n29936 = n29935 ^ n29719;
  assign n29937 = n29936 ^ n26837;
  assign n30116 = n30053 ^ n29937;
  assign n30066 = n30047 ^ n29942;
  assign n30067 = n30044 ^ n29945;
  assign n30068 = n30041 ^ n27406;
  assign n30069 = n30068 ^ n29946;
  assign n30070 = n30038 ^ n27359;
  assign n30071 = n30031 ^ n29955;
  assign n30072 = n30028 ^ n29957;
  assign n30073 = n30015 ^ n29966;
  assign n30074 = n30012 ^ n26676;
  assign n30075 = n29991 ^ n26691;
  assign n30076 = n30075 ^ n29989;
  assign n30077 = n29986 ^ n26695;
  assign n30078 = n30077 ^ n29977;
  assign n29602 = n29601 ^ n29567;
  assign n29603 = n29561 ^ n26712;
  assign n29604 = n29603 ^ n29552;
  assign n29605 = n29564 ^ n26706;
  assign n29606 = n29605 ^ n29550;
  assign n29607 = ~n29604 & ~n29606;
  assign n29608 = n29602 & n29607;
  assign n29623 = n29622 ^ n29618;
  assign n29624 = ~n29608 & ~n29623;
  assign n29639 = n29638 ^ n29627;
  assign n30079 = ~n29624 & ~n29639;
  assign n30080 = n29983 ^ n29980;
  assign n30081 = n30079 & ~n30080;
  assign n30082 = ~n30078 & ~n30081;
  assign n30083 = n30076 & n30082;
  assign n30084 = n29995 ^ n26890;
  assign n30085 = ~n30083 & n30084;
  assign n30086 = n29998 ^ n29975;
  assign n30087 = n30085 & ~n30086;
  assign n30088 = n30002 ^ n26681;
  assign n30089 = n30087 & ~n30088;
  assign n30090 = n30005 ^ n29972;
  assign n30091 = n30089 & n30090;
  assign n30092 = n30008 ^ n29970;
  assign n30093 = ~n30091 & n30092;
  assign n30094 = n30074 & ~n30093;
  assign n30095 = n30073 & n30094;
  assign n30096 = n29963 ^ n27096;
  assign n30097 = n30096 ^ n30018;
  assign n30098 = n30095 & n30097;
  assign n30099 = n30022 ^ n29961;
  assign n30100 = ~n30098 & ~n30099;
  assign n30101 = n30025 ^ n27339;
  assign n30102 = n30101 ^ n29958;
  assign n30103 = ~n30100 & n30102;
  assign n30104 = n30072 & n30103;
  assign n30105 = n30071 & ~n30104;
  assign n30106 = n30034 ^ n27326;
  assign n30107 = n30106 ^ n29951;
  assign n30108 = n30105 & n30107;
  assign n30109 = ~n30070 & n30108;
  assign n30110 = ~n30069 & ~n30109;
  assign n30111 = ~n30067 & n30110;
  assign n30112 = n30066 & n30111;
  assign n30113 = n30050 ^ n26819;
  assign n30114 = n30113 ^ n29939;
  assign n30115 = n30112 & ~n30114;
  assign n30132 = n30116 ^ n30115;
  assign n1752 = n1751 ^ n1731;
  assign n1762 = n1761 ^ n1752;
  assign n1766 = n1765 ^ n1762;
  assign n30133 = n30132 ^ n1766;
  assign n30137 = n30114 ^ n30112;
  assign n30134 = n28161 ^ n21119;
  assign n30135 = n30134 ^ n1696;
  assign n30136 = n30135 ^ n1756;
  assign n30138 = n30137 ^ n30136;
  assign n30140 = n30110 ^ n30067;
  assign n30141 = n30140 ^ n3009;
  assign n30142 = n30109 ^ n30069;
  assign n2989 = n2921 ^ n1508;
  assign n2990 = n2989 ^ n2975;
  assign n2994 = n2993 ^ n2990;
  assign n30143 = n30142 ^ n2994;
  assign n30144 = n30108 ^ n30070;
  assign n30145 = n30144 ^ n2984;
  assign n30146 = n30107 ^ n30105;
  assign n30150 = n30149 ^ n30146;
  assign n30151 = n30104 ^ n30071;
  assign n30152 = n30151 ^ n3089;
  assign n30153 = n30103 ^ n30072;
  assign n2580 = n2579 ^ n2546;
  assign n2587 = n2586 ^ n2580;
  assign n2588 = n2587 ^ n1559;
  assign n30154 = n30153 ^ n2588;
  assign n30156 = n30099 ^ n30098;
  assign n2506 = n2502 ^ n2484;
  assign n2519 = n2518 ^ n2506;
  assign n2523 = n2522 ^ n2519;
  assign n30157 = n30156 ^ n2523;
  assign n30160 = n30093 ^ n30074;
  assign n1390 = n1383 ^ n1293;
  assign n1397 = n1396 ^ n1390;
  assign n1401 = n1400 ^ n1397;
  assign n30161 = n30160 ^ n1401;
  assign n30163 = n30090 ^ n30089;
  assign n1196 = n1183 ^ n1107;
  assign n1197 = n1196 ^ n1077;
  assign n1201 = n1200 ^ n1197;
  assign n30164 = n30163 ^ n1201;
  assign n30165 = n30088 ^ n30087;
  assign n1062 = n1025 ^ n983;
  assign n1063 = n1062 ^ n1059;
  assign n1067 = n1066 ^ n1063;
  assign n30166 = n30165 ^ n1067;
  assign n30167 = n30086 ^ n30085;
  assign n30168 = n30167 ^ n1052;
  assign n30169 = n30084 ^ n30083;
  assign n30170 = n30169 ^ n3321;
  assign n30172 = n30081 ^ n30078;
  assign n30176 = n30175 ^ n30172;
  assign n30178 = n27747 ^ n20839;
  assign n30179 = n30178 ^ n24741;
  assign n30180 = n30179 ^ n587;
  assign n30177 = n30080 ^ n30079;
  assign n30181 = n30180 ^ n30177;
  assign n29644 = n29623 ^ n29608;
  assign n29641 = n27753 ^ n20845;
  assign n29642 = n29641 ^ n24748;
  assign n29643 = n29642 ^ n558;
  assign n29645 = n29644 ^ n29643;
  assign n29668 = n27759 ^ n536;
  assign n29669 = n29668 ^ n24243;
  assign n29670 = n29669 ^ n3281;
  assign n29646 = n29606 ^ n29604;
  assign n29650 = n29649 ^ n29646;
  assign n29658 = n20856 ^ n2351;
  assign n29659 = n29658 ^ n24193;
  assign n29660 = n29659 ^ n19668;
  assign n2275 = n2236 ^ n2170;
  assign n2276 = n2275 ^ n2272;
  assign n2280 = n2279 ^ n2276;
  assign n29651 = n29554 ^ n26721;
  assign n29652 = n2280 & ~n29651;
  assign n2293 = n2251 ^ n2202;
  assign n2294 = n2293 ^ n2287;
  assign n2298 = n2297 ^ n2294;
  assign n29653 = n29652 ^ n2298;
  assign n29654 = n29558 ^ n29556;
  assign n29655 = n29654 ^ n2298;
  assign n29656 = n29653 & ~n29655;
  assign n29657 = n29656 ^ n29652;
  assign n29661 = n29660 ^ n29657;
  assign n29662 = n29657 ^ n29604;
  assign n29663 = n29661 & n29662;
  assign n29664 = n29663 ^ n29660;
  assign n29665 = n29664 ^ n29646;
  assign n29666 = ~n29650 & n29665;
  assign n29667 = n29666 ^ n29649;
  assign n29671 = n29670 ^ n29667;
  assign n29672 = n29607 ^ n29602;
  assign n29673 = n29672 ^ n29667;
  assign n29674 = n29671 & n29673;
  assign n29675 = n29674 ^ n29670;
  assign n29676 = n29675 ^ n29643;
  assign n29677 = n29645 & ~n29676;
  assign n29678 = n29677 ^ n29644;
  assign n29640 = n29639 ^ n29624;
  assign n29679 = n29678 ^ n29640;
  assign n712 = n711 ^ n708;
  assign n713 = n712 ^ n563;
  assign n714 = n713 ^ n644;
  assign n30182 = n29640 ^ n714;
  assign n30183 = n29679 & ~n30182;
  assign n30184 = n30183 ^ n714;
  assign n30185 = n30184 ^ n30177;
  assign n30186 = n30181 & ~n30185;
  assign n30187 = n30186 ^ n30180;
  assign n30188 = n30187 ^ n30172;
  assign n30189 = n30176 & ~n30188;
  assign n30190 = n30189 ^ n30175;
  assign n30171 = n30082 ^ n30076;
  assign n30191 = n30190 ^ n30171;
  assign n30195 = n30194 ^ n30171;
  assign n30196 = ~n30191 & n30195;
  assign n30197 = n30196 ^ n30194;
  assign n30198 = n30197 ^ n30169;
  assign n30199 = n30170 & ~n30198;
  assign n30200 = n30199 ^ n3321;
  assign n30201 = n30200 ^ n30167;
  assign n30202 = n30168 & ~n30201;
  assign n30203 = n30202 ^ n1052;
  assign n30204 = n30203 ^ n30165;
  assign n30205 = n30166 & ~n30204;
  assign n30206 = n30205 ^ n1067;
  assign n30207 = n30206 ^ n30163;
  assign n30208 = ~n30164 & n30207;
  assign n30209 = n30208 ^ n1201;
  assign n30162 = n30092 ^ n30091;
  assign n30210 = n30209 ^ n30162;
  assign n1211 = n1192 ^ n1123;
  assign n1212 = n1211 ^ n1208;
  assign n1216 = n1215 ^ n1212;
  assign n30211 = n30209 ^ n1216;
  assign n30212 = n30210 & n30211;
  assign n30213 = n30212 ^ n1216;
  assign n30214 = n30213 ^ n30160;
  assign n30215 = n30161 & ~n30214;
  assign n30216 = n30215 ^ n1401;
  assign n30159 = n30094 ^ n30073;
  assign n30217 = n30216 ^ n30159;
  assign n30218 = n27724 ^ n2443;
  assign n30219 = n30218 ^ n1408;
  assign n30220 = n30219 ^ n3151;
  assign n30221 = n30220 ^ n30159;
  assign n30222 = n30217 & ~n30221;
  assign n30223 = n30222 ^ n30220;
  assign n30158 = n30097 ^ n30095;
  assign n30224 = n30223 ^ n30158;
  assign n3147 = n3146 ^ n2452;
  assign n3154 = n3153 ^ n3147;
  assign n3155 = n3154 ^ n2513;
  assign n30225 = n30158 ^ n3155;
  assign n30226 = n30224 & ~n30225;
  assign n30227 = n30226 ^ n3155;
  assign n30228 = n30227 ^ n30156;
  assign n30229 = n30157 & ~n30228;
  assign n30230 = n30229 ^ n2523;
  assign n30155 = n30102 ^ n30100;
  assign n30231 = n30230 ^ n30155;
  assign n3067 = n3062 ^ n3053;
  assign n3068 = n3067 ^ n2530;
  assign n3069 = n3068 ^ n2584;
  assign n30232 = n30155 ^ n3069;
  assign n30233 = ~n30231 & n30232;
  assign n30234 = n30233 ^ n3069;
  assign n30235 = n30234 ^ n30153;
  assign n30236 = ~n30154 & n30235;
  assign n30237 = n30236 ^ n2588;
  assign n30238 = n30237 ^ n3089;
  assign n30239 = ~n30152 & ~n30238;
  assign n30240 = n30239 ^ n30151;
  assign n30241 = n30240 ^ n30146;
  assign n30242 = n30150 & n30241;
  assign n30243 = n30242 ^ n30149;
  assign n30244 = n30243 ^ n30144;
  assign n30245 = ~n30145 & n30244;
  assign n30246 = n30245 ^ n2984;
  assign n30247 = n30246 ^ n30142;
  assign n30248 = ~n30143 & n30247;
  assign n30249 = n30248 ^ n2994;
  assign n30250 = n30249 ^ n30140;
  assign n30251 = n30141 & ~n30250;
  assign n30252 = n30251 ^ n3009;
  assign n30139 = n30111 ^ n30066;
  assign n30253 = n30252 ^ n30139;
  assign n1672 = n1665 ^ n1647;
  assign n1685 = n1684 ^ n1672;
  assign n1689 = n1688 ^ n1685;
  assign n30254 = n30139 ^ n1689;
  assign n30255 = n30253 & ~n30254;
  assign n30256 = n30255 ^ n1689;
  assign n30257 = n30256 ^ n30137;
  assign n30258 = n30138 & ~n30257;
  assign n30259 = n30258 ^ n30136;
  assign n30260 = n30259 ^ n30132;
  assign n30261 = n30133 & ~n30260;
  assign n30262 = n30261 ^ n1766;
  assign n30117 = ~n30115 & ~n30116;
  assign n30054 = n30053 ^ n29936;
  assign n30055 = n29937 & n30054;
  assign n30056 = n30055 ^ n26837;
  assign n30064 = n30056 ^ n26815;
  assign n29724 = n29723 ^ n29719;
  assign n29913 = n29912 ^ n29719;
  assign n29914 = ~n29724 & n29913;
  assign n29915 = n29914 ^ n29723;
  assign n29713 = n28207 ^ n27452;
  assign n29714 = n28799 ^ n28207;
  assign n29715 = ~n29713 & ~n29714;
  assign n29716 = n29715 ^ n27452;
  assign n29932 = n29915 ^ n29716;
  assign n29711 = n29464 ^ n1601;
  assign n29712 = n29711 ^ n29393;
  assign n29933 = n29932 ^ n29712;
  assign n30065 = n30064 ^ n29933;
  assign n30127 = n30117 ^ n30065;
  assign n30131 = n30130 ^ n30127;
  assign n30296 = n30262 ^ n30131;
  assign n30284 = n28921 ^ n27949;
  assign n30285 = n29612 ^ n28921;
  assign n30286 = n30284 & ~n30285;
  assign n30287 = n30286 ^ n27949;
  assign n30288 = n30256 ^ n30138;
  assign n30289 = n30287 & n30288;
  assign n30280 = n28832 ^ n27948;
  assign n30281 = n29632 ^ n28832;
  assign n30282 = n30280 & ~n30281;
  assign n30283 = n30282 ^ n27948;
  assign n30290 = n30289 ^ n30283;
  assign n30291 = n30259 ^ n30133;
  assign n30292 = n30291 ^ n30289;
  assign n30293 = n30290 & ~n30292;
  assign n30294 = n30293 ^ n30283;
  assign n30276 = n28821 ^ n27946;
  assign n30277 = n28821 ^ n28811;
  assign n30278 = ~n30276 & ~n30277;
  assign n30279 = n30278 ^ n27946;
  assign n30295 = n30294 ^ n30279;
  assign n30376 = n30296 ^ n30295;
  assign n30368 = n30288 ^ n30287;
  assign n30369 = n27315 & n30368;
  assign n30370 = n30369 ^ n27309;
  assign n30371 = n30291 ^ n30290;
  assign n30372 = n30371 ^ n30369;
  assign n30373 = n30370 & ~n30372;
  assign n30374 = n30373 ^ n27309;
  assign n30375 = n30374 ^ n27308;
  assign n30441 = n30376 ^ n30375;
  assign n30684 = n30526 ^ n30441;
  assign n2133 = n2132 ^ n2045;
  assign n2134 = n2133 ^ n2126;
  assign n2135 = n2134 ^ n2117;
  assign n30514 = n30368 ^ n27315;
  assign n30515 = n2135 & n30514;
  assign n30519 = n30518 ^ n30515;
  assign n30520 = n30371 ^ n30370;
  assign n30521 = n30520 ^ n30518;
  assign n30522 = n30519 & ~n30521;
  assign n30523 = n30522 ^ n30515;
  assign n30685 = n30684 ^ n30523;
  assign n29703 = n29661 ^ n29604;
  assign n32434 = n30685 ^ n29703;
  assign n30728 = n29480 ^ n28789;
  assign n30729 = n29729 ^ n29480;
  assign n30730 = ~n30728 & n30729;
  assign n30731 = n30730 ^ n28789;
  assign n30603 = n30223 ^ n3155;
  assign n30604 = n30603 ^ n30158;
  assign n30732 = n30731 ^ n30604;
  assign n30733 = n29360 ^ n28750;
  assign n30734 = n29735 ^ n29360;
  assign n30735 = ~n30733 & ~n30734;
  assign n30736 = n30735 ^ n28750;
  assign n30616 = n30220 ^ n30217;
  assign n30737 = n30736 ^ n30616;
  assign n30738 = n29314 ^ n28484;
  assign n30739 = n29741 ^ n29314;
  assign n30740 = ~n30738 & ~n30739;
  assign n30741 = n30740 ^ n28484;
  assign n30623 = n30213 ^ n30161;
  assign n30742 = n30741 ^ n30623;
  assign n30743 = n29111 ^ n27856;
  assign n30744 = n29884 ^ n29111;
  assign n30745 = n30743 & n30744;
  assign n30746 = n30745 ^ n27856;
  assign n30647 = n30203 ^ n30166;
  assign n30747 = n30746 ^ n30647;
  assign n30748 = n29207 ^ n27864;
  assign n30749 = n29875 ^ n29207;
  assign n30750 = n30748 & ~n30749;
  assign n30751 = n30750 ^ n27864;
  assign n30655 = n30200 ^ n1052;
  assign n30656 = n30655 ^ n30167;
  assign n30752 = n30751 ^ n30656;
  assign n30426 = n30187 ^ n30175;
  assign n30427 = n30426 ^ n30172;
  assign n30422 = n29126 ^ n28308;
  assign n30423 = n29762 ^ n29126;
  assign n30424 = n30422 & n30423;
  assign n30425 = n30424 ^ n28308;
  assign n30428 = n30427 ^ n30425;
  assign n30351 = n30184 ^ n30181;
  assign n29680 = n29679 ^ n714;
  assign n29102 = n29101 ^ n27893;
  assign n29104 = n29103 ^ n29101;
  assign n29105 = ~n29102 & n29104;
  assign n29106 = n29105 ^ n27893;
  assign n29681 = n29680 ^ n29106;
  assign n29687 = n29675 ^ n29645;
  assign n29682 = n29178 ^ n27902;
  assign n29684 = n29683 ^ n29178;
  assign n29685 = n29682 & ~n29684;
  assign n29686 = n29685 ^ n27902;
  assign n29688 = n29687 ^ n29686;
  assign n29694 = n29672 ^ n29670;
  assign n29695 = n29694 ^ n29667;
  assign n29689 = n29136 ^ n28290;
  assign n29691 = n29690 ^ n29136;
  assign n29692 = ~n29689 & n29691;
  assign n29693 = n29692 ^ n28290;
  assign n29696 = n29695 ^ n29693;
  assign n30333 = n29142 ^ n27909;
  assign n30334 = n29787 ^ n29142;
  assign n30335 = n30333 & n30334;
  assign n30336 = n30335 ^ n27909;
  assign n29697 = n29148 ^ n27915;
  assign n29700 = n29699 ^ n29148;
  assign n29701 = n29697 & n29700;
  assign n29702 = n29701 ^ n27915;
  assign n29704 = n29703 ^ n29702;
  assign n30321 = n29654 ^ n29653;
  assign n30312 = n29651 ^ n2280;
  assign n30271 = n28986 ^ n27930;
  assign n30272 = n29810 ^ n28986;
  assign n30273 = n30271 & n30272;
  assign n30274 = n30273 ^ n27930;
  assign n29934 = n29933 ^ n26815;
  assign n30057 = n30056 ^ n29933;
  assign n30058 = n29934 & n30057;
  assign n30059 = n30058 ^ n26815;
  assign n29921 = n28246 ^ n27323;
  assign n29922 = n28900 ^ n28246;
  assign n29923 = ~n29921 & n29922;
  assign n29924 = n29923 ^ n27323;
  assign n29919 = n29467 ^ n29392;
  assign n29717 = n29716 ^ n29712;
  assign n29916 = n29915 ^ n29712;
  assign n29917 = n29717 & n29916;
  assign n29918 = n29917 ^ n29716;
  assign n29920 = n29919 ^ n29918;
  assign n29930 = n29924 ^ n29920;
  assign n29931 = n29930 ^ n26729;
  assign n30119 = n30059 ^ n29931;
  assign n30118 = n30065 & n30117;
  assign n30122 = n30119 ^ n30118;
  assign n30126 = n30125 ^ n30122;
  assign n30263 = n30262 ^ n30127;
  assign n30264 = n30131 & ~n30263;
  assign n30265 = n30264 ^ n30130;
  assign n30266 = n30265 ^ n30122;
  assign n30267 = ~n30126 & n30266;
  assign n30268 = n30267 ^ n30125;
  assign n30269 = n30268 ^ n2268;
  assign n30120 = n30118 & ~n30119;
  assign n30060 = n30059 ^ n29930;
  assign n30061 = n29931 & ~n30060;
  assign n30062 = n30061 ^ n26729;
  assign n29925 = n29924 ^ n29919;
  assign n29926 = ~n29920 & ~n29925;
  assign n29927 = n29926 ^ n29924;
  assign n29709 = n29470 ^ n29387;
  assign n29705 = n27955 ^ n27317;
  assign n29706 = n28894 ^ n27955;
  assign n29707 = n29705 & ~n29706;
  assign n29708 = n29707 ^ n27317;
  assign n29710 = n29709 ^ n29708;
  assign n29928 = n29927 ^ n29710;
  assign n29929 = n29928 ^ n26725;
  assign n30063 = n30062 ^ n29929;
  assign n30121 = n30120 ^ n30063;
  assign n30270 = n30269 ^ n30121;
  assign n30275 = n30274 ^ n30270;
  assign n30300 = n30265 ^ n30126;
  assign n30297 = n30296 ^ n30294;
  assign n30298 = n30295 & ~n30297;
  assign n30299 = n30298 ^ n30279;
  assign n30301 = n30300 ^ n30299;
  assign n30302 = n28819 ^ n27936;
  assign n30303 = n29817 ^ n28819;
  assign n30304 = n30302 & n30303;
  assign n30305 = n30304 ^ n27936;
  assign n30306 = n30305 ^ n30299;
  assign n30307 = ~n30301 & ~n30306;
  assign n30308 = n30307 ^ n30300;
  assign n30309 = n30308 ^ n30270;
  assign n30310 = n30275 & ~n30309;
  assign n30311 = n30310 ^ n30274;
  assign n30313 = n30312 ^ n30311;
  assign n30314 = n29087 ^ n27923;
  assign n30315 = n29804 ^ n29087;
  assign n30316 = ~n30314 & ~n30315;
  assign n30317 = n30316 ^ n27923;
  assign n30318 = n30317 ^ n30312;
  assign n30319 = ~n30313 & ~n30318;
  assign n30320 = n30319 ^ n30317;
  assign n30322 = n30321 ^ n30320;
  assign n30323 = n29154 ^ n27917;
  assign n30324 = n29794 ^ n29154;
  assign n30325 = ~n30323 & n30324;
  assign n30326 = n30325 ^ n27917;
  assign n30327 = n30326 ^ n30321;
  assign n30328 = ~n30322 & n30327;
  assign n30329 = n30328 ^ n30326;
  assign n30330 = n30329 ^ n29702;
  assign n30331 = ~n29704 & ~n30330;
  assign n30332 = n30331 ^ n29703;
  assign n30337 = n30336 ^ n30332;
  assign n30338 = n29664 ^ n29650;
  assign n30339 = n30338 ^ n30332;
  assign n30340 = ~n30337 & n30339;
  assign n30341 = n30340 ^ n30338;
  assign n30342 = n30341 ^ n29693;
  assign n30343 = n29696 & ~n30342;
  assign n30344 = n30343 ^ n29695;
  assign n30345 = n30344 ^ n29687;
  assign n30346 = n29688 & n30345;
  assign n30347 = n30346 ^ n29686;
  assign n30348 = n30347 ^ n29106;
  assign n30349 = n29681 & n30348;
  assign n30350 = n30349 ^ n29680;
  assign n30352 = n30351 ^ n30350;
  assign n28814 = n28813 ^ n27886;
  assign n29098 = n29097 ^ n28813;
  assign n29099 = ~n28814 & ~n29098;
  assign n29100 = n29099 ^ n27886;
  assign n30419 = n30351 ^ n29100;
  assign n30420 = n30352 & ~n30419;
  assign n30421 = n30420 ^ n29100;
  assign n30575 = n30427 ^ n30421;
  assign n30576 = ~n30428 & n30575;
  assign n30577 = n30576 ^ n30425;
  assign n30573 = n30194 ^ n30191;
  assign n30753 = n30577 ^ n30573;
  assign n30569 = n29124 ^ n27879;
  assign n30570 = n29756 ^ n29124;
  assign n30571 = ~n30569 & ~n30570;
  assign n30572 = n30571 ^ n27879;
  assign n30754 = n30577 ^ n30572;
  assign n30755 = ~n30753 & ~n30754;
  assign n30756 = n30755 ^ n30573;
  assign n30662 = n30197 ^ n30170;
  assign n30757 = n30756 ^ n30662;
  assign n30758 = n29113 ^ n27872;
  assign n30759 = n29751 ^ n29113;
  assign n30760 = n30758 & n30759;
  assign n30761 = n30760 ^ n27872;
  assign n30762 = n30761 ^ n30662;
  assign n30763 = ~n30757 & n30762;
  assign n30764 = n30763 ^ n30761;
  assign n30765 = n30764 ^ n30656;
  assign n30766 = ~n30752 & ~n30765;
  assign n30767 = n30766 ^ n30751;
  assign n30768 = n30767 ^ n30647;
  assign n30769 = n30747 & n30768;
  assign n30770 = n30769 ^ n30746;
  assign n30641 = n30206 ^ n30164;
  assign n30771 = n30770 ^ n30641;
  assign n30772 = n29224 ^ n27848;
  assign n30773 = n29745 ^ n29224;
  assign n30774 = ~n30772 & n30773;
  assign n30775 = n30774 ^ n27848;
  assign n30776 = n30775 ^ n30641;
  assign n30777 = n30771 & n30776;
  assign n30778 = n30777 ^ n30775;
  assign n30634 = n30210 ^ n1216;
  assign n30779 = n30778 ^ n30634;
  assign n30780 = n29307 ^ n28338;
  assign n30781 = n29743 ^ n29307;
  assign n30782 = n30780 & ~n30781;
  assign n30783 = n30782 ^ n28338;
  assign n30784 = n30783 ^ n30634;
  assign n30785 = ~n30779 & ~n30784;
  assign n30786 = n30785 ^ n30783;
  assign n30787 = n30786 ^ n30623;
  assign n30788 = n30742 & ~n30787;
  assign n30789 = n30788 ^ n30741;
  assign n30790 = n30789 ^ n30736;
  assign n30791 = ~n30737 & ~n30790;
  assign n30792 = n30791 ^ n30616;
  assign n30793 = n30792 ^ n30604;
  assign n30794 = ~n30732 & ~n30793;
  assign n30795 = n30794 ^ n30731;
  assign n30723 = n29532 ^ n28850;
  assign n30724 = n29719 ^ n29532;
  assign n30725 = n30723 & n30724;
  assign n30726 = n30725 ^ n28850;
  assign n30596 = n30227 ^ n30157;
  assign n30727 = n30726 ^ n30596;
  assign n30837 = n30795 ^ n30727;
  assign n30838 = n30837 ^ n27269;
  assign n30839 = n30792 ^ n30731;
  assign n30840 = n30839 ^ n30604;
  assign n30841 = n30840 ^ n27852;
  assign n30842 = n30789 ^ n30737;
  assign n30843 = n30842 ^ n27859;
  assign n30844 = n30786 ^ n30742;
  assign n30845 = n30844 ^ n27867;
  assign n30846 = n30783 ^ n30779;
  assign n30847 = n30846 ^ n27875;
  assign n30848 = n30775 ^ n30771;
  assign n30849 = n30848 ^ n27985;
  assign n30850 = n30767 ^ n30747;
  assign n30851 = n30850 ^ n27882;
  assign n30852 = n30764 ^ n30752;
  assign n30853 = n30852 ^ n27889;
  assign n30854 = n30761 ^ n30757;
  assign n30855 = n30854 ^ n27897;
  assign n30574 = n30573 ^ n30572;
  assign n30578 = n30577 ^ n30574;
  assign n30579 = n30578 ^ n28002;
  assign n30429 = n30428 ^ n30421;
  assign n30430 = n30429 ^ n27837;
  assign n30357 = n30341 ^ n29696;
  assign n30358 = n30357 ^ n27274;
  assign n30359 = n30329 ^ n29704;
  assign n30360 = n30359 ^ n27276;
  assign n30361 = n30326 ^ n30322;
  assign n30362 = n30361 ^ n27282;
  assign n30363 = n30317 ^ n30313;
  assign n30364 = n30363 ^ n27289;
  assign n30365 = n30308 ^ n30274;
  assign n30366 = n30365 ^ n30270;
  assign n30367 = n30366 ^ n27295;
  assign n30377 = n30376 ^ n30374;
  assign n30378 = n30375 & ~n30377;
  assign n30379 = n30378 ^ n27308;
  assign n30380 = n30379 ^ n27301;
  assign n30381 = n30305 ^ n30300;
  assign n30382 = n30381 ^ n30299;
  assign n30383 = n30382 ^ n30379;
  assign n30384 = ~n30380 & n30383;
  assign n30385 = n30384 ^ n27301;
  assign n30386 = n30385 ^ n30366;
  assign n30387 = n30367 & ~n30386;
  assign n30388 = n30387 ^ n27295;
  assign n30389 = n30388 ^ n30363;
  assign n30390 = n30364 & n30389;
  assign n30391 = n30390 ^ n27289;
  assign n30392 = n30391 ^ n30361;
  assign n30393 = ~n30362 & ~n30392;
  assign n30394 = n30393 ^ n27282;
  assign n30395 = n30394 ^ n30359;
  assign n30396 = ~n30360 & ~n30395;
  assign n30397 = n30396 ^ n27276;
  assign n30398 = n30397 ^ n27275;
  assign n30399 = n30338 ^ n30336;
  assign n30400 = n30399 ^ n30332;
  assign n30401 = n30400 ^ n30397;
  assign n30402 = ~n30398 & n30401;
  assign n30403 = n30402 ^ n27275;
  assign n30404 = n30403 ^ n30357;
  assign n30405 = ~n30358 & ~n30404;
  assign n30406 = n30405 ^ n27274;
  assign n30355 = n30344 ^ n29686;
  assign n30356 = n30355 ^ n29687;
  assign n30407 = n30406 ^ n30356;
  assign n30408 = n30356 ^ n27273;
  assign n30409 = n30407 & n30408;
  assign n30410 = n30409 ^ n27273;
  assign n30354 = n30347 ^ n29681;
  assign n30411 = n30410 ^ n30354;
  assign n30412 = n30354 ^ n27681;
  assign n30413 = n30411 & ~n30412;
  assign n30414 = n30413 ^ n27681;
  assign n30353 = n30352 ^ n29100;
  assign n30415 = n30414 ^ n30353;
  assign n30416 = n30353 ^ n27697;
  assign n30417 = n30415 & n30416;
  assign n30418 = n30417 ^ n27697;
  assign n30566 = n30429 ^ n30418;
  assign n30567 = n30430 & ~n30566;
  assign n30568 = n30567 ^ n27837;
  assign n30856 = n30578 ^ n30568;
  assign n30857 = n30579 & ~n30856;
  assign n30858 = n30857 ^ n28002;
  assign n30859 = n30858 ^ n30854;
  assign n30860 = ~n30855 & ~n30859;
  assign n30861 = n30860 ^ n27897;
  assign n30862 = n30861 ^ n30852;
  assign n30863 = ~n30853 & ~n30862;
  assign n30864 = n30863 ^ n27889;
  assign n30865 = n30864 ^ n30850;
  assign n30866 = n30851 & n30865;
  assign n30867 = n30866 ^ n27882;
  assign n30868 = n30867 ^ n30848;
  assign n30869 = n30849 & n30868;
  assign n30870 = n30869 ^ n27985;
  assign n30871 = n30870 ^ n30846;
  assign n30872 = n30847 & ~n30871;
  assign n30873 = n30872 ^ n27875;
  assign n30874 = n30873 ^ n30844;
  assign n30875 = ~n30845 & ~n30874;
  assign n30876 = n30875 ^ n27867;
  assign n30877 = n30876 ^ n30842;
  assign n30878 = n30843 & ~n30877;
  assign n30879 = n30878 ^ n27859;
  assign n30880 = n30879 ^ n30840;
  assign n30881 = ~n30841 & n30880;
  assign n30882 = n30881 ^ n27852;
  assign n30883 = n30882 ^ n30837;
  assign n30884 = ~n30838 & ~n30883;
  assign n30885 = n30884 ^ n27269;
  assign n30796 = n30795 ^ n30596;
  assign n30797 = ~n30727 & ~n30796;
  assign n30798 = n30797 ^ n30726;
  assign n30718 = n29577 ^ n28864;
  assign n30719 = n29712 ^ n29577;
  assign n30720 = ~n30718 & n30719;
  assign n30721 = n30720 ^ n28864;
  assign n30835 = n30798 ^ n30721;
  assign n30585 = n30231 ^ n3069;
  assign n30836 = n30835 ^ n30585;
  assign n30886 = n30885 ^ n30836;
  assign n30887 = n30836 ^ n28128;
  assign n30888 = n30886 & ~n30887;
  assign n30889 = n30888 ^ n28128;
  assign n30722 = n30721 ^ n30585;
  assign n30799 = n30798 ^ n30585;
  assign n30800 = n30722 & n30799;
  assign n30801 = n30800 ^ n30721;
  assign n30713 = n28727 ^ n28226;
  assign n30714 = n29919 ^ n28727;
  assign n30715 = n30713 & n30714;
  assign n30716 = n30715 ^ n28226;
  assign n30712 = n30234 ^ n30154;
  assign n30717 = n30716 ^ n30712;
  assign n30833 = n30801 ^ n30717;
  assign n30834 = n30833 ^ n27469;
  assign n30919 = n30889 ^ n30834;
  assign n30920 = n30882 ^ n27269;
  assign n30921 = n30920 ^ n30837;
  assign n30922 = n30879 ^ n30841;
  assign n30923 = n30876 ^ n30843;
  assign n30924 = n30873 ^ n30845;
  assign n30925 = n30858 ^ n30855;
  assign n30431 = n30430 ^ n30418;
  assign n30432 = n30415 ^ n27697;
  assign n30433 = n30403 ^ n30358;
  assign n30434 = n30400 ^ n27275;
  assign n30435 = n30434 ^ n30397;
  assign n30436 = n30394 ^ n30360;
  assign n30437 = n30391 ^ n27282;
  assign n30438 = n30437 ^ n30361;
  assign n30439 = n30385 ^ n27295;
  assign n30440 = n30439 ^ n30366;
  assign n30442 = n30382 ^ n27301;
  assign n30443 = n30442 ^ n30379;
  assign n30444 = ~n30441 & ~n30443;
  assign n30445 = n30440 & n30444;
  assign n30446 = n30388 ^ n27289;
  assign n30447 = n30446 ^ n30363;
  assign n30448 = ~n30445 & ~n30447;
  assign n30449 = n30438 & ~n30448;
  assign n30450 = ~n30436 & n30449;
  assign n30451 = n30435 & ~n30450;
  assign n30452 = n30433 & n30451;
  assign n30453 = n30407 ^ n27273;
  assign n30454 = ~n30452 & ~n30453;
  assign n30455 = n30411 ^ n27681;
  assign n30456 = n30454 & ~n30455;
  assign n30457 = n30432 & n30456;
  assign n30565 = ~n30431 & n30457;
  assign n30580 = n30579 ^ n30568;
  assign n30926 = ~n30565 & n30580;
  assign n30927 = n30925 & ~n30926;
  assign n30928 = n30861 ^ n30853;
  assign n30929 = n30927 & ~n30928;
  assign n30930 = n30864 ^ n30851;
  assign n30931 = n30929 & ~n30930;
  assign n30932 = n30867 ^ n30849;
  assign n30933 = ~n30931 & ~n30932;
  assign n30934 = n30870 ^ n30847;
  assign n30935 = ~n30933 & ~n30934;
  assign n30936 = n30924 & n30935;
  assign n30937 = ~n30923 & ~n30936;
  assign n30938 = n30922 & n30937;
  assign n30939 = n30921 & n30938;
  assign n30940 = n30886 ^ n28128;
  assign n30941 = ~n30939 & n30940;
  assign n30942 = ~n30919 & n30941;
  assign n30890 = n30889 ^ n30833;
  assign n30891 = n30834 & ~n30890;
  assign n30892 = n30891 ^ n27469;
  assign n30802 = n30801 ^ n30716;
  assign n30803 = n30717 & n30802;
  assign n30804 = n30803 ^ n30712;
  assign n30707 = n28757 ^ n28233;
  assign n30708 = n29709 ^ n28757;
  assign n30709 = n30707 & n30708;
  assign n30710 = n30709 ^ n28233;
  assign n30706 = n30237 ^ n30152;
  assign n30711 = n30710 ^ n30706;
  assign n30831 = n30804 ^ n30711;
  assign n30832 = n30831 ^ n27476;
  assign n30918 = n30892 ^ n30832;
  assign n31066 = n30942 ^ n30918;
  assign n31068 = n31066 ^ n31065;
  assign n31053 = n30940 ^ n30939;
  assign n31055 = n2885 & n31053;
  assign n31051 = n30941 ^ n30919;
  assign n31074 = n31051 ^ n31050;
  assign n31075 = ~n31055 & n31074;
  assign n31052 = ~n31050 & ~n31051;
  assign n31076 = n31075 ^ n31052;
  assign n30979 = n30926 ^ n30925;
  assign n1366 = n1323 ^ n1263;
  assign n1367 = n1366 ^ n1360;
  assign n1371 = n1370 ^ n1367;
  assign n30980 = n30979 ^ n1371;
  assign n30581 = n30580 ^ n30565;
  assign n1348 = n1308 ^ n1245;
  assign n1349 = n1348 ^ n1345;
  assign n1353 = n1352 ^ n1349;
  assign n30582 = n30581 ^ n1353;
  assign n1330 = n1230 ^ n1156;
  assign n1337 = n1336 ^ n1330;
  assign n1338 = n1337 ^ n1085;
  assign n30458 = n30457 ^ n30431;
  assign n30459 = ~n1338 & ~n30458;
  assign n30460 = n30456 ^ n30432;
  assign n30462 = n30460 ^ n3347;
  assign n30461 = n3347 & ~n30460;
  assign n30463 = n30462 ^ n30461;
  assign n30464 = ~n30459 & ~n30463;
  assign n30465 = n30453 ^ n30452;
  assign n30466 = n30465 ^ n812;
  assign n30470 = n30451 ^ n30433;
  assign n30467 = n28604 ^ n21410;
  assign n30468 = n30467 ^ n668;
  assign n30469 = n30468 ^ n802;
  assign n30472 = n30470 ^ n30469;
  assign n30473 = n30450 ^ n30435;
  assign n615 = n614 ^ n605;
  assign n628 = n627 ^ n615;
  assign n632 = n631 ^ n628;
  assign n30475 = n30473 ^ n632;
  assign n30474 = ~n632 & n30473;
  assign n30476 = n30475 ^ n30474;
  assign n30477 = n30472 & ~n30476;
  assign n30471 = ~n30469 & ~n30470;
  assign n30478 = n30477 ^ n30471;
  assign n30479 = n30478 ^ n30465;
  assign n30480 = ~n30466 & ~n30479;
  assign n30481 = n30480 ^ n812;
  assign n30485 = n30455 ^ n30454;
  assign n30487 = n30485 ^ n30484;
  assign n30486 = ~n30484 & ~n30485;
  assign n30488 = n30487 ^ n30486;
  assign n30489 = ~n30481 & n30488;
  assign n30493 = n30449 ^ n30436;
  assign n30497 = n30496 ^ n30493;
  assign n30499 = n28616 ^ n576;
  assign n30500 = n30499 ^ n25004;
  assign n30501 = n30500 ^ n3260;
  assign n30498 = n30448 ^ n30438;
  assign n30502 = n30501 ^ n30498;
  assign n30503 = n30447 ^ n30445;
  assign n30507 = n30506 ^ n30503;
  assign n30509 = n28621 ^ n21375;
  assign n30510 = n30509 ^ n25010;
  assign n30511 = n30510 ^ n20274;
  assign n30508 = n30444 ^ n30440;
  assign n30512 = n30511 ^ n30508;
  assign n30527 = n30526 ^ n30523;
  assign n30528 = n30523 ^ n30441;
  assign n30529 = n30527 & n30528;
  assign n30530 = n30529 ^ n30526;
  assign n30513 = n30443 ^ n30441;
  assign n30531 = n30530 ^ n30513;
  assign n30532 = n28639 ^ n21380;
  assign n30533 = n30532 ^ n25015;
  assign n30534 = n30533 ^ n20279;
  assign n30535 = n30534 ^ n30513;
  assign n30536 = n30531 & ~n30535;
  assign n30537 = n30536 ^ n30534;
  assign n30538 = n30537 ^ n30508;
  assign n30539 = ~n30512 & n30538;
  assign n30540 = n30539 ^ n30511;
  assign n30541 = n30540 ^ n30503;
  assign n30542 = n30507 & ~n30541;
  assign n30543 = n30542 ^ n30506;
  assign n30544 = n30543 ^ n30498;
  assign n30545 = n30502 & ~n30544;
  assign n30546 = n30545 ^ n30501;
  assign n30547 = n30546 ^ n30493;
  assign n30548 = n30497 & ~n30547;
  assign n30549 = n30548 ^ n30496;
  assign n30490 = ~n812 & n30465;
  assign n30491 = ~n30471 & ~n30474;
  assign n30492 = ~n30490 & n30491;
  assign n30550 = n30549 ^ n30492;
  assign n30551 = n30492 ^ n30486;
  assign n30552 = n30492 & ~n30551;
  assign n30553 = n30552 ^ n30492;
  assign n30554 = n30550 & n30553;
  assign n30555 = n30554 ^ n30552;
  assign n30556 = n30555 ^ n30492;
  assign n30557 = n30556 ^ n30486;
  assign n30558 = n30489 & ~n30557;
  assign n30559 = n30558 ^ n30486;
  assign n30560 = n30464 & ~n30559;
  assign n30561 = n30458 ^ n1338;
  assign n30562 = ~n30461 & n30561;
  assign n30563 = n30562 ^ n30459;
  assign n30564 = ~n30560 & n30563;
  assign n30981 = n30581 ^ n30564;
  assign n30982 = ~n30582 & ~n30981;
  assign n30983 = n30982 ^ n1353;
  assign n30984 = n30983 ^ n30979;
  assign n30985 = n30980 & ~n30984;
  assign n30986 = n30985 ^ n1371;
  assign n2675 = n2623 ^ n1565;
  assign n2676 = n2675 ^ n2672;
  assign n2680 = n2679 ^ n2676;
  assign n30987 = n30936 ^ n30923;
  assign n30988 = ~n2680 & ~n30987;
  assign n2648 = n2641 ^ n2614;
  assign n2661 = n2660 ^ n2648;
  assign n2665 = n2664 ^ n2661;
  assign n30989 = n30935 ^ n30924;
  assign n30991 = n2665 & ~n30989;
  assign n30990 = n30989 ^ n2665;
  assign n30992 = n30991 ^ n30990;
  assign n30993 = ~n30988 & ~n30992;
  assign n30997 = n30932 ^ n30931;
  assign n30998 = ~n30996 & ~n30997;
  assign n30999 = n21352 ^ n1427;
  assign n31000 = n30999 ^ n3017;
  assign n31001 = n31000 ^ n2414;
  assign n31002 = n30928 ^ n30927;
  assign n31003 = ~n31001 & ~n31002;
  assign n31004 = n28588 ^ n3163;
  assign n31005 = n31004 ^ n25449;
  assign n31006 = n31005 ^ n3029;
  assign n31007 = n30930 ^ n30929;
  assign n31008 = ~n31006 & ~n31007;
  assign n31009 = ~n31003 & ~n31008;
  assign n3181 = n3177 ^ n2564;
  assign n3188 = n3187 ^ n3181;
  assign n3189 = n3188 ^ n2657;
  assign n31010 = n30934 ^ n30933;
  assign n31011 = ~n3189 & n31010;
  assign n31012 = n31009 & ~n31011;
  assign n31013 = ~n30998 & n31012;
  assign n31014 = n30938 ^ n30921;
  assign n31015 = ~n3125 & ~n31014;
  assign n31016 = n31013 & ~n31015;
  assign n31017 = n30937 ^ n30922;
  assign n2755 = n2747 ^ n2700;
  assign n2759 = n2758 ^ n2755;
  assign n2760 = n2759 ^ n1527;
  assign n31019 = n31017 ^ n2760;
  assign n31018 = n2760 & n31017;
  assign n31020 = n31019 ^ n31018;
  assign n31021 = n31016 & n31020;
  assign n31022 = n30993 & n31021;
  assign n31023 = n30986 & n31022;
  assign n31024 = n31014 ^ n3125;
  assign n31025 = n31010 ^ n3189;
  assign n31026 = n30997 ^ n30996;
  assign n31027 = n31007 ^ n31006;
  assign n31028 = n31002 ^ n31001;
  assign n31029 = n31028 ^ n31003;
  assign n31030 = n31027 & n31029;
  assign n31031 = n31030 ^ n31008;
  assign n31032 = n31031 ^ n30997;
  assign n31033 = n31026 & n31032;
  assign n31034 = n31033 ^ n30996;
  assign n31035 = ~n31025 & ~n31034;
  assign n31036 = n31035 ^ n31011;
  assign n31037 = n30993 & ~n31036;
  assign n31038 = n30987 ^ n2680;
  assign n31039 = ~n30991 & n31038;
  assign n31040 = n31039 ^ n30988;
  assign n31041 = ~n31037 & n31040;
  assign n31042 = n31019 & ~n31041;
  assign n31043 = n31042 ^ n31018;
  assign n31044 = n31043 ^ n31014;
  assign n31045 = n31024 & ~n31044;
  assign n31046 = n31045 ^ n3125;
  assign n31047 = ~n31023 & ~n31046;
  assign n31054 = n31053 ^ n2885;
  assign n31056 = n31055 ^ n31054;
  assign n31057 = ~n31052 & n31056;
  assign n31114 = ~n31047 & n31057;
  assign n31115 = n31076 & ~n31114;
  assign n31116 = n31068 & ~n31115;
  assign n31067 = n31065 & n31066;
  assign n31117 = n31116 ^ n31067;
  assign n30893 = n30892 ^ n30831;
  assign n30894 = n30832 & ~n30893;
  assign n30895 = n30894 ^ n27476;
  assign n30809 = n28799 ^ n28220;
  assign n30810 = n29510 ^ n28799;
  assign n30811 = ~n30809 & n30810;
  assign n30812 = n30811 ^ n28220;
  assign n30805 = n30804 ^ n30710;
  assign n30806 = ~n30711 & n30805;
  assign n30807 = n30806 ^ n30706;
  assign n30705 = n30240 ^ n30150;
  assign n30808 = n30807 ^ n30705;
  assign n30829 = n30812 ^ n30808;
  assign n30830 = n30829 ^ n27464;
  assign n30944 = n30895 ^ n30830;
  assign n30943 = ~n30918 & n30942;
  assign n31058 = n30944 ^ n30943;
  assign n31073 = n31061 ^ n31058;
  assign n31118 = n31117 ^ n31073;
  assign n31110 = n28921 ^ n28811;
  assign n31111 = n30312 ^ n28811;
  assign n31112 = ~n31110 & ~n31111;
  assign n31113 = n31112 ^ n28921;
  assign n31227 = n31118 ^ n31113;
  assign n31411 = n31227 ^ n27949;
  assign n2244 = n2220 ^ n2143;
  assign n2245 = n2244 ^ n2108;
  assign n2246 = n2245 ^ n2236;
  assign n31602 = n31411 ^ n2246;
  assign n32435 = n31602 ^ n30685;
  assign n32436 = n32434 & ~n32435;
  assign n32437 = n32436 ^ n29703;
  assign n30615 = n29745 ^ n29207;
  assign n30617 = n30616 ^ n29745;
  assign n30618 = n30615 & ~n30617;
  assign n30619 = n30618 ^ n29207;
  assign n30609 = n30491 & n30549;
  assign n30610 = n30478 & ~n30609;
  assign n30611 = n30610 ^ n30465;
  assign n30612 = ~n30466 & ~n30611;
  assign n30613 = n30612 ^ n812;
  assign n30614 = n30613 ^ n30487;
  assign n30620 = n30619 ^ n30614;
  assign n30622 = n29884 ^ n29113;
  assign n30624 = n30623 ^ n29884;
  assign n30625 = ~n30622 & n30624;
  assign n30626 = n30625 ^ n29113;
  assign n30621 = n30610 ^ n30466;
  assign n30627 = n30626 ^ n30621;
  assign n30633 = n29875 ^ n29124;
  assign n30635 = n30634 ^ n29875;
  assign n30636 = ~n30633 & ~n30635;
  assign n30637 = n30636 ^ n29124;
  assign n30628 = n30549 ^ n30473;
  assign n30629 = ~n30475 & n30628;
  assign n30630 = n30629 ^ n632;
  assign n30631 = n30630 ^ n30469;
  assign n30632 = n30631 ^ n30470;
  assign n30638 = n30637 ^ n30632;
  assign n30640 = n29751 ^ n29126;
  assign n30642 = n30641 ^ n29751;
  assign n30643 = n30640 & ~n30642;
  assign n30644 = n30643 ^ n29126;
  assign n30639 = n30549 ^ n30475;
  assign n30645 = n30644 ^ n30639;
  assign n30651 = n30546 ^ n30497;
  assign n30646 = n29756 ^ n28813;
  assign n30648 = n30647 ^ n29756;
  assign n30649 = n30646 & ~n30648;
  assign n30650 = n30649 ^ n28813;
  assign n30652 = n30651 ^ n30650;
  assign n30654 = n29762 ^ n29101;
  assign n30657 = n30656 ^ n29762;
  assign n30658 = n30654 & ~n30657;
  assign n30659 = n30658 ^ n29101;
  assign n30653 = n30543 ^ n30502;
  assign n30660 = n30659 ^ n30653;
  assign n30666 = n30540 ^ n30507;
  assign n30661 = n29178 ^ n29097;
  assign n30663 = n30662 ^ n29097;
  assign n30664 = n30661 & ~n30663;
  assign n30665 = n30664 ^ n29178;
  assign n30667 = n30666 ^ n30665;
  assign n30672 = n30537 ^ n30512;
  assign n30668 = n29136 ^ n29103;
  assign n30669 = n30573 ^ n29103;
  assign n30670 = ~n30668 & n30669;
  assign n30671 = n30670 ^ n29136;
  assign n30673 = n30672 ^ n30671;
  assign n30678 = n30534 ^ n30531;
  assign n30674 = n29683 ^ n29142;
  assign n30675 = n30427 ^ n29683;
  assign n30676 = ~n30674 & ~n30675;
  assign n30677 = n30676 ^ n29142;
  assign n30679 = n30678 ^ n30677;
  assign n30680 = n29690 ^ n29148;
  assign n30681 = n30351 ^ n29690;
  assign n30682 = ~n30680 & n30681;
  assign n30683 = n30682 ^ n29148;
  assign n30686 = n30685 ^ n30683;
  assign n30688 = n29787 ^ n29154;
  assign n30689 = n29787 ^ n29680;
  assign n30690 = ~n30688 & n30689;
  assign n30691 = n30690 ^ n29154;
  assign n30687 = n30520 ^ n30519;
  assign n30692 = n30691 ^ n30687;
  assign n30694 = n29699 ^ n29087;
  assign n30695 = n29699 ^ n29687;
  assign n30696 = n30694 & n30695;
  assign n30697 = n30696 ^ n29087;
  assign n30693 = n30514 ^ n2135;
  assign n30698 = n30697 ^ n30693;
  assign n31093 = n29794 ^ n28986;
  assign n31094 = n29794 ^ n29695;
  assign n31095 = ~n31093 & n31094;
  assign n31096 = n31095 ^ n28986;
  assign n30945 = n30943 & n30944;
  assign n30896 = n30895 ^ n30829;
  assign n30897 = ~n30830 & ~n30896;
  assign n30898 = n30897 ^ n27464;
  assign n30813 = n30812 ^ n30705;
  assign n30814 = ~n30808 & ~n30813;
  assign n30815 = n30814 ^ n30812;
  assign n30700 = n28900 ^ n28213;
  assign n30701 = n29504 ^ n28900;
  assign n30702 = n30700 & n30701;
  assign n30703 = n30702 ^ n28213;
  assign n30699 = n30243 ^ n30145;
  assign n30704 = n30703 ^ n30699;
  assign n30827 = n30815 ^ n30704;
  assign n30828 = n30827 ^ n27458;
  assign n30946 = n30898 ^ n30828;
  assign n30947 = ~n30945 & n30946;
  assign n30899 = n30898 ^ n30827;
  assign n30900 = ~n30828 & n30899;
  assign n30901 = n30900 ^ n27458;
  assign n30820 = n28894 ^ n28207;
  assign n30821 = n29498 ^ n28894;
  assign n30822 = ~n30820 & ~n30821;
  assign n30823 = n30822 ^ n28207;
  assign n30819 = n30246 ^ n30143;
  assign n30824 = n30823 ^ n30819;
  assign n30816 = n30815 ^ n30703;
  assign n30817 = n30704 & n30816;
  assign n30818 = n30817 ^ n30699;
  assign n30825 = n30824 ^ n30818;
  assign n30826 = n30825 ^ n27452;
  assign n30948 = n30901 ^ n30826;
  assign n30949 = n30947 & n30948;
  assign n30913 = n30249 ^ n3009;
  assign n30914 = n30913 ^ n30140;
  assign n30909 = n30819 ^ n30818;
  assign n30910 = n30824 & ~n30909;
  assign n30911 = n30910 ^ n30823;
  assign n30905 = n28844 ^ n28246;
  assign n30906 = n29544 ^ n28844;
  assign n30907 = ~n30905 & ~n30906;
  assign n30908 = n30907 ^ n28246;
  assign n30912 = n30911 ^ n30908;
  assign n30915 = n30914 ^ n30912;
  assign n30916 = n30915 ^ n27323;
  assign n30902 = n30901 ^ n30825;
  assign n30903 = ~n30826 & ~n30902;
  assign n30904 = n30903 ^ n27452;
  assign n30917 = n30916 ^ n30904;
  assign n30973 = n30949 ^ n30917;
  assign n1973 = n1952 ^ n1896;
  assign n1977 = n1976 ^ n1973;
  assign n1978 = n1977 ^ n1966;
  assign n30974 = n30973 ^ n1978;
  assign n30975 = n30948 ^ n30947;
  assign n1862 = n1831 ^ n1801;
  assign n1863 = n1862 ^ n1859;
  assign n1867 = n1866 ^ n1863;
  assign n30976 = n30975 ^ n1867;
  assign n30977 = n30946 ^ n30945;
  assign n1850 = n1822 ^ n1786;
  assign n1851 = n1850 ^ n1849;
  assign n1852 = n1851 ^ n1840;
  assign n30978 = n30977 ^ n1852;
  assign n31062 = n31058 & ~n31061;
  assign n31069 = n31068 ^ n31067;
  assign n31070 = ~n31062 & n31069;
  assign n31071 = n31057 & n31070;
  assign n31072 = ~n31047 & n31071;
  assign n31077 = n31068 & n31076;
  assign n31078 = n31077 ^ n31069;
  assign n31079 = n31078 ^ n31058;
  assign n31080 = ~n31073 & n31079;
  assign n31081 = n31080 ^ n31061;
  assign n31082 = ~n31072 & ~n31081;
  assign n31083 = n31082 ^ n30977;
  assign n31084 = ~n30978 & ~n31083;
  assign n31085 = n31084 ^ n1852;
  assign n31086 = n31085 ^ n30975;
  assign n31087 = n30976 & ~n31086;
  assign n31088 = n31087 ^ n1867;
  assign n31089 = n31088 ^ n30973;
  assign n31090 = n30974 & ~n31089;
  assign n31091 = n31090 ^ n1978;
  assign n30969 = n28885 ^ n2375;
  assign n30970 = n30969 ^ n1971;
  assign n30971 = n30970 ^ n2124;
  assign n30962 = n30904 ^ n27323;
  assign n30963 = n30915 ^ n30904;
  assign n30964 = ~n30962 & n30963;
  assign n30965 = n30964 ^ n27323;
  assign n30966 = n30965 ^ n27317;
  assign n30960 = n30253 ^ n1689;
  assign n30955 = n30914 ^ n30908;
  assign n30956 = n30914 ^ n30911;
  assign n30957 = n30955 & n30956;
  assign n30958 = n30957 ^ n30908;
  assign n30951 = n28838 ^ n27955;
  assign n30952 = n29595 ^ n28838;
  assign n30953 = n30951 & ~n30952;
  assign n30954 = n30953 ^ n27955;
  assign n30959 = n30958 ^ n30954;
  assign n30961 = n30960 ^ n30959;
  assign n30967 = n30966 ^ n30961;
  assign n30950 = n30917 & n30949;
  assign n30968 = n30967 ^ n30950;
  assign n30972 = n30971 ^ n30968;
  assign n31092 = n31091 ^ n30972;
  assign n31097 = n31096 ^ n31092;
  assign n31102 = n31088 ^ n30974;
  assign n31098 = n29804 ^ n28819;
  assign n31099 = n30338 ^ n29804;
  assign n31100 = ~n31098 & ~n31099;
  assign n31101 = n31100 ^ n28819;
  assign n31103 = n31102 ^ n31101;
  assign n31108 = n31085 ^ n30976;
  assign n31104 = n29810 ^ n28821;
  assign n31105 = n29810 ^ n29703;
  assign n31106 = ~n31104 & n31105;
  assign n31107 = n31106 ^ n28821;
  assign n31109 = n31108 ^ n31107;
  assign n31120 = n29817 ^ n28832;
  assign n31121 = n30321 ^ n29817;
  assign n31122 = ~n31120 & n31121;
  assign n31123 = n31122 ^ n28832;
  assign n31119 = n31113 & ~n31118;
  assign n31124 = n31123 ^ n31119;
  assign n31125 = n31082 ^ n30978;
  assign n31126 = n31125 ^ n31123;
  assign n31127 = n31124 & ~n31126;
  assign n31128 = n31127 ^ n31119;
  assign n31129 = n31128 ^ n31108;
  assign n31130 = ~n31109 & ~n31129;
  assign n31131 = n31130 ^ n31107;
  assign n31132 = n31131 ^ n31102;
  assign n31133 = n31103 & n31132;
  assign n31134 = n31133 ^ n31101;
  assign n31135 = n31134 ^ n31092;
  assign n31136 = n31097 & n31135;
  assign n31137 = n31136 ^ n31096;
  assign n31138 = n31137 ^ n30693;
  assign n31139 = ~n30698 & n31138;
  assign n31140 = n31139 ^ n30697;
  assign n31141 = n31140 ^ n30687;
  assign n31142 = ~n30692 & n31141;
  assign n31143 = n31142 ^ n30691;
  assign n31144 = n31143 ^ n30685;
  assign n31145 = ~n30686 & ~n31144;
  assign n31146 = n31145 ^ n30683;
  assign n31147 = n31146 ^ n30678;
  assign n31148 = n30679 & n31147;
  assign n31149 = n31148 ^ n30677;
  assign n31150 = n31149 ^ n30672;
  assign n31151 = ~n30673 & ~n31150;
  assign n31152 = n31151 ^ n30671;
  assign n31153 = n31152 ^ n30666;
  assign n31154 = n30667 & ~n31153;
  assign n31155 = n31154 ^ n30665;
  assign n31156 = n31155 ^ n30653;
  assign n31157 = n30660 & ~n31156;
  assign n31158 = n31157 ^ n30659;
  assign n31159 = n31158 ^ n30651;
  assign n31160 = n30652 & ~n31159;
  assign n31161 = n31160 ^ n30650;
  assign n31162 = n31161 ^ n30639;
  assign n31163 = n30645 & n31162;
  assign n31164 = n31163 ^ n30644;
  assign n31165 = n31164 ^ n30632;
  assign n31166 = n30638 & n31165;
  assign n31167 = n31166 ^ n30637;
  assign n31168 = n31167 ^ n30621;
  assign n31169 = n30627 & ~n31168;
  assign n31170 = n31169 ^ n30626;
  assign n31171 = n31170 ^ n30614;
  assign n31172 = ~n30620 & ~n31171;
  assign n31173 = n31172 ^ n30619;
  assign n30602 = n29743 ^ n29111;
  assign n30605 = n30604 ^ n29743;
  assign n30606 = n30602 & n30605;
  assign n30607 = n30606 ^ n29111;
  assign n30601 = n30559 ^ n30462;
  assign n30608 = n30607 ^ n30601;
  assign n31195 = n31173 ^ n30608;
  assign n31196 = n31195 ^ n27856;
  assign n31197 = n31170 ^ n30620;
  assign n31198 = n31197 ^ n27864;
  assign n31199 = n31167 ^ n30627;
  assign n31200 = n31199 ^ n27872;
  assign n31201 = n31164 ^ n30638;
  assign n31202 = n31201 ^ n27879;
  assign n31203 = n31161 ^ n30645;
  assign n31204 = n31203 ^ n28308;
  assign n31205 = n31158 ^ n30652;
  assign n31206 = n31205 ^ n27886;
  assign n31207 = n31155 ^ n30660;
  assign n31208 = n31207 ^ n27893;
  assign n31209 = n31152 ^ n30667;
  assign n31210 = n31209 ^ n27902;
  assign n31211 = n31149 ^ n30673;
  assign n31212 = n31211 ^ n28290;
  assign n31213 = n31146 ^ n30679;
  assign n31214 = n31213 ^ n27909;
  assign n31215 = n31143 ^ n30686;
  assign n31216 = n31215 ^ n27915;
  assign n31217 = n31140 ^ n30692;
  assign n31218 = n31217 ^ n27917;
  assign n31219 = n31137 ^ n30698;
  assign n31220 = n31219 ^ n27923;
  assign n31221 = n31134 ^ n31097;
  assign n31222 = n31221 ^ n27930;
  assign n31223 = n31131 ^ n31103;
  assign n31224 = n31223 ^ n27936;
  assign n31225 = n31128 ^ n31109;
  assign n31226 = n31225 ^ n27946;
  assign n31228 = n27949 & ~n31227;
  assign n31229 = n31228 ^ n27948;
  assign n31230 = n31125 ^ n31124;
  assign n31231 = n31230 ^ n31228;
  assign n31232 = n31229 & ~n31231;
  assign n31233 = n31232 ^ n27948;
  assign n31234 = n31233 ^ n31225;
  assign n31235 = ~n31226 & n31234;
  assign n31236 = n31235 ^ n27946;
  assign n31237 = n31236 ^ n31223;
  assign n31238 = ~n31224 & n31237;
  assign n31239 = n31238 ^ n27936;
  assign n31240 = n31239 ^ n31221;
  assign n31241 = ~n31222 & ~n31240;
  assign n31242 = n31241 ^ n27930;
  assign n31243 = n31242 ^ n31219;
  assign n31244 = n31220 & n31243;
  assign n31245 = n31244 ^ n27923;
  assign n31246 = n31245 ^ n31217;
  assign n31247 = n31218 & ~n31246;
  assign n31248 = n31247 ^ n27917;
  assign n31249 = n31248 ^ n31215;
  assign n31250 = n31216 & ~n31249;
  assign n31251 = n31250 ^ n27915;
  assign n31252 = n31251 ^ n31213;
  assign n31253 = ~n31214 & ~n31252;
  assign n31254 = n31253 ^ n27909;
  assign n31255 = n31254 ^ n31211;
  assign n31256 = ~n31212 & n31255;
  assign n31257 = n31256 ^ n28290;
  assign n31258 = n31257 ^ n31209;
  assign n31259 = n31210 & n31258;
  assign n31260 = n31259 ^ n27902;
  assign n31261 = n31260 ^ n31207;
  assign n31262 = ~n31208 & ~n31261;
  assign n31263 = n31262 ^ n27893;
  assign n31264 = n31263 ^ n31205;
  assign n31265 = ~n31206 & n31264;
  assign n31266 = n31265 ^ n27886;
  assign n31267 = n31266 ^ n31203;
  assign n31268 = ~n31204 & n31267;
  assign n31269 = n31268 ^ n28308;
  assign n31270 = n31269 ^ n31201;
  assign n31271 = n31202 & ~n31270;
  assign n31272 = n31271 ^ n27879;
  assign n31273 = n31272 ^ n31199;
  assign n31274 = n31200 & n31273;
  assign n31275 = n31274 ^ n27872;
  assign n31276 = n31275 ^ n31197;
  assign n31277 = n31198 & n31276;
  assign n31278 = n31277 ^ n27864;
  assign n31279 = n31278 ^ n31195;
  assign n31280 = ~n31196 & ~n31279;
  assign n31281 = n31280 ^ n27856;
  assign n31174 = n31173 ^ n30601;
  assign n31175 = n30608 & n31174;
  assign n31176 = n31175 ^ n30607;
  assign n30595 = n29741 ^ n29224;
  assign n30597 = n30596 ^ n29741;
  assign n30598 = ~n30595 & n30597;
  assign n30599 = n30598 ^ n29224;
  assign n30590 = n30559 ^ n30460;
  assign n30591 = ~n30462 & ~n30590;
  assign n30592 = n30591 ^ n3347;
  assign n30593 = n30592 ^ n1338;
  assign n30594 = n30593 ^ n30458;
  assign n30600 = n30599 ^ n30594;
  assign n31193 = n31176 ^ n30600;
  assign n31194 = n31193 ^ n27848;
  assign n31334 = n31281 ^ n31194;
  assign n31303 = n31275 ^ n31198;
  assign n31304 = n31272 ^ n31200;
  assign n31305 = n31254 ^ n31212;
  assign n31306 = n31248 ^ n31216;
  assign n31307 = n31245 ^ n31218;
  assign n31308 = n31233 ^ n31226;
  assign n31309 = n31236 ^ n31224;
  assign n31310 = n31308 & n31309;
  assign n31311 = n31239 ^ n31222;
  assign n31312 = n31310 & n31311;
  assign n31313 = n31242 ^ n31220;
  assign n31314 = ~n31312 & ~n31313;
  assign n31315 = ~n31307 & ~n31314;
  assign n31316 = ~n31306 & n31315;
  assign n31317 = n31251 ^ n31214;
  assign n31318 = ~n31316 & ~n31317;
  assign n31319 = n31305 & n31318;
  assign n31320 = n31257 ^ n31210;
  assign n31321 = ~n31319 & n31320;
  assign n31322 = n31260 ^ n31208;
  assign n31323 = n31321 & n31322;
  assign n31324 = n31263 ^ n31206;
  assign n31325 = n31323 & ~n31324;
  assign n31326 = n31266 ^ n31204;
  assign n31327 = n31325 & ~n31326;
  assign n31328 = n31269 ^ n31202;
  assign n31329 = ~n31327 & ~n31328;
  assign n31330 = n31304 & ~n31329;
  assign n31331 = ~n31303 & n31330;
  assign n31332 = n31278 ^ n31196;
  assign n31333 = n31331 & ~n31332;
  assign n31352 = n31334 ^ n31333;
  assign n3042 = n3041 ^ n3035;
  assign n3046 = n3045 ^ n3042;
  assign n3047 = n3046 ^ n2502;
  assign n31353 = n31352 ^ n3047;
  assign n31354 = n31332 ^ n31331;
  assign n2439 = n2438 ^ n2429;
  assign n2449 = n2448 ^ n2439;
  assign n2453 = n2452 ^ n2449;
  assign n31355 = n31354 ^ n2453;
  assign n31359 = n31330 ^ n31303;
  assign n31356 = n29418 ^ n1484;
  assign n31357 = n31356 ^ n1388;
  assign n31358 = n31357 ^ n2443;
  assign n31360 = n31359 ^ n31358;
  assign n31362 = n29424 ^ n1466;
  assign n31363 = n31362 ^ n25835;
  assign n31364 = n31363 ^ n1383;
  assign n31361 = n31329 ^ n31304;
  assign n31365 = n31364 ^ n31361;
  assign n31366 = n31328 ^ n31327;
  assign n1179 = n1178 ^ n1100;
  assign n1189 = n1188 ^ n1179;
  assign n1193 = n1192 ^ n1189;
  assign n31367 = n31366 ^ n1193;
  assign n31369 = n29095 ^ n1448;
  assign n31370 = n31369 ^ n1033;
  assign n31371 = n31370 ^ n1183;
  assign n31368 = n31326 ^ n31325;
  assign n31372 = n31371 ^ n31368;
  assign n31373 = n31324 ^ n31323;
  assign n1015 = n1008 ^ n942;
  assign n1022 = n1021 ^ n1015;
  assign n1026 = n1025 ^ n1022;
  assign n31374 = n31373 ^ n1026;
  assign n31375 = n31322 ^ n31321;
  assign n31376 = n31375 ^ n913;
  assign n31377 = n31320 ^ n31319;
  assign n881 = n868 ^ n832;
  assign n894 = n893 ^ n881;
  assign n898 = n897 ^ n894;
  assign n31378 = n31377 ^ n898;
  assign n31379 = n31318 ^ n31305;
  assign n31380 = n31379 ^ n3305;
  assign n31381 = n31317 ^ n31316;
  assign n31385 = n31384 ^ n31381;
  assign n31386 = n31315 ^ n31306;
  assign n31390 = n31389 ^ n31386;
  assign n31392 = n29031 ^ n22158;
  assign n31393 = n31392 ^ n25791;
  assign n31394 = n31393 ^ n711;
  assign n31391 = n31314 ^ n31307;
  assign n31395 = n31394 ^ n31391;
  assign n31399 = n31313 ^ n31312;
  assign n31396 = n29035 ^ n22128;
  assign n31397 = n31396 ^ n702;
  assign n31398 = n31397 ^ n20845;
  assign n31400 = n31399 ^ n31398;
  assign n31402 = n29039 ^ n22133;
  assign n31403 = n31402 ^ n25763;
  assign n31404 = n31403 ^ n536;
  assign n31401 = n31311 ^ n31310;
  assign n31405 = n31404 ^ n31401;
  assign n31407 = n28809 ^ n693;
  assign n31408 = n31407 ^ n25768;
  assign n31409 = n31408 ^ n20851;
  assign n31406 = n31309 ^ n31308;
  assign n31410 = n31409 ^ n31406;
  assign n31412 = n2246 & ~n31411;
  assign n2252 = n2210 ^ n2158;
  assign n2253 = n2252 ^ n2242;
  assign n2254 = n2253 ^ n2251;
  assign n31413 = n31412 ^ n2254;
  assign n31414 = n31230 ^ n31229;
  assign n31415 = n31414 ^ n2254;
  assign n31416 = n31413 & ~n31415;
  assign n31417 = n31416 ^ n31412;
  assign n31418 = n31417 ^ n31308;
  assign n31419 = n22140 ^ n2324;
  assign n31420 = n31419 ^ n25773;
  assign n31421 = n31420 ^ n20856;
  assign n31422 = n31421 ^ n31417;
  assign n31423 = n31418 & ~n31422;
  assign n31424 = n31423 ^ n31308;
  assign n31425 = n31424 ^ n31406;
  assign n31426 = ~n31410 & n31425;
  assign n31427 = n31426 ^ n31409;
  assign n31428 = n31427 ^ n31401;
  assign n31429 = ~n31405 & n31428;
  assign n31430 = n31429 ^ n31404;
  assign n31431 = n31430 ^ n31399;
  assign n31432 = n31400 & ~n31431;
  assign n31433 = n31432 ^ n31398;
  assign n31434 = n31433 ^ n31391;
  assign n31435 = ~n31395 & n31434;
  assign n31436 = n31435 ^ n31394;
  assign n31437 = n31436 ^ n31386;
  assign n31438 = n31390 & ~n31437;
  assign n31439 = n31438 ^ n31389;
  assign n31440 = n31439 ^ n31381;
  assign n31441 = n31385 & ~n31440;
  assign n31442 = n31441 ^ n31384;
  assign n31443 = n31442 ^ n31379;
  assign n31444 = n31380 & ~n31443;
  assign n31445 = n31444 ^ n3305;
  assign n31446 = n31445 ^ n31377;
  assign n31447 = n31378 & ~n31446;
  assign n31448 = n31447 ^ n898;
  assign n31449 = n31448 ^ n31375;
  assign n31450 = ~n31376 & n31449;
  assign n31451 = n31450 ^ n913;
  assign n31452 = n31451 ^ n31373;
  assign n31453 = n31374 & ~n31452;
  assign n31454 = n31453 ^ n1026;
  assign n31455 = n31454 ^ n31368;
  assign n31456 = n31372 & ~n31455;
  assign n31457 = n31456 ^ n31371;
  assign n31458 = n31457 ^ n31366;
  assign n31459 = n31367 & ~n31458;
  assign n31460 = n31459 ^ n1193;
  assign n31461 = n31460 ^ n31361;
  assign n31462 = n31365 & ~n31461;
  assign n31463 = n31462 ^ n31364;
  assign n31464 = n31463 ^ n31359;
  assign n31465 = n31360 & ~n31464;
  assign n31466 = n31465 ^ n31358;
  assign n31467 = n31466 ^ n2453;
  assign n31468 = n31355 & ~n31467;
  assign n31469 = n31468 ^ n31354;
  assign n31470 = n31469 ^ n31352;
  assign n31471 = n31353 & ~n31470;
  assign n31472 = n31471 ^ n3047;
  assign n31348 = n29410 ^ n3197;
  assign n31349 = n31348 ^ n2504;
  assign n31350 = n31349 ^ n3062;
  assign n31282 = n31281 ^ n31193;
  assign n31283 = ~n31194 & ~n31282;
  assign n31284 = n31283 ^ n27848;
  assign n31177 = n31176 ^ n30594;
  assign n31178 = n30600 & ~n31177;
  assign n31179 = n31178 ^ n30599;
  assign n30584 = n29735 ^ n29307;
  assign n30586 = n30585 ^ n29735;
  assign n30587 = ~n30584 & n30586;
  assign n30588 = n30587 ^ n29307;
  assign n30583 = n30582 ^ n30564;
  assign n30589 = n30588 ^ n30583;
  assign n31191 = n31179 ^ n30589;
  assign n31192 = n31191 ^ n28338;
  assign n31336 = n31284 ^ n31192;
  assign n31335 = ~n31333 & ~n31334;
  assign n31347 = n31336 ^ n31335;
  assign n31351 = n31350 ^ n31347;
  assign n31527 = n31472 ^ n31351;
  assign n31528 = n30960 ^ n29709;
  assign n31529 = n31054 ^ n31047;
  assign n31530 = n31529 ^ n30960;
  assign n31531 = n31528 & ~n31530;
  assign n31532 = n31531 ^ n29709;
  assign n31533 = n31527 & ~n31532;
  assign n31541 = n31445 ^ n31378;
  assign n31537 = n30604 ^ n29884;
  assign n31187 = n30983 ^ n30980;
  assign n31538 = n31187 ^ n30604;
  assign n31539 = n31537 & n31538;
  assign n31540 = n31539 ^ n29884;
  assign n31542 = n31541 ^ n31540;
  assign n31544 = n30616 ^ n29875;
  assign n31545 = n30616 ^ n30583;
  assign n31546 = n31544 & n31545;
  assign n31547 = n31546 ^ n29875;
  assign n31543 = n31442 ^ n31380;
  assign n31548 = n31547 ^ n31543;
  assign n31550 = n30623 ^ n29751;
  assign n31551 = n30623 ^ n30594;
  assign n31552 = ~n31550 & ~n31551;
  assign n31553 = n31552 ^ n29751;
  assign n31549 = n31439 ^ n31385;
  assign n31554 = n31553 ^ n31549;
  assign n31556 = n30634 ^ n29756;
  assign n31557 = n30634 ^ n30601;
  assign n31558 = ~n31556 & n31557;
  assign n31559 = n31558 ^ n29756;
  assign n31555 = n31436 ^ n31390;
  assign n31560 = n31559 ^ n31555;
  assign n31562 = n30641 ^ n29762;
  assign n31563 = n30641 ^ n30614;
  assign n31564 = ~n31562 & n31563;
  assign n31565 = n31564 ^ n29762;
  assign n31561 = n31433 ^ n31395;
  assign n31566 = n31565 ^ n31561;
  assign n31568 = n30647 ^ n29097;
  assign n31569 = n30647 ^ n30621;
  assign n31570 = n31568 & ~n31569;
  assign n31571 = n31570 ^ n29097;
  assign n31567 = n31430 ^ n31400;
  assign n31572 = n31571 ^ n31567;
  assign n31574 = n30656 ^ n29103;
  assign n31575 = n30656 ^ n30632;
  assign n31576 = ~n31574 & ~n31575;
  assign n31577 = n31576 ^ n29103;
  assign n31573 = n31427 ^ n31405;
  assign n31578 = n31577 ^ n31573;
  assign n31583 = n31424 ^ n31410;
  assign n31579 = n30662 ^ n29683;
  assign n31580 = n30662 ^ n30639;
  assign n31581 = n31579 & n31580;
  assign n31582 = n31581 ^ n29683;
  assign n31584 = n31583 ^ n31582;
  assign n31587 = n30573 ^ n29690;
  assign n31588 = n30651 ^ n30573;
  assign n31589 = ~n31587 & ~n31588;
  assign n31590 = n31589 ^ n29690;
  assign n31585 = n31421 ^ n31308;
  assign n31586 = n31585 ^ n31417;
  assign n31591 = n31590 ^ n31586;
  assign n31596 = n31414 ^ n31413;
  assign n31592 = n30427 ^ n29787;
  assign n31593 = n30653 ^ n30427;
  assign n31594 = n31592 & ~n31593;
  assign n31595 = n31594 ^ n29787;
  assign n31597 = n31596 ^ n31595;
  assign n31598 = n30351 ^ n29699;
  assign n31599 = n30666 ^ n30351;
  assign n31600 = ~n31598 & ~n31599;
  assign n31601 = n31600 ^ n29699;
  assign n31603 = n31602 ^ n31601;
  assign n31613 = n30986 & n31013;
  assign n31614 = n31036 & ~n31613;
  assign n31636 = n31614 ^ n30989;
  assign n31637 = ~n30990 & ~n31636;
  assign n31638 = n31637 ^ n2665;
  assign n31639 = n31638 ^ n31038;
  assign n31632 = n29504 ^ n28757;
  assign n31633 = n30960 ^ n29504;
  assign n31634 = n31632 & n31633;
  assign n31635 = n31634 ^ n28757;
  assign n31640 = n31639 ^ n31635;
  assign n31642 = n29510 ^ n28727;
  assign n31643 = n30914 ^ n29510;
  assign n31644 = ~n31642 & ~n31643;
  assign n31645 = n31644 ^ n28727;
  assign n31641 = n31614 ^ n30990;
  assign n31646 = n31645 ^ n31641;
  assign n31654 = n29709 ^ n29577;
  assign n31655 = n30819 ^ n29709;
  assign n31656 = n31654 & ~n31655;
  assign n31657 = n31656 ^ n29577;
  assign n31647 = n30986 & n31009;
  assign n31648 = n31031 & ~n31647;
  assign n31649 = n31648 ^ n30997;
  assign n31650 = n31026 & n31649;
  assign n31651 = n31650 ^ n30996;
  assign n31652 = n31651 ^ n3189;
  assign n31653 = n31652 ^ n31010;
  assign n31658 = n31657 ^ n31653;
  assign n31660 = n29919 ^ n29532;
  assign n31661 = n30699 ^ n29919;
  assign n31662 = ~n31660 & n31661;
  assign n31663 = n31662 ^ n29532;
  assign n31659 = n31648 ^ n31026;
  assign n31664 = n31663 ^ n31659;
  assign n31492 = n29712 ^ n29480;
  assign n31493 = n30705 ^ n29712;
  assign n31494 = ~n31492 & n31493;
  assign n31495 = n31494 ^ n29480;
  assign n31488 = n31002 ^ n30986;
  assign n31489 = n31028 & ~n31488;
  assign n31490 = n31489 ^ n31001;
  assign n31491 = n31490 ^ n31027;
  assign n31496 = n31495 ^ n31491;
  assign n31295 = n29719 ^ n29360;
  assign n31296 = n30706 ^ n29719;
  assign n31297 = ~n31295 & n31296;
  assign n31298 = n31297 ^ n29360;
  assign n31294 = n31028 ^ n30986;
  assign n31299 = n31298 ^ n31294;
  assign n31183 = n29729 ^ n29314;
  assign n31184 = n30712 ^ n29729;
  assign n31185 = ~n31183 & n31184;
  assign n31186 = n31185 ^ n29314;
  assign n31188 = n31187 ^ n31186;
  assign n31180 = n31179 ^ n30583;
  assign n31181 = n30589 & ~n31180;
  assign n31182 = n31181 ^ n30588;
  assign n31291 = n31187 ^ n31182;
  assign n31292 = ~n31188 & ~n31291;
  assign n31293 = n31292 ^ n31186;
  assign n31485 = n31294 ^ n31293;
  assign n31486 = ~n31299 & n31485;
  assign n31487 = n31486 ^ n31298;
  assign n31665 = n31491 ^ n31487;
  assign n31666 = ~n31496 & n31665;
  assign n31667 = n31666 ^ n31495;
  assign n31668 = n31667 ^ n31659;
  assign n31669 = n31664 & ~n31668;
  assign n31670 = n31669 ^ n31663;
  assign n31671 = n31670 ^ n31653;
  assign n31672 = n31658 & ~n31671;
  assign n31673 = n31672 ^ n31657;
  assign n31674 = n31673 ^ n31641;
  assign n31675 = ~n31646 & n31674;
  assign n31676 = n31675 ^ n31645;
  assign n31677 = n31676 ^ n31639;
  assign n31678 = n31640 & n31677;
  assign n31679 = n31678 ^ n31635;
  assign n31615 = n30993 & ~n31614;
  assign n31616 = n31040 & ~n31615;
  assign n31629 = n31616 ^ n2760;
  assign n31630 = n31629 ^ n31017;
  assign n31625 = n29498 ^ n28799;
  assign n31626 = n30288 ^ n29498;
  assign n31627 = ~n31625 & ~n31626;
  assign n31628 = n31627 ^ n28799;
  assign n31631 = n31630 ^ n31628;
  assign n31700 = n31679 ^ n31631;
  assign n31701 = n31700 ^ n28220;
  assign n31702 = n31676 ^ n31640;
  assign n31703 = n31702 ^ n28233;
  assign n31704 = n31673 ^ n31646;
  assign n31705 = n31704 ^ n28226;
  assign n31706 = n31670 ^ n31658;
  assign n31707 = n31706 ^ n28864;
  assign n31708 = n31667 ^ n31664;
  assign n31709 = n31708 ^ n28850;
  assign n31497 = n31496 ^ n31487;
  assign n31498 = n31497 ^ n28789;
  assign n31300 = n31299 ^ n31293;
  assign n31301 = n31300 ^ n28750;
  assign n31189 = n31188 ^ n31182;
  assign n31190 = n31189 ^ n28484;
  assign n31285 = n31284 ^ n31191;
  assign n31286 = n31192 & n31285;
  assign n31287 = n31286 ^ n28338;
  assign n31288 = n31287 ^ n31189;
  assign n31289 = ~n31190 & n31288;
  assign n31290 = n31289 ^ n28484;
  assign n31482 = n31300 ^ n31290;
  assign n31483 = n31301 & ~n31482;
  assign n31484 = n31483 ^ n28750;
  assign n31710 = n31497 ^ n31484;
  assign n31711 = n31498 & ~n31710;
  assign n31712 = n31711 ^ n28789;
  assign n31713 = n31712 ^ n31708;
  assign n31714 = n31709 & n31713;
  assign n31715 = n31714 ^ n28850;
  assign n31716 = n31715 ^ n31706;
  assign n31717 = ~n31707 & ~n31716;
  assign n31718 = n31717 ^ n28864;
  assign n31719 = n31718 ^ n31704;
  assign n31720 = ~n31705 & ~n31719;
  assign n31721 = n31720 ^ n28226;
  assign n31722 = n31721 ^ n31702;
  assign n31723 = ~n31703 & ~n31722;
  assign n31724 = n31723 ^ n28233;
  assign n31725 = n31724 ^ n31700;
  assign n31726 = n31701 & ~n31725;
  assign n31727 = n31726 ^ n28220;
  assign n31680 = n31679 ^ n31630;
  assign n31681 = n31631 & n31680;
  assign n31682 = n31681 ^ n31628;
  assign n31620 = n29544 ^ n28900;
  assign n31621 = n30291 ^ n29544;
  assign n31622 = n31620 & n31621;
  assign n31623 = n31622 ^ n28900;
  assign n31617 = n31019 & ~n31616;
  assign n31618 = n31617 ^ n31018;
  assign n31619 = n31618 ^ n31024;
  assign n31624 = n31623 ^ n31619;
  assign n31698 = n31682 ^ n31624;
  assign n31699 = n31698 ^ n28213;
  assign n31735 = n31727 ^ n31699;
  assign n31736 = n31712 ^ n31709;
  assign n31499 = n31498 ^ n31484;
  assign n31302 = n31301 ^ n31290;
  assign n31337 = ~n31335 & n31336;
  assign n31338 = n31287 ^ n31190;
  assign n31339 = n31337 & n31338;
  assign n31500 = n31302 & ~n31339;
  assign n31737 = n31499 & n31500;
  assign n31738 = n31736 & n31737;
  assign n31739 = n31715 ^ n31707;
  assign n31740 = ~n31738 & ~n31739;
  assign n31741 = n31718 ^ n31705;
  assign n31742 = n31740 & n31741;
  assign n31743 = n31721 ^ n31703;
  assign n31744 = n31742 & ~n31743;
  assign n31745 = n31724 ^ n31701;
  assign n31746 = n31744 & ~n31745;
  assign n31747 = ~n31735 & ~n31746;
  assign n31728 = n31727 ^ n31698;
  assign n31729 = ~n31699 & ~n31728;
  assign n31730 = n31729 ^ n28213;
  assign n31683 = n31682 ^ n31619;
  assign n31684 = ~n31624 & n31683;
  assign n31685 = n31684 ^ n31623;
  assign n31608 = n29595 ^ n28894;
  assign n31609 = n30296 ^ n29595;
  assign n31610 = n31608 & ~n31609;
  assign n31611 = n31610 ^ n28894;
  assign n31612 = n31611 ^ n31529;
  assign n31696 = n31685 ^ n31612;
  assign n31697 = n31696 ^ n28207;
  assign n31748 = n31730 ^ n31697;
  assign n31749 = n31747 & n31748;
  assign n31731 = n31730 ^ n31696;
  assign n31732 = ~n31697 & n31731;
  assign n31733 = n31732 ^ n28207;
  assign n31689 = n29612 ^ n28844;
  assign n31690 = n30300 ^ n29612;
  assign n31691 = ~n31689 & n31690;
  assign n31692 = n31691 ^ n28844;
  assign n31519 = n31053 ^ n31047;
  assign n31520 = n31054 & n31519;
  assign n31521 = n31520 ^ n2885;
  assign n31522 = n31521 ^ n31074;
  assign n31693 = n31692 ^ n31522;
  assign n31686 = n31685 ^ n31529;
  assign n31687 = ~n31612 & ~n31686;
  assign n31688 = n31687 ^ n31611;
  assign n31694 = n31693 ^ n31688;
  assign n31695 = n31694 ^ n28246;
  assign n31734 = n31733 ^ n31695;
  assign n31768 = n31749 ^ n31734;
  assign n31769 = n31768 ^ n2083;
  assign n31770 = n31748 ^ n31747;
  assign n31774 = n31773 ^ n31770;
  assign n31775 = n31746 ^ n31735;
  assign n31779 = n31778 ^ n31775;
  assign n31780 = n31745 ^ n31744;
  assign n31784 = n31783 ^ n31780;
  assign n31785 = n31743 ^ n31742;
  assign n31789 = n31788 ^ n31785;
  assign n31790 = n31741 ^ n31740;
  assign n31791 = n31790 ^ n1613;
  assign n31792 = n31739 ^ n31738;
  assign n2960 = n2953 ^ n2890;
  assign n2961 = n2960 ^ n2868;
  assign n2962 = n2961 ^ n1508;
  assign n31793 = n31792 ^ n2962;
  assign n31794 = n31737 ^ n31736;
  assign n2856 = n2795 ^ n1529;
  assign n2857 = n2856 ^ n2853;
  assign n2861 = n2860 ^ n2857;
  assign n31795 = n31794 ^ n2861;
  assign n31501 = n31500 ^ n31499;
  assign n31502 = n31501 ^ n2846;
  assign n31340 = n31339 ^ n31302;
  assign n3218 = n3211 ^ n2721;
  assign n3222 = n3221 ^ n3218;
  assign n3223 = n3222 ^ n2840;
  assign n31341 = n31340 ^ n3223;
  assign n31342 = n31338 ^ n31337;
  assign n31346 = n31345 ^ n31342;
  assign n31473 = n31472 ^ n31347;
  assign n31474 = n31351 & ~n31473;
  assign n31475 = n31474 ^ n31350;
  assign n31476 = n31475 ^ n31342;
  assign n31477 = ~n31346 & n31476;
  assign n31478 = n31477 ^ n31345;
  assign n31479 = n31478 ^ n31340;
  assign n31480 = ~n31341 & n31479;
  assign n31481 = n31480 ^ n3223;
  assign n31796 = n31501 ^ n31481;
  assign n31797 = n31502 & ~n31796;
  assign n31798 = n31797 ^ n2846;
  assign n31799 = n31798 ^ n31794;
  assign n31800 = n31795 & ~n31799;
  assign n31801 = n31800 ^ n2861;
  assign n31802 = n31801 ^ n31792;
  assign n31803 = ~n31793 & n31802;
  assign n31804 = n31803 ^ n2962;
  assign n31805 = n31804 ^ n31790;
  assign n31806 = ~n31791 & n31805;
  assign n31807 = n31806 ^ n1613;
  assign n31808 = n31807 ^ n31785;
  assign n31809 = n31789 & ~n31808;
  assign n31810 = n31809 ^ n31788;
  assign n31811 = n31810 ^ n31780;
  assign n31812 = n31784 & ~n31811;
  assign n31813 = n31812 ^ n31783;
  assign n31814 = n31813 ^ n31775;
  assign n31815 = n31779 & ~n31814;
  assign n31816 = n31815 ^ n31778;
  assign n31817 = n31816 ^ n31770;
  assign n31818 = n31774 & ~n31817;
  assign n31819 = n31818 ^ n31773;
  assign n31820 = n31819 ^ n31768;
  assign n31821 = n31769 & ~n31820;
  assign n31822 = n31821 ^ n2083;
  assign n31761 = n31733 ^ n28246;
  assign n31762 = n31733 ^ n31694;
  assign n31763 = ~n31761 & ~n31762;
  assign n31764 = n31763 ^ n28246;
  assign n31756 = n31688 ^ n31522;
  assign n31757 = ~n31693 & ~n31756;
  assign n31758 = n31757 ^ n31692;
  assign n31751 = n29632 ^ n28838;
  assign n31752 = n30270 ^ n29632;
  assign n31753 = n31751 & n31752;
  assign n31754 = n31753 ^ n28838;
  assign n31511 = n31115 ^ n31065;
  assign n31512 = n31511 ^ n31066;
  assign n31755 = n31754 ^ n31512;
  assign n31759 = n31758 ^ n31755;
  assign n31760 = n31759 ^ n27955;
  assign n31765 = n31764 ^ n31760;
  assign n31750 = n31734 & n31749;
  assign n31766 = n31765 ^ n31750;
  assign n31767 = n31766 ^ n2099;
  assign n31823 = n31822 ^ n31767;
  assign n31604 = n29794 ^ n29680;
  assign n31605 = n30672 ^ n29680;
  assign n31606 = ~n31604 & ~n31605;
  assign n31607 = n31606 ^ n29794;
  assign n31824 = n31823 ^ n31607;
  assign n31826 = n29804 ^ n29687;
  assign n31827 = n30678 ^ n29687;
  assign n31828 = ~n31826 & n31827;
  assign n31829 = n31828 ^ n29804;
  assign n31825 = n31819 ^ n31769;
  assign n31830 = n31829 ^ n31825;
  assign n31835 = n31816 ^ n31774;
  assign n31831 = n29810 ^ n29695;
  assign n31832 = n30685 ^ n29695;
  assign n31833 = ~n31831 & ~n31832;
  assign n31834 = n31833 ^ n29810;
  assign n31836 = n31835 ^ n31834;
  assign n31841 = n31813 ^ n31779;
  assign n31837 = n30338 ^ n29817;
  assign n31838 = n30687 ^ n30338;
  assign n31839 = n31837 & n31838;
  assign n31840 = n31839 ^ n29817;
  assign n31842 = n31841 ^ n31840;
  assign n31843 = n29703 ^ n28811;
  assign n31844 = n30693 ^ n29703;
  assign n31845 = n31843 & n31844;
  assign n31846 = n31845 ^ n28811;
  assign n31847 = n31810 ^ n31784;
  assign n31848 = ~n31846 & n31847;
  assign n31849 = n31848 ^ n31841;
  assign n31850 = n31842 & n31849;
  assign n31851 = n31850 ^ n31848;
  assign n31852 = n31851 ^ n31835;
  assign n31853 = n31836 & ~n31852;
  assign n31854 = n31853 ^ n31834;
  assign n31855 = n31854 ^ n31825;
  assign n31856 = ~n31830 & ~n31855;
  assign n31857 = n31856 ^ n31829;
  assign n31858 = n31857 ^ n31823;
  assign n31859 = ~n31824 & ~n31858;
  assign n31860 = n31859 ^ n31607;
  assign n31861 = n31860 ^ n31602;
  assign n31862 = n31603 & n31861;
  assign n31863 = n31862 ^ n31601;
  assign n31864 = n31863 ^ n31596;
  assign n31865 = n31597 & n31864;
  assign n31866 = n31865 ^ n31595;
  assign n31867 = n31866 ^ n31586;
  assign n31868 = ~n31591 & ~n31867;
  assign n31869 = n31868 ^ n31590;
  assign n31870 = n31869 ^ n31583;
  assign n31871 = ~n31584 & ~n31870;
  assign n31872 = n31871 ^ n31582;
  assign n31873 = n31872 ^ n31573;
  assign n31874 = n31578 & n31873;
  assign n31875 = n31874 ^ n31577;
  assign n31876 = n31875 ^ n31567;
  assign n31877 = n31572 & n31876;
  assign n31878 = n31877 ^ n31571;
  assign n31879 = n31878 ^ n31561;
  assign n31880 = ~n31566 & n31879;
  assign n31881 = n31880 ^ n31565;
  assign n31882 = n31881 ^ n31555;
  assign n31883 = n31560 & ~n31882;
  assign n31884 = n31883 ^ n31559;
  assign n31885 = n31884 ^ n31549;
  assign n31886 = ~n31554 & ~n31885;
  assign n31887 = n31886 ^ n31553;
  assign n31888 = n31887 ^ n31543;
  assign n31889 = ~n31548 & n31888;
  assign n31890 = n31889 ^ n31547;
  assign n31891 = n31890 ^ n31541;
  assign n31892 = ~n31542 & n31891;
  assign n31893 = n31892 ^ n31540;
  assign n31894 = n30712 ^ n29741;
  assign n31895 = n31659 ^ n30712;
  assign n31896 = n31894 & ~n31895;
  assign n31897 = n31896 ^ n29741;
  assign n31898 = n31454 ^ n31372;
  assign n31899 = n31897 & ~n31898;
  assign n31900 = n30585 ^ n29743;
  assign n31901 = n31491 ^ n30585;
  assign n31902 = n31900 & ~n31901;
  assign n31903 = n31902 ^ n29743;
  assign n31904 = n31451 ^ n31374;
  assign n31905 = ~n31903 & ~n31904;
  assign n31907 = n30596 ^ n29745;
  assign n31908 = n31294 ^ n30596;
  assign n31909 = ~n31907 & ~n31908;
  assign n31910 = n31909 ^ n29745;
  assign n31906 = n31448 ^ n31376;
  assign n31912 = n31910 ^ n31906;
  assign n31911 = ~n31906 & ~n31910;
  assign n31913 = n31912 ^ n31911;
  assign n31914 = ~n31905 & n31913;
  assign n31915 = n30706 ^ n29735;
  assign n31916 = n31653 ^ n30706;
  assign n31917 = n31915 & ~n31916;
  assign n31918 = n31917 ^ n29735;
  assign n31919 = n31457 ^ n31367;
  assign n31920 = n31918 & ~n31919;
  assign n31921 = n31914 & ~n31920;
  assign n31922 = ~n31899 & n31921;
  assign n31927 = n31460 ^ n31365;
  assign n31923 = n30705 ^ n29729;
  assign n31924 = n31641 ^ n30705;
  assign n31925 = ~n31923 & n31924;
  assign n31926 = n31925 ^ n29729;
  assign n31929 = n31927 ^ n31926;
  assign n31928 = n31926 & n31927;
  assign n31930 = n31929 ^ n31928;
  assign n31931 = n30699 ^ n29719;
  assign n31932 = n31639 ^ n30699;
  assign n31933 = ~n31931 & n31932;
  assign n31934 = n31933 ^ n29719;
  assign n31935 = n31463 ^ n31360;
  assign n31936 = ~n31934 & ~n31935;
  assign n31937 = n30914 ^ n29919;
  assign n31938 = n31619 ^ n30914;
  assign n31939 = n31937 & ~n31938;
  assign n31940 = n31939 ^ n29919;
  assign n31941 = n31469 ^ n31353;
  assign n31942 = ~n31940 & ~n31941;
  assign n31943 = ~n31936 & ~n31942;
  assign n31944 = n31930 & n31943;
  assign n31945 = n31466 ^ n31355;
  assign n31946 = n30819 ^ n29712;
  assign n31947 = n31630 ^ n30819;
  assign n31948 = ~n31946 & ~n31947;
  assign n31949 = n31948 ^ n29712;
  assign n31951 = n31945 & n31949;
  assign n31950 = n31949 ^ n31945;
  assign n31952 = n31951 ^ n31950;
  assign n31953 = n31944 & n31952;
  assign n31954 = n31922 & n31953;
  assign n31955 = ~n31893 & n31954;
  assign n31956 = n31919 ^ n31918;
  assign n31957 = n31898 ^ n31897;
  assign n31958 = n31904 ^ n31903;
  assign n31959 = n31911 ^ n31903;
  assign n31960 = ~n31958 & n31959;
  assign n31961 = n31960 ^ n31911;
  assign n31962 = n31961 ^ n31898;
  assign n31963 = ~n31957 & ~n31962;
  assign n31964 = n31963 ^ n31897;
  assign n31965 = n31964 ^ n31918;
  assign n31966 = ~n31956 & ~n31965;
  assign n31967 = n31966 ^ n31919;
  assign n31968 = n31953 & n31967;
  assign n31969 = n31941 ^ n31940;
  assign n31970 = n31935 ^ n31934;
  assign n31971 = ~n31928 & n31970;
  assign n31972 = n31971 ^ n31936;
  assign n31973 = n31950 & ~n31972;
  assign n31974 = n31973 ^ n31951;
  assign n31975 = n31974 ^ n31941;
  assign n31976 = n31969 & n31975;
  assign n31977 = n31976 ^ n31941;
  assign n31978 = ~n31968 & ~n31977;
  assign n31979 = ~n31955 & n31978;
  assign n31980 = n31532 ^ n31527;
  assign n31981 = n31980 ^ n31533;
  assign n31982 = ~n31979 & ~n31981;
  assign n31992 = ~n31533 & ~n31982;
  assign n31518 = n30288 ^ n29510;
  assign n31523 = n31522 ^ n30288;
  assign n31524 = n31518 & ~n31523;
  assign n31525 = n31524 ^ n29510;
  assign n31517 = n31475 ^ n31346;
  assign n31534 = n31525 ^ n31517;
  assign n31993 = n31992 ^ n31534;
  assign n31994 = n31993 ^ n28727;
  assign n31995 = n31980 ^ n31979;
  assign n31996 = ~n29577 & n31995;
  assign n31997 = n31996 ^ n31993;
  assign n31998 = ~n31994 & ~n31997;
  assign n31999 = n31998 ^ n28727;
  assign n32000 = ~n31893 & n31922;
  assign n32001 = ~n31967 & ~n32000;
  assign n32002 = n31930 & ~n32001;
  assign n32003 = ~n31936 & n32002;
  assign n32004 = n31972 & ~n32003;
  assign n32006 = n32004 ^ n31945;
  assign n32007 = n31950 & n32006;
  assign n32008 = n32007 ^ n31949;
  assign n32009 = n32008 ^ n31969;
  assign n32010 = n32009 ^ n29532;
  assign n32013 = ~n31928 & ~n32002;
  assign n32014 = n32013 ^ n31970;
  assign n32015 = n29360 & n32014;
  assign n32016 = n32001 ^ n31929;
  assign n32018 = n32016 ^ n29314;
  assign n32017 = ~n29314 & ~n32016;
  assign n32019 = n32018 ^ n32017;
  assign n32020 = ~n31893 & n31914;
  assign n32021 = ~n31961 & ~n32020;
  assign n32022 = n32021 ^ n31898;
  assign n32023 = ~n31957 & n32022;
  assign n32024 = n32023 ^ n31897;
  assign n32025 = n32024 ^ n31956;
  assign n32026 = n32025 ^ n29307;
  assign n32027 = n32021 ^ n31957;
  assign n32028 = n32027 ^ n29224;
  assign n32029 = n31906 ^ n31893;
  assign n32030 = n31912 & ~n32029;
  assign n32031 = n32030 ^ n31910;
  assign n32032 = n32031 ^ n31958;
  assign n32034 = n32032 ^ n29111;
  assign n32035 = n31912 ^ n31893;
  assign n32036 = ~n29207 & ~n32035;
  assign n32037 = ~n32034 & ~n32036;
  assign n32033 = ~n29111 & n32032;
  assign n32038 = n32037 ^ n32033;
  assign n32039 = n32038 ^ n32027;
  assign n32040 = n32028 & n32039;
  assign n32041 = n32040 ^ n29224;
  assign n32042 = n32041 ^ n32025;
  assign n32043 = n32026 & ~n32042;
  assign n32044 = n32043 ^ n29307;
  assign n32045 = n31890 ^ n31542;
  assign n32046 = n32045 ^ n29113;
  assign n32047 = n31887 ^ n31548;
  assign n32048 = n32047 ^ n29124;
  assign n32049 = n31884 ^ n31554;
  assign n32050 = n32049 ^ n29126;
  assign n32051 = n31881 ^ n31560;
  assign n32052 = n32051 ^ n28813;
  assign n32053 = n31878 ^ n31566;
  assign n32054 = n32053 ^ n29101;
  assign n32055 = n31875 ^ n31572;
  assign n32056 = n32055 ^ n29178;
  assign n32057 = n31872 ^ n31578;
  assign n32058 = n32057 ^ n29136;
  assign n32059 = n31869 ^ n31584;
  assign n32060 = n32059 ^ n29142;
  assign n32061 = n31866 ^ n31591;
  assign n32062 = n32061 ^ n29148;
  assign n32063 = n31863 ^ n31597;
  assign n32064 = n32063 ^ n29154;
  assign n32065 = n31860 ^ n31603;
  assign n32066 = n32065 ^ n29087;
  assign n32067 = n31857 ^ n31824;
  assign n32068 = n32067 ^ n28986;
  assign n32069 = n31854 ^ n31830;
  assign n32070 = n32069 ^ n28819;
  assign n32071 = n31851 ^ n31836;
  assign n32072 = n32071 ^ n28821;
  assign n32073 = n31847 ^ n31846;
  assign n32074 = n28921 & ~n32073;
  assign n32075 = n32074 ^ n28832;
  assign n32076 = n31848 ^ n31840;
  assign n32077 = n32076 ^ n31841;
  assign n32078 = n32077 ^ n32074;
  assign n32079 = n32075 & n32078;
  assign n32080 = n32079 ^ n28832;
  assign n32081 = n32080 ^ n32071;
  assign n32082 = ~n32072 & ~n32081;
  assign n32083 = n32082 ^ n28821;
  assign n32084 = n32083 ^ n32069;
  assign n32085 = ~n32070 & ~n32084;
  assign n32086 = n32085 ^ n28819;
  assign n32087 = n32086 ^ n32067;
  assign n32088 = ~n32068 & ~n32087;
  assign n32089 = n32088 ^ n28986;
  assign n32090 = n32089 ^ n32065;
  assign n32091 = ~n32066 & n32090;
  assign n32092 = n32091 ^ n29087;
  assign n32093 = n32092 ^ n32063;
  assign n32094 = n32064 & ~n32093;
  assign n32095 = n32094 ^ n29154;
  assign n32096 = n32095 ^ n32061;
  assign n32097 = ~n32062 & ~n32096;
  assign n32098 = n32097 ^ n29148;
  assign n32099 = n32098 ^ n32059;
  assign n32100 = ~n32060 & ~n32099;
  assign n32101 = n32100 ^ n29142;
  assign n32102 = n32101 ^ n32057;
  assign n32103 = n32058 & n32102;
  assign n32104 = n32103 ^ n29136;
  assign n32105 = n32104 ^ n32055;
  assign n32106 = ~n32056 & n32105;
  assign n32107 = n32106 ^ n29178;
  assign n32108 = n32107 ^ n32053;
  assign n32109 = ~n32054 & n32108;
  assign n32110 = n32109 ^ n29101;
  assign n32111 = n32110 ^ n32051;
  assign n32112 = n32052 & ~n32111;
  assign n32113 = n32112 ^ n28813;
  assign n32114 = n32113 ^ n32049;
  assign n32115 = n32050 & n32114;
  assign n32116 = n32115 ^ n29126;
  assign n32117 = n32116 ^ n32047;
  assign n32118 = n32048 & n32117;
  assign n32119 = n32118 ^ n29124;
  assign n32120 = n32119 ^ n32045;
  assign n32121 = n32046 & ~n32120;
  assign n32122 = n32121 ^ n29113;
  assign n32123 = ~n29224 & ~n32027;
  assign n32124 = n32035 ^ n29207;
  assign n32125 = n32124 ^ n32036;
  assign n32126 = ~n32033 & n32125;
  assign n32127 = ~n29307 & ~n32025;
  assign n32128 = n32126 & ~n32127;
  assign n32129 = ~n32123 & n32128;
  assign n32130 = n32122 & n32129;
  assign n32131 = ~n32044 & ~n32130;
  assign n32132 = n32019 & ~n32131;
  assign n32133 = ~n32015 & n32132;
  assign n32134 = n32014 ^ n29360;
  assign n32135 = n32017 ^ n32014;
  assign n32136 = n32134 & n32135;
  assign n32137 = n32136 ^ n29360;
  assign n32005 = n32004 ^ n31950;
  assign n32138 = n32005 ^ n29480;
  assign n32139 = n32137 & n32138;
  assign n32140 = n32139 ^ n32009;
  assign n32141 = n32140 ^ n32009;
  assign n32142 = ~n32133 & n32141;
  assign n32143 = n32142 ^ n32009;
  assign n32144 = ~n32010 & n32143;
  assign n32145 = n32144 ^ n29532;
  assign n32011 = n29480 & ~n32010;
  assign n32012 = n32005 & n32011;
  assign n32146 = n32145 ^ n32012;
  assign n32147 = n31995 ^ n29577;
  assign n32148 = n32147 ^ n31996;
  assign n32149 = ~n32146 & ~n32148;
  assign n32150 = n28727 & ~n31993;
  assign n32151 = n32149 & ~n32150;
  assign n32152 = n31999 & ~n32151;
  assign n31535 = ~n31533 & ~n31534;
  assign n31526 = n31517 & ~n31525;
  assign n31536 = n31535 ^ n31526;
  assign n31983 = ~n31526 & n31982;
  assign n31984 = n31536 & ~n31983;
  assign n31510 = n30291 ^ n29504;
  assign n31513 = n31512 ^ n30291;
  assign n31514 = n31510 & n31513;
  assign n31515 = n31514 ^ n29504;
  assign n31509 = n31478 ^ n31341;
  assign n31516 = n31515 ^ n31509;
  assign n31990 = n31984 ^ n31516;
  assign n31991 = n31990 ^ n28757;
  assign n32226 = n32152 ^ n31991;
  assign n32157 = ~n31996 & ~n32149;
  assign n32158 = n32157 ^ n31994;
  assign n32159 = n32147 ^ n32146;
  assign n32160 = n32131 ^ n32018;
  assign n32161 = n32122 & n32126;
  assign n32162 = n32038 & ~n32161;
  assign n32163 = n32162 ^ n32027;
  assign n32164 = n32028 & n32163;
  assign n32165 = n32164 ^ n29224;
  assign n32166 = n32165 ^ n32026;
  assign n32167 = n32162 ^ n32028;
  assign n32168 = n32122 ^ n32035;
  assign n32169 = n32124 & n32168;
  assign n32170 = n32169 ^ n29207;
  assign n32171 = n32170 ^ n32034;
  assign n32172 = n32124 ^ n32122;
  assign n32173 = ~n32171 & ~n32172;
  assign n32174 = ~n32167 & ~n32173;
  assign n32175 = ~n32166 & ~n32174;
  assign n32176 = n32160 & n32175;
  assign n32177 = n32119 ^ n32046;
  assign n32178 = n32110 ^ n32052;
  assign n32179 = n32107 ^ n32054;
  assign n32180 = n32101 ^ n32058;
  assign n32181 = n32098 ^ n32060;
  assign n32182 = n32095 ^ n32062;
  assign n32183 = n32089 ^ n32066;
  assign n32184 = n32080 ^ n32072;
  assign n32185 = n32083 ^ n32070;
  assign n32186 = n32184 & ~n32185;
  assign n32187 = n32086 ^ n32068;
  assign n32188 = n32186 & n32187;
  assign n32189 = n32183 & ~n32188;
  assign n32190 = n32092 ^ n32064;
  assign n32191 = ~n32189 & n32190;
  assign n32192 = ~n32182 & n32191;
  assign n32193 = ~n32181 & ~n32192;
  assign n32194 = ~n32180 & n32193;
  assign n32195 = n32104 ^ n32056;
  assign n32196 = ~n32194 & n32195;
  assign n32197 = n32179 & n32196;
  assign n32198 = ~n32178 & n32197;
  assign n32199 = n32113 ^ n32050;
  assign n32200 = n32198 & ~n32199;
  assign n32201 = n32116 ^ n32048;
  assign n32202 = ~n32200 & ~n32201;
  assign n32203 = ~n32177 & ~n32202;
  assign n32204 = n32203 ^ n32167;
  assign n32205 = ~n32133 & n32137;
  assign n32206 = n32205 ^ n32138;
  assign n32207 = ~n32017 & ~n32132;
  assign n32208 = n32207 ^ n32134;
  assign n32209 = n32205 ^ n32005;
  assign n32210 = n32138 & ~n32209;
  assign n32211 = n32210 ^ n29480;
  assign n32212 = n32211 ^ n32010;
  assign n32213 = ~n32208 & n32212;
  assign n32214 = ~n32206 & n32213;
  assign n32215 = n32214 ^ n32167;
  assign n32216 = ~n32167 & ~n32215;
  assign n32217 = n32216 ^ n32167;
  assign n32218 = n32204 & ~n32217;
  assign n32219 = n32218 ^ n32216;
  assign n32220 = n32219 ^ n32167;
  assign n32221 = n32220 ^ n32214;
  assign n32222 = n32176 & ~n32221;
  assign n32223 = n32222 ^ n32214;
  assign n32224 = ~n32159 & ~n32223;
  assign n32225 = ~n32158 & n32224;
  assign n32230 = n32226 ^ n32225;
  assign n32234 = n32233 ^ n32230;
  assign n32236 = n2994 ^ n1642;
  assign n32237 = n32236 ^ n26498;
  assign n32238 = n32237 ^ n21697;
  assign n32235 = n32224 ^ n32158;
  assign n32239 = n32238 ^ n32235;
  assign n32243 = n32223 ^ n32159;
  assign n32244 = n32242 & ~n32243;
  assign n32245 = n32244 ^ n32235;
  assign n32246 = n32239 & ~n32245;
  assign n32247 = n32246 ^ n32238;
  assign n32248 = n32247 ^ n32230;
  assign n32249 = ~n32234 & n32248;
  assign n32250 = n32249 ^ n32233;
  assign n32251 = n32230 & ~n32233;
  assign n32252 = ~n32172 & n32203;
  assign n32253 = ~n32171 & n32252;
  assign n32254 = ~n32167 & ~n32253;
  assign n32255 = ~n32166 & ~n32254;
  assign n32256 = n32160 & n32255;
  assign n32257 = ~n32208 & ~n32256;
  assign n32258 = ~n32206 & n32257;
  assign n32259 = n32258 ^ n32212;
  assign n32263 = n32262 ^ n32259;
  assign n32264 = n32257 ^ n32206;
  assign n32265 = n32264 ^ n3101;
  assign n32266 = n32256 ^ n32208;
  assign n2637 = n2636 ^ n2588;
  assign n2644 = n2643 ^ n2637;
  assign n2645 = n2644 ^ n1565;
  assign n32267 = n32266 ^ n2645;
  assign n3079 = n3074 ^ n3069;
  assign n3080 = n3079 ^ n2572;
  assign n3081 = n3080 ^ n2641;
  assign n32268 = n32255 ^ n32160;
  assign n32269 = n3081 & ~n32268;
  assign n32270 = n32269 ^ n32266;
  assign n32271 = n32267 & ~n32270;
  assign n32272 = n32271 ^ n2645;
  assign n32273 = n32272 ^ n32264;
  assign n32274 = ~n32265 & n32273;
  assign n32275 = n32274 ^ n3101;
  assign n32276 = n32275 ^ n32259;
  assign n32277 = n32263 & n32276;
  assign n32278 = n32277 ^ n32259;
  assign n32391 = n32254 ^ n32166;
  assign n2548 = n2544 ^ n2523;
  assign n2561 = n2560 ^ n2548;
  assign n2565 = n2564 ^ n2561;
  assign n32396 = n32391 ^ n2565;
  assign n32376 = n32253 ^ n32167;
  assign n3156 = n3155 ^ n2465;
  assign n3166 = n3165 ^ n3156;
  assign n3167 = n3166 ^ n2555;
  assign n32397 = n32376 ^ n3167;
  assign n32381 = n32252 ^ n32171;
  assign n32378 = n30220 ^ n2482;
  assign n32379 = n32378 ^ n26511;
  assign n32380 = n32379 ^ n3163;
  assign n32398 = n32381 ^ n32380;
  assign n32383 = n32203 ^ n32172;
  assign n32384 = n3144 ^ n1401;
  assign n32385 = n32384 ^ n26606;
  assign n32386 = n32385 ^ n21352;
  assign n32388 = n32383 & n32386;
  assign n32399 = n32388 ^ n32381;
  assign n32400 = n32398 & ~n32399;
  assign n32401 = n32400 ^ n32380;
  assign n32402 = n32401 ^ n32376;
  assign n32403 = n32397 & ~n32402;
  assign n32404 = n32403 ^ n3167;
  assign n32405 = n32404 ^ n32391;
  assign n32406 = ~n32396 & n32405;
  assign n32407 = n32406 ^ n2565;
  assign n32279 = n32202 ^ n32177;
  assign n1319 = n1300 ^ n1216;
  assign n1320 = n1319 ^ n1316;
  assign n1324 = n1323 ^ n1320;
  assign n32280 = n32279 ^ n1324;
  assign n32281 = n32201 ^ n32200;
  assign n1304 = n1288 ^ n1201;
  assign n1305 = n1304 ^ n1167;
  assign n1309 = n1308 ^ n1305;
  assign n32282 = n32281 ^ n1309;
  assign n32283 = n32199 ^ n32198;
  assign n1152 = n1136 ^ n1115;
  assign n1153 = n1152 ^ n1067;
  assign n1157 = n1156 ^ n1153;
  assign n32284 = n32283 ^ n1157;
  assign n32285 = n32197 ^ n32178;
  assign n32286 = n32285 ^ n1149;
  assign n32287 = n32196 ^ n32179;
  assign n32288 = n32287 ^ n3330;
  assign n32289 = n32195 ^ n32194;
  assign n32293 = n32292 ^ n32289;
  assign n32294 = n32193 ^ n32180;
  assign n32298 = n32297 ^ n32294;
  assign n32302 = n32192 ^ n32181;
  assign n32299 = n30180 ^ n22833;
  assign n32300 = n32299 ^ n26531;
  assign n32301 = n32300 ^ n614;
  assign n32303 = n32302 ^ n32301;
  assign n32304 = n32191 ^ n32182;
  assign n721 = n720 ^ n714;
  assign n722 = n721 ^ n581;
  assign n723 = n722 ^ n650;
  assign n32305 = n32304 ^ n723;
  assign n32309 = n32190 ^ n32189;
  assign n32306 = n29643 ^ n22856;
  assign n32307 = n32306 ^ n26539;
  assign n32308 = n32307 ^ n576;
  assign n32310 = n32309 ^ n32308;
  assign n32314 = n32188 ^ n32183;
  assign n32311 = n29670 ^ n548;
  assign n32312 = n32311 ^ n26544;
  assign n32313 = n32312 ^ n3284;
  assign n32315 = n32314 ^ n32313;
  assign n32316 = n32187 ^ n32186;
  assign n32320 = n32319 ^ n32316;
  assign n32322 = n29660 ^ n22327;
  assign n32323 = n32322 ^ n26556;
  assign n32324 = n32323 ^ n21380;
  assign n32321 = n32185 ^ n32184;
  assign n32325 = n32324 ^ n32321;
  assign n2401 = n2359 ^ n2298;
  assign n2402 = n2401 ^ n2393;
  assign n2406 = n2405 ^ n2402;
  assign n32326 = n32184 ^ n2406;
  assign n2378 = n2377 ^ n2268;
  assign n2379 = n2378 ^ n2191;
  assign n2380 = n2379 ^ n2132;
  assign n32327 = n32073 ^ n28921;
  assign n32328 = n2380 & ~n32327;
  assign n2383 = n2343 ^ n2280;
  assign n2384 = n2383 ^ n2370;
  assign n2388 = n2387 ^ n2384;
  assign n32329 = n32328 ^ n2388;
  assign n32330 = n32077 ^ n32075;
  assign n32331 = n32330 ^ n2388;
  assign n32332 = n32329 & n32331;
  assign n32333 = n32332 ^ n32328;
  assign n32334 = n32333 ^ n32184;
  assign n32335 = n32326 & ~n32334;
  assign n32336 = n32335 ^ n2406;
  assign n32337 = n32336 ^ n32321;
  assign n32338 = n32325 & ~n32337;
  assign n32339 = n32338 ^ n32324;
  assign n32340 = n32339 ^ n32316;
  assign n32341 = ~n32320 & n32340;
  assign n32342 = n32341 ^ n32319;
  assign n32343 = n32342 ^ n32314;
  assign n32344 = ~n32315 & n32343;
  assign n32345 = n32344 ^ n32313;
  assign n32346 = n32345 ^ n32309;
  assign n32347 = n32310 & ~n32346;
  assign n32348 = n32347 ^ n32308;
  assign n32349 = n32348 ^ n32304;
  assign n32350 = n32305 & ~n32349;
  assign n32351 = n32350 ^ n723;
  assign n32352 = n32351 ^ n32302;
  assign n32353 = n32303 & ~n32352;
  assign n32354 = n32353 ^ n32301;
  assign n32355 = n32354 ^ n32294;
  assign n32356 = ~n32298 & n32355;
  assign n32357 = n32356 ^ n32297;
  assign n32358 = n32357 ^ n32289;
  assign n32359 = n32293 & ~n32358;
  assign n32360 = n32359 ^ n32292;
  assign n32361 = n32360 ^ n32287;
  assign n32362 = ~n32288 & n32361;
  assign n32363 = n32362 ^ n3330;
  assign n32364 = n32363 ^ n32285;
  assign n32365 = n32286 & ~n32364;
  assign n32366 = n32365 ^ n1149;
  assign n32367 = n32366 ^ n32283;
  assign n32368 = n32284 & ~n32367;
  assign n32369 = n32368 ^ n1157;
  assign n32370 = n32369 ^ n32281;
  assign n32371 = n32282 & ~n32370;
  assign n32372 = n32371 ^ n1309;
  assign n32373 = n32372 ^ n32279;
  assign n32374 = ~n32280 & n32373;
  assign n32375 = n32374 ^ n1324;
  assign n32377 = ~n3167 & ~n32376;
  assign n32382 = ~n32380 & ~n32381;
  assign n32387 = n32386 ^ n32383;
  assign n32389 = n32388 ^ n32387;
  assign n32390 = ~n32382 & n32389;
  assign n32392 = ~n2565 & n32391;
  assign n32393 = n32390 & ~n32392;
  assign n32394 = ~n32377 & n32393;
  assign n32395 = n32375 & n32394;
  assign n32408 = n32407 ^ n32395;
  assign n32409 = ~n3101 & n32264;
  assign n32410 = ~n2645 & ~n32266;
  assign n32411 = n32268 ^ n3081;
  assign n32412 = n32411 ^ n32269;
  assign n32413 = ~n32410 & ~n32412;
  assign n32414 = ~n32259 & ~n32262;
  assign n32415 = n32413 & ~n32414;
  assign n32416 = ~n32409 & n32415;
  assign n32417 = n32416 ^ n32395;
  assign n32418 = ~n32395 & ~n32417;
  assign n32419 = n32418 ^ n32395;
  assign n32420 = n32408 & ~n32419;
  assign n32421 = n32420 ^ n32418;
  assign n32422 = n32421 ^ n32395;
  assign n32423 = n32422 ^ n32416;
  assign n32424 = ~n32278 & ~n32423;
  assign n32425 = n32424 ^ n32278;
  assign n32426 = ~n32235 & ~n32238;
  assign n32427 = n32243 ^ n32242;
  assign n32428 = n32427 ^ n32244;
  assign n32429 = ~n32426 & ~n32428;
  assign n32430 = n32425 & n32429;
  assign n32431 = ~n32251 & n32430;
  assign n32432 = ~n32250 & ~n32431;
  assign n32227 = n32225 & n32226;
  assign n32153 = n32152 ^ n31990;
  assign n32154 = n31991 & n32153;
  assign n32155 = n32154 ^ n28757;
  assign n31985 = n31984 ^ n31509;
  assign n31986 = ~n31516 & ~n31985;
  assign n31987 = n31986 ^ n31515;
  assign n31504 = n30296 ^ n29498;
  assign n31505 = n31118 ^ n30296;
  assign n31506 = n31504 & n31505;
  assign n31507 = n31506 ^ n29498;
  assign n31503 = n31502 ^ n31481;
  assign n31508 = n31507 ^ n31503;
  assign n31988 = n31987 ^ n31508;
  assign n31989 = n31988 ^ n28799;
  assign n32156 = n32155 ^ n31989;
  assign n32228 = n32227 ^ n32156;
  assign n1733 = n1729 ^ n1689;
  assign n1743 = n1742 ^ n1733;
  assign n1744 = n1743 ^ n1710;
  assign n32229 = n32228 ^ n1744;
  assign n32433 = n32432 ^ n32229;
  assign n32438 = n32437 ^ n32433;
  assign n32439 = ~n28811 & ~n32438;
  assign n32440 = n32439 ^ n29817;
  assign n32486 = ~n1744 & n32228;
  assign n32487 = n32429 & ~n32486;
  assign n32488 = ~n32251 & n32487;
  assign n32489 = n32425 & n32488;
  assign n32490 = n32250 ^ n32228;
  assign n32491 = ~n32229 & n32490;
  assign n32492 = n32491 ^ n1744;
  assign n32493 = ~n32489 & ~n32492;
  assign n32483 = n30136 ^ n22801;
  assign n32484 = n32483 ^ n1715;
  assign n32485 = n32484 ^ n1822;
  assign n32494 = n32493 ^ n32485;
  assign n32481 = n32156 & ~n32228;
  assign n32474 = n30300 ^ n29544;
  assign n32475 = n31125 ^ n30300;
  assign n32476 = n32474 & n32475;
  assign n32477 = n32476 ^ n29544;
  assign n32460 = ~n31503 & ~n31507;
  assign n32461 = ~n31526 & ~n32460;
  assign n32462 = ~n31981 & n32461;
  assign n32463 = ~n31509 & n31515;
  assign n32464 = n32463 ^ n31516;
  assign n32465 = n32462 & ~n32464;
  assign n32466 = ~n31979 & n32465;
  assign n32467 = ~n31516 & ~n31536;
  assign n32468 = n32467 ^ n32463;
  assign n32469 = n32468 ^ n31507;
  assign n32470 = n31508 & ~n32469;
  assign n32471 = n32470 ^ n31503;
  assign n32472 = ~n32466 & ~n32471;
  assign n32459 = n31798 ^ n31795;
  assign n32473 = n32472 ^ n32459;
  assign n32478 = n32477 ^ n32473;
  assign n32479 = n32478 ^ n28900;
  assign n32447 = n31999 ^ n31990;
  assign n32448 = n31991 & n32447;
  assign n32449 = n32448 ^ n28757;
  assign n32450 = n32449 ^ n31988;
  assign n32451 = ~n31989 & ~n32450;
  assign n32452 = n32451 ^ n28799;
  assign n32453 = ~n28757 & ~n31990;
  assign n32454 = n28799 & ~n31988;
  assign n32455 = ~n32453 & ~n32454;
  assign n32456 = ~n32150 & n32455;
  assign n32457 = n32149 & n32456;
  assign n32458 = n32452 & ~n32457;
  assign n32480 = n32479 ^ n32458;
  assign n32482 = n32481 ^ n32480;
  assign n32495 = n32494 ^ n32482;
  assign n32442 = n31596 ^ n30678;
  assign n32443 = n30678 ^ n30338;
  assign n32444 = n32442 & n32443;
  assign n32445 = n32444 ^ n30338;
  assign n32441 = n32433 & ~n32437;
  assign n32446 = n32445 ^ n32441;
  assign n32496 = n32495 ^ n32446;
  assign n32955 = n32496 ^ n32439;
  assign n32956 = ~n32440 & n32955;
  assign n32957 = n32956 ^ n29817;
  assign n32780 = n32495 ^ n32445;
  assign n32781 = ~n32446 & n32780;
  assign n32782 = n32781 ^ n32441;
  assign n32775 = n30672 ^ n29695;
  assign n32776 = n31586 ^ n30672;
  assign n32777 = n32775 & n32776;
  assign n32778 = n32777 ^ n29695;
  assign n32752 = n32485 ^ n32482;
  assign n32753 = n32493 ^ n32482;
  assign n32754 = ~n32752 & ~n32753;
  assign n32755 = n32754 ^ n32485;
  assign n32703 = n32477 ^ n32459;
  assign n32704 = n32473 & ~n32703;
  assign n32705 = n32704 ^ n32477;
  assign n32698 = n30270 ^ n29595;
  assign n32699 = n31108 ^ n30270;
  assign n32700 = ~n32698 & n32699;
  assign n32701 = n32700 ^ n29595;
  assign n32572 = n31801 ^ n31793;
  assign n32702 = n32701 ^ n32572;
  assign n32726 = n32705 ^ n32702;
  assign n32735 = n32726 ^ n28894;
  assign n32721 = n32458 ^ n28900;
  assign n32722 = n32478 ^ n32458;
  assign n32723 = n32721 & n32722;
  assign n32724 = n32723 ^ n28900;
  assign n32736 = n32735 ^ n32724;
  assign n32734 = n32480 & ~n32481;
  assign n32750 = n32736 ^ n32734;
  assign n1818 = n1817 ^ n1766;
  assign n1828 = n1827 ^ n1818;
  assign n1832 = n1831 ^ n1828;
  assign n32751 = n32750 ^ n1832;
  assign n32774 = n32755 ^ n32751;
  assign n32779 = n32778 ^ n32774;
  assign n32953 = n32782 ^ n32779;
  assign n32954 = n32953 ^ n29810;
  assign n33050 = n32957 ^ n32954;
  assign n33257 = n33256 ^ n33050;
  assign n32498 = n23152 ^ n2065;
  assign n32499 = n32498 ^ n30971;
  assign n32500 = n32499 ^ n2220;
  assign n32501 = n32438 ^ n28811;
  assign n32502 = n32500 & n32501;
  assign n2229 = n2228 ^ n2135;
  assign n2230 = n2229 ^ n2222;
  assign n2231 = n2230 ^ n2210;
  assign n32503 = n32502 ^ n2231;
  assign n32497 = n32496 ^ n32440;
  assign n33258 = n32497 ^ n2231;
  assign n33259 = n32503 & ~n33258;
  assign n33260 = n33259 ^ n32502;
  assign n33261 = n33260 ^ n33050;
  assign n33262 = n33257 & ~n33261;
  assign n33263 = n33262 ^ n33256;
  assign n32958 = n32957 ^ n32953;
  assign n32959 = n32954 & n32958;
  assign n32960 = n32959 ^ n29810;
  assign n32783 = n32782 ^ n32774;
  assign n32784 = ~n32779 & ~n32783;
  assign n32785 = n32784 ^ n32782;
  assign n32769 = n30666 ^ n29687;
  assign n32770 = n31583 ^ n30666;
  assign n32771 = n32769 & n32770;
  assign n32772 = n32771 ^ n29687;
  assign n32756 = n32755 ^ n32750;
  assign n32757 = ~n32751 & n32756;
  assign n32758 = n32757 ^ n1832;
  assign n32725 = n32724 ^ n28894;
  assign n32727 = n32726 ^ n32724;
  assign n32728 = ~n32725 & n32727;
  assign n32729 = n32728 ^ n28894;
  assign n32706 = n32705 ^ n32701;
  assign n32707 = n32702 & ~n32706;
  assign n32708 = n32707 ^ n32705;
  assign n32693 = n30312 ^ n29612;
  assign n32694 = n31102 ^ n30312;
  assign n32695 = ~n32693 & n32694;
  assign n32696 = n32695 ^ n29612;
  assign n32560 = n31804 ^ n31791;
  assign n32697 = n32696 ^ n32560;
  assign n32719 = n32708 ^ n32697;
  assign n32720 = n32719 ^ n28844;
  assign n32738 = n32729 ^ n32720;
  assign n32737 = n32734 & ~n32736;
  assign n32745 = n32738 ^ n32737;
  assign n32749 = n32748 ^ n32745;
  assign n32768 = n32758 ^ n32749;
  assign n32773 = n32772 ^ n32768;
  assign n32951 = n32785 ^ n32773;
  assign n32952 = n32951 ^ n29804;
  assign n33051 = n32960 ^ n32952;
  assign n33252 = n33051 ^ n33050;
  assign n33249 = n30526 ^ n23097;
  assign n33250 = n33249 ^ n27142;
  assign n33251 = n33250 ^ n693;
  assign n33253 = n33252 ^ n33251;
  assign n33442 = n33263 ^ n33253;
  assign n32663 = n32336 ^ n32325;
  assign n34859 = n33442 ^ n32663;
  assign n32578 = n31522 ^ n30914;
  assign n32579 = n32459 ^ n31522;
  assign n32580 = n32578 & ~n32579;
  assign n32581 = n32580 ^ n30914;
  assign n32565 = n32375 & n32390;
  assign n32566 = ~n32401 & ~n32565;
  assign n32577 = n32566 ^ n32397;
  assign n32582 = n32581 ^ n32577;
  assign n32587 = n31529 ^ n30819;
  assign n32588 = n31529 ^ n31503;
  assign n32589 = n32587 & n32588;
  assign n32590 = n32589 ^ n30819;
  assign n32583 = n32383 ^ n32375;
  assign n32584 = n32387 & ~n32583;
  assign n32585 = n32584 ^ n32386;
  assign n32586 = n32585 ^ n32398;
  assign n32591 = n32590 ^ n32586;
  assign n32593 = n31619 ^ n30699;
  assign n32594 = n31619 ^ n31509;
  assign n32595 = ~n32593 & n32594;
  assign n32596 = n32595 ^ n30699;
  assign n32592 = n32387 ^ n32375;
  assign n32597 = n32596 ^ n32592;
  assign n32599 = n31630 ^ n30705;
  assign n32600 = n31630 ^ n31517;
  assign n32601 = n32599 & ~n32600;
  assign n32602 = n32601 ^ n30705;
  assign n32598 = n32372 ^ n32280;
  assign n32603 = n32602 ^ n32598;
  assign n32605 = n31639 ^ n30706;
  assign n32606 = n31639 ^ n31527;
  assign n32607 = ~n32605 & ~n32606;
  assign n32608 = n32607 ^ n30706;
  assign n32604 = n32369 ^ n32282;
  assign n32609 = n32608 ^ n32604;
  assign n32611 = n31641 ^ n30712;
  assign n32612 = n31941 ^ n31641;
  assign n32613 = ~n32611 & ~n32612;
  assign n32614 = n32613 ^ n30712;
  assign n32610 = n32366 ^ n32284;
  assign n32615 = n32614 ^ n32610;
  assign n32620 = n32363 ^ n32286;
  assign n32616 = n31653 ^ n30585;
  assign n32617 = n31945 ^ n31653;
  assign n32618 = ~n32616 & n32617;
  assign n32619 = n32618 ^ n30585;
  assign n32621 = n32620 ^ n32619;
  assign n32623 = n31659 ^ n30596;
  assign n32624 = n31935 ^ n31659;
  assign n32625 = ~n32623 & n32624;
  assign n32626 = n32625 ^ n30596;
  assign n32622 = n32360 ^ n32288;
  assign n32627 = n32626 ^ n32622;
  assign n32629 = n31491 ^ n30604;
  assign n32630 = n31927 ^ n31491;
  assign n32631 = ~n32629 & ~n32630;
  assign n32632 = n32631 ^ n30604;
  assign n32628 = n32357 ^ n32293;
  assign n32633 = n32632 ^ n32628;
  assign n32638 = n32354 ^ n32298;
  assign n32634 = n31294 ^ n30616;
  assign n32635 = n31919 ^ n31294;
  assign n32636 = ~n32634 & ~n32635;
  assign n32637 = n32636 ^ n30616;
  assign n32639 = n32638 ^ n32637;
  assign n32641 = n31187 ^ n30623;
  assign n32642 = n31898 ^ n31187;
  assign n32643 = n32641 & ~n32642;
  assign n32644 = n32643 ^ n30623;
  assign n32640 = n32351 ^ n32303;
  assign n32645 = n32644 ^ n32640;
  assign n32650 = n32348 ^ n32305;
  assign n32646 = n30634 ^ n30583;
  assign n32647 = n31904 ^ n30583;
  assign n32648 = ~n32646 & ~n32647;
  assign n32649 = n32648 ^ n30634;
  assign n32652 = n32650 ^ n32649;
  assign n32651 = n32649 & ~n32650;
  assign n32653 = n32652 ^ n32651;
  assign n32654 = n32653 ^ n32644;
  assign n32655 = n32645 & ~n32654;
  assign n32656 = n32655 ^ n32640;
  assign n32657 = n32656 ^ n32637;
  assign n32658 = ~n32639 & ~n32657;
  assign n32659 = n32658 ^ n32656;
  assign n32660 = n32659 ^ n32628;
  assign n32661 = ~n32633 & ~n32660;
  assign n32662 = n32661 ^ n32632;
  assign n32664 = n30662 ^ n30621;
  assign n32665 = n31549 ^ n30621;
  assign n32666 = n32664 & ~n32665;
  assign n32667 = n32666 ^ n30662;
  assign n32668 = ~n32663 & ~n32667;
  assign n32519 = n32339 ^ n32320;
  assign n32669 = n30656 ^ n30614;
  assign n32670 = n31543 ^ n30614;
  assign n32671 = n32669 & ~n32670;
  assign n32672 = n32671 ^ n30656;
  assign n32673 = n32519 & ~n32672;
  assign n32674 = ~n32668 & ~n32673;
  assign n32679 = n32333 ^ n32326;
  assign n32675 = n30632 ^ n30573;
  assign n32676 = n31555 ^ n30632;
  assign n32677 = n32675 & ~n32676;
  assign n32678 = n32677 ^ n30573;
  assign n32680 = n32679 ^ n32678;
  assign n32682 = n30639 ^ n30427;
  assign n32683 = n31561 ^ n30639;
  assign n32684 = ~n32682 & ~n32683;
  assign n32685 = n32684 ^ n30427;
  assign n32681 = n32330 ^ n32329;
  assign n32686 = n32685 ^ n32681;
  assign n32688 = n30651 ^ n30351;
  assign n32689 = n31567 ^ n30651;
  assign n32690 = n32688 & ~n32689;
  assign n32691 = n32690 ^ n30351;
  assign n32687 = n32327 ^ n2380;
  assign n32692 = n32691 ^ n32687;
  assign n32763 = n30653 ^ n29680;
  assign n32764 = n31573 ^ n30653;
  assign n32765 = ~n32763 & n32764;
  assign n32766 = n32765 ^ n29680;
  assign n32759 = n32758 ^ n32745;
  assign n32760 = ~n32749 & n32759;
  assign n32761 = n32760 ^ n32748;
  assign n32739 = n32737 & ~n32738;
  assign n32730 = n32729 ^ n32719;
  assign n32731 = ~n32720 & ~n32730;
  assign n32732 = n32731 ^ n28844;
  assign n32712 = n30321 ^ n29632;
  assign n32713 = n31092 ^ n30321;
  assign n32714 = n32712 & n32713;
  assign n32715 = n32714 ^ n29632;
  assign n32549 = n31807 ^ n31789;
  assign n32716 = n32715 ^ n32549;
  assign n32709 = n32708 ^ n32560;
  assign n32710 = ~n32697 & ~n32709;
  assign n32711 = n32710 ^ n32696;
  assign n32717 = n32716 ^ n32711;
  assign n32718 = n32717 ^ n28838;
  assign n32733 = n32732 ^ n32718;
  assign n32740 = n32739 ^ n32733;
  assign n32744 = n32743 ^ n32740;
  assign n32762 = n32761 ^ n32744;
  assign n32767 = n32766 ^ n32762;
  assign n32786 = n32785 ^ n32768;
  assign n32787 = ~n32773 & n32786;
  assign n32788 = n32787 ^ n32772;
  assign n32789 = n32788 ^ n32762;
  assign n32790 = ~n32767 & ~n32789;
  assign n32791 = n32790 ^ n32766;
  assign n32792 = n32791 ^ n32687;
  assign n32793 = ~n32692 & ~n32792;
  assign n32794 = n32793 ^ n32691;
  assign n32795 = n32794 ^ n32685;
  assign n32796 = n32686 & n32795;
  assign n32797 = n32796 ^ n32794;
  assign n32798 = n32797 ^ n32679;
  assign n32799 = ~n32680 & n32798;
  assign n32800 = n32799 ^ n32797;
  assign n32801 = n32674 & n32800;
  assign n32513 = n32342 ^ n32315;
  assign n32802 = n30647 ^ n30601;
  assign n32803 = n31541 ^ n30601;
  assign n32804 = n32802 & ~n32803;
  assign n32805 = n32804 ^ n30647;
  assign n32806 = n32513 & ~n32805;
  assign n32807 = n32801 & ~n32806;
  assign n32506 = n32345 ^ n32310;
  assign n32808 = n30641 ^ n30594;
  assign n32809 = n31906 ^ n30594;
  assign n32810 = ~n32808 & n32809;
  assign n32811 = n32810 ^ n30641;
  assign n32812 = ~n32506 & n32811;
  assign n32813 = n32807 & ~n32812;
  assign n32814 = n32811 ^ n32506;
  assign n32815 = n32805 ^ n32513;
  assign n32816 = n32672 ^ n32519;
  assign n32817 = n32667 ^ n32663;
  assign n32818 = n32817 ^ n32668;
  assign n32819 = ~n32816 & n32818;
  assign n32820 = n32819 ^ n32673;
  assign n32821 = n32820 ^ n32513;
  assign n32822 = ~n32815 & ~n32821;
  assign n32823 = n32822 ^ n32805;
  assign n32824 = n32823 ^ n32506;
  assign n32825 = ~n32814 & ~n32824;
  assign n32826 = n32825 ^ n32811;
  assign n32827 = ~n32813 & n32826;
  assign n32828 = ~n32640 & ~n32644;
  assign n32829 = n32637 & n32638;
  assign n32830 = ~n32628 & n32632;
  assign n32831 = ~n32651 & ~n32830;
  assign n32832 = ~n32829 & n32831;
  assign n32833 = ~n32828 & n32832;
  assign n32834 = n32827 & n32833;
  assign n32835 = n32834 ^ n32833;
  assign n32836 = n32662 & n32835;
  assign n32837 = n32836 ^ n32662;
  assign n32838 = n32837 ^ n32622;
  assign n32839 = ~n32627 & ~n32838;
  assign n32840 = n32839 ^ n32626;
  assign n32841 = n32840 ^ n32619;
  assign n32842 = n32621 & ~n32841;
  assign n32843 = n32842 ^ n32620;
  assign n32844 = n32843 ^ n32610;
  assign n32845 = ~n32615 & ~n32844;
  assign n32846 = n32845 ^ n32614;
  assign n32847 = n32846 ^ n32604;
  assign n32848 = ~n32609 & n32847;
  assign n32849 = n32848 ^ n32608;
  assign n32850 = n32849 ^ n32598;
  assign n32851 = n32603 & ~n32850;
  assign n32852 = n32851 ^ n32602;
  assign n32853 = n32852 ^ n32592;
  assign n32854 = ~n32597 & n32853;
  assign n32855 = n32854 ^ n32596;
  assign n32856 = n32855 ^ n32586;
  assign n32857 = ~n32591 & n32856;
  assign n32858 = n32857 ^ n32590;
  assign n32859 = n32858 ^ n32577;
  assign n32860 = ~n32582 & ~n32859;
  assign n32861 = n32860 ^ n32581;
  assign n32571 = n31512 ^ n30960;
  assign n32573 = n32572 ^ n31512;
  assign n32574 = n32571 & ~n32573;
  assign n32575 = n32574 ^ n30960;
  assign n32567 = n32566 ^ n32376;
  assign n32568 = n32397 & n32567;
  assign n32569 = n32568 ^ n3167;
  assign n32570 = n32569 ^ n32396;
  assign n32576 = n32575 ^ n32570;
  assign n32887 = n32861 ^ n32576;
  assign n32888 = n32887 ^ n29709;
  assign n32889 = n32858 ^ n32582;
  assign n32890 = n32889 ^ n29919;
  assign n32891 = n32855 ^ n32591;
  assign n32892 = n32891 ^ n29712;
  assign n32893 = n32852 ^ n32597;
  assign n32894 = n32893 ^ n29719;
  assign n32895 = n32849 ^ n32603;
  assign n32896 = n32895 ^ n29729;
  assign n32897 = n32846 ^ n32609;
  assign n32898 = n32897 ^ n29735;
  assign n32899 = n32843 ^ n32615;
  assign n32900 = n32899 ^ n29741;
  assign n32901 = n32840 ^ n32621;
  assign n32902 = n32901 ^ n29743;
  assign n32903 = n32837 ^ n32627;
  assign n32904 = n32903 ^ n29745;
  assign n32906 = ~n32651 & ~n32826;
  assign n32905 = ~n32651 & n32813;
  assign n32907 = n32906 ^ n32905;
  assign n32908 = n32905 ^ n32656;
  assign n32909 = ~n32905 & n32908;
  assign n32910 = n32909 ^ n32905;
  assign n32911 = n32907 & ~n32910;
  assign n32912 = n32911 ^ n32909;
  assign n32913 = n32912 ^ n32905;
  assign n32914 = n32913 ^ n32656;
  assign n32915 = ~n32828 & n32914;
  assign n32916 = n32915 ^ n32656;
  assign n32917 = n32916 ^ n32638;
  assign n32918 = n32639 & n32917;
  assign n32919 = n32918 ^ n32637;
  assign n32920 = n32919 ^ n32633;
  assign n32921 = n32920 ^ n29884;
  assign n32922 = n32916 ^ n32639;
  assign n32923 = n32922 ^ n29875;
  assign n32924 = ~n32653 & ~n32906;
  assign n32925 = ~n32905 & n32924;
  assign n32926 = n32925 ^ n32645;
  assign n32927 = n32926 ^ n29751;
  assign n32928 = n32827 ^ n32652;
  assign n32929 = n32928 ^ n29756;
  assign n32930 = ~n32807 & ~n32823;
  assign n32931 = n32930 ^ n32814;
  assign n32932 = n32931 ^ n29762;
  assign n32933 = ~n32801 & n32820;
  assign n32934 = n32933 ^ n32815;
  assign n32935 = n32934 ^ n29097;
  assign n32936 = n32800 ^ n32663;
  assign n32937 = n32817 & ~n32936;
  assign n32938 = n32937 ^ n32667;
  assign n32939 = n32938 ^ n32816;
  assign n32940 = n32939 ^ n29103;
  assign n32941 = n32817 ^ n32800;
  assign n32942 = n32941 ^ n29683;
  assign n32943 = n32797 ^ n32680;
  assign n32944 = n32943 ^ n29690;
  assign n32945 = n32794 ^ n32686;
  assign n32946 = n32945 ^ n29787;
  assign n32947 = n32791 ^ n32692;
  assign n32948 = n32947 ^ n29699;
  assign n32949 = n32788 ^ n32767;
  assign n32950 = n32949 ^ n29794;
  assign n32961 = n32960 ^ n32951;
  assign n32962 = n32952 & n32961;
  assign n32963 = n32962 ^ n29804;
  assign n32964 = n32963 ^ n32949;
  assign n32965 = ~n32950 & ~n32964;
  assign n32966 = n32965 ^ n29794;
  assign n32967 = n32966 ^ n32947;
  assign n32968 = ~n32948 & ~n32967;
  assign n32969 = n32968 ^ n29699;
  assign n32970 = n32969 ^ n32945;
  assign n32971 = ~n32946 & ~n32970;
  assign n32972 = n32971 ^ n29787;
  assign n32973 = n32972 ^ n32943;
  assign n32974 = ~n32944 & ~n32973;
  assign n32975 = n32974 ^ n29690;
  assign n32976 = n32975 ^ n32941;
  assign n32977 = n32942 & n32976;
  assign n32978 = n32977 ^ n29683;
  assign n32979 = n32978 ^ n32939;
  assign n32980 = n32940 & n32979;
  assign n32981 = n32980 ^ n29103;
  assign n32982 = n32981 ^ n32934;
  assign n32983 = n32935 & n32982;
  assign n32984 = n32983 ^ n29097;
  assign n32985 = n32984 ^ n32931;
  assign n32986 = n32932 & ~n32985;
  assign n32987 = n32986 ^ n29762;
  assign n32988 = n32987 ^ n32928;
  assign n32989 = n32929 & ~n32988;
  assign n32990 = n32989 ^ n29756;
  assign n32991 = n32990 ^ n32926;
  assign n32992 = n32927 & n32991;
  assign n32993 = n32992 ^ n29751;
  assign n32994 = n32993 ^ n32922;
  assign n32995 = ~n32923 & n32994;
  assign n32996 = n32995 ^ n29875;
  assign n32997 = n32996 ^ n32920;
  assign n32998 = ~n32921 & n32997;
  assign n32999 = n32998 ^ n29884;
  assign n33000 = n32999 ^ n32903;
  assign n33001 = ~n32904 & n33000;
  assign n33002 = n33001 ^ n29745;
  assign n33003 = n33002 ^ n32901;
  assign n33004 = n32902 & n33003;
  assign n33005 = n33004 ^ n29743;
  assign n33006 = n33005 ^ n32899;
  assign n33007 = n32900 & n33006;
  assign n33008 = n33007 ^ n29741;
  assign n33009 = n33008 ^ n32897;
  assign n33010 = ~n32898 & n33009;
  assign n33011 = n33010 ^ n29735;
  assign n33012 = n33011 ^ n32895;
  assign n33013 = ~n32896 & ~n33012;
  assign n33014 = n33013 ^ n29729;
  assign n33015 = n33014 ^ n32893;
  assign n33016 = n32894 & ~n33015;
  assign n33017 = n33016 ^ n29719;
  assign n33018 = n33017 ^ n32891;
  assign n33019 = n32892 & ~n33018;
  assign n33020 = n33019 ^ n29712;
  assign n33021 = n33020 ^ n32889;
  assign n33022 = n32890 & ~n33021;
  assign n33023 = n33022 ^ n29919;
  assign n33024 = n33023 ^ n32887;
  assign n33025 = ~n32888 & ~n33024;
  assign n33026 = n33025 ^ n29709;
  assign n32862 = n32861 ^ n32570;
  assign n32863 = n32576 & n32862;
  assign n32864 = n32863 ^ n32575;
  assign n32559 = n31118 ^ n30288;
  assign n32561 = n32560 ^ n31118;
  assign n32562 = ~n32559 & ~n32561;
  assign n32563 = n32562 ^ n30288;
  assign n32530 = ~n32395 & ~n32407;
  assign n32558 = n32530 ^ n32411;
  assign n32564 = n32563 ^ n32558;
  assign n32885 = n32864 ^ n32564;
  assign n32886 = n32885 ^ n29510;
  assign n33042 = n33026 ^ n32886;
  assign n33043 = n33023 ^ n32888;
  assign n33044 = n33017 ^ n32892;
  assign n33045 = n33014 ^ n32894;
  assign n33046 = n32996 ^ n32921;
  assign n33047 = n32984 ^ n32932;
  assign n33048 = n32969 ^ n32946;
  assign n33049 = n32963 ^ n32950;
  assign n33052 = n33050 & ~n33051;
  assign n33053 = ~n33049 & n33052;
  assign n33054 = n32966 ^ n32948;
  assign n33055 = ~n33053 & ~n33054;
  assign n33056 = ~n33048 & ~n33055;
  assign n33057 = n32972 ^ n32944;
  assign n33058 = n33056 & n33057;
  assign n33059 = n32975 ^ n32942;
  assign n33060 = ~n33058 & ~n33059;
  assign n33061 = n32978 ^ n32940;
  assign n33062 = n33060 & n33061;
  assign n33063 = n32981 ^ n32935;
  assign n33064 = ~n33062 & n33063;
  assign n33065 = ~n33047 & n33064;
  assign n33066 = n32987 ^ n32929;
  assign n33067 = n33065 & ~n33066;
  assign n33068 = n32990 ^ n32927;
  assign n33069 = n33067 & ~n33068;
  assign n33070 = n32993 ^ n32923;
  assign n33071 = ~n33069 & n33070;
  assign n33072 = ~n33046 & ~n33071;
  assign n33073 = n32999 ^ n32904;
  assign n33074 = n33072 & ~n33073;
  assign n33075 = n33002 ^ n32902;
  assign n33076 = n33074 & n33075;
  assign n33077 = n33005 ^ n32900;
  assign n33078 = ~n33076 & n33077;
  assign n33079 = n33008 ^ n32898;
  assign n33080 = ~n33078 & ~n33079;
  assign n33081 = n33011 ^ n32896;
  assign n33082 = n33080 & ~n33081;
  assign n33083 = n33045 & ~n33082;
  assign n33084 = n33044 & n33083;
  assign n33085 = n33020 ^ n32890;
  assign n33086 = n33084 & n33085;
  assign n33087 = n33043 & ~n33086;
  assign n33088 = ~n33042 & n33087;
  assign n33027 = n33026 ^ n32885;
  assign n33028 = ~n32886 & ~n33027;
  assign n33029 = n33028 ^ n29510;
  assign n32865 = n32864 ^ n32558;
  assign n32866 = n32564 & n32865;
  assign n32867 = n32866 ^ n32563;
  assign n32553 = n32530 ^ n32268;
  assign n32554 = ~n32411 & ~n32553;
  assign n32555 = n32554 ^ n3081;
  assign n32556 = n32555 ^ n32267;
  assign n32548 = n31125 ^ n30291;
  assign n32550 = n32549 ^ n31125;
  assign n32551 = n32548 & ~n32550;
  assign n32552 = n32551 ^ n30291;
  assign n32557 = n32556 ^ n32552;
  assign n32883 = n32867 ^ n32557;
  assign n32884 = n32883 ^ n29504;
  assign n33041 = n33029 ^ n32884;
  assign n33146 = n33088 ^ n33041;
  assign n33150 = n33149 ^ n33146;
  assign n33151 = n33087 ^ n33042;
  assign n33152 = n33151 ^ n2957;
  assign n33153 = n33086 ^ n33043;
  assign n33157 = n33156 ^ n33153;
  assign n33158 = n33085 ^ n33084;
  assign n2821 = n2817 ^ n2760;
  assign n2825 = n2824 ^ n2821;
  assign n2826 = n2825 ^ n1529;
  assign n33159 = n33158 ^ n2826;
  assign n33160 = n33083 ^ n33044;
  assign n2732 = n2680 ^ n1574;
  assign n2733 = n2732 ^ n2729;
  assign n2737 = n2736 ^ n2733;
  assign n33161 = n33160 ^ n2737;
  assign n33162 = n33082 ^ n33045;
  assign n2705 = n2698 ^ n2665;
  assign n2718 = n2717 ^ n2705;
  assign n2722 = n2721 ^ n2718;
  assign n33163 = n33162 ^ n2722;
  assign n3193 = n3189 ^ n2601;
  assign n3200 = n3199 ^ n3193;
  assign n3201 = n3200 ^ n2714;
  assign n33164 = n33081 ^ n33080;
  assign n33165 = n3201 & n33164;
  assign n33166 = n33165 ^ n33162;
  assign n33167 = ~n33163 & n33166;
  assign n33168 = n33167 ^ n2722;
  assign n33169 = n33168 ^ n2737;
  assign n33170 = n33161 & ~n33169;
  assign n33171 = n33170 ^ n33160;
  assign n33172 = n33171 ^ n33158;
  assign n33173 = n33159 & ~n33172;
  assign n33174 = n33173 ^ n2826;
  assign n33201 = n33071 ^ n33046;
  assign n1462 = n1419 ^ n1353;
  assign n1463 = n1462 ^ n1459;
  assign n1467 = n1466 ^ n1463;
  assign n33202 = n33201 ^ n1467;
  assign n33203 = n33070 ^ n33069;
  assign n1444 = n1338 ^ n1252;
  assign n1451 = n1450 ^ n1444;
  assign n1452 = n1451 ^ n1178;
  assign n33204 = n33203 ^ n1452;
  assign n33206 = n3347 ^ n1237;
  assign n33207 = n33206 ^ n1013;
  assign n33208 = n33207 ^ n1448;
  assign n33205 = n33068 ^ n33067;
  assign n33209 = n33208 ^ n33205;
  assign n33211 = n30484 ^ n1228;
  assign n33212 = n33211 ^ n27130;
  assign n33213 = n33212 ^ n1008;
  assign n33210 = n33066 ^ n33065;
  assign n33214 = n33213 ^ n33210;
  assign n33215 = n33064 ^ n33047;
  assign n864 = n863 ^ n812;
  assign n874 = n873 ^ n864;
  assign n878 = n877 ^ n874;
  assign n33216 = n33215 ^ n878;
  assign n33218 = n30469 ^ n23070;
  assign n33219 = n33218 ^ n787;
  assign n33220 = n33219 ^ n868;
  assign n33217 = n33063 ^ n33062;
  assign n33221 = n33220 ^ n33217;
  assign n33222 = n33061 ^ n33060;
  assign n775 = n774 ^ n756;
  assign n776 = n775 ^ n632;
  assign n780 = n779 ^ n776;
  assign n33223 = n33222 ^ n780;
  assign n33224 = n33059 ^ n33058;
  assign n33228 = n33227 ^ n33224;
  assign n33230 = n30501 ^ n600;
  assign n33231 = n33230 ^ n27181;
  assign n33232 = n33231 ^ n3266;
  assign n33229 = n33057 ^ n33056;
  assign n33233 = n33232 ^ n33229;
  assign n33234 = n33055 ^ n33048;
  assign n33238 = n33237 ^ n33234;
  assign n33240 = n30511 ^ n23106;
  assign n33241 = n33240 ^ n27167;
  assign n33242 = n33241 ^ n22128;
  assign n33239 = n33054 ^ n33053;
  assign n33243 = n33242 ^ n33239;
  assign n33245 = n30534 ^ n23082;
  assign n33246 = n33245 ^ n27158;
  assign n33247 = n33246 ^ n22133;
  assign n33244 = n33052 ^ n33049;
  assign n33248 = n33247 ^ n33244;
  assign n33264 = n33263 ^ n33252;
  assign n33265 = n33253 & ~n33264;
  assign n33266 = n33265 ^ n33251;
  assign n33267 = n33266 ^ n33244;
  assign n33268 = n33248 & ~n33267;
  assign n33269 = n33268 ^ n33247;
  assign n33270 = n33269 ^ n33242;
  assign n33271 = n33243 & ~n33270;
  assign n33272 = n33271 ^ n33239;
  assign n33273 = n33272 ^ n33234;
  assign n33274 = ~n33238 & n33273;
  assign n33275 = n33274 ^ n33237;
  assign n33276 = n33275 ^ n33229;
  assign n33277 = ~n33233 & n33276;
  assign n33278 = n33277 ^ n33232;
  assign n33279 = n33278 ^ n33224;
  assign n33280 = n33228 & ~n33279;
  assign n33281 = n33280 ^ n33227;
  assign n33282 = n33281 ^ n33222;
  assign n33283 = n33223 & ~n33282;
  assign n33284 = n33283 ^ n780;
  assign n33285 = n33284 ^ n33217;
  assign n33286 = n33221 & ~n33285;
  assign n33287 = n33286 ^ n33220;
  assign n33288 = n33287 ^ n33215;
  assign n33289 = n33216 & ~n33288;
  assign n33290 = n33289 ^ n878;
  assign n33291 = n33290 ^ n33210;
  assign n33292 = n33214 & ~n33291;
  assign n33293 = n33292 ^ n33213;
  assign n33294 = n33293 ^ n33205;
  assign n33295 = n33209 & ~n33294;
  assign n33296 = n33295 ^ n33208;
  assign n33297 = n33296 ^ n33203;
  assign n33298 = ~n33204 & n33297;
  assign n33299 = n33298 ^ n1452;
  assign n33300 = n33299 ^ n33201;
  assign n33301 = ~n33202 & n33300;
  assign n33302 = n33301 ^ n1467;
  assign n33180 = n33077 ^ n33076;
  assign n33181 = n31006 ^ n3175;
  assign n33182 = n33181 ^ n27116;
  assign n33183 = n33182 ^ n3041;
  assign n33303 = n33180 & ~n33183;
  assign n33187 = n33075 ^ n33074;
  assign n33188 = n31001 ^ n23486;
  assign n33189 = n33188 ^ n3023;
  assign n33190 = n33189 ^ n2438;
  assign n33193 = n33187 & ~n33190;
  assign n33185 = n33073 ^ n33072;
  assign n1480 = n1435 ^ n1371;
  assign n1481 = n1480 ^ n1474;
  assign n1485 = n1484 ^ n1481;
  assign n33304 = n33185 ^ n1485;
  assign n33186 = n1485 & n33185;
  assign n33305 = n33304 ^ n33186;
  assign n33175 = n33079 ^ n33078;
  assign n33306 = n33175 & ~n33178;
  assign n33307 = n33305 & ~n33306;
  assign n33308 = ~n33193 & n33307;
  assign n33309 = ~n33303 & n33308;
  assign n33310 = n33302 & n33309;
  assign n33179 = n33178 ^ n33175;
  assign n33184 = n33183 ^ n33180;
  assign n33191 = n33190 ^ n33187;
  assign n33192 = ~n33186 & ~n33191;
  assign n33194 = n33193 ^ n33192;
  assign n33195 = n33194 ^ n33180;
  assign n33196 = ~n33184 & ~n33195;
  assign n33197 = n33196 ^ n33183;
  assign n33198 = n33197 ^ n33175;
  assign n33199 = ~n33179 & n33198;
  assign n33200 = n33199 ^ n33178;
  assign n33311 = n33310 ^ n33200;
  assign n33312 = ~n2737 & ~n33160;
  assign n33313 = ~n2722 & n33162;
  assign n33314 = n33164 ^ n3201;
  assign n33315 = n33314 ^ n33165;
  assign n33316 = ~n33313 & n33315;
  assign n33317 = ~n2826 & ~n33158;
  assign n33318 = n33316 & ~n33317;
  assign n33319 = ~n33312 & n33318;
  assign n33320 = n33319 ^ n33310;
  assign n33321 = ~n33310 & ~n33320;
  assign n33322 = n33321 ^ n33310;
  assign n33323 = n33311 & ~n33322;
  assign n33324 = n33323 ^ n33321;
  assign n33325 = n33324 ^ n33310;
  assign n33326 = n33325 ^ n33319;
  assign n33327 = ~n33174 & ~n33326;
  assign n33328 = n33327 ^ n33174;
  assign n33329 = n33328 ^ n33153;
  assign n33330 = n33157 & ~n33329;
  assign n33331 = n33330 ^ n33156;
  assign n33332 = n33331 ^ n33151;
  assign n33333 = n33152 & ~n33332;
  assign n33334 = n33333 ^ n2957;
  assign n33335 = n33334 ^ n33146;
  assign n33336 = n33150 & ~n33335;
  assign n33337 = n33336 ^ n33149;
  assign n33089 = ~n33041 & n33088;
  assign n33030 = n33029 ^ n32883;
  assign n33031 = n32884 & ~n33030;
  assign n33032 = n33031 ^ n29504;
  assign n32868 = n32867 ^ n32556;
  assign n32869 = n32557 & ~n32868;
  assign n32870 = n32869 ^ n32552;
  assign n32543 = n31108 ^ n30296;
  assign n32544 = n31847 ^ n31108;
  assign n32545 = n32543 & ~n32544;
  assign n32546 = n32545 ^ n30296;
  assign n32531 = n32413 & ~n32530;
  assign n32532 = ~n32272 & ~n32531;
  assign n32542 = n32532 ^ n32265;
  assign n32547 = n32546 ^ n32542;
  assign n32881 = n32870 ^ n32547;
  assign n32882 = n32881 ^ n29498;
  assign n33040 = n33032 ^ n32882;
  assign n33141 = n33089 ^ n33040;
  assign n33145 = n33144 ^ n33141;
  assign n33370 = n33337 ^ n33145;
  assign n33371 = n31586 ^ n30685;
  assign n33372 = n32687 ^ n31586;
  assign n33373 = ~n33371 & n33372;
  assign n33374 = n33373 ^ n30685;
  assign n33375 = n33370 & ~n33374;
  assign n33364 = n31583 ^ n30678;
  assign n33365 = n32681 ^ n31583;
  assign n33366 = n33364 & ~n33365;
  assign n33367 = n33366 ^ n30678;
  assign n33415 = n33375 ^ n33367;
  assign n33338 = n33337 ^ n33141;
  assign n33339 = n33145 & ~n33338;
  assign n33340 = n33339 ^ n33144;
  assign n33033 = n33032 ^ n32881;
  assign n33034 = n32882 & ~n33033;
  assign n33035 = n33034 ^ n29498;
  assign n32871 = n32870 ^ n32542;
  assign n32872 = n32547 & ~n32871;
  assign n32873 = n32872 ^ n32546;
  assign n32537 = n31102 ^ n30300;
  assign n32538 = n31841 ^ n31102;
  assign n32539 = ~n32537 & ~n32538;
  assign n32540 = n32539 ^ n30300;
  assign n32533 = n32532 ^ n32264;
  assign n32534 = ~n32265 & ~n32533;
  assign n32535 = n32534 ^ n3101;
  assign n32536 = n32535 ^ n32263;
  assign n32541 = n32540 ^ n32536;
  assign n32879 = n32873 ^ n32541;
  assign n32880 = n32879 ^ n29544;
  assign n33091 = n33035 ^ n32880;
  assign n33090 = ~n33040 & n33089;
  assign n33136 = n33091 ^ n33090;
  assign n33140 = n33139 ^ n33136;
  assign n33368 = n33340 ^ n33140;
  assign n33416 = n33415 ^ n33368;
  assign n33412 = n33374 ^ n33370;
  assign n33413 = ~n29703 & ~n33412;
  assign n33414 = n33413 ^ n30338;
  assign n33495 = n33416 ^ n33414;
  assign n2187 = n2150 ^ n2099;
  assign n2188 = n2187 ^ n2170;
  assign n2192 = n2191 ^ n2188;
  assign n33492 = n33412 ^ n29703;
  assign n33493 = n2192 & n33492;
  assign n2336 = n2246 ^ n2202;
  assign n2337 = n2336 ^ n2318;
  assign n2344 = n2343 ^ n2337;
  assign n33494 = n33493 ^ n2344;
  assign n34228 = n33495 ^ n33494;
  assign n34860 = n34228 ^ n33442;
  assign n34861 = n34859 & n34860;
  assign n34862 = n34861 ^ n32663;
  assign n33398 = n33260 ^ n33257;
  assign n34853 = n33398 ^ n32679;
  assign n34200 = n33492 ^ n2192;
  assign n34854 = n34200 ^ n33398;
  assign n34855 = n34853 & ~n34854;
  assign n34856 = n34855 ^ n32679;
  assign n34714 = n32238 ^ n1684;
  assign n34715 = n34714 ^ n28561;
  assign n34716 = n34715 ^ n23468;
  assign n33672 = n33287 ^ n33216;
  assign n33668 = n31941 ^ n31659;
  assign n33669 = n32592 ^ n31941;
  assign n33670 = ~n33668 & ~n33669;
  assign n33671 = n33670 ^ n31659;
  assign n33674 = n33672 ^ n33671;
  assign n33600 = n33284 ^ n33221;
  assign n33596 = n31945 ^ n31491;
  assign n33597 = n32598 ^ n31945;
  assign n33598 = n33596 & n33597;
  assign n33599 = n33598 ^ n31491;
  assign n33601 = n33600 ^ n33599;
  assign n33602 = n31935 ^ n31294;
  assign n33603 = n32604 ^ n31935;
  assign n33604 = n33602 & ~n33603;
  assign n33605 = n33604 ^ n31294;
  assign n33542 = n33281 ^ n33223;
  assign n33606 = n33605 ^ n33542;
  assign n33611 = n33278 ^ n33228;
  assign n33607 = n31927 ^ n31187;
  assign n33608 = n32610 ^ n31927;
  assign n33609 = n33607 & ~n33608;
  assign n33610 = n33609 ^ n31187;
  assign n33612 = n33611 ^ n33610;
  assign n33617 = n33275 ^ n33233;
  assign n33613 = n31919 ^ n30583;
  assign n33614 = n32620 ^ n31919;
  assign n33615 = n33613 & ~n33614;
  assign n33616 = n33615 ^ n30583;
  assign n33618 = n33617 ^ n33616;
  assign n33394 = n31543 ^ n30632;
  assign n33395 = n32650 ^ n31543;
  assign n33396 = n33394 & ~n33395;
  assign n33397 = n33396 ^ n30632;
  assign n33399 = n33398 ^ n33397;
  assign n32505 = n31549 ^ n30639;
  assign n32507 = n32506 ^ n31549;
  assign n32508 = ~n32505 & ~n32507;
  assign n32509 = n32508 ^ n30639;
  assign n32504 = n32503 ^ n32497;
  assign n32510 = n32509 ^ n32504;
  assign n32512 = n31555 ^ n30651;
  assign n32514 = n32513 ^ n31555;
  assign n32515 = n32512 & n32514;
  assign n32516 = n32515 ^ n30651;
  assign n32511 = n32501 ^ n32500;
  assign n32517 = n32516 ^ n32511;
  assign n32874 = n32873 ^ n32536;
  assign n32875 = ~n32541 & ~n32874;
  assign n32876 = n32875 ^ n32540;
  assign n32525 = n31092 ^ n30270;
  assign n32526 = n31835 ^ n31092;
  assign n32527 = n32525 & n32526;
  assign n32528 = n32527 ^ n30270;
  assign n32523 = n32425 ^ n32242;
  assign n32524 = n32523 ^ n32243;
  assign n32529 = n32528 ^ n32524;
  assign n32877 = n32876 ^ n32529;
  assign n32878 = n32877 ^ n29595;
  assign n33036 = n33035 ^ n32879;
  assign n33037 = n32880 & n33036;
  assign n33038 = n33037 ^ n29544;
  assign n33108 = n33038 ^ n32877;
  assign n33109 = ~n32878 & ~n33108;
  assign n33110 = n33109 ^ n29595;
  assign n33101 = n30693 ^ n30312;
  assign n33102 = n31825 ^ n30693;
  assign n33103 = ~n33101 & ~n33102;
  assign n33104 = n33103 ^ n30312;
  assign n33097 = n32425 ^ n32243;
  assign n33098 = ~n32427 & n33097;
  assign n33099 = n33098 ^ n32242;
  assign n33100 = n33099 ^ n32239;
  assign n33105 = n33104 ^ n33100;
  assign n33094 = n32876 ^ n32524;
  assign n33095 = n32529 & ~n33094;
  assign n33096 = n33095 ^ n32528;
  assign n33106 = n33105 ^ n33096;
  assign n33107 = n33106 ^ n29612;
  assign n33111 = n33110 ^ n33107;
  assign n33039 = n33038 ^ n32878;
  assign n33092 = ~n33090 & n33091;
  assign n33093 = n33039 & n33092;
  assign n33132 = n33111 ^ n33093;
  assign n1934 = n1903 ^ n1867;
  assign n1935 = n1934 ^ n1931;
  assign n1939 = n1938 ^ n1935;
  assign n33133 = n33132 ^ n1939;
  assign n33134 = n33092 ^ n33039;
  assign n1922 = n1891 ^ n1852;
  assign n1923 = n1922 ^ n1921;
  assign n1924 = n1923 ^ n1912;
  assign n33135 = n33134 ^ n1924;
  assign n33341 = n33340 ^ n33136;
  assign n33342 = ~n33140 & n33341;
  assign n33343 = n33342 ^ n33139;
  assign n33344 = n33343 ^ n33134;
  assign n33345 = n33135 & ~n33344;
  assign n33346 = n33345 ^ n1924;
  assign n33347 = n33346 ^ n33132;
  assign n33348 = n33133 & ~n33347;
  assign n33349 = n33348 ^ n1939;
  assign n33125 = n33110 ^ n29612;
  assign n33126 = n33110 ^ n33106;
  assign n33127 = n33125 & ~n33126;
  assign n33128 = n33127 ^ n29612;
  assign n33120 = n33100 ^ n33096;
  assign n33121 = ~n33105 & n33120;
  assign n33122 = n33121 ^ n33104;
  assign n33117 = ~n32247 & ~n32430;
  assign n33118 = n33117 ^ n32234;
  assign n33113 = n30687 ^ n30321;
  assign n33114 = n31823 ^ n30687;
  assign n33115 = n33113 & n33114;
  assign n33116 = n33115 ^ n30321;
  assign n33119 = n33118 ^ n33116;
  assign n33123 = n33122 ^ n33119;
  assign n33124 = n33123 ^ n29632;
  assign n33129 = n33128 ^ n33124;
  assign n33112 = n33093 & n33111;
  assign n33130 = n33129 ^ n33112;
  assign n2047 = n2039 ^ n1978;
  assign n2054 = n2053 ^ n2047;
  assign n2058 = n2057 ^ n2054;
  assign n33131 = n33130 ^ n2058;
  assign n33350 = n33349 ^ n33131;
  assign n32518 = n31561 ^ n30653;
  assign n32520 = n32519 ^ n31561;
  assign n32521 = ~n32518 & ~n32520;
  assign n32522 = n32521 ^ n30653;
  assign n33351 = n33350 ^ n32522;
  assign n33356 = n33346 ^ n33133;
  assign n33352 = n32663 ^ n31567;
  assign n33353 = n31567 ^ n30666;
  assign n33354 = ~n33352 & n33353;
  assign n33355 = n33354 ^ n30666;
  assign n33357 = n33356 ^ n33355;
  assign n33359 = n32679 ^ n31573;
  assign n33360 = n31573 ^ n30672;
  assign n33361 = n33359 & n33360;
  assign n33362 = n33361 ^ n30672;
  assign n33358 = n33343 ^ n33135;
  assign n33363 = n33362 ^ n33358;
  assign n33369 = n33368 ^ n33367;
  assign n33376 = n33375 ^ n33368;
  assign n33377 = ~n33369 & ~n33376;
  assign n33378 = n33377 ^ n33375;
  assign n33379 = n33378 ^ n33358;
  assign n33380 = ~n33363 & ~n33379;
  assign n33381 = n33380 ^ n33362;
  assign n33382 = n33381 ^ n33356;
  assign n33383 = n33357 & n33382;
  assign n33384 = n33383 ^ n33355;
  assign n33385 = n33384 ^ n33350;
  assign n33386 = n33351 & ~n33385;
  assign n33387 = n33386 ^ n32522;
  assign n33388 = n33387 ^ n32511;
  assign n33389 = n32517 & n33388;
  assign n33390 = n33389 ^ n32511;
  assign n33391 = n33390 ^ n32504;
  assign n33392 = ~n32510 & ~n33391;
  assign n33393 = n33392 ^ n32509;
  assign n33444 = n33398 ^ n33393;
  assign n33445 = n33399 & n33444;
  assign n33446 = n33445 ^ n33397;
  assign n33527 = n31906 ^ n30614;
  assign n33528 = n32638 ^ n31906;
  assign n33529 = ~n33527 & ~n33528;
  assign n33530 = n33529 ^ n30614;
  assign n33531 = n33266 ^ n33248;
  assign n33619 = ~n33530 & ~n33531;
  assign n33438 = n31541 ^ n30621;
  assign n33439 = n32640 ^ n31541;
  assign n33440 = n33438 & ~n33439;
  assign n33441 = n33440 ^ n30621;
  assign n33620 = n33441 & n33442;
  assign n33443 = n33442 ^ n33441;
  assign n33621 = n33620 ^ n33443;
  assign n33622 = ~n33619 & n33621;
  assign n33623 = n31904 ^ n30601;
  assign n33624 = n32628 ^ n31904;
  assign n33625 = n33623 & ~n33624;
  assign n33626 = n33625 ^ n30601;
  assign n33627 = n33269 ^ n33243;
  assign n33628 = ~n33626 & ~n33627;
  assign n33629 = n33622 & ~n33628;
  assign n33630 = n31898 ^ n30594;
  assign n33631 = n32622 ^ n31898;
  assign n33632 = n33630 & n33631;
  assign n33633 = n33632 ^ n30594;
  assign n33634 = n33272 ^ n33238;
  assign n33635 = ~n33633 & n33634;
  assign n33636 = n33629 & ~n33635;
  assign n33637 = n33446 & n33636;
  assign n33638 = n33634 ^ n33633;
  assign n33639 = n33627 ^ n33626;
  assign n33532 = n33531 ^ n33530;
  assign n33640 = n33620 ^ n33530;
  assign n33641 = n33532 & ~n33640;
  assign n33642 = n33641 ^ n33531;
  assign n33643 = n33642 ^ n33627;
  assign n33644 = n33639 & ~n33643;
  assign n33645 = n33644 ^ n33626;
  assign n33646 = n33645 ^ n33633;
  assign n33647 = ~n33638 & ~n33646;
  assign n33648 = n33647 ^ n33634;
  assign n33649 = ~n33637 & n33648;
  assign n33650 = n33649 ^ n33617;
  assign n33651 = ~n33618 & ~n33650;
  assign n33652 = n33651 ^ n33616;
  assign n33653 = n33652 ^ n33610;
  assign n33654 = ~n33612 & n33653;
  assign n33655 = n33654 ^ n33652;
  assign n33656 = n33655 ^ n33542;
  assign n33657 = n33606 & ~n33656;
  assign n33658 = n33657 ^ n33605;
  assign n33659 = n33658 ^ n33600;
  assign n33660 = n33601 & ~n33659;
  assign n33661 = n33660 ^ n33599;
  assign n33808 = n33672 ^ n33661;
  assign n33809 = ~n33674 & ~n33808;
  assign n33810 = n33809 ^ n33671;
  assign n33666 = n33290 ^ n33214;
  assign n33662 = n31653 ^ n31527;
  assign n33663 = n32586 ^ n31527;
  assign n33664 = ~n33662 & ~n33663;
  assign n33665 = n33664 ^ n31653;
  assign n33729 = n33666 ^ n33665;
  assign n33811 = n33810 ^ n33729;
  assign n33812 = n33811 ^ n30585;
  assign n33813 = n33674 ^ n33661;
  assign n33814 = n33813 ^ n30596;
  assign n33815 = n33658 ^ n33601;
  assign n33816 = n33815 ^ n30604;
  assign n33817 = n33655 ^ n33606;
  assign n33818 = n33817 ^ n30616;
  assign n33819 = n33652 ^ n33612;
  assign n33820 = n33819 ^ n30623;
  assign n33821 = n33649 ^ n33618;
  assign n33822 = n33821 ^ n30634;
  assign n33823 = n33446 & n33622;
  assign n33824 = ~n33642 & ~n33823;
  assign n33825 = n33824 ^ n33627;
  assign n33826 = n33639 & n33825;
  assign n33827 = n33826 ^ n33626;
  assign n33828 = n33827 ^ n33638;
  assign n33829 = n33828 ^ n30641;
  assign n33830 = n33824 ^ n33639;
  assign n33831 = n33830 ^ n30647;
  assign n33524 = n33446 ^ n33442;
  assign n33525 = n33443 & ~n33524;
  assign n33526 = n33525 ^ n33441;
  assign n33533 = n33532 ^ n33526;
  assign n33534 = n33533 ^ n30656;
  assign n33447 = n33446 ^ n33443;
  assign n33448 = n33447 ^ n30662;
  assign n33400 = n33399 ^ n33393;
  assign n33401 = n33400 ^ n30573;
  assign n33402 = n33390 ^ n32510;
  assign n33403 = n33402 ^ n30427;
  assign n33404 = n33387 ^ n32517;
  assign n33405 = n33404 ^ n30351;
  assign n33406 = n33384 ^ n33351;
  assign n33407 = n33406 ^ n29680;
  assign n33408 = n33381 ^ n33357;
  assign n33409 = n33408 ^ n29687;
  assign n33410 = n33378 ^ n33363;
  assign n33411 = n33410 ^ n29695;
  assign n33417 = n33416 ^ n33413;
  assign n33418 = ~n33414 & ~n33417;
  assign n33419 = n33418 ^ n30338;
  assign n33420 = n33419 ^ n33410;
  assign n33421 = n33411 & ~n33420;
  assign n33422 = n33421 ^ n29695;
  assign n33423 = n33422 ^ n33408;
  assign n33424 = ~n33409 & ~n33423;
  assign n33425 = n33424 ^ n29687;
  assign n33426 = n33425 ^ n33406;
  assign n33427 = ~n33407 & ~n33426;
  assign n33428 = n33427 ^ n29680;
  assign n33429 = n33428 ^ n33404;
  assign n33430 = n33405 & n33429;
  assign n33431 = n33430 ^ n30351;
  assign n33432 = n33431 ^ n33402;
  assign n33433 = ~n33403 & n33432;
  assign n33434 = n33433 ^ n30427;
  assign n33435 = n33434 ^ n33400;
  assign n33436 = ~n33401 & n33435;
  assign n33437 = n33436 ^ n30573;
  assign n33521 = n33447 ^ n33437;
  assign n33522 = n33448 & ~n33521;
  assign n33523 = n33522 ^ n30662;
  assign n33832 = n33533 ^ n33523;
  assign n33833 = n33534 & ~n33832;
  assign n33834 = n33833 ^ n30656;
  assign n33835 = n33834 ^ n33830;
  assign n33836 = ~n33831 & n33835;
  assign n33837 = n33836 ^ n30647;
  assign n33838 = n33837 ^ n33828;
  assign n33839 = n33829 & n33838;
  assign n33840 = n33839 ^ n30641;
  assign n33841 = n33840 ^ n33821;
  assign n33842 = ~n33822 & n33841;
  assign n33843 = n33842 ^ n30634;
  assign n33844 = n33843 ^ n33819;
  assign n33845 = n33820 & n33844;
  assign n33846 = n33845 ^ n30623;
  assign n33847 = n33846 ^ n33817;
  assign n33848 = ~n33818 & ~n33847;
  assign n33849 = n33848 ^ n30616;
  assign n33850 = n33849 ^ n33815;
  assign n33851 = ~n33816 & n33850;
  assign n33852 = n33851 ^ n30604;
  assign n33853 = n33852 ^ n33813;
  assign n33854 = ~n33814 & ~n33853;
  assign n33855 = n33854 ^ n30596;
  assign n33856 = n33855 ^ n33811;
  assign n33857 = n33812 & ~n33856;
  assign n33858 = n33857 ^ n30585;
  assign n33673 = ~n33671 & n33672;
  assign n33730 = n33673 ^ n33665;
  assign n33731 = ~n33729 & n33730;
  assign n33732 = n33731 ^ n33666;
  assign n33667 = n33665 & ~n33666;
  assign n33675 = n33674 ^ n33673;
  assign n33676 = ~n33667 & ~n33675;
  assign n33799 = n33661 & n33676;
  assign n33800 = ~n33732 & ~n33799;
  assign n33688 = n33293 ^ n33209;
  assign n33684 = n31641 ^ n31517;
  assign n33685 = n32577 ^ n31517;
  assign n33686 = ~n33684 & ~n33685;
  assign n33687 = n33686 ^ n31641;
  assign n33690 = n33688 ^ n33687;
  assign n33806 = n33800 ^ n33690;
  assign n33807 = n33806 ^ n30712;
  assign n33918 = n33858 ^ n33807;
  assign n33901 = n33855 ^ n33812;
  assign n33902 = n33837 ^ n33829;
  assign n33903 = n33834 ^ n33831;
  assign n33449 = n33448 ^ n33437;
  assign n33450 = n33431 ^ n33403;
  assign n33451 = n33425 ^ n33407;
  assign n33452 = n33422 ^ n33409;
  assign n33453 = n33419 ^ n33411;
  assign n33454 = ~n33452 & n33453;
  assign n33455 = n33451 & n33454;
  assign n33456 = n33428 ^ n33405;
  assign n33457 = ~n33455 & ~n33456;
  assign n33458 = n33450 & ~n33457;
  assign n33459 = n33434 ^ n33401;
  assign n33460 = n33458 & n33459;
  assign n33520 = n33449 & ~n33460;
  assign n33535 = n33534 ^ n33523;
  assign n33904 = n33520 & n33535;
  assign n33905 = n33903 & ~n33904;
  assign n33906 = ~n33902 & n33905;
  assign n33907 = n33840 ^ n33822;
  assign n33908 = n33906 & ~n33907;
  assign n33909 = n33843 ^ n33820;
  assign n33910 = n33908 & n33909;
  assign n33911 = n33846 ^ n33818;
  assign n33912 = ~n33910 & ~n33911;
  assign n33913 = n33849 ^ n33816;
  assign n33914 = ~n33912 & ~n33913;
  assign n33915 = n33852 ^ n33814;
  assign n33916 = n33914 & ~n33915;
  assign n33917 = ~n33901 & n33916;
  assign n34013 = n33918 ^ n33917;
  assign n2466 = n2465 ^ n2453;
  assign n2485 = n2484 ^ n2466;
  assign n2492 = n2491 ^ n2485;
  assign n34048 = n34013 ^ n2492;
  assign n34016 = n31358 ^ n3033;
  assign n34017 = n34016 ^ n3146;
  assign n34018 = n34017 ^ n2482;
  assign n34015 = n33916 ^ n33901;
  assign n34049 = n34018 ^ n34015;
  assign n34020 = n33915 ^ n33914;
  assign n34021 = n31364 ^ n2424;
  assign n34022 = n34021 ^ n27724;
  assign n34023 = n34022 ^ n3144;
  assign n34025 = n34020 & n34023;
  assign n34050 = n34025 ^ n34015;
  assign n34051 = n34049 & ~n34050;
  assign n34052 = n34051 ^ n34018;
  assign n33956 = n33913 ^ n33912;
  assign n1281 = n1280 ^ n1193;
  assign n1294 = n1293 ^ n1281;
  assign n1301 = n1300 ^ n1294;
  assign n33957 = n33956 ^ n1301;
  assign n33959 = n31371 ^ n24072;
  assign n33960 = n33959 ^ n1123;
  assign n33961 = n33960 ^ n1288;
  assign n33958 = n33911 ^ n33910;
  assign n33962 = n33961 ^ n33958;
  assign n33963 = n33909 ^ n33908;
  assign n1108 = n1107 ^ n1095;
  assign n1109 = n1108 ^ n1026;
  assign n1116 = n1115 ^ n1109;
  assign n33964 = n33963 ^ n1116;
  assign n33965 = n33907 ^ n33906;
  assign n33966 = n33965 ^ n994;
  assign n33467 = n31394 ^ n23678;
  assign n33468 = n33467 ^ n27747;
  assign n33469 = n33468 ^ n720;
  assign n33466 = n33459 ^ n33458;
  assign n33470 = n33469 ^ n33466;
  assign n33474 = n33457 ^ n33450;
  assign n33471 = n31398 ^ n23683;
  assign n33472 = n33471 ^ n708;
  assign n33473 = n33472 ^ n22856;
  assign n33475 = n33474 ^ n33473;
  assign n33479 = n33456 ^ n33455;
  assign n33476 = n31404 ^ n23688;
  assign n33477 = n33476 ^ n27753;
  assign n33478 = n33477 ^ n548;
  assign n33480 = n33479 ^ n33478;
  assign n33484 = n33454 ^ n33451;
  assign n33481 = n31409 ^ n696;
  assign n33482 = n33481 ^ n27759;
  assign n33483 = n33482 ^ n22842;
  assign n33485 = n33484 ^ n33483;
  assign n33487 = n31421 ^ n23700;
  assign n33488 = n33487 ^ n27763;
  assign n33489 = n33488 ^ n22327;
  assign n33486 = n33453 ^ n33452;
  assign n33490 = n33489 ^ n33486;
  assign n2360 = n2312 ^ n2254;
  assign n2361 = n2360 ^ n2351;
  assign n2362 = n2361 ^ n2359;
  assign n33491 = n33453 ^ n2362;
  assign n33496 = n33495 ^ n2344;
  assign n33497 = n33494 & n33496;
  assign n33498 = n33497 ^ n33493;
  assign n33499 = n33498 ^ n33453;
  assign n33500 = n33491 & ~n33499;
  assign n33501 = n33500 ^ n2362;
  assign n33502 = n33501 ^ n33486;
  assign n33503 = n33490 & ~n33502;
  assign n33504 = n33503 ^ n33489;
  assign n33505 = n33504 ^ n33484;
  assign n33506 = ~n33485 & n33505;
  assign n33507 = n33506 ^ n33483;
  assign n33508 = n33507 ^ n33479;
  assign n33509 = n33480 & ~n33508;
  assign n33510 = n33509 ^ n33478;
  assign n33511 = n33510 ^ n33474;
  assign n33512 = n33475 & ~n33511;
  assign n33513 = n33512 ^ n33473;
  assign n33514 = n33513 ^ n33466;
  assign n33515 = ~n33470 & n33514;
  assign n33516 = n33515 ^ n33469;
  assign n33536 = n33535 ^ n33520;
  assign n33967 = ~n33536 & ~n33539;
  assign n33461 = n33460 ^ n33449;
  assign n33968 = ~n33461 & n33464;
  assign n33465 = n33464 ^ n33461;
  assign n33969 = n33968 ^ n33465;
  assign n33970 = ~n33967 & ~n33969;
  assign n33971 = n33904 ^ n33903;
  assign n33972 = ~n3314 & ~n33971;
  assign n33973 = n33970 & ~n33972;
  assign n968 = n967 ^ n898;
  assign n975 = n974 ^ n968;
  assign n976 = n975 ^ n940;
  assign n33974 = n33905 ^ n33902;
  assign n33975 = ~n976 & ~n33974;
  assign n33976 = n33973 & ~n33975;
  assign n33977 = n33516 & n33976;
  assign n33978 = n33974 ^ n976;
  assign n33979 = n33971 ^ n3314;
  assign n33540 = n33539 ^ n33536;
  assign n33980 = n33540 & ~n33968;
  assign n33981 = n33980 ^ n33967;
  assign n33982 = n33979 & n33981;
  assign n33983 = n33982 ^ n33972;
  assign n33984 = n33983 ^ n33974;
  assign n33985 = n33978 & n33984;
  assign n33986 = n33985 ^ n976;
  assign n33987 = ~n33977 & ~n33986;
  assign n33988 = n33987 ^ n33965;
  assign n33989 = n33966 & n33988;
  assign n33990 = n33989 ^ n994;
  assign n33991 = n33990 ^ n1116;
  assign n33992 = ~n33964 & ~n33991;
  assign n33993 = n33992 ^ n33963;
  assign n33994 = n33993 ^ n33958;
  assign n33995 = n33962 & n33994;
  assign n33996 = n33995 ^ n33961;
  assign n33997 = n33996 ^ n33956;
  assign n33998 = ~n33957 & n33997;
  assign n33999 = n33998 ^ n1301;
  assign n34019 = ~n34015 & ~n34018;
  assign n34024 = n34023 ^ n34020;
  assign n34026 = n34025 ^ n34024;
  assign n34027 = ~n34019 & n34026;
  assign n34354 = n33999 & n34027;
  assign n34355 = ~n34052 & ~n34354;
  assign n34356 = n34355 ^ n34013;
  assign n34357 = ~n34048 & ~n34356;
  assign n34358 = n34357 ^ n2492;
  assign n33919 = ~n33917 & n33918;
  assign n33859 = n33858 ^ n33806;
  assign n33860 = n33807 & n33859;
  assign n33861 = n33860 ^ n30712;
  assign n33801 = n33800 ^ n33688;
  assign n33802 = n33690 & n33801;
  assign n33803 = n33802 ^ n33687;
  assign n33678 = n31639 ^ n31509;
  assign n33679 = n32570 ^ n31509;
  assign n33680 = ~n33678 & ~n33679;
  assign n33681 = n33680 ^ n31639;
  assign n33677 = n33296 ^ n33204;
  assign n33728 = n33681 ^ n33677;
  assign n33804 = n33803 ^ n33728;
  assign n33805 = n33804 ^ n30706;
  assign n33900 = n33861 ^ n33805;
  assign n34028 = n33919 ^ n33900;
  assign n3054 = n3053 ^ n3047;
  assign n3055 = n3054 ^ n2544;
  assign n3059 = n3058 ^ n3055;
  assign n34047 = n34028 ^ n3059;
  assign n34359 = n34358 ^ n34047;
  assign n34350 = n33118 ^ n32549;
  assign n33544 = n33328 ^ n33156;
  assign n33545 = n33544 ^ n33153;
  assign n34351 = n33545 ^ n33118;
  assign n34352 = n34350 & ~n34351;
  assign n34353 = n34352 ^ n32549;
  assign n34360 = n34359 ^ n34353;
  assign n34509 = n34355 ^ n34048;
  assign n34365 = n34020 ^ n33999;
  assign n34366 = n34024 & ~n34365;
  assign n34367 = n34366 ^ n34023;
  assign n34368 = n34367 ^ n34049;
  assign n33555 = ~n33200 & ~n33310;
  assign n33556 = n33316 & ~n33555;
  assign n33557 = ~n33168 & ~n33556;
  assign n33567 = n33557 ^ n33161;
  assign n34361 = n33567 ^ n32524;
  assign n34362 = n32572 ^ n32524;
  assign n34363 = ~n34361 & n34362;
  assign n34364 = n34363 ^ n32572;
  assign n34369 = n34368 ^ n34364;
  assign n34374 = n34024 ^ n33999;
  assign n33573 = n33555 ^ n33164;
  assign n33574 = n33314 & n33573;
  assign n33575 = n33574 ^ n3201;
  assign n33576 = n33575 ^ n33163;
  assign n34370 = n33576 ^ n32536;
  assign n34371 = n32536 ^ n32459;
  assign n34372 = n34370 & n34371;
  assign n34373 = n34372 ^ n32459;
  assign n34375 = n34374 ^ n34373;
  assign n34380 = n33996 ^ n33957;
  assign n33582 = n33555 ^ n33314;
  assign n34376 = n33582 ^ n32542;
  assign n34377 = n32542 ^ n31503;
  assign n34378 = n34376 & n34377;
  assign n34379 = n34378 ^ n31503;
  assign n34381 = n34380 ^ n34379;
  assign n34386 = n33993 ^ n33962;
  assign n33588 = n33302 & n33305;
  assign n33589 = ~n33193 & n33588;
  assign n33590 = n33194 & ~n33589;
  assign n33591 = n33590 ^ n33180;
  assign n33592 = ~n33184 & ~n33591;
  assign n33593 = n33592 ^ n33183;
  assign n33594 = n33593 ^ n33179;
  assign n34382 = n33594 ^ n32556;
  assign n34383 = n32556 ^ n31509;
  assign n34384 = n34382 & ~n34383;
  assign n34385 = n34384 ^ n31509;
  assign n34387 = n34386 ^ n34385;
  assign n33718 = n33590 ^ n33184;
  assign n34389 = n33718 ^ n32558;
  assign n34390 = n32558 ^ n31517;
  assign n34391 = ~n34389 & ~n34390;
  assign n34392 = n34391 ^ n31517;
  assign n34388 = n33990 ^ n33964;
  assign n34393 = n34392 ^ n34388;
  assign n34400 = n33516 & n33970;
  assign n34401 = n33981 & ~n34400;
  assign n34402 = n34401 ^ n33971;
  assign n34403 = n33979 & n34402;
  assign n34404 = n34403 ^ n3314;
  assign n34405 = n34404 ^ n33978;
  assign n33693 = n33304 ^ n33302;
  assign n34396 = n33693 ^ n32577;
  assign n34397 = n32577 ^ n31941;
  assign n34398 = n34396 & ~n34397;
  assign n34399 = n34398 ^ n31941;
  assign n34406 = n34405 ^ n34399;
  assign n34411 = n34401 ^ n33979;
  assign n33703 = n33299 ^ n33202;
  assign n34407 = n33703 ^ n32586;
  assign n34408 = n32586 ^ n31945;
  assign n34409 = n34407 & n34408;
  assign n34410 = n34409 ^ n31945;
  assign n34412 = n34411 ^ n34410;
  assign n34413 = n33677 ^ n32592;
  assign n34414 = n32592 ^ n31935;
  assign n34415 = n34413 & n34414;
  assign n34416 = n34415 ^ n31935;
  assign n33517 = n33516 ^ n33461;
  assign n33518 = ~n33465 & n33517;
  assign n33519 = n33518 ^ n33464;
  assign n33541 = n33540 ^ n33519;
  assign n34417 = n34416 ^ n33541;
  assign n34422 = n33516 ^ n33465;
  assign n34418 = n32598 ^ n31927;
  assign n34419 = n33688 ^ n32598;
  assign n34420 = ~n34418 & n34419;
  assign n34421 = n34420 ^ n31927;
  assign n34423 = n34422 ^ n34421;
  assign n34428 = n33513 ^ n33470;
  assign n34424 = n33666 ^ n32604;
  assign n34425 = n32604 ^ n31919;
  assign n34426 = ~n34424 & n34425;
  assign n34427 = n34426 ^ n31919;
  assign n34429 = n34428 ^ n34427;
  assign n34434 = n33510 ^ n33475;
  assign n34430 = n32610 ^ n31898;
  assign n34431 = n33672 ^ n32610;
  assign n34432 = n34430 & ~n34431;
  assign n34433 = n34432 ^ n31898;
  assign n34435 = n34434 ^ n34433;
  assign n34437 = n32620 ^ n31904;
  assign n34438 = n33600 ^ n32620;
  assign n34439 = n34437 & ~n34438;
  assign n34440 = n34439 ^ n31904;
  assign n34436 = n33507 ^ n33480;
  assign n34441 = n34440 ^ n34436;
  assign n34442 = n33504 ^ n33485;
  assign n34443 = n32622 ^ n31906;
  assign n34444 = n33542 ^ n32622;
  assign n34445 = n34443 & n34444;
  assign n34446 = n34445 ^ n31906;
  assign n34457 = n34442 & n34446;
  assign n34447 = n34446 ^ n34442;
  assign n34449 = n32628 ^ n31541;
  assign n34450 = n33611 ^ n32628;
  assign n34451 = n34449 & ~n34450;
  assign n34452 = n34451 ^ n31541;
  assign n34448 = n33501 ^ n33490;
  assign n34454 = n34452 ^ n34448;
  assign n34453 = ~n34448 & ~n34452;
  assign n34455 = n34454 ^ n34453;
  assign n34456 = n34447 & n34455;
  assign n34458 = n34457 ^ n34456;
  assign n34293 = n32638 ^ n31543;
  assign n34294 = n33617 ^ n32638;
  assign n34295 = ~n34293 & ~n34294;
  assign n34296 = n34295 ^ n31543;
  assign n34292 = n33498 ^ n33491;
  assign n34297 = n34296 ^ n34292;
  assign n34224 = n32640 ^ n31549;
  assign n34225 = n33634 ^ n32640;
  assign n34226 = n34224 & n34225;
  assign n34227 = n34226 ^ n31549;
  assign n34229 = n34228 ^ n34227;
  assign n34196 = n32650 ^ n31555;
  assign n34197 = n33627 ^ n32650;
  assign n34198 = n34196 & ~n34197;
  assign n34199 = n34198 ^ n31555;
  assign n34201 = n34200 ^ n34199;
  assign n34141 = n32506 ^ n31561;
  assign n34142 = n33531 ^ n32506;
  assign n34143 = ~n34141 & ~n34142;
  assign n34144 = n34143 ^ n31561;
  assign n33563 = n31835 ^ n31108;
  assign n33564 = n32433 ^ n31835;
  assign n33565 = n33563 & ~n33564;
  assign n33566 = n33565 ^ n31108;
  assign n33568 = n33567 ^ n33566;
  assign n33569 = n31841 ^ n31125;
  assign n33570 = n33118 ^ n31841;
  assign n33571 = n33569 & ~n33570;
  assign n33572 = n33571 ^ n31125;
  assign n33577 = n33576 ^ n33572;
  assign n33578 = n31847 ^ n31118;
  assign n33579 = n33100 ^ n31847;
  assign n33580 = ~n33578 & ~n33579;
  assign n33581 = n33580 ^ n31118;
  assign n33583 = n33582 ^ n33581;
  assign n33584 = n32549 ^ n31512;
  assign n33585 = n32549 ^ n32524;
  assign n33586 = ~n33584 & n33585;
  assign n33587 = n33586 ^ n31512;
  assign n33595 = n33594 ^ n33587;
  assign n33682 = n33677 & ~n33681;
  assign n33683 = n33676 & ~n33682;
  assign n33689 = n33687 & n33688;
  assign n33691 = n33690 ^ n33689;
  assign n33692 = n33683 & n33691;
  assign n33694 = n32459 ^ n31619;
  assign n33695 = n32556 ^ n32459;
  assign n33696 = n33694 & ~n33695;
  assign n33697 = n33696 ^ n31619;
  assign n33698 = ~n33693 & ~n33697;
  assign n33699 = n31630 ^ n31503;
  assign n33700 = n32558 ^ n31503;
  assign n33701 = ~n33699 & ~n33700;
  assign n33702 = n33701 ^ n31630;
  assign n33705 = ~n33702 & ~n33703;
  assign n33704 = n33703 ^ n33702;
  assign n33706 = n33705 ^ n33704;
  assign n33707 = ~n33698 & n33706;
  assign n33708 = n32572 ^ n31529;
  assign n33709 = n32572 ^ n32542;
  assign n33710 = n33708 & n33709;
  assign n33711 = n33710 ^ n31529;
  assign n33712 = ~n33186 & ~n33588;
  assign n33713 = n33712 ^ n33191;
  assign n33715 = ~n33711 & n33713;
  assign n33714 = n33713 ^ n33711;
  assign n33716 = n33715 ^ n33714;
  assign n33717 = n33707 & ~n33716;
  assign n33719 = n32560 ^ n31522;
  assign n33720 = n32560 ^ n32536;
  assign n33721 = ~n33719 & n33720;
  assign n33722 = n33721 ^ n31522;
  assign n33723 = ~n33718 & ~n33722;
  assign n33724 = n33717 & ~n33723;
  assign n33725 = n33692 & n33724;
  assign n33726 = n33661 & n33725;
  assign n33727 = n33722 ^ n33718;
  assign n33733 = n33690 & n33732;
  assign n33734 = n33733 ^ n33689;
  assign n33735 = n33734 ^ n33677;
  assign n33736 = ~n33728 & n33735;
  assign n33737 = n33736 ^ n33681;
  assign n33738 = n33717 & n33737;
  assign n33739 = n33738 ^ n33722;
  assign n33740 = n33739 ^ n33722;
  assign n33741 = n33697 ^ n33693;
  assign n33742 = n33705 ^ n33697;
  assign n33743 = n33741 & ~n33742;
  assign n33744 = n33743 ^ n33693;
  assign n33745 = ~n33714 & n33744;
  assign n33746 = n33745 ^ n33715;
  assign n33747 = n33746 ^ n33722;
  assign n33748 = n33747 ^ n33722;
  assign n33749 = ~n33740 & ~n33748;
  assign n33750 = n33749 ^ n33722;
  assign n33751 = n33727 & n33750;
  assign n33752 = n33751 ^ n33718;
  assign n33753 = ~n33726 & ~n33752;
  assign n33754 = n33753 ^ n33594;
  assign n33755 = n33595 & ~n33754;
  assign n33756 = n33755 ^ n33587;
  assign n33757 = n33756 ^ n33582;
  assign n33758 = n33583 & ~n33757;
  assign n33759 = n33758 ^ n33581;
  assign n33760 = n33759 ^ n33576;
  assign n33761 = ~n33577 & ~n33760;
  assign n33762 = n33761 ^ n33572;
  assign n33763 = n33762 ^ n33567;
  assign n33764 = ~n33568 & n33763;
  assign n33765 = n33764 ^ n33566;
  assign n33558 = n33557 ^ n33160;
  assign n33559 = n33161 & n33558;
  assign n33560 = n33559 ^ n2737;
  assign n33561 = n33560 ^ n33159;
  assign n33551 = n31825 ^ n31102;
  assign n33552 = n32495 ^ n31825;
  assign n33553 = n33551 & ~n33552;
  assign n33554 = n33553 ^ n31102;
  assign n33562 = n33561 ^ n33554;
  assign n33771 = n33765 ^ n33562;
  assign n33772 = n33771 ^ n30300;
  assign n33773 = n33762 ^ n33568;
  assign n33774 = n33773 ^ n30296;
  assign n33775 = n33759 ^ n33577;
  assign n33776 = n33775 ^ n30291;
  assign n33777 = n33756 ^ n33583;
  assign n33778 = n33777 ^ n30288;
  assign n33779 = n33753 ^ n33595;
  assign n33780 = n33779 ^ n30960;
  assign n33781 = n33661 & n33692;
  assign n33782 = ~n33737 & ~n33781;
  assign n33783 = n33707 & ~n33782;
  assign n33784 = ~n33744 & ~n33783;
  assign n33785 = n33784 ^ n33713;
  assign n33786 = ~n33714 & n33785;
  assign n33787 = n33786 ^ n33711;
  assign n33788 = n33787 ^ n33727;
  assign n33789 = n33788 ^ n30914;
  assign n33790 = n33784 ^ n33714;
  assign n33791 = n33790 ^ n30819;
  assign n33792 = n33782 ^ n33703;
  assign n33793 = n33704 & ~n33792;
  assign n33794 = n33793 ^ n33702;
  assign n33795 = n33794 ^ n33741;
  assign n33796 = n33795 ^ n30699;
  assign n33797 = n33782 ^ n33704;
  assign n33798 = n33797 ^ n30705;
  assign n33862 = n33861 ^ n33804;
  assign n33863 = n33805 & ~n33862;
  assign n33864 = n33863 ^ n30706;
  assign n33865 = n33864 ^ n33797;
  assign n33866 = n33798 & ~n33865;
  assign n33867 = n33866 ^ n30705;
  assign n33868 = n33867 ^ n33795;
  assign n33869 = n33796 & ~n33868;
  assign n33870 = n33869 ^ n30699;
  assign n33871 = n33870 ^ n33790;
  assign n33872 = ~n33791 & n33871;
  assign n33873 = n33872 ^ n30819;
  assign n33874 = n33873 ^ n33788;
  assign n33875 = ~n33789 & ~n33874;
  assign n33876 = n33875 ^ n30914;
  assign n33877 = n33876 ^ n33779;
  assign n33878 = n33780 & n33877;
  assign n33879 = n33878 ^ n30960;
  assign n33880 = n33879 ^ n33777;
  assign n33881 = ~n33778 & ~n33880;
  assign n33882 = n33881 ^ n30288;
  assign n33883 = n33882 ^ n33775;
  assign n33884 = n33776 & ~n33883;
  assign n33885 = n33884 ^ n30291;
  assign n33886 = n33885 ^ n33773;
  assign n33887 = ~n33774 & n33886;
  assign n33888 = n33887 ^ n30296;
  assign n33889 = n33888 ^ n33771;
  assign n33890 = ~n33772 & ~n33889;
  assign n33891 = n33890 ^ n30300;
  assign n33766 = n33765 ^ n33561;
  assign n33767 = n33562 & ~n33766;
  assign n33768 = n33767 ^ n33554;
  assign n33546 = n31823 ^ n31092;
  assign n33547 = n32774 ^ n31823;
  assign n33548 = n33546 & ~n33547;
  assign n33549 = n33548 ^ n31092;
  assign n33550 = n33549 ^ n33545;
  assign n33769 = n33768 ^ n33550;
  assign n33770 = n33769 ^ n30270;
  assign n33892 = n33891 ^ n33770;
  assign n33893 = n33888 ^ n33772;
  assign n33894 = n33882 ^ n33776;
  assign n33895 = n33879 ^ n33778;
  assign n33896 = n33876 ^ n33780;
  assign n33897 = n33873 ^ n33789;
  assign n33898 = n33867 ^ n33796;
  assign n33899 = n33864 ^ n33798;
  assign n33920 = n33900 & ~n33919;
  assign n33921 = n33899 & n33920;
  assign n33922 = ~n33898 & ~n33921;
  assign n33923 = n33870 ^ n33791;
  assign n33924 = n33922 & n33923;
  assign n33925 = n33897 & n33924;
  assign n33926 = ~n33896 & ~n33925;
  assign n33927 = ~n33895 & n33926;
  assign n33928 = ~n33894 & n33927;
  assign n33929 = n33885 ^ n33774;
  assign n33930 = n33928 & n33929;
  assign n33931 = ~n33893 & ~n33930;
  assign n34102 = ~n33892 & n33931;
  assign n34098 = n33891 ^ n33769;
  assign n34099 = n33770 & ~n34098;
  assign n34100 = n34099 ^ n30270;
  assign n34091 = n31602 ^ n30693;
  assign n34092 = n32768 ^ n31602;
  assign n34093 = ~n34091 & ~n34092;
  assign n34094 = n34093 ^ n30693;
  assign n34090 = n33331 ^ n33152;
  assign n34095 = n34094 ^ n34090;
  assign n34087 = n33768 ^ n33545;
  assign n34088 = ~n33550 & ~n34087;
  assign n34089 = n34088 ^ n33549;
  assign n34096 = n34095 ^ n34089;
  assign n34097 = n34096 ^ n30312;
  assign n34101 = n34100 ^ n34097;
  assign n34103 = n34102 ^ n34101;
  assign n34107 = n34106 ^ n34103;
  assign n33932 = n33931 ^ n33892;
  assign n33936 = n33935 ^ n33932;
  assign n33938 = n31783 ^ n22801;
  assign n33939 = n33938 ^ n1731;
  assign n33940 = n33939 ^ n24121;
  assign n33937 = n33930 ^ n33893;
  assign n33941 = n33940 ^ n33937;
  assign n33945 = n33929 ^ n33928;
  assign n33942 = n31788 ^ n24019;
  assign n33943 = n33942 ^ n28161;
  assign n33944 = n33943 ^ n1729;
  assign n33946 = n33945 ^ n33944;
  assign n33947 = n33927 ^ n33894;
  assign n1629 = n1628 ^ n1613;
  assign n1648 = n1647 ^ n1629;
  assign n1655 = n1654 ^ n1648;
  assign n33948 = n33947 ^ n1655;
  assign n33952 = n33926 ^ n33895;
  assign n33949 = n24026 ^ n2962;
  assign n33950 = n33949 ^ n2937;
  assign n33951 = n33950 ^ n1642;
  assign n33953 = n33952 ^ n33951;
  assign n33954 = n33925 ^ n33896;
  assign n2928 = n2927 ^ n2861;
  assign n2929 = n2928 ^ n2921;
  assign n2930 = n2929 ^ n1538;
  assign n33955 = n33954 ^ n2930;
  assign n34003 = n33921 ^ n33898;
  assign n34004 = ~n34002 & ~n34003;
  assign n34008 = n33920 ^ n33899;
  assign n34005 = n31350 ^ n2546;
  assign n34006 = n34005 ^ n3209;
  assign n34007 = n34006 ^ n3074;
  assign n34010 = n34008 ^ n34007;
  assign n34009 = n34007 & ~n34008;
  assign n34011 = n34010 ^ n34009;
  assign n34012 = ~n34004 & ~n34011;
  assign n34014 = ~n2492 & n34013;
  assign n34029 = ~n3059 & ~n34028;
  assign n34030 = n34027 & ~n34029;
  assign n34031 = ~n34014 & n34030;
  assign n34032 = n33924 ^ n33897;
  assign n34033 = ~n2914 & ~n34032;
  assign n3230 = n3223 ^ n2787;
  assign n3234 = n3233 ^ n3230;
  assign n3235 = n3234 ^ n2908;
  assign n34034 = n33923 ^ n33922;
  assign n34036 = n3235 & n34034;
  assign n34035 = n34034 ^ n3235;
  assign n34037 = n34036 ^ n34035;
  assign n34038 = ~n34033 & n34037;
  assign n34039 = n34031 & n34038;
  assign n34040 = n34012 & n34039;
  assign n34041 = n33999 & n34040;
  assign n34042 = n34032 ^ n2914;
  assign n34043 = n34003 ^ n34002;
  assign n34044 = n34009 ^ n34003;
  assign n34045 = n34043 & ~n34044;
  assign n34046 = n34045 ^ n34002;
  assign n34053 = n34052 ^ n2492;
  assign n34054 = ~n34048 & n34053;
  assign n34055 = n34054 ^ n2492;
  assign n34056 = n34047 & n34055;
  assign n34057 = n34056 ^ n34047;
  assign n34058 = n34057 ^ n34029;
  assign n34059 = n34012 & ~n34058;
  assign n34060 = ~n34036 & ~n34059;
  assign n34061 = ~n34046 & n34060;
  assign n34062 = n34061 ^ n34032;
  assign n34063 = n34062 ^ n34032;
  assign n34064 = n34037 & ~n34063;
  assign n34065 = n34064 ^ n34032;
  assign n34066 = n34042 & ~n34065;
  assign n34067 = n34066 ^ n2914;
  assign n34068 = ~n34041 & ~n34067;
  assign n34069 = n34068 ^ n33954;
  assign n34070 = ~n33955 & ~n34069;
  assign n34071 = n34070 ^ n2930;
  assign n34072 = n34071 ^ n33951;
  assign n34073 = n33953 & ~n34072;
  assign n34074 = n34073 ^ n33952;
  assign n34075 = n34074 ^ n33947;
  assign n34076 = n33948 & ~n34075;
  assign n34077 = n34076 ^ n1655;
  assign n34078 = n34077 ^ n33945;
  assign n34079 = ~n33946 & n34078;
  assign n34080 = n34079 ^ n33944;
  assign n34081 = n34080 ^ n33937;
  assign n34082 = n33941 & ~n34081;
  assign n34083 = n34082 ^ n33940;
  assign n34084 = n34083 ^ n33932;
  assign n34085 = ~n33936 & n34084;
  assign n34086 = n34085 ^ n33935;
  assign n34164 = n34103 ^ n34086;
  assign n34165 = ~n34107 & n34164;
  assign n34166 = n34165 ^ n34106;
  assign n34157 = n34100 ^ n30312;
  assign n34158 = n34100 ^ n34096;
  assign n34159 = n34157 & ~n34158;
  assign n34160 = n34159 ^ n30312;
  assign n34150 = n31596 ^ n30687;
  assign n34151 = n32762 ^ n31596;
  assign n34152 = n34150 & ~n34151;
  assign n34153 = n34152 ^ n30687;
  assign n34149 = n33334 ^ n33150;
  assign n34154 = n34153 ^ n34149;
  assign n34146 = n34090 ^ n34089;
  assign n34147 = n34095 & n34146;
  assign n34148 = n34147 ^ n34094;
  assign n34155 = n34154 ^ n34148;
  assign n34156 = n34155 ^ n30321;
  assign n34161 = n34160 ^ n34156;
  assign n34145 = ~n34101 & n34102;
  assign n34162 = n34161 ^ n34145;
  assign n34163 = n34162 ^ n2182;
  assign n34167 = n34166 ^ n34163;
  assign n34193 = n34144 & ~n34167;
  assign n34168 = n34167 ^ n34144;
  assign n34194 = n34193 ^ n34168;
  assign n34215 = n34200 ^ n34194;
  assign n34216 = n34215 ^ n34199;
  assign n34109 = n32513 ^ n31567;
  assign n34110 = n33442 ^ n32513;
  assign n34111 = ~n34109 & n34110;
  assign n34112 = n34111 ^ n31567;
  assign n34108 = n34107 ^ n34086;
  assign n34113 = n34112 ^ n34108;
  assign n34115 = n32519 ^ n31573;
  assign n34116 = n33398 ^ n32519;
  assign n34117 = n34115 & n34116;
  assign n34118 = n34117 ^ n31573;
  assign n34114 = n34083 ^ n33936;
  assign n34119 = n34118 ^ n34114;
  assign n34121 = n32663 ^ n31583;
  assign n34122 = n32663 ^ n32504;
  assign n34123 = ~n34121 & ~n34122;
  assign n34124 = n34123 ^ n31583;
  assign n34120 = n34080 ^ n33941;
  assign n34125 = n34124 ^ n34120;
  assign n34126 = n32679 ^ n31586;
  assign n34127 = n32679 ^ n32511;
  assign n34128 = n34126 & ~n34127;
  assign n34129 = n34128 ^ n31586;
  assign n34130 = n34077 ^ n33946;
  assign n34131 = n34129 & ~n34130;
  assign n34132 = n34131 ^ n34120;
  assign n34133 = n34125 & n34132;
  assign n34134 = n34133 ^ n34131;
  assign n34135 = n34134 ^ n34118;
  assign n34136 = n34119 & n34135;
  assign n34137 = n34136 ^ n34114;
  assign n34138 = n34137 ^ n34112;
  assign n34139 = ~n34113 & n34138;
  assign n34140 = n34139 ^ n34108;
  assign n34217 = ~n34140 & ~n34193;
  assign n34218 = n34217 ^ n34199;
  assign n34219 = n34218 ^ n34199;
  assign n34220 = n34216 & ~n34219;
  assign n34221 = n34220 ^ n34199;
  assign n34222 = n34201 & n34221;
  assign n34223 = n34222 ^ n34200;
  assign n34289 = n34228 ^ n34223;
  assign n34290 = ~n34229 & n34289;
  assign n34291 = n34290 ^ n34227;
  assign n34459 = n34296 ^ n34291;
  assign n34460 = n34297 & ~n34459;
  assign n34461 = n34460 ^ n34292;
  assign n34462 = ~n34453 & ~n34457;
  assign n34463 = n34461 & n34462;
  assign n34464 = n34458 & ~n34463;
  assign n34465 = n34464 ^ n34440;
  assign n34466 = n34441 & n34465;
  assign n34467 = n34466 ^ n34436;
  assign n34468 = n34467 ^ n34434;
  assign n34469 = n34435 & ~n34468;
  assign n34470 = n34469 ^ n34433;
  assign n34471 = n34470 ^ n34428;
  assign n34472 = n34429 & ~n34471;
  assign n34473 = n34472 ^ n34470;
  assign n34474 = n34473 ^ n34421;
  assign n34475 = ~n34423 & ~n34474;
  assign n34476 = n34475 ^ n34422;
  assign n34477 = n34476 ^ n33541;
  assign n34478 = n34417 & n34477;
  assign n34479 = n34478 ^ n34416;
  assign n34480 = n34479 ^ n34411;
  assign n34481 = ~n34412 & n34480;
  assign n34482 = n34481 ^ n34410;
  assign n34483 = n34482 ^ n34405;
  assign n34484 = n34406 & ~n34483;
  assign n34485 = n34484 ^ n34399;
  assign n34394 = n33987 ^ n994;
  assign n34395 = n34394 ^ n33965;
  assign n34486 = n34485 ^ n34395;
  assign n34487 = n33713 ^ n32570;
  assign n34488 = n32570 ^ n31527;
  assign n34489 = n34487 & ~n34488;
  assign n34490 = n34489 ^ n31527;
  assign n34491 = n34490 ^ n34395;
  assign n34492 = n34486 & ~n34491;
  assign n34493 = n34492 ^ n34490;
  assign n34494 = n34493 ^ n34388;
  assign n34495 = n34393 & n34494;
  assign n34496 = n34495 ^ n34392;
  assign n34497 = n34496 ^ n34386;
  assign n34498 = n34387 & ~n34497;
  assign n34499 = n34498 ^ n34385;
  assign n34500 = n34499 ^ n34380;
  assign n34501 = ~n34381 & ~n34500;
  assign n34502 = n34501 ^ n34379;
  assign n34503 = n34502 ^ n34374;
  assign n34504 = n34375 & ~n34503;
  assign n34505 = n34504 ^ n34373;
  assign n34506 = n34505 ^ n34368;
  assign n34507 = ~n34369 & ~n34506;
  assign n34508 = n34507 ^ n34364;
  assign n34510 = n34509 ^ n34508;
  assign n34511 = n33561 ^ n33100;
  assign n34512 = n33100 ^ n32560;
  assign n34513 = ~n34511 & ~n34512;
  assign n34514 = n34513 ^ n32560;
  assign n34515 = n34514 ^ n34509;
  assign n34516 = n34510 & ~n34515;
  assign n34517 = n34516 ^ n34514;
  assign n34518 = n34517 ^ n34359;
  assign n34519 = n34360 & n34518;
  assign n34520 = n34519 ^ n34353;
  assign n34316 = n33999 & n34031;
  assign n34317 = n34058 & ~n34316;
  assign n34348 = n34317 ^ n34010;
  assign n34344 = n32433 ^ n31847;
  assign n34345 = n34090 ^ n32433;
  assign n34346 = n34344 & ~n34345;
  assign n34347 = n34346 ^ n31847;
  assign n34349 = n34348 ^ n34347;
  assign n34542 = n34520 ^ n34349;
  assign n34543 = n34542 ^ n31118;
  assign n34544 = n34517 ^ n34360;
  assign n34545 = n34544 ^ n31512;
  assign n34546 = n34514 ^ n34510;
  assign n34547 = n34546 ^ n31522;
  assign n34548 = n34505 ^ n34364;
  assign n34549 = n34548 ^ n34368;
  assign n34550 = n34549 ^ n31529;
  assign n34551 = n34502 ^ n34375;
  assign n34552 = n34551 ^ n31619;
  assign n34553 = n34499 ^ n34381;
  assign n34554 = n34553 ^ n31630;
  assign n34555 = n34496 ^ n34387;
  assign n34556 = n34555 ^ n31639;
  assign n34557 = n34493 ^ n34393;
  assign n34558 = n34557 ^ n31641;
  assign n34559 = n34490 ^ n34486;
  assign n34560 = n34559 ^ n31653;
  assign n34561 = n34482 ^ n34399;
  assign n34562 = n34561 ^ n34405;
  assign n34563 = n34562 ^ n31659;
  assign n34564 = n34479 ^ n34410;
  assign n34565 = n34564 ^ n34411;
  assign n34566 = n34565 ^ n31491;
  assign n34567 = n34476 ^ n34417;
  assign n34568 = n34567 ^ n31294;
  assign n34569 = n34473 ^ n34423;
  assign n34570 = n34569 ^ n31187;
  assign n34571 = n34470 ^ n34429;
  assign n34572 = n34571 ^ n30583;
  assign n34573 = n34467 ^ n34435;
  assign n34574 = n34573 ^ n30594;
  assign n34575 = n34464 ^ n34441;
  assign n34576 = n34575 ^ n30601;
  assign n34577 = n34461 ^ n34452;
  assign n34578 = n34454 & ~n34577;
  assign n34579 = n34578 ^ n34448;
  assign n34580 = n34579 ^ n34447;
  assign n34581 = n34580 ^ n30614;
  assign n34582 = n34461 ^ n34454;
  assign n34583 = n34582 ^ n30621;
  assign n34230 = n34229 ^ n34223;
  assign n34231 = n34230 ^ n30639;
  assign n34192 = ~n34140 & ~n34168;
  assign n34195 = n34194 ^ n34192;
  assign n34202 = n34201 ^ n34195;
  assign n34203 = n34202 ^ n30651;
  assign n34169 = n34168 ^ n34140;
  assign n34170 = n34169 ^ n30653;
  assign n34171 = n34137 ^ n34113;
  assign n34172 = n34171 ^ n30666;
  assign n34173 = n34134 ^ n34119;
  assign n34174 = n34173 ^ n30672;
  assign n34175 = n34130 ^ n34129;
  assign n34176 = ~n30685 & ~n34175;
  assign n34177 = n34176 ^ n30678;
  assign n34178 = n34131 ^ n34124;
  assign n34179 = n34178 ^ n34120;
  assign n34180 = n34179 ^ n34176;
  assign n34181 = ~n34177 & n34180;
  assign n34182 = n34181 ^ n30678;
  assign n34183 = n34182 ^ n34173;
  assign n34184 = ~n34174 & n34183;
  assign n34185 = n34184 ^ n30672;
  assign n34186 = n34185 ^ n34171;
  assign n34187 = n34172 & n34186;
  assign n34188 = n34187 ^ n30666;
  assign n34189 = n34188 ^ n34169;
  assign n34190 = n34170 & ~n34189;
  assign n34191 = n34190 ^ n30653;
  assign n34212 = n34202 ^ n34191;
  assign n34213 = n34203 & ~n34212;
  assign n34214 = n34213 ^ n30651;
  assign n34299 = n34230 ^ n34214;
  assign n34300 = n34231 & n34299;
  assign n34301 = n34300 ^ n30639;
  assign n34298 = n34297 ^ n34291;
  assign n34302 = n34301 ^ n34298;
  assign n34584 = n34298 ^ n30632;
  assign n34585 = n34302 & n34584;
  assign n34586 = n34585 ^ n30632;
  assign n34587 = n34586 ^ n34582;
  assign n34588 = n34583 & ~n34587;
  assign n34589 = n34588 ^ n30621;
  assign n34590 = n34589 ^ n34580;
  assign n34591 = n34581 & ~n34590;
  assign n34592 = n34591 ^ n30614;
  assign n34593 = n34592 ^ n34575;
  assign n34594 = ~n34576 & n34593;
  assign n34595 = n34594 ^ n30601;
  assign n34596 = n34595 ^ n34573;
  assign n34597 = n34574 & ~n34596;
  assign n34598 = n34597 ^ n30594;
  assign n34599 = n34598 ^ n34571;
  assign n34600 = ~n34572 & n34599;
  assign n34601 = n34600 ^ n30583;
  assign n34602 = n34601 ^ n34569;
  assign n34603 = ~n34570 & n34602;
  assign n34604 = n34603 ^ n31187;
  assign n34605 = n34604 ^ n34567;
  assign n34606 = ~n34568 & n34605;
  assign n34607 = n34606 ^ n31294;
  assign n34608 = n34607 ^ n34565;
  assign n34609 = ~n34566 & n34608;
  assign n34610 = n34609 ^ n31491;
  assign n34611 = n34610 ^ n34562;
  assign n34612 = ~n34563 & ~n34611;
  assign n34613 = n34612 ^ n31659;
  assign n34614 = n34613 ^ n34559;
  assign n34615 = n34560 & ~n34614;
  assign n34616 = n34615 ^ n31653;
  assign n34617 = n34616 ^ n34557;
  assign n34618 = n34558 & n34617;
  assign n34619 = n34618 ^ n31641;
  assign n34620 = n34619 ^ n34555;
  assign n34621 = ~n34556 & n34620;
  assign n34622 = n34621 ^ n31639;
  assign n34623 = n34622 ^ n34553;
  assign n34624 = ~n34554 & ~n34623;
  assign n34625 = n34624 ^ n31630;
  assign n34626 = n34625 ^ n34551;
  assign n34627 = n34552 & n34626;
  assign n34628 = n34627 ^ n31619;
  assign n34629 = n34628 ^ n34549;
  assign n34630 = n34550 & n34629;
  assign n34631 = n34630 ^ n31529;
  assign n34632 = n34631 ^ n34546;
  assign n34633 = n34547 & n34632;
  assign n34634 = n34633 ^ n31522;
  assign n34635 = n34634 ^ n34544;
  assign n34636 = n34545 & n34635;
  assign n34637 = n34636 ^ n31512;
  assign n34638 = n34637 ^ n34542;
  assign n34639 = ~n34543 & n34638;
  assign n34640 = n34639 ^ n31118;
  assign n34521 = n34520 ^ n34348;
  assign n34522 = n34349 & ~n34521;
  assign n34523 = n34522 ^ n34347;
  assign n34339 = n34317 ^ n34008;
  assign n34340 = ~n34010 & ~n34339;
  assign n34341 = n34340 ^ n34007;
  assign n34342 = n34341 ^ n34043;
  assign n34335 = n32495 ^ n31841;
  assign n34336 = n34149 ^ n32495;
  assign n34337 = n34335 & ~n34336;
  assign n34338 = n34337 ^ n31841;
  assign n34343 = n34342 ^ n34338;
  assign n34540 = n34523 ^ n34343;
  assign n34541 = n34540 ^ n31125;
  assign n34701 = n34640 ^ n34541;
  assign n34654 = n34637 ^ n31118;
  assign n34655 = n34654 ^ n34542;
  assign n34656 = n34625 ^ n31619;
  assign n34657 = n34656 ^ n34551;
  assign n34658 = n34616 ^ n34558;
  assign n34659 = n34613 ^ n31653;
  assign n34660 = n34659 ^ n34559;
  assign n34661 = n34610 ^ n34563;
  assign n34662 = n34604 ^ n31294;
  assign n34663 = n34662 ^ n34567;
  assign n34664 = n34595 ^ n30594;
  assign n34665 = n34664 ^ n34573;
  assign n34666 = n34589 ^ n30614;
  assign n34667 = n34666 ^ n34580;
  assign n34303 = n34302 ^ n30632;
  assign n34204 = n34203 ^ n34191;
  assign n34205 = n34182 ^ n34174;
  assign n34206 = n34185 ^ n34172;
  assign n34207 = ~n34205 & n34206;
  assign n34208 = n34188 ^ n30653;
  assign n34209 = n34208 ^ n34169;
  assign n34210 = n34207 & ~n34209;
  assign n34211 = n34204 & ~n34210;
  assign n34232 = n34231 ^ n34214;
  assign n34304 = ~n34211 & ~n34232;
  assign n34668 = n34303 & n34304;
  assign n34669 = n34586 ^ n34583;
  assign n34670 = ~n34668 & n34669;
  assign n34671 = n34667 & n34670;
  assign n34672 = n34592 ^ n34576;
  assign n34673 = ~n34671 & n34672;
  assign n34674 = ~n34665 & n34673;
  assign n34675 = n34598 ^ n34572;
  assign n34676 = n34674 & n34675;
  assign n34677 = n34601 ^ n31187;
  assign n34678 = n34677 ^ n34569;
  assign n34679 = n34676 & n34678;
  assign n34680 = ~n34663 & ~n34679;
  assign n34681 = n34607 ^ n31491;
  assign n34682 = n34681 ^ n34565;
  assign n34683 = ~n34680 & n34682;
  assign n34684 = n34661 & n34683;
  assign n34685 = n34660 & n34684;
  assign n34686 = ~n34658 & ~n34685;
  assign n34687 = n34619 ^ n31639;
  assign n34688 = n34687 ^ n34555;
  assign n34689 = ~n34686 & n34688;
  assign n34690 = n34622 ^ n34554;
  assign n34691 = n34689 & n34690;
  assign n34692 = ~n34657 & ~n34691;
  assign n34693 = n34628 ^ n34550;
  assign n34694 = n34692 & n34693;
  assign n34695 = n34631 ^ n31522;
  assign n34696 = n34695 ^ n34546;
  assign n34697 = n34694 & ~n34696;
  assign n34698 = n34634 ^ n34545;
  assign n34699 = ~n34697 & ~n34698;
  assign n34700 = ~n34655 & n34699;
  assign n34713 = n34701 ^ n34700;
  assign n34717 = n34716 ^ n34713;
  assign n34718 = n34699 ^ n34655;
  assign n34722 = n34721 ^ n34718;
  assign n34723 = n34698 ^ n34697;
  assign n34727 = n34726 ^ n34723;
  assign n34728 = n34696 ^ n34694;
  assign n34729 = n34728 ^ n3113;
  assign n34730 = n34693 ^ n34692;
  assign n2694 = n2693 ^ n2645;
  assign n2701 = n2700 ^ n2694;
  assign n2702 = n2701 ^ n1574;
  assign n34731 = n34730 ^ n2702;
  assign n34732 = n34691 ^ n34657;
  assign n3091 = n3086 ^ n3081;
  assign n3092 = n3091 ^ n2623;
  assign n3093 = n3092 ^ n2698;
  assign n34733 = n34732 ^ n3093;
  assign n34734 = n34690 ^ n34689;
  assign n2602 = n2601 ^ n2565;
  assign n2615 = n2614 ^ n2602;
  assign n2616 = n2615 ^ n2586;
  assign n34735 = n34734 ^ n2616;
  assign n34736 = n34688 ^ n34686;
  assign n3168 = n3167 ^ n2530;
  assign n3178 = n3177 ^ n3168;
  assign n3179 = n3178 ^ n2612;
  assign n34737 = n34736 ^ n3179;
  assign n34739 = n32380 ^ n2518;
  assign n34740 = n34739 ^ n28583;
  assign n34741 = n34740 ^ n3175;
  assign n34738 = n34685 ^ n34658;
  assign n34742 = n34741 ^ n34738;
  assign n34744 = n32386 ^ n3153;
  assign n34745 = n34744 ^ n28588;
  assign n34746 = n34745 ^ n23486;
  assign n34743 = n34684 ^ n34660;
  assign n34747 = n34746 ^ n34743;
  assign n34749 = n34682 ^ n34680;
  assign n1412 = n1396 ^ n1309;
  assign n1413 = n1412 ^ n1263;
  assign n1420 = n1419 ^ n1413;
  assign n34750 = n34749 ^ n1420;
  assign n34751 = n34679 ^ n34663;
  assign n1248 = n1245 ^ n1157;
  assign n1249 = n1248 ^ n1208;
  assign n1253 = n1252 ^ n1249;
  assign n34752 = n34751 ^ n1253;
  assign n34753 = n34678 ^ n34676;
  assign n1221 = n1149 ^ n1077;
  assign n1231 = n1230 ^ n1221;
  assign n1238 = n1237 ^ n1231;
  assign n34754 = n34753 ^ n1238;
  assign n34755 = n34675 ^ n34674;
  assign n3334 = n3330 ^ n1059;
  assign n3338 = n3337 ^ n3334;
  assign n3339 = n3338 ^ n1228;
  assign n34756 = n34755 ^ n3339;
  assign n34757 = n34673 ^ n34665;
  assign n34761 = n34760 ^ n34757;
  assign n34762 = n34672 ^ n34671;
  assign n34766 = n34765 ^ n34762;
  assign n34770 = n34670 ^ n34667;
  assign n34767 = n32301 ^ n24769;
  assign n34768 = n34767 ^ n28604;
  assign n34769 = n34768 ^ n756;
  assign n34771 = n34770 ^ n34769;
  assign n34772 = n34669 ^ n34668;
  assign n730 = n729 ^ n723;
  assign n731 = n730 ^ n605;
  assign n732 = n731 ^ n659;
  assign n34773 = n34772 ^ n732;
  assign n34305 = n34304 ^ n34303;
  assign n34285 = n32308 ^ n24741;
  assign n34286 = n34285 ^ n28611;
  assign n34287 = n34286 ^ n600;
  assign n34774 = n34305 ^ n34287;
  assign n34234 = n32313 ^ n563;
  assign n34235 = n34234 ^ n28616;
  assign n34236 = n34235 ^ n3287;
  assign n34233 = n34232 ^ n34211;
  assign n34237 = n34236 ^ n34233;
  assign n34238 = n34210 ^ n34204;
  assign n34242 = n34241 ^ n34238;
  assign n34244 = n28621 ^ n24243;
  assign n34245 = n34244 ^ n32324;
  assign n34246 = n34245 ^ n23082;
  assign n34243 = n34209 ^ n34207;
  assign n34247 = n34246 ^ n34243;
  assign n34251 = n34206 ^ n34205;
  assign n34248 = n24202 ^ n2406;
  assign n34249 = n34248 ^ n28639;
  assign n34250 = n34249 ^ n23097;
  assign n34252 = n34251 ^ n34250;
  assign n34253 = n24193 ^ n2388;
  assign n34254 = n34253 ^ n28625;
  assign n34255 = n34254 ^ n23088;
  assign n34256 = n34255 ^ n34205;
  assign n34262 = n2380 ^ n2287;
  assign n34263 = n34262 ^ n28628;
  assign n34264 = n34263 ^ n2228;
  assign n34257 = n32743 ^ n2272;
  assign n34258 = n34257 ^ n2045;
  assign n34259 = n34258 ^ n23152;
  assign n34260 = n34175 ^ n30685;
  assign n34261 = n34259 & n34260;
  assign n34265 = n34264 ^ n34261;
  assign n34266 = n34179 ^ n34177;
  assign n34267 = n34266 ^ n34264;
  assign n34268 = n34265 & ~n34267;
  assign n34269 = n34268 ^ n34261;
  assign n34270 = n34269 ^ n34205;
  assign n34271 = ~n34256 & n34270;
  assign n34272 = n34271 ^ n34255;
  assign n34273 = n34272 ^ n34251;
  assign n34274 = n34252 & ~n34273;
  assign n34275 = n34274 ^ n34250;
  assign n34276 = n34275 ^ n34243;
  assign n34277 = n34247 & ~n34276;
  assign n34278 = n34277 ^ n34246;
  assign n34279 = n34278 ^ n34238;
  assign n34280 = ~n34242 & n34279;
  assign n34281 = n34280 ^ n34241;
  assign n34282 = n34281 ^ n34233;
  assign n34283 = ~n34237 & n34282;
  assign n34284 = n34283 ^ n34236;
  assign n34775 = n34305 ^ n34284;
  assign n34776 = ~n34774 & n34775;
  assign n34777 = n34776 ^ n34287;
  assign n34778 = n34777 ^ n34772;
  assign n34779 = ~n34773 & n34778;
  assign n34780 = n34779 ^ n732;
  assign n34781 = n34780 ^ n34770;
  assign n34782 = n34771 & ~n34781;
  assign n34783 = n34782 ^ n34769;
  assign n34784 = n34783 ^ n34762;
  assign n34785 = n34766 & ~n34784;
  assign n34786 = n34785 ^ n34765;
  assign n34787 = n34786 ^ n34757;
  assign n34788 = n34761 & ~n34787;
  assign n34789 = n34788 ^ n34760;
  assign n34790 = n34789 ^ n34755;
  assign n34791 = ~n34756 & n34790;
  assign n34792 = n34791 ^ n3339;
  assign n34793 = n34792 ^ n34753;
  assign n34794 = ~n34754 & n34793;
  assign n34795 = n34794 ^ n1238;
  assign n34796 = n34795 ^ n34751;
  assign n34797 = n34752 & ~n34796;
  assign n34798 = n34797 ^ n1253;
  assign n34799 = n34798 ^ n34749;
  assign n34800 = n34750 & ~n34799;
  assign n34801 = n34800 ^ n1420;
  assign n34748 = n34683 ^ n34661;
  assign n34802 = n34801 ^ n34748;
  assign n1436 = n1435 ^ n1324;
  assign n1437 = n1436 ^ n1427;
  assign n1438 = n1437 ^ n1408;
  assign n34803 = n34748 ^ n1438;
  assign n34804 = n34802 & ~n34803;
  assign n34805 = n34804 ^ n1438;
  assign n34806 = n34805 ^ n34743;
  assign n34807 = ~n34747 & n34806;
  assign n34808 = n34807 ^ n34746;
  assign n34809 = n34808 ^ n34738;
  assign n34810 = n34742 & ~n34809;
  assign n34811 = n34810 ^ n34741;
  assign n34812 = n34811 ^ n34736;
  assign n34813 = n34737 & ~n34812;
  assign n34814 = n34813 ^ n3179;
  assign n34815 = n34814 ^ n34734;
  assign n34816 = ~n34735 & n34815;
  assign n34817 = n34816 ^ n2616;
  assign n34818 = n34817 ^ n34732;
  assign n34819 = n34733 & ~n34818;
  assign n34820 = n34819 ^ n3093;
  assign n34821 = n34820 ^ n34730;
  assign n34822 = n34731 & ~n34821;
  assign n34823 = n34822 ^ n2702;
  assign n34824 = n34823 ^ n34728;
  assign n34825 = ~n34729 & n34824;
  assign n34826 = n34825 ^ n3113;
  assign n34827 = n34826 ^ n34723;
  assign n34828 = ~n34727 & n34827;
  assign n34829 = n34828 ^ n34726;
  assign n34830 = n34829 ^ n34718;
  assign n34831 = n34722 & ~n34830;
  assign n34832 = n34831 ^ n34721;
  assign n34833 = n34832 ^ n34713;
  assign n34834 = ~n34717 & n34833;
  assign n34835 = n34834 ^ n34716;
  assign n34702 = n34700 & n34701;
  assign n34641 = n34640 ^ n34540;
  assign n34642 = n34541 & n34641;
  assign n34643 = n34642 ^ n31125;
  assign n34652 = n34643 ^ n31108;
  assign n34524 = n34523 ^ n34342;
  assign n34525 = n34343 & ~n34524;
  assign n34526 = n34525 ^ n34338;
  assign n34318 = n34012 & ~n34317;
  assign n34319 = ~n34046 & ~n34318;
  assign n34333 = n34319 ^ n34035;
  assign n34329 = n32774 ^ n31835;
  assign n34330 = n33370 ^ n32774;
  assign n34331 = ~n34329 & n34330;
  assign n34332 = n34331 ^ n31835;
  assign n34334 = n34333 ^ n34332;
  assign n34538 = n34526 ^ n34334;
  assign n34653 = n34652 ^ n34538;
  assign n34712 = n34702 ^ n34653;
  assign n34836 = n34835 ^ n34712;
  assign n34857 = n34839 ^ n34836;
  assign n34858 = n34856 & ~n34857;
  assign n34863 = n34862 ^ n34858;
  assign n34840 = n34839 ^ n34712;
  assign n34841 = n34836 & ~n34840;
  assign n34842 = n34841 ^ n34839;
  assign n34539 = n34538 ^ n31108;
  assign n34644 = n34643 ^ n34538;
  assign n34645 = ~n34539 & n34644;
  assign n34646 = n34645 ^ n31108;
  assign n34527 = n34526 ^ n34333;
  assign n34528 = ~n34334 & n34527;
  assign n34529 = n34528 ^ n34332;
  assign n34324 = n32768 ^ n31825;
  assign n34325 = n33368 ^ n32768;
  assign n34326 = ~n34324 & ~n34325;
  assign n34327 = n34326 ^ n31825;
  assign n34535 = n34529 ^ n34327;
  assign n34320 = n34319 ^ n34034;
  assign n34321 = n34035 & n34320;
  assign n34322 = n34321 ^ n3235;
  assign n34323 = n34322 ^ n34042;
  assign n34536 = n34535 ^ n34323;
  assign n34537 = n34536 ^ n31102;
  assign n34704 = n34646 ^ n34537;
  assign n34703 = n34653 & n34702;
  assign n34710 = n34704 ^ n34703;
  assign n1768 = n1761 ^ n1744;
  assign n1787 = n1786 ^ n1768;
  assign n1794 = n1793 ^ n1787;
  assign n34711 = n34710 ^ n1794;
  assign n34864 = n34842 ^ n34711;
  assign n34865 = n34864 ^ n34862;
  assign n34866 = n34863 & n34865;
  assign n34867 = n34866 ^ n34858;
  assign n34848 = n33531 ^ n32519;
  assign n34849 = n34292 ^ n33531;
  assign n34850 = ~n34848 & ~n34849;
  assign n34851 = n34850 ^ n32519;
  assign n34843 = n34842 ^ n34710;
  assign n34844 = ~n34711 & n34843;
  assign n34845 = n34844 ^ n1794;
  assign n34707 = n32485 ^ n24699;
  assign n34708 = n34707 ^ n1801;
  assign n34709 = n34708 ^ n1891;
  assign n34846 = n34845 ^ n34709;
  assign n34705 = ~n34703 & n34704;
  assign n34647 = n34646 ^ n34536;
  assign n34648 = n34537 & ~n34647;
  assign n34649 = n34648 ^ n31102;
  assign n34650 = n34649 ^ n31092;
  assign n34328 = n34327 ^ n34323;
  assign n34530 = n34529 ^ n34323;
  assign n34531 = n34328 & ~n34530;
  assign n34532 = n34531 ^ n34327;
  assign n34312 = n32762 ^ n31823;
  assign n34313 = n33358 ^ n32762;
  assign n34314 = ~n34312 & ~n34313;
  assign n34315 = n34314 ^ n31823;
  assign n34533 = n34532 ^ n34315;
  assign n34310 = n34068 ^ n2930;
  assign n34311 = n34310 ^ n33954;
  assign n34534 = n34533 ^ n34311;
  assign n34651 = n34650 ^ n34534;
  assign n34706 = n34705 ^ n34651;
  assign n34847 = n34846 ^ n34706;
  assign n34852 = n34851 ^ n34847;
  assign n34868 = n34867 ^ n34852;
  assign n35274 = n34868 ^ n31573;
  assign n34869 = n34857 ^ n34856;
  assign n34870 = n31586 & ~n34869;
  assign n34871 = n34870 ^ n31583;
  assign n34872 = n34864 ^ n34863;
  assign n34873 = n34872 ^ n34870;
  assign n34874 = ~n34871 & n34873;
  assign n34875 = n34874 ^ n31583;
  assign n35275 = n34875 ^ n34868;
  assign n35276 = n35274 & ~n35275;
  assign n35277 = n35276 ^ n31573;
  assign n35115 = n34867 ^ n34847;
  assign n35116 = ~n34852 & ~n35115;
  assign n35117 = n35116 ^ n34851;
  assign n35110 = n33627 ^ n32513;
  assign n35111 = n34448 ^ n33627;
  assign n35112 = ~n35110 & ~n35111;
  assign n35113 = n35112 ^ n32513;
  assign n35092 = n34709 ^ n34706;
  assign n35093 = n34845 ^ n34706;
  assign n35094 = n35092 & ~n35093;
  assign n35095 = n35094 ^ n34709;
  assign n35066 = n34534 ^ n31092;
  assign n35067 = n34649 ^ n34534;
  assign n35068 = n35066 & n35067;
  assign n35069 = n35068 ^ n31092;
  assign n35070 = n35069 ^ n30693;
  assign n35060 = n34315 ^ n34311;
  assign n35061 = n34532 ^ n34311;
  assign n35062 = ~n35060 & ~n35061;
  assign n35063 = n35062 ^ n34315;
  assign n35056 = n32687 ^ n31602;
  assign n35057 = n33356 ^ n32687;
  assign n35058 = n35056 & n35057;
  assign n35059 = n35058 ^ n31602;
  assign n35064 = n35063 ^ n35059;
  assign n34929 = n34071 ^ n33953;
  assign n35065 = n35064 ^ n34929;
  assign n35071 = n35070 ^ n35065;
  assign n35055 = n34651 & n34705;
  assign n35090 = n35071 ^ n35055;
  assign n1884 = n1883 ^ n1832;
  assign n1897 = n1896 ^ n1884;
  assign n1904 = n1903 ^ n1897;
  assign n35091 = n35090 ^ n1904;
  assign n35109 = n35095 ^ n35091;
  assign n35114 = n35113 ^ n35109;
  assign n35272 = n35117 ^ n35114;
  assign n35273 = n35272 ^ n31567;
  assign n35377 = n35277 ^ n35273;
  assign n34876 = n34875 ^ n31573;
  assign n34877 = n34876 ^ n34868;
  assign n35561 = n35377 ^ n34877;
  assign n35565 = n35564 ^ n35561;
  assign n2331 = n2330 ^ n2231;
  assign n2332 = n2331 ^ n2324;
  assign n2333 = n2332 ^ n2312;
  assign n34878 = n34877 ^ n2333;
  assign n34881 = n32500 ^ n25019;
  assign n34882 = n34881 ^ n2158;
  assign n34883 = n34882 ^ n2318;
  assign n2137 = n2126 ^ n2058;
  assign n2144 = n2143 ^ n2137;
  assign n2151 = n2150 ^ n2144;
  assign n34879 = n34869 ^ n31586;
  assign n34880 = n2151 & ~n34879;
  assign n34884 = n34883 ^ n34880;
  assign n34885 = n34872 ^ n34871;
  assign n34886 = n34885 ^ n34883;
  assign n34887 = n34884 & ~n34886;
  assign n34888 = n34887 ^ n34880;
  assign n35566 = n34888 ^ n34877;
  assign n35567 = n34878 & ~n35566;
  assign n35568 = n35567 ^ n2333;
  assign n35569 = n35568 ^ n35561;
  assign n35570 = n35565 & ~n35569;
  assign n35571 = n35570 ^ n35564;
  assign n35556 = n33251 ^ n25010;
  assign n35557 = n35556 ^ n29039;
  assign n35558 = n35557 ^ n696;
  assign n35769 = n35571 ^ n35558;
  assign n35278 = n35277 ^ n35272;
  assign n35279 = ~n35273 & ~n35278;
  assign n35280 = n35279 ^ n31567;
  assign n35379 = n35280 ^ n31561;
  assign n35118 = n35117 ^ n35109;
  assign n35119 = n35114 & ~n35118;
  assign n35120 = n35119 ^ n35113;
  assign n35104 = n33634 ^ n32506;
  assign n35105 = n34442 ^ n33634;
  assign n35106 = ~n35104 & ~n35105;
  assign n35107 = n35106 ^ n32506;
  assign n35099 = n32748 ^ n2266;
  assign n35100 = n35099 ^ n28885;
  assign n35101 = n35100 ^ n2039;
  assign n35096 = n35095 ^ n35090;
  assign n35097 = ~n35091 & n35096;
  assign n35098 = n35097 ^ n1904;
  assign n35102 = n35101 ^ n35098;
  assign n35082 = n35059 ^ n34929;
  assign n35083 = n35063 ^ n34929;
  assign n35084 = ~n35082 & n35083;
  assign n35085 = n35084 ^ n35059;
  assign n35078 = n32681 ^ n31596;
  assign n35079 = n33350 ^ n32681;
  assign n35080 = ~n35078 & n35079;
  assign n35081 = n35080 ^ n31596;
  assign n35086 = n35085 ^ n35081;
  assign n34922 = n34074 ^ n33948;
  assign n35087 = n35086 ^ n34922;
  assign n35073 = n35065 ^ n30693;
  assign n35074 = n35069 ^ n35065;
  assign n35075 = n35073 & n35074;
  assign n35076 = n35075 ^ n30693;
  assign n35077 = n35076 ^ n30687;
  assign n35088 = n35087 ^ n35077;
  assign n35072 = n35055 & ~n35071;
  assign n35089 = n35088 ^ n35072;
  assign n35103 = n35102 ^ n35089;
  assign n35108 = n35107 ^ n35103;
  assign n35270 = n35120 ^ n35108;
  assign n35380 = n35379 ^ n35270;
  assign n35378 = n34877 & ~n35377;
  assign n35559 = n35380 ^ n35378;
  assign n35770 = n35769 ^ n35559;
  assign n35764 = n34405 ^ n33672;
  assign n35001 = n34780 ^ n34769;
  assign n35002 = n35001 ^ n34770;
  assign n35765 = n35002 ^ n34405;
  assign n35766 = n35764 & ~n35765;
  assign n35767 = n35766 ^ n33672;
  assign n35716 = n35568 ^ n35565;
  assign n35712 = n34411 ^ n33600;
  assign n35008 = n34777 ^ n34773;
  assign n35713 = n35008 ^ n34411;
  assign n35714 = ~n35712 & ~n35713;
  assign n35715 = n35714 ^ n33600;
  assign n35717 = n35716 ^ n35715;
  assign n34889 = n34888 ^ n34878;
  assign n33543 = n33542 ^ n33541;
  assign n34288 = n34287 ^ n34284;
  assign n34306 = n34305 ^ n34288;
  assign n34307 = n34306 ^ n33541;
  assign n34308 = n33543 & n34307;
  assign n34309 = n34308 ^ n33542;
  assign n34890 = n34889 ^ n34309;
  assign n34898 = n34879 ^ n2151;
  assign n34892 = n34428 ^ n33617;
  assign n34893 = n34278 ^ n34241;
  assign n34894 = n34893 ^ n34238;
  assign n34895 = n34894 ^ n34428;
  assign n34896 = n34892 & ~n34895;
  assign n34897 = n34896 ^ n33617;
  assign n34899 = n34898 ^ n34897;
  assign n35655 = n34434 ^ n33634;
  assign n35136 = n34275 ^ n34246;
  assign n35137 = n35136 ^ n34243;
  assign n35656 = n35137 ^ n34434;
  assign n35657 = ~n35655 & ~n35656;
  assign n35658 = n35657 ^ n33634;
  assign n34918 = n34820 ^ n2702;
  assign n34919 = n34918 ^ n34730;
  assign n34914 = n33358 ^ n32774;
  assign n34915 = n34130 ^ n33358;
  assign n34916 = ~n34914 & n34915;
  assign n34917 = n34916 ^ n32774;
  assign n34920 = n34919 ^ n34917;
  assign n34926 = n34817 ^ n34733;
  assign n34921 = n33368 ^ n32495;
  assign n34923 = n34922 ^ n33368;
  assign n34924 = ~n34921 & n34923;
  assign n34925 = n34924 ^ n32495;
  assign n34927 = n34926 ^ n34925;
  assign n34933 = n34814 ^ n2616;
  assign n34934 = n34933 ^ n34734;
  assign n34928 = n33370 ^ n32433;
  assign n34930 = n34929 ^ n33370;
  assign n34931 = n34928 & ~n34930;
  assign n34932 = n34931 ^ n32433;
  assign n34935 = n34934 ^ n34932;
  assign n34940 = n34811 ^ n3179;
  assign n34941 = n34940 ^ n34736;
  assign n34936 = n34149 ^ n33118;
  assign n34937 = n34311 ^ n34149;
  assign n34938 = n34936 & ~n34937;
  assign n34939 = n34938 ^ n33118;
  assign n34942 = n34941 ^ n34939;
  assign n34947 = n34808 ^ n34742;
  assign n34943 = n34090 ^ n33100;
  assign n34944 = n34323 ^ n34090;
  assign n34945 = n34943 & ~n34944;
  assign n34946 = n34945 ^ n33100;
  assign n34948 = n34947 ^ n34946;
  assign n34953 = n34805 ^ n34747;
  assign n34949 = n33545 ^ n32524;
  assign n34950 = n34333 ^ n33545;
  assign n34951 = ~n34949 & n34950;
  assign n34952 = n34951 ^ n32524;
  assign n34954 = n34953 ^ n34952;
  assign n34959 = n34802 ^ n1438;
  assign n34955 = n33561 ^ n32536;
  assign n34956 = n34342 ^ n33561;
  assign n34957 = n34955 & ~n34956;
  assign n34958 = n34957 ^ n32536;
  assign n34960 = n34959 ^ n34958;
  assign n34965 = n34798 ^ n1420;
  assign n34966 = n34965 ^ n34749;
  assign n34961 = n33567 ^ n32542;
  assign n34962 = n34348 ^ n33567;
  assign n34963 = ~n34961 & n34962;
  assign n34964 = n34963 ^ n32542;
  assign n34967 = n34966 ^ n34964;
  assign n34972 = n34795 ^ n34752;
  assign n34968 = n33576 ^ n32556;
  assign n34969 = n34359 ^ n33576;
  assign n34970 = ~n34968 & n34969;
  assign n34971 = n34970 ^ n32556;
  assign n34973 = n34972 ^ n34971;
  assign n34976 = n33582 ^ n32558;
  assign n34977 = n34509 ^ n33582;
  assign n34978 = ~n34976 & n34977;
  assign n34979 = n34978 ^ n32558;
  assign n34974 = n34792 ^ n1238;
  assign n34975 = n34974 ^ n34753;
  assign n34980 = n34979 ^ n34975;
  assign n34983 = n33594 ^ n32570;
  assign n34984 = n34368 ^ n33594;
  assign n34985 = n34983 & n34984;
  assign n34986 = n34985 ^ n32570;
  assign n34981 = n34789 ^ n3339;
  assign n34982 = n34981 ^ n34755;
  assign n34987 = n34986 ^ n34982;
  assign n34990 = n33718 ^ n32577;
  assign n34991 = n34374 ^ n33718;
  assign n34992 = ~n34990 & ~n34991;
  assign n34993 = n34992 ^ n32577;
  assign n34988 = n34786 ^ n34760;
  assign n34989 = n34988 ^ n34757;
  assign n34994 = n34993 ^ n34989;
  assign n34996 = n33713 ^ n32586;
  assign n34997 = n34380 ^ n33713;
  assign n34998 = n34996 & n34997;
  assign n34999 = n34998 ^ n32586;
  assign n34995 = n34783 ^ n34766;
  assign n35000 = n34999 ^ n34995;
  assign n35003 = n33693 ^ n32592;
  assign n35004 = n34386 ^ n33693;
  assign n35005 = n35003 & n35004;
  assign n35006 = n35005 ^ n32592;
  assign n35007 = n35006 ^ n35002;
  assign n35009 = n33703 ^ n32598;
  assign n35010 = n34388 ^ n33703;
  assign n35011 = n35009 & ~n35010;
  assign n35012 = n35011 ^ n32598;
  assign n35013 = n35012 ^ n35008;
  assign n35014 = n33677 ^ n32604;
  assign n35015 = n34395 ^ n33677;
  assign n35016 = ~n35014 & ~n35015;
  assign n35017 = n35016 ^ n32604;
  assign n35018 = n35017 ^ n34306;
  assign n35023 = n34281 ^ n34237;
  assign n35019 = n33688 ^ n32610;
  assign n35020 = n34405 ^ n33688;
  assign n35021 = n35019 & ~n35020;
  assign n35022 = n35021 ^ n32610;
  assign n35024 = n35023 ^ n35022;
  assign n35025 = n33666 ^ n32620;
  assign n35026 = n34411 ^ n33666;
  assign n35027 = n35025 & n35026;
  assign n35028 = n35027 ^ n32620;
  assign n35029 = n35028 ^ n34894;
  assign n35034 = n34272 ^ n34250;
  assign n35035 = n35034 ^ n34251;
  assign n35030 = n33600 ^ n32628;
  assign n35031 = n34422 ^ n33600;
  assign n35032 = n35030 & n35031;
  assign n35033 = n35032 ^ n32628;
  assign n35036 = n35035 ^ n35033;
  assign n35041 = n34269 ^ n34256;
  assign n35037 = n33542 ^ n32638;
  assign n35038 = n34428 ^ n33542;
  assign n35039 = ~n35037 & n35038;
  assign n35040 = n35039 ^ n32638;
  assign n35042 = n35041 ^ n35040;
  assign n35047 = n34266 ^ n34265;
  assign n35043 = n33611 ^ n32640;
  assign n35044 = n34434 ^ n33611;
  assign n35045 = n35043 & ~n35044;
  assign n35046 = n35045 ^ n32640;
  assign n35048 = n35047 ^ n35046;
  assign n35050 = n33617 ^ n32650;
  assign n35051 = n34436 ^ n33617;
  assign n35052 = ~n35050 & n35051;
  assign n35053 = n35052 ^ n32650;
  assign n35049 = n34260 ^ n34259;
  assign n35054 = n35053 ^ n35049;
  assign n35121 = n35120 ^ n35103;
  assign n35122 = n35108 & n35121;
  assign n35123 = n35122 ^ n35107;
  assign n35124 = n35123 ^ n35049;
  assign n35125 = n35054 & ~n35124;
  assign n35126 = n35125 ^ n35053;
  assign n35127 = n35126 ^ n35047;
  assign n35128 = n35048 & ~n35127;
  assign n35129 = n35128 ^ n35046;
  assign n35130 = n35129 ^ n35041;
  assign n35131 = n35042 & n35130;
  assign n35132 = n35131 ^ n35040;
  assign n35133 = n35132 ^ n35035;
  assign n35134 = n35036 & n35133;
  assign n35135 = n35134 ^ n35033;
  assign n35138 = n35137 ^ n35135;
  assign n35139 = n33672 ^ n32622;
  assign n35140 = n33672 ^ n33541;
  assign n35141 = ~n35139 & ~n35140;
  assign n35142 = n35141 ^ n32622;
  assign n35143 = n35142 ^ n35137;
  assign n35144 = ~n35138 & ~n35143;
  assign n35145 = n35144 ^ n35142;
  assign n35146 = n35145 ^ n34894;
  assign n35147 = ~n35029 & ~n35146;
  assign n35148 = n35147 ^ n35028;
  assign n35149 = n35148 ^ n35023;
  assign n35150 = ~n35024 & n35149;
  assign n35151 = n35150 ^ n35022;
  assign n35152 = n35151 ^ n34306;
  assign n35153 = ~n35018 & n35152;
  assign n35154 = n35153 ^ n35017;
  assign n35155 = n35154 ^ n35008;
  assign n35156 = n35013 & n35155;
  assign n35157 = n35156 ^ n35012;
  assign n35158 = n35157 ^ n35002;
  assign n35159 = n35007 & n35158;
  assign n35160 = n35159 ^ n35006;
  assign n35161 = n35160 ^ n34995;
  assign n35162 = n35000 & ~n35161;
  assign n35163 = n35162 ^ n34999;
  assign n35164 = n35163 ^ n34989;
  assign n35165 = ~n34994 & ~n35164;
  assign n35166 = n35165 ^ n34993;
  assign n35167 = n35166 ^ n34982;
  assign n35168 = n34987 & ~n35167;
  assign n35169 = n35168 ^ n34986;
  assign n35170 = n35169 ^ n34975;
  assign n35171 = ~n34980 & ~n35170;
  assign n35172 = n35171 ^ n34979;
  assign n35173 = n35172 ^ n34972;
  assign n35174 = n34973 & ~n35173;
  assign n35175 = n35174 ^ n34971;
  assign n35176 = n35175 ^ n34966;
  assign n35177 = n34967 & ~n35176;
  assign n35178 = n35177 ^ n34964;
  assign n35179 = n35178 ^ n34959;
  assign n35180 = ~n34960 & n35179;
  assign n35181 = n35180 ^ n34958;
  assign n35182 = n35181 ^ n34953;
  assign n35183 = n34954 & n35182;
  assign n35184 = n35183 ^ n34952;
  assign n35185 = n35184 ^ n34947;
  assign n35186 = n34948 & n35185;
  assign n35187 = n35186 ^ n34946;
  assign n35188 = n35187 ^ n34941;
  assign n35189 = n34942 & ~n35188;
  assign n35190 = n35189 ^ n34939;
  assign n35191 = n35190 ^ n34934;
  assign n35192 = ~n34935 & n35191;
  assign n35193 = n35192 ^ n34932;
  assign n35194 = n35193 ^ n34926;
  assign n35195 = n34927 & ~n35194;
  assign n35196 = n35195 ^ n34925;
  assign n35197 = n35196 ^ n34919;
  assign n35198 = ~n34920 & ~n35197;
  assign n35199 = n35198 ^ n34917;
  assign n34908 = n33356 ^ n32768;
  assign n34909 = n34120 ^ n33356;
  assign n34910 = ~n34908 & ~n34909;
  assign n34911 = n34910 ^ n32768;
  assign n35215 = n35199 ^ n34911;
  assign n34912 = n34823 ^ n34729;
  assign n35216 = n35215 ^ n34912;
  assign n35217 = n35216 ^ n31825;
  assign n35218 = n35196 ^ n34917;
  assign n35219 = n35218 ^ n34919;
  assign n35220 = n35219 ^ n31835;
  assign n35221 = n35193 ^ n34927;
  assign n35222 = n35221 ^ n31841;
  assign n35223 = n35190 ^ n34935;
  assign n35224 = n35223 ^ n31847;
  assign n35225 = n35187 ^ n34942;
  assign n35226 = n35225 ^ n32549;
  assign n35227 = n35184 ^ n34948;
  assign n35228 = n35227 ^ n32560;
  assign n35229 = n35181 ^ n34954;
  assign n35230 = n35229 ^ n32572;
  assign n35231 = n35178 ^ n34960;
  assign n35232 = n35231 ^ n32459;
  assign n35233 = n35175 ^ n34967;
  assign n35234 = n35233 ^ n31503;
  assign n35235 = n35172 ^ n34973;
  assign n35236 = n35235 ^ n31509;
  assign n35237 = n35169 ^ n34980;
  assign n35238 = n35237 ^ n31517;
  assign n35239 = n35166 ^ n34987;
  assign n35240 = n35239 ^ n31527;
  assign n35241 = n35163 ^ n34994;
  assign n35242 = n35241 ^ n31941;
  assign n35243 = n35160 ^ n35000;
  assign n35244 = n35243 ^ n31945;
  assign n35245 = n35157 ^ n35007;
  assign n35246 = n35245 ^ n31935;
  assign n35247 = n35154 ^ n35012;
  assign n35248 = n35247 ^ n35008;
  assign n35249 = n35248 ^ n31927;
  assign n35250 = n35151 ^ n35018;
  assign n35251 = n35250 ^ n31919;
  assign n35252 = n35148 ^ n35024;
  assign n35253 = n35252 ^ n31898;
  assign n35254 = n35145 ^ n35029;
  assign n35255 = n35254 ^ n31904;
  assign n35256 = n35142 ^ n35138;
  assign n35257 = n35256 ^ n31906;
  assign n35258 = n35132 ^ n35033;
  assign n35259 = n35258 ^ n35035;
  assign n35260 = n35259 ^ n31541;
  assign n35261 = n35129 ^ n35040;
  assign n35262 = n35261 ^ n35041;
  assign n35263 = n35262 ^ n31543;
  assign n35264 = n35126 ^ n35046;
  assign n35265 = n35264 ^ n35047;
  assign n35266 = n35265 ^ n31549;
  assign n35267 = n35123 ^ n35053;
  assign n35268 = n35267 ^ n35049;
  assign n35269 = n35268 ^ n31555;
  assign n35271 = n35270 ^ n31561;
  assign n35281 = n35280 ^ n35270;
  assign n35282 = n35271 & n35281;
  assign n35283 = n35282 ^ n31561;
  assign n35284 = n35283 ^ n35268;
  assign n35285 = n35269 & n35284;
  assign n35286 = n35285 ^ n31555;
  assign n35287 = n35286 ^ n35265;
  assign n35288 = n35266 & ~n35287;
  assign n35289 = n35288 ^ n31549;
  assign n35290 = n35289 ^ n35262;
  assign n35291 = n35263 & ~n35290;
  assign n35292 = n35291 ^ n31543;
  assign n35293 = n35292 ^ n35259;
  assign n35294 = ~n35260 & n35293;
  assign n35295 = n35294 ^ n31541;
  assign n35296 = n35295 ^ n35256;
  assign n35297 = n35257 & n35296;
  assign n35298 = n35297 ^ n31906;
  assign n35299 = n35298 ^ n35254;
  assign n35300 = n35255 & n35299;
  assign n35301 = n35300 ^ n31904;
  assign n35302 = n35301 ^ n35252;
  assign n35303 = ~n35253 & n35302;
  assign n35304 = n35303 ^ n31898;
  assign n35305 = n35304 ^ n35250;
  assign n35306 = ~n35251 & n35305;
  assign n35307 = n35306 ^ n31919;
  assign n35308 = n35307 ^ n35248;
  assign n35309 = n35249 & ~n35308;
  assign n35310 = n35309 ^ n31927;
  assign n35311 = n35310 ^ n35245;
  assign n35312 = ~n35246 & n35311;
  assign n35313 = n35312 ^ n31935;
  assign n35314 = n35313 ^ n35243;
  assign n35315 = n35244 & ~n35314;
  assign n35316 = n35315 ^ n31945;
  assign n35317 = n35316 ^ n35241;
  assign n35318 = ~n35242 & n35317;
  assign n35319 = n35318 ^ n31941;
  assign n35320 = n35319 ^ n35239;
  assign n35321 = ~n35240 & n35320;
  assign n35322 = n35321 ^ n31527;
  assign n35323 = n35322 ^ n35237;
  assign n35324 = ~n35238 & ~n35323;
  assign n35325 = n35324 ^ n31517;
  assign n35326 = n35325 ^ n35235;
  assign n35327 = ~n35236 & n35326;
  assign n35328 = n35327 ^ n31509;
  assign n35329 = n35328 ^ n35233;
  assign n35330 = n35234 & n35329;
  assign n35331 = n35330 ^ n31503;
  assign n35332 = n35331 ^ n35231;
  assign n35333 = ~n35232 & n35332;
  assign n35334 = n35333 ^ n32459;
  assign n35335 = n35334 ^ n35229;
  assign n35336 = ~n35230 & ~n35335;
  assign n35337 = n35336 ^ n32572;
  assign n35338 = n35337 ^ n35227;
  assign n35339 = n35228 & ~n35338;
  assign n35340 = n35339 ^ n32560;
  assign n35341 = n35340 ^ n35225;
  assign n35342 = n35226 & n35341;
  assign n35343 = n35342 ^ n32549;
  assign n35344 = n35343 ^ n35223;
  assign n35345 = ~n35224 & n35344;
  assign n35346 = n35345 ^ n31847;
  assign n35347 = n35346 ^ n35221;
  assign n35348 = n35222 & ~n35347;
  assign n35349 = n35348 ^ n31841;
  assign n35350 = n35349 ^ n35219;
  assign n35351 = ~n35220 & n35350;
  assign n35352 = n35351 ^ n31835;
  assign n35353 = n35352 ^ n35216;
  assign n35354 = ~n35217 & n35353;
  assign n35355 = n35354 ^ n31825;
  assign n35361 = n35355 ^ n31823;
  assign n34913 = n34912 ^ n34911;
  assign n35200 = n35199 ^ n34912;
  assign n35201 = n34913 & ~n35200;
  assign n35202 = n35201 ^ n34911;
  assign n34903 = n33350 ^ n32762;
  assign n34904 = n34114 ^ n33350;
  assign n34905 = n34903 & n34904;
  assign n34906 = n34905 ^ n32762;
  assign n35212 = n35202 ^ n34906;
  assign n34901 = n34826 ^ n34726;
  assign n34902 = n34901 ^ n34723;
  assign n35213 = n35212 ^ n34902;
  assign n35362 = n35361 ^ n35213;
  assign n35363 = n35349 ^ n35220;
  assign n35364 = n35337 ^ n35228;
  assign n35365 = n35331 ^ n35232;
  assign n35366 = n35325 ^ n35236;
  assign n35367 = n35319 ^ n35240;
  assign n35368 = n35316 ^ n35242;
  assign n35369 = n35307 ^ n35249;
  assign n35370 = n35304 ^ n31919;
  assign n35371 = n35370 ^ n35250;
  assign n35372 = n35292 ^ n31541;
  assign n35373 = n35372 ^ n35259;
  assign n35374 = n35289 ^ n31543;
  assign n35375 = n35374 ^ n35262;
  assign n35376 = n35283 ^ n35269;
  assign n35381 = n35378 & ~n35380;
  assign n35382 = ~n35376 & ~n35381;
  assign n35383 = n35286 ^ n31549;
  assign n35384 = n35383 ^ n35265;
  assign n35385 = ~n35382 & ~n35384;
  assign n35386 = ~n35375 & n35385;
  assign n35387 = ~n35373 & ~n35386;
  assign n35388 = n35295 ^ n31906;
  assign n35389 = n35388 ^ n35256;
  assign n35390 = n35387 & n35389;
  assign n35391 = n35298 ^ n31904;
  assign n35392 = n35391 ^ n35254;
  assign n35393 = ~n35390 & n35392;
  assign n35394 = n35301 ^ n35253;
  assign n35395 = n35393 & n35394;
  assign n35396 = n35371 & n35395;
  assign n35397 = ~n35369 & n35396;
  assign n35398 = n35310 ^ n31935;
  assign n35399 = n35398 ^ n35245;
  assign n35400 = ~n35397 & ~n35399;
  assign n35401 = n35313 ^ n35244;
  assign n35402 = ~n35400 & ~n35401;
  assign n35403 = n35368 & n35402;
  assign n35404 = n35367 & n35403;
  assign n35405 = n35322 ^ n31517;
  assign n35406 = n35405 ^ n35237;
  assign n35407 = ~n35404 & ~n35406;
  assign n35408 = ~n35366 & ~n35407;
  assign n35409 = n35328 ^ n31503;
  assign n35410 = n35409 ^ n35233;
  assign n35411 = n35408 & n35410;
  assign n35412 = ~n35365 & ~n35411;
  assign n35413 = n35334 ^ n32572;
  assign n35414 = n35413 ^ n35229;
  assign n35415 = n35412 & ~n35414;
  assign n35416 = ~n35364 & n35415;
  assign n35417 = n35340 ^ n35226;
  assign n35418 = ~n35416 & n35417;
  assign n35419 = n35343 ^ n35224;
  assign n35420 = n35418 & n35419;
  assign n35421 = n35346 ^ n31841;
  assign n35422 = n35421 ^ n35221;
  assign n35423 = n35420 & ~n35422;
  assign n35424 = n35363 & n35423;
  assign n35425 = n35352 ^ n31825;
  assign n35426 = n35425 ^ n35216;
  assign n35427 = ~n35424 & ~n35426;
  assign n35428 = ~n35362 & n35427;
  assign n35214 = n35213 ^ n31823;
  assign n35356 = n35355 ^ n35213;
  assign n35357 = ~n35214 & ~n35356;
  assign n35358 = n35357 ^ n31823;
  assign n35359 = n35358 ^ n31602;
  assign n35207 = n32687 ^ n32511;
  assign n35208 = n34108 ^ n32511;
  assign n35209 = ~n35207 & n35208;
  assign n35210 = n35209 ^ n32687;
  assign n34907 = n34906 ^ n34902;
  assign n35203 = n35202 ^ n34902;
  assign n35204 = ~n34907 & ~n35203;
  assign n35205 = n35204 ^ n34906;
  assign n34900 = n34829 ^ n34722;
  assign n35206 = n35205 ^ n34900;
  assign n35211 = n35210 ^ n35206;
  assign n35360 = n35359 ^ n35211;
  assign n35447 = n35428 ^ n35360;
  assign n2003 = n1976 ^ n1924;
  assign n2004 = n2003 ^ n2002;
  assign n2005 = n2004 ^ n1990;
  assign n35448 = n35447 ^ n2005;
  assign n35449 = n35427 ^ n35362;
  assign n35453 = n35452 ^ n35449;
  assign n35454 = n35426 ^ n35424;
  assign n35458 = n35457 ^ n35454;
  assign n35460 = n33149 ^ n25427;
  assign n35461 = n35460 ^ n29386;
  assign n35462 = n35461 ^ n24019;
  assign n35459 = n35423 ^ n35363;
  assign n35463 = n35462 ^ n35459;
  assign n35464 = n35422 ^ n35420;
  assign n35468 = n35467 ^ n35464;
  assign n35469 = n35419 ^ n35418;
  assign n35473 = n35472 ^ n35469;
  assign n35474 = n35417 ^ n35416;
  assign n2887 = n2883 ^ n2826;
  assign n2891 = n2890 ^ n2887;
  assign n2892 = n2891 ^ n1538;
  assign n35475 = n35474 ^ n2892;
  assign n35476 = n35415 ^ n35364;
  assign n2798 = n2737 ^ n1583;
  assign n2799 = n2798 ^ n2795;
  assign n2803 = n2802 ^ n2799;
  assign n35477 = n35476 ^ n2803;
  assign n35478 = n35414 ^ n35412;
  assign n2765 = n2758 ^ n2722;
  assign n2781 = n2780 ^ n2765;
  assign n2788 = n2787 ^ n2781;
  assign n35479 = n35478 ^ n2788;
  assign n35480 = n35411 ^ n35365;
  assign n3205 = n3201 ^ n2672;
  assign n3212 = n3211 ^ n3205;
  assign n3213 = n3212 ^ n2777;
  assign n35481 = n35480 ^ n3213;
  assign n35482 = n35410 ^ n35408;
  assign n35486 = n35485 ^ n35482;
  assign n35490 = n35407 ^ n35366;
  assign n35487 = n29410 ^ n3187;
  assign n35488 = n35487 ^ n33183;
  assign n35489 = n35488 ^ n3058;
  assign n35491 = n35490 ^ n35489;
  assign n35495 = n35406 ^ n35404;
  assign n35492 = n33190 ^ n25444;
  assign n35493 = n35492 ^ n3035;
  assign n35494 = n35493 ^ n2491;
  assign n35496 = n35495 ^ n35494;
  assign n35500 = n35403 ^ n35367;
  assign n35497 = n25449 ^ n1485;
  assign n35498 = n35497 ^ n2429;
  assign n35499 = n35498 ^ n3033;
  assign n35501 = n35500 ^ n35499;
  assign n35505 = n35402 ^ n35368;
  assign n35502 = n3017 ^ n1467;
  assign n35503 = n35502 ^ n29418;
  assign n35504 = n35503 ^ n2424;
  assign n35506 = n35505 ^ n35504;
  assign n35510 = n35401 ^ n35400;
  assign n35507 = n1452 ^ n1360;
  assign n35508 = n35507 ^ n29424;
  assign n35509 = n35508 ^ n1280;
  assign n35511 = n35510 ^ n35509;
  assign n35513 = n33208 ^ n1345;
  assign n35514 = n35513 ^ n1100;
  assign n35515 = n35514 ^ n24072;
  assign n35512 = n35399 ^ n35397;
  assign n35516 = n35515 ^ n35512;
  assign n35518 = n33213 ^ n1336;
  assign n35519 = n35518 ^ n29095;
  assign n35520 = n35519 ^ n1095;
  assign n35517 = n35396 ^ n35369;
  assign n35521 = n35520 ^ n35517;
  assign n35522 = n35395 ^ n35371;
  assign n930 = n929 ^ n878;
  assign n943 = n942 ^ n930;
  assign n950 = n949 ^ n943;
  assign n35523 = n35522 ^ n950;
  assign n35525 = n33220 ^ n25058;
  assign n35526 = n35525 ^ n847;
  assign n35527 = n35526 ^ n940;
  assign n35524 = n35394 ^ n35393;
  assign n35528 = n35527 ^ n35524;
  assign n35529 = n35392 ^ n35390;
  assign n814 = n807 ^ n780;
  assign n833 = n832 ^ n814;
  assign n840 = n839 ^ n833;
  assign n35530 = n35529 ^ n840;
  assign n35531 = n35389 ^ n35387;
  assign n35535 = n35534 ^ n35531;
  assign n35537 = n33232 ^ n627;
  assign n35538 = n35537 ^ n29021;
  assign n35539 = n35538 ^ n3272;
  assign n35536 = n35386 ^ n35373;
  assign n35540 = n35539 ^ n35536;
  assign n35541 = n35385 ^ n35375;
  assign n35545 = n35544 ^ n35541;
  assign n35547 = n33242 ^ n25004;
  assign n35548 = n35547 ^ n29031;
  assign n35549 = n35548 ^ n23683;
  assign n35546 = n35384 ^ n35382;
  assign n35550 = n35549 ^ n35546;
  assign n35554 = n35381 ^ n35376;
  assign n35551 = n33247 ^ n25035;
  assign n35552 = n35551 ^ n29035;
  assign n35553 = n35552 ^ n23688;
  assign n35555 = n35554 ^ n35553;
  assign n35560 = n35559 ^ n35558;
  assign n35572 = n35571 ^ n35559;
  assign n35573 = n35560 & ~n35572;
  assign n35574 = n35573 ^ n35558;
  assign n35575 = n35574 ^ n35554;
  assign n35576 = n35555 & ~n35575;
  assign n35577 = n35576 ^ n35553;
  assign n35578 = n35577 ^ n35546;
  assign n35579 = ~n35550 & n35578;
  assign n35580 = n35579 ^ n35549;
  assign n35581 = n35580 ^ n35541;
  assign n35582 = n35545 & ~n35581;
  assign n35583 = n35582 ^ n35544;
  assign n35584 = n35583 ^ n35536;
  assign n35585 = n35540 & ~n35584;
  assign n35586 = n35585 ^ n35539;
  assign n35587 = n35586 ^ n35531;
  assign n35588 = n35535 & ~n35587;
  assign n35589 = n35588 ^ n35534;
  assign n35590 = n35589 ^ n35529;
  assign n35591 = n35530 & ~n35590;
  assign n35592 = n35591 ^ n840;
  assign n35593 = n35592 ^ n35524;
  assign n35594 = ~n35528 & n35593;
  assign n35595 = n35594 ^ n35527;
  assign n35596 = n35595 ^ n35522;
  assign n35597 = ~n35523 & n35596;
  assign n35598 = n35597 ^ n950;
  assign n35599 = n35598 ^ n35517;
  assign n35600 = n35521 & ~n35599;
  assign n35601 = n35600 ^ n35520;
  assign n35602 = n35601 ^ n35512;
  assign n35603 = n35516 & ~n35602;
  assign n35604 = n35603 ^ n35515;
  assign n35605 = n35604 ^ n35510;
  assign n35606 = ~n35511 & n35605;
  assign n35607 = n35606 ^ n35509;
  assign n35608 = n35607 ^ n35505;
  assign n35609 = ~n35506 & n35608;
  assign n35610 = n35609 ^ n35504;
  assign n35611 = n35610 ^ n35500;
  assign n35612 = ~n35501 & n35611;
  assign n35613 = n35612 ^ n35499;
  assign n35614 = n35613 ^ n35495;
  assign n35615 = n35496 & ~n35614;
  assign n35616 = n35615 ^ n35494;
  assign n35617 = n35616 ^ n35490;
  assign n35618 = ~n35491 & n35617;
  assign n35619 = n35618 ^ n35489;
  assign n35620 = n35619 ^ n35482;
  assign n35621 = ~n35486 & n35620;
  assign n35622 = n35621 ^ n35485;
  assign n35623 = n35622 ^ n35480;
  assign n35624 = n35481 & ~n35623;
  assign n35625 = n35624 ^ n3213;
  assign n35626 = n35625 ^ n35478;
  assign n35627 = ~n35479 & n35626;
  assign n35628 = n35627 ^ n2788;
  assign n35629 = n35628 ^ n35476;
  assign n35630 = ~n35477 & n35629;
  assign n35631 = n35630 ^ n2803;
  assign n35632 = n35631 ^ n35474;
  assign n35633 = n35475 & ~n35632;
  assign n35634 = n35633 ^ n2892;
  assign n35635 = n35634 ^ n35469;
  assign n35636 = ~n35473 & n35635;
  assign n35637 = n35636 ^ n35472;
  assign n35638 = n35637 ^ n35464;
  assign n35639 = n35468 & ~n35638;
  assign n35640 = n35639 ^ n35467;
  assign n35641 = n35640 ^ n35459;
  assign n35642 = ~n35463 & n35641;
  assign n35643 = n35642 ^ n35462;
  assign n35644 = n35643 ^ n35454;
  assign n35645 = n35458 & ~n35644;
  assign n35646 = n35645 ^ n35457;
  assign n35647 = n35646 ^ n35449;
  assign n35648 = ~n35453 & n35647;
  assign n35649 = n35648 ^ n35452;
  assign n35650 = n35649 ^ n35447;
  assign n35651 = ~n35448 & n35650;
  assign n35652 = n35651 ^ n2005;
  assign n2015 = n1971 ^ n1939;
  assign n2016 = n2015 ^ n2012;
  assign n2023 = n2022 ^ n2016;
  assign n35653 = n35652 ^ n2023;
  assign n35440 = n35211 ^ n31602;
  assign n35441 = n35358 ^ n35211;
  assign n35442 = n35440 & ~n35441;
  assign n35443 = n35442 ^ n31602;
  assign n35444 = n35443 ^ n31596;
  assign n35435 = n35210 ^ n34900;
  assign n35436 = ~n35206 & ~n35435;
  assign n35437 = n35436 ^ n35210;
  assign n35431 = n32681 ^ n32504;
  assign n35432 = n34167 ^ n32504;
  assign n35433 = ~n35431 & ~n35432;
  assign n35434 = n35433 ^ n32681;
  assign n35438 = n35437 ^ n35434;
  assign n35430 = n34832 ^ n34717;
  assign n35439 = n35438 ^ n35430;
  assign n35445 = n35444 ^ n35439;
  assign n35429 = ~n35360 & n35428;
  assign n35446 = n35445 ^ n35429;
  assign n35654 = n35653 ^ n35446;
  assign n35659 = n35658 ^ n35654;
  assign n35661 = n34436 ^ n33627;
  assign n35662 = n35035 ^ n34436;
  assign n35663 = n35661 & ~n35662;
  assign n35664 = n35663 ^ n33627;
  assign n35660 = n35649 ^ n35448;
  assign n35665 = n35664 ^ n35660;
  assign n35668 = n34442 ^ n33531;
  assign n35669 = n35041 ^ n34442;
  assign n35670 = ~n35668 & ~n35669;
  assign n35671 = n35670 ^ n33531;
  assign n35666 = n35646 ^ n35452;
  assign n35667 = n35666 ^ n35449;
  assign n35672 = n35671 ^ n35667;
  assign n35674 = n34448 ^ n33442;
  assign n35675 = n35047 ^ n34448;
  assign n35676 = n35674 & ~n35675;
  assign n35677 = n35676 ^ n33442;
  assign n35673 = n35643 ^ n35458;
  assign n35678 = n35677 ^ n35673;
  assign n35679 = n35640 ^ n35462;
  assign n35680 = n35679 ^ n35459;
  assign n35681 = n34292 ^ n33398;
  assign n35682 = n35049 ^ n34292;
  assign n35683 = n35681 & ~n35682;
  assign n35684 = n35683 ^ n33398;
  assign n35685 = ~n35680 & n35684;
  assign n35686 = n35685 ^ n35673;
  assign n35687 = ~n35678 & n35686;
  assign n35688 = n35687 ^ n35685;
  assign n35689 = n35688 ^ n35667;
  assign n35690 = ~n35672 & n35689;
  assign n35691 = n35690 ^ n35671;
  assign n35692 = n35691 ^ n35660;
  assign n35693 = ~n35665 & n35692;
  assign n35694 = n35693 ^ n35664;
  assign n35695 = n35694 ^ n35654;
  assign n35696 = n35659 & n35695;
  assign n35697 = n35696 ^ n35658;
  assign n35698 = n35697 ^ n34898;
  assign n35699 = n34899 & ~n35698;
  assign n35700 = n35699 ^ n34897;
  assign n34891 = n34885 ^ n34884;
  assign n35701 = n35700 ^ n34891;
  assign n35702 = n34422 ^ n33611;
  assign n35703 = n35023 ^ n34422;
  assign n35704 = ~n35702 & ~n35703;
  assign n35705 = n35704 ^ n33611;
  assign n35706 = n35705 ^ n34891;
  assign n35707 = n35701 & n35706;
  assign n35708 = n35707 ^ n35705;
  assign n35709 = n35708 ^ n34889;
  assign n35710 = n34890 & ~n35709;
  assign n35711 = n35710 ^ n34309;
  assign n35761 = n35716 ^ n35711;
  assign n35762 = n35717 & ~n35761;
  assign n35763 = n35762 ^ n35715;
  assign n35768 = n35767 ^ n35763;
  assign n35771 = n35770 ^ n35768;
  assign n35772 = n35771 ^ n32622;
  assign n35718 = n35717 ^ n35711;
  assign n35719 = n35718 ^ n32628;
  assign n35720 = n35708 ^ n34890;
  assign n35721 = n35720 ^ n32638;
  assign n35722 = n35705 ^ n35701;
  assign n35723 = n35722 ^ n32640;
  assign n35724 = n35697 ^ n34899;
  assign n35725 = n35724 ^ n32650;
  assign n35726 = n35694 ^ n35659;
  assign n35727 = n35726 ^ n32506;
  assign n35728 = n35691 ^ n35665;
  assign n35729 = n35728 ^ n32513;
  assign n35730 = n35688 ^ n35672;
  assign n35731 = n35730 ^ n32519;
  assign n35732 = n35684 ^ n35680;
  assign n35733 = n32679 & ~n35732;
  assign n35734 = n35733 ^ n32663;
  assign n35735 = n35685 ^ n35677;
  assign n35736 = n35735 ^ n35673;
  assign n35737 = n35736 ^ n35733;
  assign n35738 = n35734 & ~n35737;
  assign n35739 = n35738 ^ n32663;
  assign n35740 = n35739 ^ n35730;
  assign n35741 = n35731 & n35740;
  assign n35742 = n35741 ^ n32519;
  assign n35743 = n35742 ^ n35728;
  assign n35744 = n35729 & ~n35743;
  assign n35745 = n35744 ^ n32513;
  assign n35746 = n35745 ^ n35726;
  assign n35747 = n35727 & n35746;
  assign n35748 = n35747 ^ n32506;
  assign n35749 = n35748 ^ n35724;
  assign n35750 = ~n35725 & n35749;
  assign n35751 = n35750 ^ n32650;
  assign n35752 = n35751 ^ n35722;
  assign n35753 = ~n35723 & n35752;
  assign n35754 = n35753 ^ n32640;
  assign n35755 = n35754 ^ n35720;
  assign n35756 = ~n35721 & ~n35755;
  assign n35757 = n35756 ^ n32638;
  assign n35758 = n35757 ^ n35718;
  assign n35759 = n35719 & n35758;
  assign n35760 = n35759 ^ n32628;
  assign n35773 = n35772 ^ n35760;
  assign n35774 = n35757 ^ n32628;
  assign n35775 = n35774 ^ n35718;
  assign n35776 = n35754 ^ n35721;
  assign n35777 = n35739 ^ n32519;
  assign n35778 = n35777 ^ n35730;
  assign n35779 = n35742 ^ n35729;
  assign n35780 = ~n35778 & n35779;
  assign n35781 = n35745 ^ n32506;
  assign n35782 = n35781 ^ n35726;
  assign n35783 = n35780 & n35782;
  assign n35784 = n35748 ^ n35725;
  assign n35785 = ~n35783 & ~n35784;
  assign n35786 = n35751 ^ n32640;
  assign n35787 = n35786 ^ n35722;
  assign n35788 = ~n35785 & n35787;
  assign n35789 = n35776 & n35788;
  assign n35790 = ~n35775 & ~n35789;
  assign n35791 = ~n35773 & n35790;
  assign n35801 = n34395 ^ n33666;
  assign n35802 = n34995 ^ n34395;
  assign n35803 = ~n35801 & n35802;
  assign n35804 = n35803 ^ n33666;
  assign n35800 = n35574 ^ n35555;
  assign n35805 = n35804 ^ n35800;
  assign n35796 = n35770 ^ n35767;
  assign n35797 = n35770 ^ n35763;
  assign n35798 = n35796 & ~n35797;
  assign n35799 = n35798 ^ n35767;
  assign n35806 = n35805 ^ n35799;
  assign n35792 = n35771 ^ n35760;
  assign n35793 = ~n35772 & ~n35792;
  assign n35794 = n35793 ^ n32622;
  assign n35795 = n35794 ^ n32620;
  assign n35807 = n35806 ^ n35795;
  assign n35808 = ~n35791 & n35807;
  assign n35817 = n34388 ^ n33688;
  assign n35818 = n34989 ^ n34388;
  assign n35819 = ~n35817 & n35818;
  assign n35820 = n35819 ^ n33688;
  assign n35816 = n35577 ^ n35550;
  assign n35821 = n35820 ^ n35816;
  assign n35813 = n35800 ^ n35799;
  assign n35814 = n35805 & ~n35813;
  assign n35815 = n35814 ^ n35804;
  assign n35822 = n35821 ^ n35815;
  assign n35823 = n35822 ^ n32610;
  assign n35809 = n35806 ^ n32620;
  assign n35810 = n35806 ^ n35794;
  assign n35811 = n35809 & n35810;
  assign n35812 = n35811 ^ n32620;
  assign n35824 = n35823 ^ n35812;
  assign n35908 = n35808 & n35824;
  assign n35918 = n34386 ^ n33677;
  assign n35919 = n34982 ^ n34386;
  assign n35920 = n35918 & ~n35919;
  assign n35921 = n35920 ^ n33677;
  assign n35916 = n35580 ^ n35544;
  assign n35917 = n35916 ^ n35541;
  assign n35922 = n35921 ^ n35917;
  assign n35913 = n35816 ^ n35815;
  assign n35914 = ~n35821 & n35913;
  assign n35915 = n35914 ^ n35820;
  assign n35923 = n35922 ^ n35915;
  assign n35909 = n35822 ^ n35812;
  assign n35910 = ~n35823 & n35909;
  assign n35911 = n35910 ^ n32610;
  assign n35912 = n35911 ^ n32604;
  assign n35924 = n35923 ^ n35912;
  assign n36232 = n35908 & n35924;
  assign n36158 = n35923 ^ n32604;
  assign n36159 = n35923 ^ n35911;
  assign n36160 = ~n36158 & n36159;
  assign n36161 = n36160 ^ n32604;
  assign n36046 = n35917 ^ n35915;
  assign n36047 = ~n35922 & ~n36046;
  assign n36048 = n36047 ^ n35921;
  assign n36041 = n34380 ^ n33703;
  assign n36042 = n34975 ^ n34380;
  assign n36043 = n36041 & ~n36042;
  assign n36044 = n36043 ^ n33703;
  assign n36155 = n36048 ^ n36044;
  assign n36040 = n35583 ^ n35540;
  assign n36156 = n36155 ^ n36040;
  assign n36157 = n36156 ^ n32598;
  assign n36231 = n36161 ^ n36157;
  assign n36341 = n36232 ^ n36231;
  assign n1070 = n1033 ^ n994;
  assign n1071 = n1070 ^ n1067;
  assign n1078 = n1077 ^ n1071;
  assign n36342 = n36341 ^ n1078;
  assign n35925 = n35924 ^ n35908;
  assign n1037 = n1021 ^ n976;
  assign n1053 = n1052 ^ n1037;
  assign n1060 = n1059 ^ n1053;
  assign n35926 = n35925 ^ n1060;
  assign n35825 = n35824 ^ n35808;
  assign n35826 = n35825 ^ n3323;
  assign n35827 = n35807 ^ n35791;
  assign n35831 = n35830 ^ n35827;
  assign n35832 = n35790 ^ n35773;
  assign n35836 = n35835 ^ n35832;
  assign n35840 = n35789 ^ n35775;
  assign n35837 = n33469 ^ n25754;
  assign n35838 = n35837 ^ n30180;
  assign n35839 = n35838 ^ n729;
  assign n35841 = n35840 ^ n35839;
  assign n35845 = n35788 ^ n35776;
  assign n35842 = n33473 ^ n25798;
  assign n35843 = n35842 ^ n714;
  assign n35844 = n35843 ^ n24741;
  assign n35846 = n35845 ^ n35844;
  assign n35850 = n35787 ^ n35785;
  assign n35847 = n33478 ^ n25791;
  assign n35848 = n35847 ^ n29643;
  assign n35849 = n35848 ^ n563;
  assign n35851 = n35850 ^ n35849;
  assign n35855 = n35784 ^ n35783;
  assign n35852 = n33483 ^ n702;
  assign n35853 = n35852 ^ n29670;
  assign n35854 = n35853 ^ n24748;
  assign n35856 = n35855 ^ n35854;
  assign n35858 = n33489 ^ n25763;
  assign n35859 = n35858 ^ n29649;
  assign n35860 = n35859 ^ n24243;
  assign n35857 = n35782 ^ n35780;
  assign n35861 = n35860 ^ n35857;
  assign n35863 = n24202 ^ n2362;
  assign n35864 = n35863 ^ n29660;
  assign n35865 = n35864 ^ n25768;
  assign n35862 = n35779 ^ n35778;
  assign n35866 = n35865 ^ n35862;
  assign n35867 = n25773 ^ n2344;
  assign n35868 = n35867 ^ n2298;
  assign n35869 = n35868 ^ n24193;
  assign n35870 = n35869 ^ n35778;
  assign n2259 = n2182 ^ n2108;
  assign n2269 = n2268 ^ n2259;
  assign n2273 = n2272 ^ n2269;
  assign n35871 = n35732 ^ n32679;
  assign n35872 = n2273 & ~n35871;
  assign n2283 = n2242 ^ n2192;
  assign n2284 = n2283 ^ n2280;
  assign n2288 = n2287 ^ n2284;
  assign n35873 = n35872 ^ n2288;
  assign n35874 = n35736 ^ n35734;
  assign n35875 = n35874 ^ n2288;
  assign n35876 = n35873 & ~n35875;
  assign n35877 = n35876 ^ n35872;
  assign n35878 = n35877 ^ n35778;
  assign n35879 = ~n35870 & n35878;
  assign n35880 = n35879 ^ n35869;
  assign n35881 = n35880 ^ n35862;
  assign n35882 = n35866 & ~n35881;
  assign n35883 = n35882 ^ n35865;
  assign n35884 = n35883 ^ n35857;
  assign n35885 = ~n35861 & n35884;
  assign n35886 = n35885 ^ n35860;
  assign n35887 = n35886 ^ n35855;
  assign n35888 = n35856 & ~n35887;
  assign n35889 = n35888 ^ n35854;
  assign n35890 = n35889 ^ n35850;
  assign n35891 = n35851 & ~n35890;
  assign n35892 = n35891 ^ n35849;
  assign n35893 = n35892 ^ n35845;
  assign n35894 = ~n35846 & n35893;
  assign n35895 = n35894 ^ n35844;
  assign n35896 = n35895 ^ n35840;
  assign n35897 = n35841 & ~n35896;
  assign n35898 = n35897 ^ n35839;
  assign n35899 = n35898 ^ n35832;
  assign n35900 = ~n35836 & n35899;
  assign n35901 = n35900 ^ n35835;
  assign n35902 = n35901 ^ n35827;
  assign n35903 = n35831 & ~n35902;
  assign n35904 = n35903 ^ n35830;
  assign n35905 = n35904 ^ n35825;
  assign n35906 = ~n35826 & n35905;
  assign n35907 = n35906 ^ n3323;
  assign n36343 = n35925 ^ n35907;
  assign n36344 = ~n35926 & n36343;
  assign n36345 = n36344 ^ n1060;
  assign n36346 = n36345 ^ n36341;
  assign n36347 = ~n36342 & n36346;
  assign n36348 = n36347 ^ n1078;
  assign n36233 = n36231 & n36232;
  assign n36162 = n36161 ^ n36156;
  assign n36163 = ~n36157 & ~n36162;
  assign n36164 = n36163 ^ n32598;
  assign n36229 = n36164 ^ n32592;
  assign n36045 = n36044 ^ n36040;
  assign n36049 = n36048 ^ n36040;
  assign n36050 = ~n36045 & n36049;
  assign n36051 = n36050 ^ n36044;
  assign n36035 = n34374 ^ n33693;
  assign n36036 = n34972 ^ n34374;
  assign n36037 = n36035 & ~n36036;
  assign n36038 = n36037 ^ n33693;
  assign n36033 = n35586 ^ n35534;
  assign n36034 = n36033 ^ n35531;
  assign n36039 = n36038 ^ n36034;
  assign n36153 = n36051 ^ n36039;
  assign n36230 = n36229 ^ n36153;
  assign n36339 = n36233 ^ n36230;
  assign n1195 = n1188 ^ n1116;
  assign n1202 = n1201 ^ n1195;
  assign n1209 = n1208 ^ n1202;
  assign n36340 = n36339 ^ n1209;
  assign n36679 = n36348 ^ n36340;
  assign n36008 = n35601 ^ n35516;
  assign n38048 = n36679 ^ n36008;
  assign n36516 = n34989 ^ n34405;
  assign n36517 = n36034 ^ n34989;
  assign n36518 = n36516 & ~n36517;
  assign n36519 = n36518 ^ n34405;
  assign n36514 = n35883 ^ n35860;
  assign n36515 = n36514 ^ n35857;
  assign n36520 = n36519 ^ n36515;
  assign n36463 = n35880 ^ n35865;
  assign n36464 = n36463 ^ n35862;
  assign n36458 = n34995 ^ n34411;
  assign n36459 = n36040 ^ n34995;
  assign n36460 = ~n36458 & ~n36459;
  assign n36461 = n36460 ^ n34411;
  assign n36510 = n36464 ^ n36461;
  assign n35934 = n35877 ^ n35870;
  assign n35930 = n35002 ^ n33541;
  assign n35931 = n35917 ^ n35002;
  assign n35932 = n35930 & ~n35931;
  assign n35933 = n35932 ^ n33541;
  assign n35935 = n35934 ^ n35933;
  assign n35940 = n35874 ^ n35873;
  assign n35936 = n35008 ^ n34422;
  assign n35937 = n35816 ^ n35008;
  assign n35938 = n35936 & ~n35937;
  assign n35939 = n35938 ^ n34422;
  assign n35941 = n35940 ^ n35939;
  assign n35946 = n35871 ^ n2273;
  assign n35942 = n34428 ^ n34306;
  assign n35943 = n35800 ^ n34306;
  assign n35944 = n35942 & n35943;
  assign n35945 = n35944 ^ n34428;
  assign n35947 = n35946 ^ n35945;
  assign n36406 = n35023 ^ n34434;
  assign n36407 = n35770 ^ n35023;
  assign n36408 = ~n36406 & n36407;
  assign n36409 = n36408 ^ n34434;
  assign n35966 = n35625 ^ n35479;
  assign n35962 = n34114 ^ n33358;
  assign n35963 = n34857 ^ n34114;
  assign n35964 = ~n35962 & ~n35963;
  assign n35965 = n35964 ^ n33358;
  assign n35967 = n35966 ^ n35965;
  assign n35972 = n35622 ^ n35481;
  assign n35968 = n34120 ^ n33368;
  assign n35969 = n35430 ^ n34120;
  assign n35970 = ~n35968 & n35969;
  assign n35971 = n35970 ^ n33368;
  assign n35973 = n35972 ^ n35971;
  assign n35978 = n35619 ^ n35485;
  assign n35979 = n35978 ^ n35482;
  assign n35974 = n34130 ^ n33370;
  assign n35975 = n34900 ^ n34130;
  assign n35976 = ~n35974 & n35975;
  assign n35977 = n35976 ^ n33370;
  assign n35980 = n35979 ^ n35977;
  assign n35983 = n34922 ^ n34149;
  assign n35984 = n34922 ^ n34902;
  assign n35985 = n35983 & n35984;
  assign n35986 = n35985 ^ n34149;
  assign n35981 = n35616 ^ n35489;
  assign n35982 = n35981 ^ n35490;
  assign n35987 = n35986 ^ n35982;
  assign n35992 = n35613 ^ n35496;
  assign n35988 = n34929 ^ n34090;
  assign n35989 = n34929 ^ n34912;
  assign n35990 = n35988 & n35989;
  assign n35991 = n35990 ^ n34090;
  assign n35993 = n35992 ^ n35991;
  assign n35998 = n35610 ^ n35501;
  assign n35994 = n34311 ^ n33545;
  assign n35995 = n34919 ^ n34311;
  assign n35996 = n35994 & ~n35995;
  assign n35997 = n35996 ^ n33545;
  assign n35999 = n35998 ^ n35997;
  assign n36003 = n34333 ^ n33567;
  assign n36004 = n34934 ^ n34333;
  assign n36005 = n36003 & ~n36004;
  assign n36006 = n36005 ^ n33567;
  assign n36001 = n35604 ^ n35509;
  assign n36002 = n36001 ^ n35510;
  assign n36007 = n36006 ^ n36002;
  assign n36009 = n34342 ^ n33576;
  assign n36010 = n34941 ^ n34342;
  assign n36011 = ~n36009 & ~n36010;
  assign n36012 = n36011 ^ n33576;
  assign n36013 = n36012 ^ n36008;
  assign n36018 = n35598 ^ n35520;
  assign n36019 = n36018 ^ n35517;
  assign n36014 = n34348 ^ n33582;
  assign n36015 = n34947 ^ n34348;
  assign n36016 = ~n36014 & ~n36015;
  assign n36017 = n36016 ^ n33582;
  assign n36020 = n36019 ^ n36017;
  assign n36021 = n34359 ^ n33594;
  assign n36022 = n34953 ^ n34359;
  assign n36023 = ~n36021 & n36022;
  assign n36024 = n36023 ^ n33594;
  assign n35928 = n35595 ^ n35523;
  assign n36025 = n36024 ^ n35928;
  assign n36030 = n35592 ^ n35527;
  assign n36031 = n36030 ^ n35524;
  assign n36026 = n34509 ^ n33718;
  assign n36027 = n34959 ^ n34509;
  assign n36028 = n36026 & n36027;
  assign n36029 = n36028 ^ n33718;
  assign n36032 = n36031 ^ n36029;
  assign n36055 = n35589 ^ n35530;
  assign n36052 = n36051 ^ n36034;
  assign n36053 = n36039 & n36052;
  assign n36054 = n36053 ^ n36038;
  assign n36056 = n36055 ^ n36054;
  assign n36057 = n34368 ^ n33713;
  assign n36058 = n34966 ^ n34368;
  assign n36059 = n36057 & ~n36058;
  assign n36060 = n36059 ^ n33713;
  assign n36061 = n36060 ^ n36055;
  assign n36062 = ~n36056 & n36061;
  assign n36063 = n36062 ^ n36060;
  assign n36064 = n36063 ^ n36031;
  assign n36065 = ~n36032 & n36064;
  assign n36066 = n36065 ^ n36029;
  assign n36067 = n36066 ^ n35928;
  assign n36068 = n36025 & n36067;
  assign n36069 = n36068 ^ n36024;
  assign n36070 = n36069 ^ n36019;
  assign n36071 = ~n36020 & n36070;
  assign n36072 = n36071 ^ n36017;
  assign n36073 = n36072 ^ n36008;
  assign n36074 = ~n36013 & n36073;
  assign n36075 = n36074 ^ n36012;
  assign n36076 = n36075 ^ n36002;
  assign n36077 = n36007 & ~n36076;
  assign n36078 = n36077 ^ n36006;
  assign n36000 = n35607 ^ n35506;
  assign n36079 = n36078 ^ n36000;
  assign n36080 = n34323 ^ n33561;
  assign n36081 = n34926 ^ n34323;
  assign n36082 = n36080 & ~n36081;
  assign n36083 = n36082 ^ n33561;
  assign n36084 = n36083 ^ n36000;
  assign n36085 = ~n36079 & ~n36084;
  assign n36086 = n36085 ^ n36083;
  assign n36087 = n36086 ^ n35998;
  assign n36088 = ~n35999 & n36087;
  assign n36089 = n36088 ^ n35997;
  assign n36090 = n36089 ^ n35992;
  assign n36091 = n35993 & ~n36090;
  assign n36092 = n36091 ^ n35991;
  assign n36093 = n36092 ^ n35982;
  assign n36094 = ~n35987 & n36093;
  assign n36095 = n36094 ^ n35986;
  assign n36096 = n36095 ^ n35979;
  assign n36097 = ~n35980 & n36096;
  assign n36098 = n36097 ^ n35977;
  assign n36099 = n36098 ^ n35972;
  assign n36100 = ~n35973 & ~n36099;
  assign n36101 = n36100 ^ n35971;
  assign n36102 = n36101 ^ n35966;
  assign n36103 = ~n35967 & ~n36102;
  assign n36104 = n36103 ^ n35965;
  assign n35960 = n35628 ^ n35477;
  assign n35956 = n34108 ^ n33356;
  assign n35957 = n34864 ^ n34108;
  assign n35958 = ~n35956 & ~n35957;
  assign n35959 = n35958 ^ n33356;
  assign n35961 = n35960 ^ n35959;
  assign n36120 = n36104 ^ n35961;
  assign n36121 = n36120 ^ n32768;
  assign n36122 = n36101 ^ n35967;
  assign n36123 = n36122 ^ n32774;
  assign n36124 = n36098 ^ n35973;
  assign n36125 = n36124 ^ n32495;
  assign n36126 = n36095 ^ n35980;
  assign n36127 = n36126 ^ n32433;
  assign n36128 = n36092 ^ n35986;
  assign n36129 = n36128 ^ n35982;
  assign n36130 = n36129 ^ n33118;
  assign n36131 = n36089 ^ n35993;
  assign n36132 = n36131 ^ n33100;
  assign n36133 = n36086 ^ n35999;
  assign n36134 = n36133 ^ n32524;
  assign n36135 = n36083 ^ n36079;
  assign n36136 = n36135 ^ n32536;
  assign n36137 = n36075 ^ n36006;
  assign n36138 = n36137 ^ n36002;
  assign n36139 = n36138 ^ n32542;
  assign n36142 = n36069 ^ n36017;
  assign n36143 = n36142 ^ n36019;
  assign n36144 = n36143 ^ n32558;
  assign n36145 = n36066 ^ n36024;
  assign n36146 = n36145 ^ n35928;
  assign n36147 = n36146 ^ n32570;
  assign n36148 = n36063 ^ n36029;
  assign n36149 = n36148 ^ n36031;
  assign n36150 = n36149 ^ n32577;
  assign n36151 = n36060 ^ n36056;
  assign n36152 = n36151 ^ n32586;
  assign n36154 = n36153 ^ n32592;
  assign n36165 = n36164 ^ n36153;
  assign n36166 = ~n36154 & ~n36165;
  assign n36167 = n36166 ^ n32592;
  assign n36168 = n36167 ^ n36151;
  assign n36169 = n36152 & ~n36168;
  assign n36170 = n36169 ^ n32586;
  assign n36171 = n36170 ^ n36149;
  assign n36172 = n36150 & n36171;
  assign n36173 = n36172 ^ n32577;
  assign n36174 = n36173 ^ n36146;
  assign n36175 = ~n36147 & n36174;
  assign n36176 = n36175 ^ n32570;
  assign n36177 = n36176 ^ n36143;
  assign n36178 = n36144 & n36177;
  assign n36179 = n36178 ^ n32558;
  assign n36140 = n36072 ^ n36012;
  assign n36141 = n36140 ^ n36008;
  assign n36180 = n36179 ^ n36141;
  assign n36181 = n36141 ^ n32556;
  assign n36182 = ~n36180 & n36181;
  assign n36183 = n36182 ^ n32556;
  assign n36184 = n36183 ^ n36138;
  assign n36185 = ~n36139 & n36184;
  assign n36186 = n36185 ^ n32542;
  assign n36187 = n36186 ^ n36135;
  assign n36188 = n36136 & ~n36187;
  assign n36189 = n36188 ^ n32536;
  assign n36190 = n36189 ^ n36133;
  assign n36191 = n36134 & n36190;
  assign n36192 = n36191 ^ n32524;
  assign n36193 = n36192 ^ n36131;
  assign n36194 = n36132 & n36193;
  assign n36195 = n36194 ^ n33100;
  assign n36196 = n36195 ^ n36129;
  assign n36197 = ~n36130 & n36196;
  assign n36198 = n36197 ^ n33118;
  assign n36199 = n36198 ^ n36126;
  assign n36200 = ~n36127 & n36199;
  assign n36201 = n36200 ^ n32433;
  assign n36202 = n36201 ^ n36124;
  assign n36203 = ~n36125 & n36202;
  assign n36204 = n36203 ^ n32495;
  assign n36205 = n36204 ^ n36122;
  assign n36206 = ~n36123 & ~n36205;
  assign n36207 = n36206 ^ n32774;
  assign n36208 = n36207 ^ n36120;
  assign n36209 = n36121 & ~n36208;
  assign n36210 = n36209 ^ n32768;
  assign n36216 = n36210 ^ n32762;
  assign n36105 = n36104 ^ n35960;
  assign n36106 = ~n35961 & n36105;
  assign n36107 = n36106 ^ n35959;
  assign n35951 = n34167 ^ n33350;
  assign n35952 = n34847 ^ n34167;
  assign n35953 = n35951 & ~n35952;
  assign n35954 = n35953 ^ n33350;
  assign n36117 = n36107 ^ n35954;
  assign n35949 = n35631 ^ n2892;
  assign n35950 = n35949 ^ n35474;
  assign n36118 = n36117 ^ n35950;
  assign n36217 = n36216 ^ n36118;
  assign n36218 = n36207 ^ n32768;
  assign n36219 = n36218 ^ n36120;
  assign n36220 = n36201 ^ n32495;
  assign n36221 = n36220 ^ n36124;
  assign n36222 = n36198 ^ n36127;
  assign n36223 = n36192 ^ n36132;
  assign n36224 = n36189 ^ n32524;
  assign n36225 = n36224 ^ n36133;
  assign n36226 = n36176 ^ n32558;
  assign n36227 = n36226 ^ n36143;
  assign n36228 = n36167 ^ n36152;
  assign n36234 = n36230 & ~n36233;
  assign n36235 = ~n36228 & ~n36234;
  assign n36236 = n36170 ^ n36150;
  assign n36237 = n36235 & ~n36236;
  assign n36238 = n36173 ^ n32570;
  assign n36239 = n36238 ^ n36146;
  assign n36240 = n36237 & ~n36239;
  assign n36241 = ~n36227 & ~n36240;
  assign n36242 = n36180 ^ n32556;
  assign n36243 = ~n36241 & ~n36242;
  assign n36244 = n36183 ^ n32542;
  assign n36245 = n36244 ^ n36138;
  assign n36246 = n36243 & n36245;
  assign n36247 = n36186 ^ n32536;
  assign n36248 = n36247 ^ n36135;
  assign n36249 = ~n36246 & n36248;
  assign n36250 = n36225 & n36249;
  assign n36251 = ~n36223 & n36250;
  assign n36252 = n36195 ^ n36130;
  assign n36253 = ~n36251 & n36252;
  assign n36254 = n36222 & n36253;
  assign n36255 = n36221 & n36254;
  assign n36256 = n36204 ^ n36123;
  assign n36257 = n36255 & n36256;
  assign n36258 = ~n36219 & ~n36257;
  assign n36259 = ~n36217 & n36258;
  assign n36119 = n36118 ^ n32762;
  assign n36211 = n36210 ^ n36118;
  assign n36212 = n36119 & n36211;
  assign n36213 = n36212 ^ n32762;
  assign n36214 = n36213 ^ n32687;
  assign n36112 = n34200 ^ n32511;
  assign n36113 = n35109 ^ n34200;
  assign n36114 = n36112 & n36113;
  assign n36115 = n36114 ^ n32511;
  assign n35955 = n35954 ^ n35950;
  assign n36108 = n36107 ^ n35950;
  assign n36109 = n35955 & ~n36108;
  assign n36110 = n36109 ^ n35954;
  assign n35948 = n35634 ^ n35473;
  assign n36111 = n36110 ^ n35948;
  assign n36116 = n36115 ^ n36111;
  assign n36215 = n36214 ^ n36116;
  assign n36278 = n36259 ^ n36215;
  assign n36282 = n36281 ^ n36278;
  assign n36286 = n36258 ^ n36217;
  assign n36283 = n33940 ^ n26111;
  assign n36284 = n36283 ^ n1766;
  assign n36285 = n36284 ^ n24699;
  assign n36287 = n36286 ^ n36285;
  assign n36291 = n36257 ^ n36219;
  assign n36288 = n33944 ^ n26116;
  assign n36289 = n36288 ^ n30136;
  assign n36290 = n36289 ^ n1761;
  assign n36292 = n36291 ^ n36290;
  assign n36293 = n36256 ^ n36255;
  assign n1671 = n1670 ^ n1655;
  assign n1690 = n1689 ^ n1671;
  assign n1697 = n1696 ^ n1690;
  assign n36294 = n36293 ^ n1697;
  assign n36298 = n36254 ^ n36221;
  assign n36295 = n33951 ^ n26123;
  assign n36296 = n36295 ^ n3009;
  assign n36297 = n36296 ^ n1684;
  assign n36299 = n36298 ^ n36297;
  assign n36300 = n36253 ^ n36222;
  assign n2997 = n2930 ^ n1547;
  assign n2998 = n2997 ^ n2994;
  assign n3002 = n3001 ^ n2998;
  assign n36301 = n36300 ^ n3002;
  assign n36302 = n36252 ^ n36251;
  assign n36303 = n36302 ^ n2987;
  assign n36305 = n3235 ^ n2853;
  assign n36306 = n36305 ^ n30149;
  assign n36307 = n36306 ^ n2981;
  assign n36304 = n36250 ^ n36223;
  assign n36308 = n36307 ^ n36304;
  assign n36309 = n36249 ^ n36225;
  assign n36313 = n36312 ^ n36309;
  assign n36315 = n34007 ^ n3221;
  assign n36316 = n36315 ^ n2588;
  assign n36317 = n36316 ^ n3086;
  assign n36314 = n36248 ^ n36246;
  assign n36318 = n36317 ^ n36314;
  assign n36319 = n36245 ^ n36243;
  assign n3066 = n3065 ^ n3059;
  assign n3070 = n3069 ^ n3066;
  assign n3071 = n3070 ^ n2586;
  assign n36320 = n36319 ^ n3071;
  assign n36321 = n36242 ^ n36241;
  assign n2505 = n2504 ^ n2492;
  assign n2524 = n2523 ^ n2505;
  assign n2531 = n2530 ^ n2524;
  assign n36322 = n36321 ^ n2531;
  assign n36326 = n36240 ^ n36227;
  assign n36323 = n34018 ^ n3045;
  assign n36324 = n36323 ^ n3155;
  assign n36325 = n36324 ^ n2518;
  assign n36327 = n36326 ^ n36325;
  assign n36329 = n34023 ^ n2448;
  assign n36330 = n36329 ^ n30220;
  assign n36331 = n36330 ^ n3153;
  assign n36328 = n36239 ^ n36237;
  assign n36332 = n36331 ^ n36328;
  assign n36335 = n33961 ^ n25835;
  assign n36336 = n36335 ^ n1216;
  assign n36337 = n36336 ^ n1396;
  assign n36334 = n36234 ^ n36228;
  assign n36338 = n36337 ^ n36334;
  assign n36349 = n36348 ^ n36339;
  assign n36350 = ~n36340 & n36349;
  assign n36351 = n36350 ^ n1209;
  assign n36352 = n36351 ^ n36334;
  assign n36353 = ~n36338 & n36352;
  assign n36354 = n36353 ^ n36337;
  assign n36333 = n36236 ^ n36235;
  assign n36355 = n36354 ^ n36333;
  assign n1389 = n1388 ^ n1301;
  assign n1402 = n1401 ^ n1389;
  assign n1409 = n1408 ^ n1402;
  assign n36356 = n36333 ^ n1409;
  assign n36357 = ~n36355 & n36356;
  assign n36358 = n36357 ^ n1409;
  assign n36359 = n36358 ^ n36328;
  assign n36360 = n36332 & ~n36359;
  assign n36361 = n36360 ^ n36331;
  assign n36362 = n36361 ^ n36326;
  assign n36363 = n36327 & ~n36362;
  assign n36364 = n36363 ^ n36325;
  assign n36365 = n36364 ^ n36321;
  assign n36366 = ~n36322 & n36365;
  assign n36367 = n36366 ^ n2531;
  assign n36368 = n36367 ^ n36319;
  assign n36369 = ~n36320 & n36368;
  assign n36370 = n36369 ^ n3071;
  assign n36371 = n36370 ^ n36314;
  assign n36372 = ~n36318 & n36371;
  assign n36373 = n36372 ^ n36317;
  assign n36374 = n36373 ^ n36309;
  assign n36375 = n36313 & ~n36374;
  assign n36376 = n36375 ^ n36312;
  assign n36377 = n36376 ^ n36304;
  assign n36378 = ~n36308 & n36377;
  assign n36379 = n36378 ^ n36307;
  assign n36380 = n36379 ^ n36302;
  assign n36381 = n36303 & ~n36380;
  assign n36382 = n36381 ^ n2987;
  assign n36383 = n36382 ^ n36300;
  assign n36384 = ~n36301 & n36383;
  assign n36385 = n36384 ^ n3002;
  assign n36386 = n36385 ^ n36298;
  assign n36387 = ~n36299 & n36386;
  assign n36388 = n36387 ^ n36297;
  assign n36389 = n36388 ^ n36293;
  assign n36390 = ~n36294 & n36389;
  assign n36391 = n36390 ^ n1697;
  assign n36392 = n36391 ^ n36291;
  assign n36393 = n36292 & ~n36392;
  assign n36394 = n36393 ^ n36290;
  assign n36395 = n36394 ^ n36286;
  assign n36396 = ~n36287 & n36395;
  assign n36397 = n36396 ^ n36285;
  assign n36398 = n36397 ^ n36278;
  assign n36399 = n36282 & ~n36398;
  assign n36400 = n36399 ^ n36281;
  assign n36404 = n36403 ^ n36400;
  assign n36271 = n36116 ^ n32687;
  assign n36272 = n36213 ^ n36116;
  assign n36273 = n36271 & n36272;
  assign n36274 = n36273 ^ n32687;
  assign n36275 = n36274 ^ n32681;
  assign n36267 = n36115 ^ n35948;
  assign n36268 = n36111 & ~n36267;
  assign n36269 = n36268 ^ n36115;
  assign n36265 = n35637 ^ n35468;
  assign n36261 = n34228 ^ n32504;
  assign n36262 = n35103 ^ n34228;
  assign n36263 = ~n36261 & n36262;
  assign n36264 = n36263 ^ n32504;
  assign n36266 = n36265 ^ n36264;
  assign n36270 = n36269 ^ n36266;
  assign n36276 = n36275 ^ n36270;
  assign n36260 = n36215 & n36259;
  assign n36277 = n36276 ^ n36260;
  assign n36405 = n36404 ^ n36277;
  assign n36410 = n36409 ^ n36405;
  assign n36415 = n36397 ^ n36282;
  assign n36411 = n34894 ^ n34436;
  assign n36412 = n35716 ^ n34894;
  assign n36413 = ~n36411 & n36412;
  assign n36414 = n36413 ^ n34436;
  assign n36416 = n36415 ^ n36414;
  assign n36419 = n35137 ^ n34442;
  assign n36420 = n35137 ^ n34889;
  assign n36421 = ~n36419 & ~n36420;
  assign n36422 = n36421 ^ n34442;
  assign n36417 = n36394 ^ n36285;
  assign n36418 = n36417 ^ n36286;
  assign n36423 = n36422 ^ n36418;
  assign n36428 = n36391 ^ n36292;
  assign n36424 = n35035 ^ n34448;
  assign n36425 = n35035 ^ n34891;
  assign n36426 = n36424 & ~n36425;
  assign n36427 = n36426 ^ n34448;
  assign n36429 = n36428 ^ n36427;
  assign n36430 = n35041 ^ n34292;
  assign n36431 = n35041 ^ n34898;
  assign n36432 = ~n36430 & ~n36431;
  assign n36433 = n36432 ^ n34292;
  assign n36434 = n36388 ^ n1697;
  assign n36435 = n36434 ^ n36293;
  assign n36436 = n36433 & ~n36435;
  assign n36437 = n36436 ^ n36428;
  assign n36438 = ~n36429 & n36437;
  assign n36439 = n36438 ^ n36436;
  assign n36440 = n36439 ^ n36418;
  assign n36441 = n36423 & n36440;
  assign n36442 = n36441 ^ n36422;
  assign n36443 = n36442 ^ n36415;
  assign n36444 = n36416 & n36443;
  assign n36445 = n36444 ^ n36414;
  assign n36446 = n36445 ^ n36405;
  assign n36447 = ~n36410 & n36446;
  assign n36448 = n36447 ^ n36409;
  assign n36449 = n36448 ^ n35946;
  assign n36450 = n35947 & n36449;
  assign n36451 = n36450 ^ n35945;
  assign n36452 = n36451 ^ n35940;
  assign n36453 = ~n35941 & n36452;
  assign n36454 = n36453 ^ n35939;
  assign n36455 = n36454 ^ n35934;
  assign n36456 = ~n35935 & ~n36455;
  assign n36457 = n36456 ^ n35933;
  assign n36511 = n36464 ^ n36457;
  assign n36512 = ~n36510 & ~n36511;
  assign n36513 = n36512 ^ n36461;
  assign n36521 = n36520 ^ n36513;
  assign n36522 = n36521 ^ n33672;
  assign n36462 = n36461 ^ n36457;
  assign n36465 = n36464 ^ n36462;
  assign n36466 = n36465 ^ n33600;
  assign n36467 = n36454 ^ n35935;
  assign n36468 = n36467 ^ n33542;
  assign n36469 = n36451 ^ n35939;
  assign n36470 = n36469 ^ n35940;
  assign n36471 = n36470 ^ n33611;
  assign n36472 = n36448 ^ n35947;
  assign n36473 = n36472 ^ n33617;
  assign n36474 = n36445 ^ n36410;
  assign n36475 = n36474 ^ n33634;
  assign n36476 = n36442 ^ n36414;
  assign n36477 = n36476 ^ n36415;
  assign n36478 = n36477 ^ n33627;
  assign n36479 = n36439 ^ n36423;
  assign n36480 = n36479 ^ n33531;
  assign n36481 = n36435 ^ n36433;
  assign n36482 = n33398 & ~n36481;
  assign n36483 = n36482 ^ n33442;
  assign n36484 = n36436 ^ n36427;
  assign n36485 = n36484 ^ n36428;
  assign n36486 = n36485 ^ n36482;
  assign n36487 = n36483 & ~n36486;
  assign n36488 = n36487 ^ n33442;
  assign n36489 = n36488 ^ n36479;
  assign n36490 = n36480 & ~n36489;
  assign n36491 = n36490 ^ n33531;
  assign n36492 = n36491 ^ n36477;
  assign n36493 = ~n36478 & n36492;
  assign n36494 = n36493 ^ n33627;
  assign n36495 = n36494 ^ n36474;
  assign n36496 = n36475 & n36495;
  assign n36497 = n36496 ^ n33634;
  assign n36498 = n36497 ^ n36472;
  assign n36499 = ~n36473 & n36498;
  assign n36500 = n36499 ^ n33617;
  assign n36501 = n36500 ^ n36470;
  assign n36502 = n36471 & n36501;
  assign n36503 = n36502 ^ n33611;
  assign n36504 = n36503 ^ n36467;
  assign n36505 = n36468 & ~n36504;
  assign n36506 = n36505 ^ n33542;
  assign n36507 = n36506 ^ n36465;
  assign n36508 = ~n36466 & n36507;
  assign n36509 = n36508 ^ n33600;
  assign n36523 = n36522 ^ n36509;
  assign n36524 = n36506 ^ n33600;
  assign n36525 = n36524 ^ n36465;
  assign n36526 = n36491 ^ n36478;
  assign n36527 = n36488 ^ n33531;
  assign n36528 = n36527 ^ n36479;
  assign n36529 = n36526 & ~n36528;
  assign n36530 = n36494 ^ n33634;
  assign n36531 = n36530 ^ n36474;
  assign n36532 = n36529 & ~n36531;
  assign n36533 = n36497 ^ n36473;
  assign n36534 = ~n36532 & n36533;
  assign n36535 = n36500 ^ n33611;
  assign n36536 = n36535 ^ n36470;
  assign n36537 = ~n36534 & n36536;
  assign n36538 = n36503 ^ n36468;
  assign n36539 = n36537 & ~n36538;
  assign n36540 = ~n36525 & ~n36539;
  assign n36617 = n36523 & n36540;
  assign n36629 = n36521 ^ n36509;
  assign n36630 = n36522 & ~n36629;
  assign n36631 = n36630 ^ n33672;
  assign n36632 = n36631 ^ n33666;
  assign n36625 = n36515 ^ n36513;
  assign n36626 = ~n36520 & ~n36625;
  assign n36627 = n36626 ^ n36519;
  assign n36622 = n35886 ^ n35854;
  assign n36623 = n36622 ^ n35855;
  assign n36618 = n34982 ^ n34395;
  assign n36619 = n36055 ^ n34982;
  assign n36620 = n36618 & n36619;
  assign n36621 = n36620 ^ n34395;
  assign n36624 = n36623 ^ n36621;
  assign n36628 = n36627 ^ n36624;
  assign n36633 = n36632 ^ n36628;
  assign n36895 = ~n36617 & n36633;
  assign n36825 = n36631 ^ n36628;
  assign n36826 = n36632 & n36825;
  assign n36827 = n36826 ^ n33666;
  assign n36736 = n36627 ^ n36623;
  assign n36737 = n36627 ^ n36621;
  assign n36738 = n36736 & n36737;
  assign n36739 = n36738 ^ n36623;
  assign n36731 = n34975 ^ n34388;
  assign n36732 = n36031 ^ n34975;
  assign n36733 = n36731 & ~n36732;
  assign n36734 = n36733 ^ n34388;
  assign n36730 = n35889 ^ n35851;
  assign n36735 = n36734 ^ n36730;
  assign n36823 = n36739 ^ n36735;
  assign n36824 = n36823 ^ n33688;
  assign n36894 = n36827 ^ n36824;
  assign n36996 = n36895 ^ n36894;
  assign n37000 = n36999 ^ n36996;
  assign n36634 = n36633 ^ n36617;
  assign n36614 = n34769 ^ n26526;
  assign n36615 = n36614 ^ n30469;
  assign n36616 = n36615 ^ n807;
  assign n36635 = n36634 ^ n36616;
  assign n36541 = n36540 ^ n36523;
  assign n739 = n738 ^ n732;
  assign n669 = n668 ^ n632;
  assign n740 = n739 ^ n669;
  assign n36542 = n36541 ^ n740;
  assign n36545 = n34236 ^ n581;
  assign n36546 = n36545 ^ n30501;
  assign n36547 = n36546 ^ n3290;
  assign n36544 = n36538 ^ n36537;
  assign n36548 = n36547 ^ n36544;
  assign n36549 = n36536 ^ n36534;
  assign n36553 = n36552 ^ n36549;
  assign n36555 = n34246 ^ n26544;
  assign n36556 = n36555 ^ n30511;
  assign n36557 = n36556 ^ n25035;
  assign n36554 = n36533 ^ n36532;
  assign n36558 = n36557 ^ n36554;
  assign n36562 = n36531 ^ n36529;
  assign n36559 = n34250 ^ n26562;
  assign n36560 = n36559 ^ n30534;
  assign n36561 = n36560 ^ n25010;
  assign n36563 = n36562 ^ n36561;
  assign n36565 = n34264 ^ n2330;
  assign n36566 = n36565 ^ n2393;
  assign n36567 = n36566 ^ n30518;
  assign n36568 = n36567 ^ n36528;
  assign n36572 = n35101 ^ n2377;
  assign n36573 = n36572 ^ n2126;
  assign n36574 = n36573 ^ n30971;
  assign n36575 = n36481 ^ n33398;
  assign n36576 = n36574 & ~n36575;
  assign n36569 = n34259 ^ n2370;
  assign n36570 = n36569 ^ n25019;
  assign n36571 = n36570 ^ n2135;
  assign n36577 = n36576 ^ n36571;
  assign n36578 = n36485 ^ n36483;
  assign n36579 = n36578 ^ n36571;
  assign n36580 = n36577 & ~n36579;
  assign n36581 = n36580 ^ n36576;
  assign n36582 = n36581 ^ n36528;
  assign n36583 = ~n36568 & n36582;
  assign n36584 = n36583 ^ n36567;
  assign n36564 = n36528 ^ n36526;
  assign n36585 = n36584 ^ n36564;
  assign n36586 = n34255 ^ n26556;
  assign n36587 = n36586 ^ n25015;
  assign n36588 = n36587 ^ n30526;
  assign n36589 = n36588 ^ n36564;
  assign n36590 = ~n36585 & n36589;
  assign n36591 = n36590 ^ n36588;
  assign n36592 = n36591 ^ n36562;
  assign n36593 = n36563 & ~n36592;
  assign n36594 = n36593 ^ n36561;
  assign n36595 = n36594 ^ n36554;
  assign n36596 = ~n36558 & n36595;
  assign n36597 = n36596 ^ n36557;
  assign n36598 = n36597 ^ n36549;
  assign n36599 = n36553 & ~n36598;
  assign n36600 = n36599 ^ n36552;
  assign n36601 = n36600 ^ n36544;
  assign n36602 = n36548 & ~n36601;
  assign n36603 = n36602 ^ n36547;
  assign n36543 = n36539 ^ n36525;
  assign n36604 = n36603 ^ n36543;
  assign n36605 = n34287 ^ n26531;
  assign n36606 = n36605 ^ n30496;
  assign n36607 = n36606 ^ n627;
  assign n36608 = n36607 ^ n36543;
  assign n36609 = ~n36604 & n36608;
  assign n36610 = n36609 ^ n36607;
  assign n36611 = n36610 ^ n36541;
  assign n36612 = n36542 & ~n36611;
  assign n36613 = n36612 ^ n740;
  assign n37001 = n36634 ^ n36613;
  assign n37002 = n36635 & ~n37001;
  assign n37003 = n37002 ^ n36616;
  assign n37004 = n37003 ^ n36996;
  assign n37005 = ~n37000 & n37004;
  assign n37006 = n37005 ^ n36999;
  assign n36828 = n36827 ^ n36823;
  assign n36829 = ~n36824 & n36828;
  assign n36830 = n36829 ^ n33688;
  assign n36897 = n36830 ^ n33677;
  assign n36740 = n36739 ^ n36730;
  assign n36741 = ~n36735 & ~n36740;
  assign n36742 = n36741 ^ n36734;
  assign n36725 = n34972 ^ n34386;
  assign n36726 = n35928 ^ n34972;
  assign n36727 = ~n36725 & n36726;
  assign n36728 = n36727 ^ n34386;
  assign n36820 = n36742 ^ n36728;
  assign n36723 = n35892 ^ n35844;
  assign n36724 = n36723 ^ n35845;
  assign n36821 = n36820 ^ n36724;
  assign n36898 = n36897 ^ n36821;
  assign n36896 = n36894 & n36895;
  assign n36995 = n36898 ^ n36896;
  assign n37007 = n37006 ^ n36995;
  assign n37358 = n37010 ^ n37007;
  assign n38049 = n37358 ^ n36679;
  assign n38050 = ~n38048 & n38049;
  assign n38051 = n38050 ^ n36008;
  assign n37193 = n35816 ^ n35023;
  assign n37194 = n36515 ^ n35816;
  assign n37195 = n37193 & ~n37194;
  assign n37196 = n37195 ^ n35023;
  assign n37085 = n36379 ^ n2987;
  assign n37086 = n37085 ^ n36302;
  assign n36945 = n36376 ^ n36308;
  assign n36940 = n35109 ^ n34108;
  assign n36941 = n35673 ^ n35109;
  assign n36942 = n36940 & n36941;
  assign n36943 = n36942 ^ n34108;
  assign n37080 = n36945 ^ n36943;
  assign n36886 = n36373 ^ n36312;
  assign n36887 = n36886 ^ n36309;
  assign n36881 = n34847 ^ n34114;
  assign n36882 = n35680 ^ n34847;
  assign n36883 = ~n36881 & n36882;
  assign n36884 = n36883 ^ n34114;
  assign n36936 = n36887 ^ n36884;
  assign n36789 = n36370 ^ n36317;
  assign n36790 = n36789 ^ n36314;
  assign n36785 = n34864 ^ n34120;
  assign n36786 = n36265 ^ n34864;
  assign n36787 = ~n36785 & n36786;
  assign n36788 = n36787 ^ n34120;
  assign n36791 = n36790 ^ n36788;
  assign n36644 = n36367 ^ n3071;
  assign n36645 = n36644 ^ n36319;
  assign n36640 = n34857 ^ n34130;
  assign n36641 = n35948 ^ n34857;
  assign n36642 = n36640 & ~n36641;
  assign n36643 = n36642 ^ n34130;
  assign n36646 = n36645 ^ n36643;
  assign n36649 = n35430 ^ n34922;
  assign n36650 = n35950 ^ n35430;
  assign n36651 = ~n36649 & n36650;
  assign n36652 = n36651 ^ n34922;
  assign n36647 = n36364 ^ n2531;
  assign n36648 = n36647 ^ n36321;
  assign n36653 = n36652 ^ n36648;
  assign n36655 = n34929 ^ n34900;
  assign n36656 = n35960 ^ n34900;
  assign n36657 = n36655 & n36656;
  assign n36658 = n36657 ^ n34929;
  assign n36654 = n36361 ^ n36327;
  assign n36659 = n36658 ^ n36654;
  assign n36664 = n36358 ^ n36332;
  assign n36660 = n34902 ^ n34311;
  assign n36661 = n35966 ^ n34902;
  assign n36662 = ~n36660 & ~n36661;
  assign n36663 = n36662 ^ n34311;
  assign n36665 = n36664 ^ n36663;
  assign n36670 = n36355 ^ n1409;
  assign n36666 = n34912 ^ n34323;
  assign n36667 = n35972 ^ n34912;
  assign n36668 = ~n36666 & n36667;
  assign n36669 = n36668 ^ n34323;
  assign n36671 = n36670 ^ n36669;
  assign n36674 = n34919 ^ n34333;
  assign n36675 = n35979 ^ n34919;
  assign n36676 = ~n36674 & n36675;
  assign n36677 = n36676 ^ n34333;
  assign n36672 = n36351 ^ n36337;
  assign n36673 = n36672 ^ n36334;
  assign n36678 = n36677 ^ n36673;
  assign n36680 = n34926 ^ n34342;
  assign n36681 = n35982 ^ n34926;
  assign n36682 = n36680 & n36681;
  assign n36683 = n36682 ^ n34342;
  assign n36684 = n36683 ^ n36679;
  assign n36687 = n34934 ^ n34348;
  assign n36688 = n35992 ^ n34934;
  assign n36689 = ~n36687 & n36688;
  assign n36690 = n36689 ^ n34348;
  assign n36685 = n36345 ^ n1078;
  assign n36686 = n36685 ^ n36341;
  assign n36691 = n36690 ^ n36686;
  assign n36692 = n34941 ^ n34359;
  assign n36693 = n35998 ^ n34941;
  assign n36694 = n36692 & n36693;
  assign n36695 = n36694 ^ n34359;
  assign n35927 = n35926 ^ n35907;
  assign n36696 = n36695 ^ n35927;
  assign n36701 = n35904 ^ n3323;
  assign n36702 = n36701 ^ n35825;
  assign n36697 = n34947 ^ n34509;
  assign n36698 = n36000 ^ n34947;
  assign n36699 = n36697 & n36698;
  assign n36700 = n36699 ^ n34509;
  assign n36703 = n36702 ^ n36700;
  assign n36708 = n35901 ^ n35831;
  assign n36704 = n34953 ^ n34368;
  assign n36705 = n36002 ^ n34953;
  assign n36706 = ~n36704 & ~n36705;
  assign n36707 = n36706 ^ n34368;
  assign n36709 = n36708 ^ n36707;
  assign n36714 = n35898 ^ n35835;
  assign n36715 = n36714 ^ n35832;
  assign n36710 = n34959 ^ n34374;
  assign n36711 = n36008 ^ n34959;
  assign n36712 = ~n36710 & n36711;
  assign n36713 = n36712 ^ n34374;
  assign n36716 = n36715 ^ n36713;
  assign n36718 = n34966 ^ n34380;
  assign n36719 = n36019 ^ n34966;
  assign n36720 = ~n36718 & ~n36719;
  assign n36721 = n36720 ^ n34380;
  assign n36717 = n35895 ^ n35841;
  assign n36722 = n36721 ^ n36717;
  assign n36729 = n36728 ^ n36724;
  assign n36743 = n36742 ^ n36724;
  assign n36744 = n36729 & ~n36743;
  assign n36745 = n36744 ^ n36728;
  assign n36746 = n36745 ^ n36717;
  assign n36747 = ~n36722 & n36746;
  assign n36748 = n36747 ^ n36721;
  assign n36749 = n36748 ^ n36715;
  assign n36750 = ~n36716 & ~n36749;
  assign n36751 = n36750 ^ n36713;
  assign n36752 = n36751 ^ n36708;
  assign n36753 = n36709 & ~n36752;
  assign n36754 = n36753 ^ n36707;
  assign n36755 = n36754 ^ n36702;
  assign n36756 = ~n36703 & n36755;
  assign n36757 = n36756 ^ n36700;
  assign n36758 = n36757 ^ n35927;
  assign n36759 = ~n36696 & n36758;
  assign n36760 = n36759 ^ n36695;
  assign n36761 = n36760 ^ n36686;
  assign n36762 = ~n36691 & n36761;
  assign n36763 = n36762 ^ n36690;
  assign n36764 = n36763 ^ n36679;
  assign n36765 = ~n36684 & n36764;
  assign n36766 = n36765 ^ n36683;
  assign n36767 = n36766 ^ n36673;
  assign n36768 = n36678 & n36767;
  assign n36769 = n36768 ^ n36677;
  assign n36770 = n36769 ^ n36670;
  assign n36771 = n36671 & n36770;
  assign n36772 = n36771 ^ n36669;
  assign n36773 = n36772 ^ n36664;
  assign n36774 = n36665 & ~n36773;
  assign n36775 = n36774 ^ n36663;
  assign n36776 = n36775 ^ n36654;
  assign n36777 = n36659 & ~n36776;
  assign n36778 = n36777 ^ n36658;
  assign n36779 = n36778 ^ n36648;
  assign n36780 = ~n36653 & n36779;
  assign n36781 = n36780 ^ n36652;
  assign n36782 = n36781 ^ n36645;
  assign n36783 = n36646 & n36782;
  assign n36784 = n36783 ^ n36643;
  assign n36878 = n36790 ^ n36784;
  assign n36879 = ~n36791 & ~n36878;
  assign n36880 = n36879 ^ n36788;
  assign n36937 = n36887 ^ n36880;
  assign n36938 = ~n36936 & ~n36937;
  assign n36939 = n36938 ^ n36884;
  assign n37081 = n36945 ^ n36939;
  assign n37082 = n37080 & ~n37081;
  assign n37083 = n37082 ^ n36943;
  assign n37076 = n35103 ^ n34167;
  assign n37077 = n35667 ^ n35103;
  assign n37078 = n37076 & n37077;
  assign n37079 = n37078 ^ n34167;
  assign n37084 = n37083 ^ n37079;
  assign n37087 = n37086 ^ n37084;
  assign n37139 = n37087 ^ n33350;
  assign n36944 = n36943 ^ n36939;
  assign n36946 = n36945 ^ n36944;
  assign n37071 = n36946 ^ n33356;
  assign n36885 = n36884 ^ n36880;
  assign n36888 = n36887 ^ n36885;
  assign n36889 = n36888 ^ n33358;
  assign n36792 = n36791 ^ n36784;
  assign n36793 = n36792 ^ n33368;
  assign n36794 = n36781 ^ n36646;
  assign n36795 = n36794 ^ n33370;
  assign n36796 = n36778 ^ n36652;
  assign n36797 = n36796 ^ n36648;
  assign n36798 = n36797 ^ n34149;
  assign n36799 = n36772 ^ n36665;
  assign n36800 = n36799 ^ n33545;
  assign n36801 = n36769 ^ n36671;
  assign n36802 = n36801 ^ n33561;
  assign n36803 = n36766 ^ n36678;
  assign n36804 = n36803 ^ n33567;
  assign n36805 = n36763 ^ n36683;
  assign n36806 = n36805 ^ n36679;
  assign n36807 = n36806 ^ n33576;
  assign n36808 = n36760 ^ n36691;
  assign n36809 = n36808 ^ n33582;
  assign n36810 = n36757 ^ n36696;
  assign n36811 = n36810 ^ n33594;
  assign n36812 = n36754 ^ n36703;
  assign n36813 = n36812 ^ n33718;
  assign n36814 = n36751 ^ n36709;
  assign n36815 = n36814 ^ n33713;
  assign n36816 = n36748 ^ n36716;
  assign n36817 = n36816 ^ n33693;
  assign n36818 = n36745 ^ n36722;
  assign n36819 = n36818 ^ n33703;
  assign n36822 = n36821 ^ n33677;
  assign n36831 = n36830 ^ n36821;
  assign n36832 = n36822 & n36831;
  assign n36833 = n36832 ^ n33677;
  assign n36834 = n36833 ^ n36818;
  assign n36835 = ~n36819 & n36834;
  assign n36836 = n36835 ^ n33703;
  assign n36837 = n36836 ^ n36816;
  assign n36838 = n36817 & n36837;
  assign n36839 = n36838 ^ n33693;
  assign n36840 = n36839 ^ n36814;
  assign n36841 = n36815 & ~n36840;
  assign n36842 = n36841 ^ n33713;
  assign n36843 = n36842 ^ n36812;
  assign n36844 = ~n36813 & n36843;
  assign n36845 = n36844 ^ n33718;
  assign n36846 = n36845 ^ n36810;
  assign n36847 = n36811 & n36846;
  assign n36848 = n36847 ^ n33594;
  assign n36849 = n36848 ^ n36808;
  assign n36850 = n36809 & ~n36849;
  assign n36851 = n36850 ^ n33582;
  assign n36852 = n36851 ^ n36806;
  assign n36853 = n36807 & ~n36852;
  assign n36854 = n36853 ^ n33576;
  assign n36855 = n36854 ^ n36803;
  assign n36856 = ~n36804 & n36855;
  assign n36857 = n36856 ^ n33567;
  assign n36858 = n36857 ^ n36801;
  assign n36859 = ~n36802 & ~n36858;
  assign n36860 = n36859 ^ n33561;
  assign n36861 = n36860 ^ n36799;
  assign n36862 = n36800 & ~n36861;
  assign n36863 = n36862 ^ n33545;
  assign n36864 = n36863 ^ n34090;
  assign n36865 = n36775 ^ n36659;
  assign n36866 = n36865 ^ n36863;
  assign n36867 = n36864 & ~n36866;
  assign n36868 = n36867 ^ n34090;
  assign n36869 = n36868 ^ n36797;
  assign n36870 = ~n36798 & n36869;
  assign n36871 = n36870 ^ n34149;
  assign n36872 = n36871 ^ n36794;
  assign n36873 = n36795 & ~n36872;
  assign n36874 = n36873 ^ n33370;
  assign n36875 = n36874 ^ n36792;
  assign n36876 = ~n36793 & ~n36875;
  assign n36877 = n36876 ^ n33368;
  assign n36932 = n36888 ^ n36877;
  assign n36933 = ~n36889 & ~n36932;
  assign n36934 = n36933 ^ n33358;
  assign n37072 = n36946 ^ n36934;
  assign n37073 = ~n37071 & n37072;
  assign n37074 = n37073 ^ n33356;
  assign n37140 = n37087 ^ n37074;
  assign n37141 = ~n37139 & n37140;
  assign n37142 = n37141 ^ n33350;
  assign n37143 = n37142 ^ n32511;
  assign n37134 = n35049 ^ n34200;
  assign n37135 = n35660 ^ n35049;
  assign n37136 = n37134 & n37135;
  assign n37137 = n37136 ^ n34200;
  assign n37132 = n36382 ^ n36301;
  assign n37128 = n37086 ^ n37079;
  assign n37129 = n37086 ^ n37083;
  assign n37130 = n37128 & n37129;
  assign n37131 = n37130 ^ n37079;
  assign n37133 = n37132 ^ n37131;
  assign n37138 = n37137 ^ n37133;
  assign n37144 = n37143 ^ n37138;
  assign n37075 = n37074 ^ n33350;
  assign n37088 = n37087 ^ n37075;
  assign n36890 = n36889 ^ n36877;
  assign n36891 = n36845 ^ n36811;
  assign n36892 = n36836 ^ n33693;
  assign n36893 = n36892 ^ n36816;
  assign n36899 = n36896 & ~n36898;
  assign n36900 = n36833 ^ n36819;
  assign n36901 = n36899 & ~n36900;
  assign n36902 = ~n36893 & ~n36901;
  assign n36903 = n36839 ^ n36815;
  assign n36904 = ~n36902 & ~n36903;
  assign n36905 = n36842 ^ n36813;
  assign n36906 = n36904 & n36905;
  assign n36907 = ~n36891 & n36906;
  assign n36908 = n36848 ^ n33582;
  assign n36909 = n36908 ^ n36808;
  assign n36910 = ~n36907 & ~n36909;
  assign n36911 = n36851 ^ n36807;
  assign n36912 = ~n36910 & n36911;
  assign n36913 = n36854 ^ n33567;
  assign n36914 = n36913 ^ n36803;
  assign n36915 = n36912 & ~n36914;
  assign n36916 = n36857 ^ n36802;
  assign n36917 = ~n36915 & n36916;
  assign n36918 = n36860 ^ n33545;
  assign n36919 = n36918 ^ n36799;
  assign n36920 = n36917 & n36919;
  assign n36921 = n36865 ^ n34090;
  assign n36922 = n36921 ^ n36863;
  assign n36923 = n36920 & n36922;
  assign n36924 = n36868 ^ n36798;
  assign n36925 = ~n36923 & n36924;
  assign n36926 = n36871 ^ n36795;
  assign n36927 = n36925 & ~n36926;
  assign n36928 = n36874 ^ n33368;
  assign n36929 = n36928 ^ n36792;
  assign n36930 = n36927 & n36929;
  assign n36931 = ~n36890 & n36930;
  assign n36935 = n36934 ^ n33356;
  assign n36947 = n36946 ^ n36935;
  assign n37089 = ~n36931 & ~n36947;
  assign n37127 = ~n37088 & n37089;
  assign n37145 = n37144 ^ n37127;
  assign n37124 = n34709 ^ n26798;
  assign n37125 = n37124 ^ n1976;
  assign n37126 = n37125 ^ n1867;
  assign n37146 = n37145 ^ n37126;
  assign n37090 = n37089 ^ n37088;
  assign n1834 = n1827 ^ n1794;
  assign n1853 = n1852 ^ n1834;
  assign n1860 = n1859 ^ n1853;
  assign n37091 = n37090 ^ n1860;
  assign n36950 = n34716 ^ n1742;
  assign n36951 = n36950 ^ n31065;
  assign n36952 = n36951 ^ n25427;
  assign n36949 = n36930 ^ n36890;
  assign n36953 = n36952 ^ n36949;
  assign n36954 = n36929 ^ n36927;
  assign n36958 = n36957 ^ n36954;
  assign n36959 = n36926 ^ n36925;
  assign n36963 = n36962 ^ n36959;
  assign n36964 = n36924 ^ n36923;
  assign n36965 = n36964 ^ n3131;
  assign n36966 = n36922 ^ n36920;
  assign n2754 = n2753 ^ n2702;
  assign n2761 = n2760 ^ n2754;
  assign n2762 = n2761 ^ n1583;
  assign n36967 = n36966 ^ n2762;
  assign n36968 = n36919 ^ n36917;
  assign n3103 = n3098 ^ n3093;
  assign n3104 = n3103 ^ n2680;
  assign n3105 = n3104 ^ n2758;
  assign n36969 = n36968 ^ n3105;
  assign n36970 = n36916 ^ n36915;
  assign n2647 = n2643 ^ n2616;
  assign n2666 = n2665 ^ n2647;
  assign n2673 = n2672 ^ n2666;
  assign n36971 = n36970 ^ n2673;
  assign n36972 = n36914 ^ n36912;
  assign n3180 = n3179 ^ n2572;
  assign n3190 = n3189 ^ n3180;
  assign n3191 = n3190 ^ n2660;
  assign n36973 = n36972 ^ n3191;
  assign n36975 = n34741 ^ n2560;
  assign n36976 = n36975 ^ n30996;
  assign n36977 = n36976 ^ n3187;
  assign n36974 = n36911 ^ n36910;
  assign n36978 = n36977 ^ n36974;
  assign n36980 = n34746 ^ n3165;
  assign n36981 = n36980 ^ n31006;
  assign n36982 = n36981 ^ n25444;
  assign n36979 = n36909 ^ n36907;
  assign n36983 = n36982 ^ n36979;
  assign n36987 = n36906 ^ n36891;
  assign n36984 = n26511 ^ n1438;
  assign n36985 = n36984 ^ n31001;
  assign n36986 = n36985 ^ n25449;
  assign n36988 = n36987 ^ n36986;
  assign n36990 = n36903 ^ n36902;
  assign n1356 = n1316 ^ n1253;
  assign n1357 = n1356 ^ n1353;
  assign n1361 = n1360 ^ n1357;
  assign n36991 = n36990 ^ n1361;
  assign n36993 = n36900 ^ n36899;
  assign n3343 = n3339 ^ n1136;
  assign n3344 = n3343 ^ n1336;
  assign n3348 = n3347 ^ n3344;
  assign n36994 = n36993 ^ n3348;
  assign n37011 = n37010 ^ n36995;
  assign n37012 = ~n37007 & n37011;
  assign n37013 = n37012 ^ n37010;
  assign n37014 = n37013 ^ n36993;
  assign n37015 = n36994 & ~n37014;
  assign n37016 = n37015 ^ n3348;
  assign n36992 = n36901 ^ n36893;
  assign n37017 = n37016 ^ n36992;
  assign n1329 = n1238 ^ n1167;
  assign n1339 = n1338 ^ n1329;
  assign n1346 = n1345 ^ n1339;
  assign n37018 = n36992 ^ n1346;
  assign n37019 = ~n37017 & n37018;
  assign n37020 = n37019 ^ n1346;
  assign n37021 = n37020 ^ n36990;
  assign n37022 = ~n36991 & n37021;
  assign n37023 = n37022 ^ n1361;
  assign n36989 = n36905 ^ n36904;
  assign n37024 = n37023 ^ n36989;
  assign n37025 = n26606 ^ n1420;
  assign n37026 = n37025 ^ n1371;
  assign n37027 = n37026 ^ n3017;
  assign n37028 = n37027 ^ n36989;
  assign n37029 = n37024 & ~n37028;
  assign n37030 = n37029 ^ n37027;
  assign n37031 = n37030 ^ n36987;
  assign n37032 = n36988 & ~n37031;
  assign n37033 = n37032 ^ n36986;
  assign n37034 = n37033 ^ n36982;
  assign n37035 = n36983 & ~n37034;
  assign n37036 = n37035 ^ n36979;
  assign n37037 = n37036 ^ n36974;
  assign n37038 = n36978 & ~n37037;
  assign n37039 = n37038 ^ n36977;
  assign n37040 = n37039 ^ n36972;
  assign n37041 = n36973 & ~n37040;
  assign n37042 = n37041 ^ n3191;
  assign n37043 = n37042 ^ n36970;
  assign n37044 = ~n36971 & n37043;
  assign n37045 = n37044 ^ n2673;
  assign n37046 = n37045 ^ n36968;
  assign n37047 = n36969 & ~n37046;
  assign n37048 = n37047 ^ n3105;
  assign n37049 = n37048 ^ n36966;
  assign n37050 = n36967 & ~n37049;
  assign n37051 = n37050 ^ n2762;
  assign n37052 = n37051 ^ n36964;
  assign n37053 = n36965 & ~n37052;
  assign n37054 = n37053 ^ n3131;
  assign n37055 = n37054 ^ n36959;
  assign n37056 = n36963 & ~n37055;
  assign n37057 = n37056 ^ n36962;
  assign n37058 = n37057 ^ n36954;
  assign n37059 = ~n36958 & n37058;
  assign n37060 = n37059 ^ n36957;
  assign n37061 = n37060 ^ n36949;
  assign n37062 = n36953 & ~n37061;
  assign n37063 = n37062 ^ n36952;
  assign n36948 = n36947 ^ n36931;
  assign n37064 = n37063 ^ n36948;
  assign n37065 = n34839 ^ n1715;
  assign n37066 = n37065 ^ n1849;
  assign n37067 = n37066 ^ n31061;
  assign n37068 = n37067 ^ n36948;
  assign n37069 = ~n37064 & n37068;
  assign n37070 = n37069 ^ n37067;
  assign n37121 = n37090 ^ n37070;
  assign n37122 = ~n37091 & n37121;
  assign n37123 = n37122 ^ n1860;
  assign n37188 = n37145 ^ n37123;
  assign n37189 = ~n37146 & n37188;
  assign n37190 = n37189 ^ n37126;
  assign n1959 = n1958 ^ n1904;
  assign n1972 = n1971 ^ n1959;
  assign n1979 = n1978 ^ n1972;
  assign n37191 = n37190 ^ n1979;
  assign n37181 = n37138 ^ n32511;
  assign n37182 = n37142 ^ n37138;
  assign n37183 = ~n37181 & n37182;
  assign n37184 = n37183 ^ n32511;
  assign n37185 = n37184 ^ n32504;
  assign n37179 = n36385 ^ n36299;
  assign n37175 = n37137 ^ n37132;
  assign n37176 = n37133 & ~n37175;
  assign n37177 = n37176 ^ n37137;
  assign n37171 = n35047 ^ n34228;
  assign n37172 = n35654 ^ n35047;
  assign n37173 = ~n37171 & n37172;
  assign n37174 = n37173 ^ n34228;
  assign n37178 = n37177 ^ n37174;
  assign n37180 = n37179 ^ n37178;
  assign n37186 = n37185 ^ n37180;
  assign n37170 = n37127 & ~n37144;
  assign n37187 = n37186 ^ n37170;
  assign n37192 = n37191 ^ n37187;
  assign n37197 = n37196 ^ n37192;
  assign n37147 = n37146 ^ n37123;
  assign n37116 = n35800 ^ n34894;
  assign n37117 = n36464 ^ n35800;
  assign n37118 = ~n37116 & ~n37117;
  assign n37119 = n37118 ^ n34894;
  assign n37166 = n37147 ^ n37119;
  assign n37093 = n35770 ^ n35137;
  assign n37094 = n35934 ^ n35770;
  assign n37095 = n37093 & n37094;
  assign n37096 = n37095 ^ n35137;
  assign n37092 = n37091 ^ n37070;
  assign n37097 = n37096 ^ n37092;
  assign n37104 = n35716 ^ n35035;
  assign n37105 = n35940 ^ n35716;
  assign n37106 = n37104 & ~n37105;
  assign n37107 = n37106 ^ n35035;
  assign n37098 = n35041 ^ n34889;
  assign n37099 = n35946 ^ n34889;
  assign n37100 = ~n37098 & n37099;
  assign n37101 = n37100 ^ n35041;
  assign n37102 = n37060 ^ n36953;
  assign n37103 = ~n37101 & n37102;
  assign n37108 = n37107 ^ n37103;
  assign n37109 = n37067 ^ n37064;
  assign n37110 = n37109 ^ n37107;
  assign n37111 = n37108 & ~n37110;
  assign n37112 = n37111 ^ n37103;
  assign n37113 = n37112 ^ n37092;
  assign n37114 = ~n37097 & n37113;
  assign n37115 = n37114 ^ n37096;
  assign n37167 = n37147 ^ n37115;
  assign n37168 = n37166 & n37167;
  assign n37169 = n37168 ^ n37119;
  assign n37198 = n37197 ^ n37169;
  assign n37120 = n37119 ^ n37115;
  assign n37148 = n37147 ^ n37120;
  assign n37149 = n37148 ^ n34436;
  assign n37150 = n37112 ^ n37097;
  assign n37151 = n37150 ^ n34442;
  assign n37152 = n37102 ^ n37101;
  assign n37153 = n34292 & ~n37152;
  assign n37154 = n37153 ^ n34448;
  assign n37155 = n37109 ^ n37108;
  assign n37156 = n37155 ^ n37153;
  assign n37157 = n37154 & ~n37156;
  assign n37158 = n37157 ^ n34448;
  assign n37159 = n37158 ^ n37150;
  assign n37160 = n37151 & n37159;
  assign n37161 = n37160 ^ n34442;
  assign n37162 = n37161 ^ n37148;
  assign n37163 = n37149 & n37162;
  assign n37164 = n37163 ^ n34436;
  assign n37165 = n37164 ^ n34434;
  assign n37199 = n37198 ^ n37165;
  assign n37200 = n37161 ^ n37149;
  assign n37201 = n37158 ^ n34442;
  assign n37202 = n37201 ^ n37150;
  assign n37203 = n37200 & ~n37202;
  assign n37237 = n37199 & n37203;
  assign n37250 = n36575 ^ n36574;
  assign n37245 = n35917 ^ n34306;
  assign n37246 = n36623 ^ n35917;
  assign n37247 = ~n37245 & ~n37246;
  assign n37248 = n37247 ^ n34306;
  assign n37242 = n37192 ^ n37169;
  assign n37243 = n37197 & ~n37242;
  assign n37244 = n37243 ^ n37196;
  assign n37249 = n37248 ^ n37244;
  assign n37251 = n37250 ^ n37249;
  assign n37252 = n37251 ^ n34428;
  assign n37238 = n37198 ^ n34434;
  assign n37239 = n37198 ^ n37164;
  assign n37240 = ~n37238 & n37239;
  assign n37241 = n37240 ^ n34434;
  assign n37253 = n37252 ^ n37241;
  assign n37671 = ~n37237 & n37253;
  assign n37574 = n37251 ^ n37241;
  assign n37575 = n37252 & n37574;
  assign n37576 = n37575 ^ n34428;
  assign n37669 = n37576 ^ n34422;
  assign n37420 = n37250 ^ n37248;
  assign n37421 = n37250 ^ n37244;
  assign n37422 = n37420 & ~n37421;
  assign n37423 = n37422 ^ n37248;
  assign n37415 = n36040 ^ n35008;
  assign n37416 = n36730 ^ n36040;
  assign n37417 = ~n37415 & ~n37416;
  assign n37418 = n37417 ^ n35008;
  assign n37571 = n37423 ^ n37418;
  assign n37414 = n36578 ^ n36577;
  assign n37572 = n37571 ^ n37414;
  assign n37670 = n37669 ^ n37572;
  assign n37819 = n37671 ^ n37670;
  assign n37816 = n35553 ^ n27174;
  assign n37817 = n37816 ^ n31398;
  assign n37818 = n37817 ^ n25791;
  assign n37820 = n37819 ^ n37818;
  assign n37254 = n37253 ^ n37237;
  assign n37234 = n35558 ^ n27167;
  assign n37235 = n37234 ^ n31404;
  assign n37236 = n37235 ^ n702;
  assign n37255 = n37254 ^ n37236;
  assign n37205 = n35564 ^ n27158;
  assign n37206 = n37205 ^ n31409;
  assign n37207 = n37206 ^ n25763;
  assign n37204 = n37203 ^ n37199;
  assign n37208 = n37207 ^ n37204;
  assign n37210 = n27142 ^ n2333;
  assign n37211 = n37210 ^ n31421;
  assign n37212 = n37211 ^ n25768;
  assign n37209 = n37202 ^ n37200;
  assign n37213 = n37212 ^ n37209;
  assign n37214 = n34883 ^ n27147;
  assign n37215 = n37214 ^ n2254;
  assign n37216 = n37215 ^ n25773;
  assign n37217 = n37216 ^ n37202;
  assign n2102 = n2065 ^ n2023;
  assign n2109 = n2108 ^ n2102;
  assign n2110 = n2109 ^ n2099;
  assign n37218 = n37152 ^ n34292;
  assign n37219 = n2110 & ~n37218;
  assign n2233 = n2222 ^ n2151;
  assign n2243 = n2242 ^ n2233;
  assign n2247 = n2246 ^ n2243;
  assign n37220 = n37219 ^ n2247;
  assign n37221 = n37155 ^ n37154;
  assign n37222 = n37221 ^ n2247;
  assign n37223 = n37220 & ~n37222;
  assign n37224 = n37223 ^ n37219;
  assign n37225 = n37224 ^ n37202;
  assign n37226 = ~n37217 & n37225;
  assign n37227 = n37226 ^ n37216;
  assign n37228 = n37227 ^ n37212;
  assign n37229 = n37213 & ~n37228;
  assign n37230 = n37229 ^ n37209;
  assign n37231 = n37230 ^ n37204;
  assign n37232 = ~n37208 & n37231;
  assign n37233 = n37232 ^ n37207;
  assign n37821 = n37254 ^ n37233;
  assign n37822 = ~n37255 & n37821;
  assign n37823 = n37822 ^ n37236;
  assign n37824 = n37823 ^ n37819;
  assign n37825 = ~n37820 & n37824;
  assign n37826 = n37825 ^ n37818;
  assign n37812 = n35549 ^ n27181;
  assign n37813 = n37812 ^ n31394;
  assign n37814 = n37813 ^ n25798;
  assign n37672 = ~n37670 & ~n37671;
  assign n37573 = n37572 ^ n34422;
  assign n37577 = n37576 ^ n37572;
  assign n37578 = ~n37573 & n37577;
  assign n37579 = n37578 ^ n34422;
  assign n37667 = n37579 ^ n33541;
  assign n37419 = n37418 ^ n37414;
  assign n37424 = n37423 ^ n37414;
  assign n37425 = ~n37419 & n37424;
  assign n37426 = n37425 ^ n37418;
  assign n37408 = n36034 ^ n35002;
  assign n37409 = n36724 ^ n36034;
  assign n37410 = n37408 & n37409;
  assign n37411 = n37410 ^ n35002;
  assign n37568 = n37426 ^ n37411;
  assign n37412 = n36581 ^ n36568;
  assign n37569 = n37568 ^ n37412;
  assign n37668 = n37667 ^ n37569;
  assign n37811 = n37672 ^ n37668;
  assign n37815 = n37814 ^ n37811;
  assign n38047 = n37826 ^ n37815;
  assign n38052 = n38051 ^ n38047;
  assign n37981 = n37823 ^ n37820;
  assign n37977 = n36686 ^ n36019;
  assign n37364 = n37003 ^ n37000;
  assign n37978 = n37364 ^ n36686;
  assign n37979 = ~n37977 & ~n37978;
  assign n37980 = n37979 ^ n36019;
  assign n37982 = n37981 ^ n37980;
  assign n37256 = n37255 ^ n37233;
  assign n35929 = n35928 ^ n35927;
  assign n36636 = n36635 ^ n36613;
  assign n36637 = n36636 ^ n35927;
  assign n36638 = n35929 & n36637;
  assign n36639 = n36638 ^ n35928;
  assign n37257 = n37256 ^ n36639;
  assign n37263 = n37230 ^ n37208;
  assign n37258 = n36702 ^ n36031;
  assign n37259 = n36610 ^ n36542;
  assign n37260 = n37259 ^ n36702;
  assign n37261 = n37258 & n37260;
  assign n37262 = n37261 ^ n36031;
  assign n37264 = n37263 ^ n37262;
  assign n37270 = n37227 ^ n37213;
  assign n37265 = n36708 ^ n36055;
  assign n37266 = n36607 ^ n36604;
  assign n37267 = n37266 ^ n36708;
  assign n37268 = n37265 & ~n37267;
  assign n37269 = n37268 ^ n36055;
  assign n37271 = n37270 ^ n37269;
  assign n37277 = n37224 ^ n37217;
  assign n37272 = n36715 ^ n36034;
  assign n37273 = n36600 ^ n36548;
  assign n37274 = n37273 ^ n36715;
  assign n37275 = ~n37272 & n37274;
  assign n37276 = n37275 ^ n36034;
  assign n37278 = n37277 ^ n37276;
  assign n37284 = n37221 ^ n37220;
  assign n37279 = n36717 ^ n36040;
  assign n37280 = n36597 ^ n36553;
  assign n37281 = n37280 ^ n36717;
  assign n37282 = n37279 & ~n37281;
  assign n37283 = n37282 ^ n36040;
  assign n37285 = n37284 ^ n37283;
  assign n37291 = n37218 ^ n2110;
  assign n37286 = n36724 ^ n35917;
  assign n37287 = n36594 ^ n36558;
  assign n37288 = n37287 ^ n36724;
  assign n37289 = ~n37286 & ~n37288;
  assign n37290 = n37289 ^ n35917;
  assign n37292 = n37291 ^ n37290;
  assign n37918 = n36730 ^ n35816;
  assign n37400 = n36591 ^ n36563;
  assign n37919 = n37400 ^ n36730;
  assign n37920 = ~n37918 & ~n37919;
  assign n37921 = n37920 ^ n35816;
  assign n37304 = n37045 ^ n36969;
  assign n37300 = n35667 ^ n34847;
  assign n37301 = n36435 ^ n35667;
  assign n37302 = ~n37300 & ~n37301;
  assign n37303 = n37302 ^ n34847;
  assign n37305 = n37304 ^ n37303;
  assign n37310 = n37042 ^ n36971;
  assign n37306 = n35673 ^ n34864;
  assign n37307 = n37179 ^ n35673;
  assign n37308 = ~n37306 & n37307;
  assign n37309 = n37308 ^ n34864;
  assign n37311 = n37310 ^ n37309;
  assign n37316 = n37039 ^ n36973;
  assign n37312 = n35680 ^ n34857;
  assign n37313 = n37132 ^ n35680;
  assign n37314 = n37312 & ~n37313;
  assign n37315 = n37314 ^ n34857;
  assign n37317 = n37316 ^ n37315;
  assign n37322 = n37036 ^ n36978;
  assign n37318 = n36265 ^ n35430;
  assign n37319 = n37086 ^ n36265;
  assign n37320 = ~n37318 & ~n37319;
  assign n37321 = n37320 ^ n35430;
  assign n37323 = n37322 ^ n37321;
  assign n37328 = n37033 ^ n36983;
  assign n37324 = n35948 ^ n34900;
  assign n37325 = n36945 ^ n35948;
  assign n37326 = ~n37324 & ~n37325;
  assign n37327 = n37326 ^ n34900;
  assign n37329 = n37328 ^ n37327;
  assign n37472 = n37030 ^ n36988;
  assign n37334 = n37027 ^ n37024;
  assign n37330 = n35960 ^ n34912;
  assign n37331 = n36790 ^ n35960;
  assign n37332 = n37330 & ~n37331;
  assign n37333 = n37332 ^ n34912;
  assign n37335 = n37334 ^ n37333;
  assign n37340 = n37020 ^ n36991;
  assign n37336 = n35966 ^ n34919;
  assign n37337 = n36645 ^ n35966;
  assign n37338 = ~n37336 & ~n37337;
  assign n37339 = n37338 ^ n34919;
  assign n37341 = n37340 ^ n37339;
  assign n37343 = n35972 ^ n34926;
  assign n37344 = n36648 ^ n35972;
  assign n37345 = n37343 & n37344;
  assign n37346 = n37345 ^ n34926;
  assign n37342 = n37017 ^ n1346;
  assign n37347 = n37346 ^ n37342;
  assign n37352 = n37013 ^ n36994;
  assign n37348 = n35979 ^ n34934;
  assign n37349 = n36654 ^ n35979;
  assign n37350 = n37348 & n37349;
  assign n37351 = n37350 ^ n34934;
  assign n37353 = n37352 ^ n37351;
  assign n37354 = n35982 ^ n34941;
  assign n37355 = n36664 ^ n35982;
  assign n37356 = ~n37354 & n37355;
  assign n37357 = n37356 ^ n34941;
  assign n37359 = n37358 ^ n37357;
  assign n37360 = n35992 ^ n34947;
  assign n37361 = n36670 ^ n35992;
  assign n37362 = n37360 & ~n37361;
  assign n37363 = n37362 ^ n34947;
  assign n37365 = n37364 ^ n37363;
  assign n37366 = n35998 ^ n34953;
  assign n37367 = n36673 ^ n35998;
  assign n37368 = n37366 & ~n37367;
  assign n37369 = n37368 ^ n34953;
  assign n37370 = n37369 ^ n36636;
  assign n37371 = n36000 ^ n34959;
  assign n37372 = n36679 ^ n36000;
  assign n37373 = n37371 & ~n37372;
  assign n37374 = n37373 ^ n34959;
  assign n37375 = n37374 ^ n37259;
  assign n37376 = n36002 ^ n34966;
  assign n37377 = n36686 ^ n36002;
  assign n37378 = ~n37376 & ~n37377;
  assign n37379 = n37378 ^ n34966;
  assign n37380 = n37379 ^ n37266;
  assign n37381 = n36008 ^ n34972;
  assign n37382 = n36008 ^ n35927;
  assign n37383 = n37381 & n37382;
  assign n37384 = n37383 ^ n34972;
  assign n37385 = n37384 ^ n37273;
  assign n37386 = n36019 ^ n34975;
  assign n37387 = n36702 ^ n36019;
  assign n37388 = ~n37386 & n37387;
  assign n37389 = n37388 ^ n34975;
  assign n37390 = n37389 ^ n37280;
  assign n37391 = n35928 ^ n34982;
  assign n37392 = n36708 ^ n35928;
  assign n37393 = n37391 & n37392;
  assign n37394 = n37393 ^ n34982;
  assign n37395 = n37394 ^ n37287;
  assign n37396 = n36031 ^ n34989;
  assign n37397 = n36715 ^ n36031;
  assign n37398 = ~n37396 & ~n37397;
  assign n37399 = n37398 ^ n34989;
  assign n37401 = n37400 ^ n37399;
  assign n37406 = n36588 ^ n36585;
  assign n37402 = n36055 ^ n34995;
  assign n37403 = n36717 ^ n36055;
  assign n37404 = n37402 & ~n37403;
  assign n37405 = n37404 ^ n34995;
  assign n37407 = n37406 ^ n37405;
  assign n37413 = n37412 ^ n37411;
  assign n37427 = n37426 ^ n37412;
  assign n37428 = ~n37413 & ~n37427;
  assign n37429 = n37428 ^ n37411;
  assign n37430 = n37429 ^ n37406;
  assign n37431 = n37407 & ~n37430;
  assign n37432 = n37431 ^ n37405;
  assign n37433 = n37432 ^ n37400;
  assign n37434 = n37401 & ~n37433;
  assign n37435 = n37434 ^ n37399;
  assign n37436 = n37435 ^ n37287;
  assign n37437 = n37395 & n37436;
  assign n37438 = n37437 ^ n37394;
  assign n37439 = n37438 ^ n37280;
  assign n37440 = ~n37390 & n37439;
  assign n37441 = n37440 ^ n37389;
  assign n37442 = n37441 ^ n37273;
  assign n37443 = n37385 & n37442;
  assign n37444 = n37443 ^ n37384;
  assign n37445 = n37444 ^ n37266;
  assign n37446 = n37380 & ~n37445;
  assign n37447 = n37446 ^ n37379;
  assign n37448 = n37447 ^ n37259;
  assign n37449 = ~n37375 & ~n37448;
  assign n37450 = n37449 ^ n37374;
  assign n37451 = n37450 ^ n36636;
  assign n37452 = ~n37370 & n37451;
  assign n37453 = n37452 ^ n37369;
  assign n37454 = n37453 ^ n37364;
  assign n37455 = ~n37365 & ~n37454;
  assign n37456 = n37455 ^ n37363;
  assign n37457 = n37456 ^ n37358;
  assign n37458 = n37359 & ~n37457;
  assign n37459 = n37458 ^ n37357;
  assign n37460 = n37459 ^ n37352;
  assign n37461 = ~n37353 & ~n37460;
  assign n37462 = n37461 ^ n37351;
  assign n37463 = n37462 ^ n37342;
  assign n37464 = n37347 & n37463;
  assign n37465 = n37464 ^ n37346;
  assign n37466 = n37465 ^ n37340;
  assign n37467 = ~n37341 & n37466;
  assign n37468 = n37467 ^ n37339;
  assign n37469 = n37468 ^ n37334;
  assign n37470 = n37335 & n37469;
  assign n37471 = n37470 ^ n37333;
  assign n37473 = n37472 ^ n37471;
  assign n37474 = n35950 ^ n34902;
  assign n37475 = n36887 ^ n35950;
  assign n37476 = ~n37474 & ~n37475;
  assign n37477 = n37476 ^ n34902;
  assign n37478 = n37477 ^ n37472;
  assign n37479 = n37473 & ~n37478;
  assign n37480 = n37479 ^ n37477;
  assign n37481 = n37480 ^ n37328;
  assign n37482 = n37329 & n37481;
  assign n37483 = n37482 ^ n37327;
  assign n37484 = n37483 ^ n37322;
  assign n37485 = ~n37323 & ~n37484;
  assign n37486 = n37485 ^ n37321;
  assign n37487 = n37486 ^ n37316;
  assign n37488 = ~n37317 & n37487;
  assign n37489 = n37488 ^ n37315;
  assign n37490 = n37489 ^ n37310;
  assign n37491 = n37311 & ~n37490;
  assign n37492 = n37491 ^ n37309;
  assign n37493 = n37492 ^ n37304;
  assign n37494 = n37305 & n37493;
  assign n37495 = n37494 ^ n37303;
  assign n37294 = n35660 ^ n35109;
  assign n37295 = n36428 ^ n35660;
  assign n37296 = n37294 & n37295;
  assign n37297 = n37296 ^ n35109;
  assign n37516 = n37495 ^ n37297;
  assign n37298 = n37048 ^ n36967;
  assign n37517 = n37516 ^ n37298;
  assign n37518 = n37517 ^ n34108;
  assign n37519 = n37492 ^ n37303;
  assign n37520 = n37519 ^ n37304;
  assign n37521 = n37520 ^ n34114;
  assign n37522 = n37489 ^ n37309;
  assign n37523 = n37522 ^ n37310;
  assign n37524 = n37523 ^ n34120;
  assign n37525 = n37486 ^ n37315;
  assign n37526 = n37525 ^ n37316;
  assign n37527 = n37526 ^ n34130;
  assign n37528 = n37483 ^ n37321;
  assign n37529 = n37528 ^ n37322;
  assign n37530 = n37529 ^ n34922;
  assign n37531 = n37480 ^ n37327;
  assign n37532 = n37531 ^ n37328;
  assign n37533 = n37532 ^ n34929;
  assign n37534 = n37477 ^ n37473;
  assign n37535 = n37534 ^ n34311;
  assign n37536 = n37468 ^ n37333;
  assign n37537 = n37536 ^ n37334;
  assign n37538 = n37537 ^ n34323;
  assign n37539 = n37465 ^ n37341;
  assign n37540 = n37539 ^ n34333;
  assign n37541 = n37462 ^ n37347;
  assign n37542 = n37541 ^ n34342;
  assign n37543 = n37459 ^ n37353;
  assign n37544 = n37543 ^ n34348;
  assign n37545 = n37456 ^ n37359;
  assign n37546 = n37545 ^ n34359;
  assign n37547 = n37453 ^ n37365;
  assign n37548 = n37547 ^ n34509;
  assign n37549 = n37450 ^ n37370;
  assign n37550 = n37549 ^ n34368;
  assign n37552 = n37444 ^ n37380;
  assign n37553 = n37552 ^ n34380;
  assign n37554 = n37441 ^ n37384;
  assign n37555 = n37554 ^ n37273;
  assign n37556 = n37555 ^ n34386;
  assign n37557 = n37438 ^ n37390;
  assign n37558 = n37557 ^ n34388;
  assign n37559 = n37435 ^ n37394;
  assign n37560 = n37559 ^ n37287;
  assign n37561 = n37560 ^ n34395;
  assign n37562 = n37432 ^ n37399;
  assign n37563 = n37562 ^ n37400;
  assign n37564 = n37563 ^ n34405;
  assign n37565 = n37429 ^ n37405;
  assign n37566 = n37565 ^ n37406;
  assign n37567 = n37566 ^ n34411;
  assign n37570 = n37569 ^ n33541;
  assign n37580 = n37579 ^ n37569;
  assign n37581 = n37570 & n37580;
  assign n37582 = n37581 ^ n33541;
  assign n37583 = n37582 ^ n37566;
  assign n37584 = ~n37567 & ~n37583;
  assign n37585 = n37584 ^ n34411;
  assign n37586 = n37585 ^ n37563;
  assign n37587 = n37564 & n37586;
  assign n37588 = n37587 ^ n34405;
  assign n37589 = n37588 ^ n37560;
  assign n37590 = ~n37561 & ~n37589;
  assign n37591 = n37590 ^ n34395;
  assign n37592 = n37591 ^ n37557;
  assign n37593 = ~n37558 & n37592;
  assign n37594 = n37593 ^ n34388;
  assign n37595 = n37594 ^ n37555;
  assign n37596 = n37556 & ~n37595;
  assign n37597 = n37596 ^ n34386;
  assign n37598 = n37597 ^ n37552;
  assign n37599 = ~n37553 & n37598;
  assign n37600 = n37599 ^ n34380;
  assign n37551 = n37447 ^ n37375;
  assign n37601 = n37600 ^ n37551;
  assign n37602 = n37551 ^ n34374;
  assign n37603 = ~n37601 & ~n37602;
  assign n37604 = n37603 ^ n34374;
  assign n37605 = n37604 ^ n37549;
  assign n37606 = n37550 & ~n37605;
  assign n37607 = n37606 ^ n34368;
  assign n37608 = n37607 ^ n37547;
  assign n37609 = n37548 & ~n37608;
  assign n37610 = n37609 ^ n34509;
  assign n37611 = n37610 ^ n37545;
  assign n37612 = n37546 & ~n37611;
  assign n37613 = n37612 ^ n34359;
  assign n37614 = n37613 ^ n37543;
  assign n37615 = ~n37544 & n37614;
  assign n37616 = n37615 ^ n34348;
  assign n37617 = n37616 ^ n37541;
  assign n37618 = ~n37542 & n37617;
  assign n37619 = n37618 ^ n34342;
  assign n37620 = n37619 ^ n37539;
  assign n37621 = n37540 & n37620;
  assign n37622 = n37621 ^ n34333;
  assign n37623 = n37622 ^ n37537;
  assign n37624 = n37538 & n37623;
  assign n37625 = n37624 ^ n34323;
  assign n37626 = n37625 ^ n37534;
  assign n37627 = n37535 & ~n37626;
  assign n37628 = n37627 ^ n34311;
  assign n37629 = n37628 ^ n37532;
  assign n37630 = ~n37533 & n37629;
  assign n37631 = n37630 ^ n34929;
  assign n37632 = n37631 ^ n37529;
  assign n37633 = ~n37530 & n37632;
  assign n37634 = n37633 ^ n34922;
  assign n37635 = n37634 ^ n37526;
  assign n37636 = ~n37527 & ~n37635;
  assign n37637 = n37636 ^ n34130;
  assign n37638 = n37637 ^ n37523;
  assign n37639 = ~n37524 & ~n37638;
  assign n37640 = n37639 ^ n34120;
  assign n37641 = n37640 ^ n37520;
  assign n37642 = n37521 & n37641;
  assign n37643 = n37642 ^ n34114;
  assign n37644 = n37643 ^ n37517;
  assign n37645 = n37518 & ~n37644;
  assign n37646 = n37645 ^ n34108;
  assign n37652 = n37646 ^ n34167;
  assign n37501 = n35654 ^ n35103;
  assign n37502 = n36418 ^ n35654;
  assign n37503 = ~n37501 & ~n37502;
  assign n37504 = n37503 ^ n35103;
  assign n37499 = n37051 ^ n36965;
  assign n37299 = n37298 ^ n37297;
  assign n37496 = n37495 ^ n37298;
  assign n37497 = ~n37299 & ~n37496;
  assign n37498 = n37497 ^ n37297;
  assign n37500 = n37499 ^ n37498;
  assign n37514 = n37504 ^ n37500;
  assign n37653 = n37652 ^ n37514;
  assign n37654 = n37640 ^ n34114;
  assign n37655 = n37654 ^ n37520;
  assign n37656 = n37637 ^ n34120;
  assign n37657 = n37656 ^ n37523;
  assign n37658 = n37634 ^ n34130;
  assign n37659 = n37658 ^ n37526;
  assign n37660 = n37625 ^ n34311;
  assign n37661 = n37660 ^ n37534;
  assign n37662 = n37622 ^ n37538;
  assign n37663 = n37616 ^ n37542;
  assign n37664 = n37610 ^ n37546;
  assign n37665 = n37582 ^ n34411;
  assign n37666 = n37665 ^ n37566;
  assign n37673 = n37668 & n37672;
  assign n37674 = ~n37666 & ~n37673;
  assign n37675 = n37585 ^ n34405;
  assign n37676 = n37675 ^ n37563;
  assign n37677 = n37674 & ~n37676;
  assign n37678 = n37588 ^ n34395;
  assign n37679 = n37678 ^ n37560;
  assign n37680 = ~n37677 & n37679;
  assign n37681 = n37591 ^ n37558;
  assign n37682 = n37680 & ~n37681;
  assign n37683 = n37594 ^ n37556;
  assign n37684 = n37682 & n37683;
  assign n37685 = n37597 ^ n37553;
  assign n37686 = n37684 & ~n37685;
  assign n37687 = n37601 ^ n34374;
  assign n37688 = ~n37686 & n37687;
  assign n37689 = n37604 ^ n37550;
  assign n37690 = ~n37688 & ~n37689;
  assign n37691 = n37607 ^ n37548;
  assign n37692 = n37690 & ~n37691;
  assign n37693 = ~n37664 & n37692;
  assign n37694 = n37613 ^ n37544;
  assign n37695 = ~n37693 & ~n37694;
  assign n37696 = n37663 & ~n37695;
  assign n37697 = n37619 ^ n37540;
  assign n37698 = n37696 & ~n37697;
  assign n37699 = ~n37662 & ~n37698;
  assign n37700 = n37661 & n37699;
  assign n37701 = n37628 ^ n34929;
  assign n37702 = n37701 ^ n37532;
  assign n37703 = n37700 & ~n37702;
  assign n37704 = n37631 ^ n37530;
  assign n37705 = ~n37703 & n37704;
  assign n37706 = n37659 & n37705;
  assign n37707 = ~n37657 & n37706;
  assign n37708 = ~n37655 & n37707;
  assign n37709 = n37643 ^ n34108;
  assign n37710 = n37709 ^ n37517;
  assign n37711 = ~n37708 & ~n37710;
  assign n37712 = n37653 & n37711;
  assign n37515 = n37514 ^ n34167;
  assign n37647 = n37646 ^ n37514;
  assign n37648 = ~n37515 & ~n37647;
  assign n37649 = n37648 ^ n34167;
  assign n37650 = n37649 ^ n34200;
  assign n37509 = n35049 ^ n34898;
  assign n37510 = n36415 ^ n34898;
  assign n37511 = ~n37509 & n37510;
  assign n37512 = n37511 ^ n35049;
  assign n37505 = n37504 ^ n37499;
  assign n37506 = n37500 & n37505;
  assign n37507 = n37506 ^ n37504;
  assign n37293 = n37054 ^ n36963;
  assign n37508 = n37507 ^ n37293;
  assign n37513 = n37512 ^ n37508;
  assign n37651 = n37650 ^ n37513;
  assign n37731 = n37712 ^ n37651;
  assign n37735 = n37734 ^ n37731;
  assign n37736 = n37711 ^ n37653;
  assign n37740 = n37739 ^ n37736;
  assign n37742 = n35462 ^ n27433;
  assign n37743 = n37742 ^ n26116;
  assign n37744 = n37743 ^ n31783;
  assign n37741 = n37710 ^ n37708;
  assign n37745 = n37744 ^ n37741;
  assign n37746 = n37707 ^ n37655;
  assign n37750 = n37749 ^ n37746;
  assign n37751 = n37706 ^ n37657;
  assign n37755 = n37754 ^ n37751;
  assign n37757 = n37704 ^ n37703;
  assign n2864 = n2803 ^ n1592;
  assign n2865 = n2864 ^ n2861;
  assign n2869 = n2868 ^ n2865;
  assign n37758 = n37757 ^ n2869;
  assign n37759 = n37702 ^ n37700;
  assign n2831 = n2824 ^ n2788;
  assign n2847 = n2846 ^ n2831;
  assign n2854 = n2853 ^ n2847;
  assign n37760 = n37759 ^ n2854;
  assign n37761 = n37699 ^ n37661;
  assign n3217 = n3213 ^ n2729;
  assign n3224 = n3223 ^ n3217;
  assign n3225 = n3224 ^ n2843;
  assign n37762 = n37761 ^ n3225;
  assign n37763 = n37698 ^ n37662;
  assign n37767 = n37766 ^ n37763;
  assign n37771 = n37697 ^ n37696;
  assign n37768 = n35489 ^ n3199;
  assign n37769 = n37768 ^ n31350;
  assign n37770 = n37769 ^ n3065;
  assign n37772 = n37771 ^ n37770;
  assign n37776 = n37695 ^ n37663;
  assign n37773 = n35494 ^ n27111;
  assign n37774 = n37773 ^ n3047;
  assign n37775 = n37774 ^ n2504;
  assign n37777 = n37776 ^ n37775;
  assign n37781 = n37694 ^ n37693;
  assign n37778 = n35499 ^ n27116;
  assign n37779 = n37778 ^ n2453;
  assign n37780 = n37779 ^ n3045;
  assign n37782 = n37781 ^ n37780;
  assign n37786 = n37692 ^ n37664;
  assign n37783 = n35504 ^ n3023;
  assign n37784 = n37783 ^ n2448;
  assign n37785 = n37784 ^ n31358;
  assign n37787 = n37786 ^ n37785;
  assign n37791 = n37691 ^ n37690;
  assign n37788 = n35509 ^ n1474;
  assign n37789 = n37788 ^ n31364;
  assign n37790 = n37789 ^ n1388;
  assign n37792 = n37791 ^ n37790;
  assign n37794 = n35515 ^ n1459;
  assign n37795 = n37794 ^ n1193;
  assign n37796 = n37795 ^ n25835;
  assign n37793 = n37689 ^ n37688;
  assign n37797 = n37796 ^ n37793;
  assign n37799 = n37685 ^ n37684;
  assign n1014 = n1013 ^ n950;
  assign n1027 = n1026 ^ n1014;
  assign n1034 = n1033 ^ n1027;
  assign n37800 = n37799 ^ n1034;
  assign n37802 = n37681 ^ n37680;
  assign n880 = n873 ^ n840;
  assign n899 = n898 ^ n880;
  assign n906 = n905 ^ n899;
  assign n37803 = n37802 ^ n906;
  assign n37806 = n31384 ^ n774;
  assign n37807 = n37806 ^ n35539;
  assign n37808 = n37807 ^ n3303;
  assign n37805 = n37676 ^ n37674;
  assign n37809 = n37808 ^ n37805;
  assign n37827 = n37826 ^ n37811;
  assign n37828 = ~n37815 & n37827;
  assign n37829 = n37828 ^ n37814;
  assign n37810 = n37673 ^ n37666;
  assign n37830 = n37829 ^ n37810;
  assign n37834 = n37833 ^ n37810;
  assign n37835 = ~n37830 & n37834;
  assign n37836 = n37835 ^ n37833;
  assign n37837 = n37836 ^ n37805;
  assign n37838 = ~n37809 & n37837;
  assign n37839 = n37838 ^ n37808;
  assign n37804 = n37679 ^ n37677;
  assign n37840 = n37839 ^ n37804;
  assign n37844 = n37843 ^ n37804;
  assign n37845 = ~n37840 & n37844;
  assign n37846 = n37845 ^ n37843;
  assign n37847 = n37846 ^ n37802;
  assign n37848 = n37803 & ~n37847;
  assign n37849 = n37848 ^ n906;
  assign n37801 = n37683 ^ n37682;
  assign n37850 = n37849 ^ n37801;
  assign n37851 = n35527 ^ n27130;
  assign n37852 = n37851 ^ n913;
  assign n37853 = n37852 ^ n1021;
  assign n37854 = n37853 ^ n37801;
  assign n37855 = n37850 & ~n37854;
  assign n37856 = n37855 ^ n37853;
  assign n37857 = n37856 ^ n37799;
  assign n37858 = n37800 & ~n37857;
  assign n37859 = n37858 ^ n1034;
  assign n37798 = n37687 ^ n37686;
  assign n37860 = n37859 ^ n37798;
  assign n37861 = n35520 ^ n1450;
  assign n37862 = n37861 ^ n31371;
  assign n37863 = n37862 ^ n1188;
  assign n37864 = n37863 ^ n37798;
  assign n37865 = n37860 & ~n37864;
  assign n37866 = n37865 ^ n37863;
  assign n37867 = n37866 ^ n37793;
  assign n37868 = ~n37797 & n37867;
  assign n37869 = n37868 ^ n37796;
  assign n37870 = n37869 ^ n37791;
  assign n37871 = n37792 & ~n37870;
  assign n37872 = n37871 ^ n37790;
  assign n37873 = n37872 ^ n37786;
  assign n37874 = n37787 & ~n37873;
  assign n37875 = n37874 ^ n37785;
  assign n37876 = n37875 ^ n37781;
  assign n37877 = n37782 & ~n37876;
  assign n37878 = n37877 ^ n37780;
  assign n37879 = n37878 ^ n37776;
  assign n37880 = n37777 & ~n37879;
  assign n37881 = n37880 ^ n37775;
  assign n37882 = n37881 ^ n37771;
  assign n37883 = n37772 & ~n37882;
  assign n37884 = n37883 ^ n37770;
  assign n37885 = n37884 ^ n37763;
  assign n37886 = n37767 & ~n37885;
  assign n37887 = n37886 ^ n37766;
  assign n37888 = n37887 ^ n37761;
  assign n37889 = n37762 & ~n37888;
  assign n37890 = n37889 ^ n3225;
  assign n37891 = n37890 ^ n37759;
  assign n37892 = ~n37760 & n37891;
  assign n37893 = n37892 ^ n2854;
  assign n37894 = n37893 ^ n37757;
  assign n37895 = n37758 & ~n37894;
  assign n37896 = n37895 ^ n2869;
  assign n37756 = n37705 ^ n37659;
  assign n37897 = n37896 ^ n37756;
  assign n2959 = n2955 ^ n2892;
  assign n2963 = n2962 ^ n2959;
  assign n2964 = n2963 ^ n1547;
  assign n37898 = n37756 ^ n2964;
  assign n37899 = n37897 & ~n37898;
  assign n37900 = n37899 ^ n2964;
  assign n37901 = n37900 ^ n37751;
  assign n37902 = n37755 & ~n37901;
  assign n37903 = n37902 ^ n37754;
  assign n37904 = n37903 ^ n37746;
  assign n37905 = n37750 & ~n37904;
  assign n37906 = n37905 ^ n37749;
  assign n37907 = n37906 ^ n37744;
  assign n37908 = n37745 & ~n37907;
  assign n37909 = n37908 ^ n37741;
  assign n37910 = n37909 ^ n37736;
  assign n37911 = n37740 & ~n37910;
  assign n37912 = n37911 ^ n37739;
  assign n37913 = n37912 ^ n37731;
  assign n37914 = n37735 & ~n37913;
  assign n37915 = n37914 ^ n37734;
  assign n2090 = n2053 ^ n2005;
  assign n2091 = n2090 ^ n2089;
  assign n2092 = n2091 ^ n2083;
  assign n37916 = n37915 ^ n2092;
  assign n37724 = n37513 ^ n34200;
  assign n37725 = n37649 ^ n37513;
  assign n37726 = n37724 & ~n37725;
  assign n37727 = n37726 ^ n34200;
  assign n37728 = n37727 ^ n34228;
  assign n37719 = n35047 ^ n34891;
  assign n37720 = n36405 ^ n34891;
  assign n37721 = n37719 & n37720;
  assign n37722 = n37721 ^ n35047;
  assign n37715 = n37512 ^ n37293;
  assign n37716 = ~n37508 & n37715;
  assign n37717 = n37716 ^ n37512;
  assign n37714 = n37057 ^ n36958;
  assign n37718 = n37717 ^ n37714;
  assign n37723 = n37722 ^ n37718;
  assign n37729 = n37728 ^ n37723;
  assign n37713 = n37651 & n37712;
  assign n37730 = n37729 ^ n37713;
  assign n37917 = n37916 ^ n37730;
  assign n37922 = n37921 ^ n37917;
  assign n37927 = n37912 ^ n37735;
  assign n37923 = n36623 ^ n35800;
  assign n37924 = n37406 ^ n36623;
  assign n37925 = n37923 & ~n37924;
  assign n37926 = n37925 ^ n35800;
  assign n37928 = n37927 ^ n37926;
  assign n37930 = n36515 ^ n35770;
  assign n37931 = n37412 ^ n36515;
  assign n37932 = ~n37930 & ~n37931;
  assign n37933 = n37932 ^ n35770;
  assign n37929 = n37909 ^ n37740;
  assign n37934 = n37933 ^ n37929;
  assign n37941 = n36464 ^ n35716;
  assign n37942 = n37414 ^ n36464;
  assign n37943 = n37941 & ~n37942;
  assign n37944 = n37943 ^ n35716;
  assign n37935 = n35934 ^ n34889;
  assign n37936 = n37250 ^ n35934;
  assign n37937 = ~n37935 & ~n37936;
  assign n37938 = n37937 ^ n34889;
  assign n37939 = n37903 ^ n37750;
  assign n37940 = n37938 & n37939;
  assign n37945 = n37944 ^ n37940;
  assign n37946 = n37906 ^ n37745;
  assign n37947 = n37946 ^ n37944;
  assign n37948 = n37945 & ~n37947;
  assign n37949 = n37948 ^ n37940;
  assign n37950 = n37949 ^ n37929;
  assign n37951 = n37934 & ~n37950;
  assign n37952 = n37951 ^ n37933;
  assign n37953 = n37952 ^ n37927;
  assign n37954 = n37928 & ~n37953;
  assign n37955 = n37954 ^ n37926;
  assign n37956 = n37955 ^ n37917;
  assign n37957 = n37922 & n37956;
  assign n37958 = n37957 ^ n37921;
  assign n37959 = n37958 ^ n37291;
  assign n37960 = ~n37292 & ~n37959;
  assign n37961 = n37960 ^ n37290;
  assign n37962 = n37961 ^ n37284;
  assign n37963 = n37285 & ~n37962;
  assign n37964 = n37963 ^ n37283;
  assign n37965 = n37964 ^ n37277;
  assign n37966 = ~n37278 & n37965;
  assign n37967 = n37966 ^ n37276;
  assign n37968 = n37967 ^ n37270;
  assign n37969 = n37271 & ~n37968;
  assign n37970 = n37969 ^ n37269;
  assign n37971 = n37970 ^ n37263;
  assign n37972 = n37264 & n37971;
  assign n37973 = n37972 ^ n37262;
  assign n37974 = n37973 ^ n37256;
  assign n37975 = n37257 & ~n37974;
  assign n37976 = n37975 ^ n36639;
  assign n38044 = n37981 ^ n37976;
  assign n38045 = ~n37982 & ~n38044;
  assign n38046 = n38045 ^ n37980;
  assign n38280 = n38047 ^ n38046;
  assign n38281 = ~n38052 & n38280;
  assign n38282 = n38281 ^ n38051;
  assign n38275 = n36673 ^ n36002;
  assign n38276 = n37352 ^ n36673;
  assign n38277 = n38275 & n38276;
  assign n38278 = n38277 ^ n36002;
  assign n38168 = n37833 ^ n37830;
  assign n38279 = n38278 ^ n38168;
  assign n38380 = n38282 ^ n38279;
  assign n38381 = n38380 ^ n34966;
  assign n38053 = n38052 ^ n38046;
  assign n38054 = n38053 ^ n34972;
  assign n37983 = n37982 ^ n37976;
  assign n37984 = n37983 ^ n34975;
  assign n37985 = n37973 ^ n37257;
  assign n37986 = n37985 ^ n34982;
  assign n37987 = n37970 ^ n37264;
  assign n37988 = n37987 ^ n34989;
  assign n37989 = n37967 ^ n37269;
  assign n37990 = n37989 ^ n37270;
  assign n37991 = n37990 ^ n34995;
  assign n37992 = n37964 ^ n37278;
  assign n37993 = n37992 ^ n35002;
  assign n37994 = n37961 ^ n37283;
  assign n37995 = n37994 ^ n37284;
  assign n37996 = n37995 ^ n35008;
  assign n37997 = n37958 ^ n37292;
  assign n37998 = n37997 ^ n34306;
  assign n37999 = n37955 ^ n37922;
  assign n38000 = n37999 ^ n35023;
  assign n38001 = n37952 ^ n37926;
  assign n38002 = n38001 ^ n37927;
  assign n38003 = n38002 ^ n34894;
  assign n38004 = n37949 ^ n37933;
  assign n38005 = n38004 ^ n37929;
  assign n38006 = n38005 ^ n35137;
  assign n38007 = n37939 ^ n37938;
  assign n38008 = ~n35041 & n38007;
  assign n38009 = n38008 ^ n35035;
  assign n38010 = n37946 ^ n37945;
  assign n38011 = n38010 ^ n38008;
  assign n38012 = n38009 & ~n38011;
  assign n38013 = n38012 ^ n35035;
  assign n38014 = n38013 ^ n38005;
  assign n38015 = n38006 & ~n38014;
  assign n38016 = n38015 ^ n35137;
  assign n38017 = n38016 ^ n38002;
  assign n38018 = ~n38003 & ~n38017;
  assign n38019 = n38018 ^ n34894;
  assign n38020 = n38019 ^ n37999;
  assign n38021 = ~n38000 & n38020;
  assign n38022 = n38021 ^ n35023;
  assign n38023 = n38022 ^ n37997;
  assign n38024 = ~n37998 & n38023;
  assign n38025 = n38024 ^ n34306;
  assign n38026 = n38025 ^ n37995;
  assign n38027 = ~n37996 & n38026;
  assign n38028 = n38027 ^ n35008;
  assign n38029 = n38028 ^ n37992;
  assign n38030 = ~n37993 & ~n38029;
  assign n38031 = n38030 ^ n35002;
  assign n38032 = n38031 ^ n37990;
  assign n38033 = n37991 & ~n38032;
  assign n38034 = n38033 ^ n34995;
  assign n38035 = n38034 ^ n37987;
  assign n38036 = n37988 & ~n38035;
  assign n38037 = n38036 ^ n34989;
  assign n38038 = n38037 ^ n37985;
  assign n38039 = n37986 & n38038;
  assign n38040 = n38039 ^ n34982;
  assign n38041 = n38040 ^ n37983;
  assign n38042 = ~n37984 & n38041;
  assign n38043 = n38042 ^ n34975;
  assign n38382 = n38053 ^ n38043;
  assign n38383 = ~n38054 & ~n38382;
  assign n38384 = n38383 ^ n34972;
  assign n38385 = n38384 ^ n38380;
  assign n38386 = ~n38381 & n38385;
  assign n38387 = n38386 ^ n34966;
  assign n38283 = n38282 ^ n38168;
  assign n38284 = ~n38279 & ~n38283;
  assign n38285 = n38284 ^ n38278;
  assign n38270 = n36670 ^ n36000;
  assign n38271 = n37342 ^ n36670;
  assign n38272 = ~n38270 & ~n38271;
  assign n38273 = n38272 ^ n36000;
  assign n38269 = n37836 ^ n37809;
  assign n38274 = n38273 ^ n38269;
  assign n38378 = n38285 ^ n38274;
  assign n38379 = n38378 ^ n34959;
  assign n38447 = n38387 ^ n38379;
  assign n38448 = n38384 ^ n38381;
  assign n38055 = n38054 ^ n38043;
  assign n38056 = n38022 ^ n37998;
  assign n38057 = n38013 ^ n38006;
  assign n38058 = n38016 ^ n38003;
  assign n38059 = ~n38057 & n38058;
  assign n38060 = n38019 ^ n38000;
  assign n38061 = n38059 & ~n38060;
  assign n38062 = n38056 & ~n38061;
  assign n38063 = n38025 ^ n37996;
  assign n38064 = ~n38062 & ~n38063;
  assign n38065 = n38028 ^ n37993;
  assign n38066 = n38064 & ~n38065;
  assign n38067 = n38031 ^ n37991;
  assign n38068 = ~n38066 & n38067;
  assign n38069 = n38034 ^ n37988;
  assign n38070 = n38068 & n38069;
  assign n38071 = n38037 ^ n37986;
  assign n38072 = ~n38070 & ~n38071;
  assign n38073 = n38040 ^ n37984;
  assign n38074 = n38072 & ~n38073;
  assign n38449 = ~n38055 & n38074;
  assign n38450 = n38448 & n38449;
  assign n38451 = n38447 & ~n38450;
  assign n38388 = n38387 ^ n38378;
  assign n38389 = n38379 & n38388;
  assign n38390 = n38389 ^ n34959;
  assign n38286 = n38285 ^ n38269;
  assign n38287 = n38274 & ~n38286;
  assign n38288 = n38287 ^ n38273;
  assign n38267 = n37843 ^ n37840;
  assign n38263 = n36664 ^ n35998;
  assign n38264 = n37340 ^ n36664;
  assign n38265 = ~n38263 & n38264;
  assign n38266 = n38265 ^ n35998;
  assign n38268 = n38267 ^ n38266;
  assign n38376 = n38288 ^ n38268;
  assign n38377 = n38376 ^ n34953;
  assign n38446 = n38390 ^ n38377;
  assign n38543 = n38451 ^ n38446;
  assign n1303 = n1293 ^ n1209;
  assign n1310 = n1309 ^ n1303;
  assign n1317 = n1316 ^ n1310;
  assign n38544 = n38543 ^ n1317;
  assign n38546 = n38449 ^ n38448;
  assign n1127 = n1107 ^ n1060;
  assign n1137 = n1136 ^ n1127;
  assign n1150 = n1149 ^ n1137;
  assign n38547 = n38546 ^ n1150;
  assign n38076 = n38073 ^ n38072;
  assign n38080 = n38079 ^ n38076;
  assign n38081 = n38071 ^ n38070;
  assign n38085 = n38084 ^ n38081;
  assign n38089 = n38069 ^ n38068;
  assign n38086 = n35839 ^ n27737;
  assign n38087 = n38086 ^ n32301;
  assign n38088 = n38087 ^ n738;
  assign n38090 = n38089 ^ n38088;
  assign n38095 = n38065 ^ n38064;
  assign n38092 = n35849 ^ n27747;
  assign n38093 = n38092 ^ n32308;
  assign n38094 = n38093 ^ n581;
  assign n38096 = n38095 ^ n38094;
  assign n38100 = n38063 ^ n38062;
  assign n38097 = n35854 ^ n708;
  assign n38098 = n38097 ^ n32313;
  assign n38099 = n38098 ^ n26539;
  assign n38101 = n38100 ^ n38099;
  assign n38103 = n35860 ^ n27753;
  assign n38104 = n38103 ^ n32319;
  assign n38105 = n38104 ^ n26544;
  assign n38102 = n38061 ^ n38056;
  assign n38106 = n38105 ^ n38102;
  assign n38110 = n38060 ^ n38059;
  assign n38107 = n35865 ^ n27759;
  assign n38108 = n38107 ^ n32324;
  assign n38109 = n38108 ^ n26562;
  assign n38111 = n38110 ^ n38109;
  assign n2394 = n2393 ^ n2288;
  assign n2395 = n2394 ^ n2351;
  assign n2396 = n2395 ^ n2388;
  assign n38113 = n38057 ^ n2396;
  assign n38114 = n36403 ^ n2170;
  assign n38115 = n38114 ^ n2377;
  assign n38116 = n38115 ^ n32743;
  assign n38117 = n38007 ^ n35041;
  assign n38118 = n38116 & ~n38117;
  assign n2367 = n2273 ^ n2202;
  assign n2371 = n2370 ^ n2367;
  assign n2381 = n2380 ^ n2371;
  assign n38119 = n38118 ^ n2381;
  assign n38120 = n38010 ^ n38009;
  assign n38121 = n38120 ^ n2381;
  assign n38122 = n38119 & ~n38121;
  assign n38123 = n38122 ^ n38118;
  assign n38124 = n38123 ^ n38057;
  assign n38125 = ~n38113 & n38124;
  assign n38126 = n38125 ^ n2396;
  assign n38112 = n38058 ^ n38057;
  assign n38127 = n38126 ^ n38112;
  assign n38128 = n35869 ^ n27763;
  assign n38129 = n38128 ^ n26556;
  assign n38130 = n38129 ^ n2406;
  assign n38131 = n38130 ^ n38112;
  assign n38132 = ~n38127 & n38131;
  assign n38133 = n38132 ^ n38130;
  assign n38134 = n38133 ^ n38110;
  assign n38135 = n38111 & ~n38134;
  assign n38136 = n38135 ^ n38109;
  assign n38137 = n38136 ^ n38102;
  assign n38138 = ~n38106 & n38137;
  assign n38139 = n38138 ^ n38105;
  assign n38140 = n38139 ^ n38100;
  assign n38141 = ~n38101 & n38140;
  assign n38142 = n38141 ^ n38099;
  assign n38143 = n38142 ^ n38095;
  assign n38144 = n38096 & ~n38143;
  assign n38145 = n38144 ^ n38094;
  assign n38091 = n38067 ^ n38066;
  assign n38146 = n38145 ^ n38091;
  assign n38147 = n35844 ^ n27742;
  assign n38148 = n38147 ^ n723;
  assign n38149 = n38148 ^ n26531;
  assign n38150 = n38149 ^ n38091;
  assign n38151 = n38146 & ~n38150;
  assign n38152 = n38151 ^ n38149;
  assign n38153 = n38152 ^ n38089;
  assign n38154 = n38090 & ~n38153;
  assign n38155 = n38154 ^ n38088;
  assign n38156 = n38155 ^ n38081;
  assign n38157 = ~n38085 & n38156;
  assign n38158 = n38157 ^ n38084;
  assign n38159 = n38158 ^ n38076;
  assign n38160 = n38080 & ~n38159;
  assign n38161 = n38160 ^ n38079;
  assign n38075 = n38074 ^ n38055;
  assign n38162 = n38161 ^ n38075;
  assign n38548 = n38075 ^ n3332;
  assign n38549 = ~n38162 & n38548;
  assign n38550 = n38549 ^ n3332;
  assign n38551 = n38550 ^ n38546;
  assign n38552 = ~n38547 & n38551;
  assign n38553 = n38552 ^ n1150;
  assign n38545 = n38450 ^ n38447;
  assign n38554 = n38553 ^ n38545;
  assign n1160 = n1123 ^ n1078;
  assign n1161 = n1160 ^ n1157;
  assign n1168 = n1167 ^ n1161;
  assign n38555 = n38545 ^ n1168;
  assign n38556 = n38554 & ~n38555;
  assign n38557 = n38556 ^ n1168;
  assign n38558 = n38557 ^ n38543;
  assign n38559 = ~n38544 & n38558;
  assign n38560 = n38559 ^ n1317;
  assign n38452 = ~n38446 & ~n38451;
  assign n38391 = n38390 ^ n38376;
  assign n38392 = ~n38377 & n38391;
  assign n38393 = n38392 ^ n34953;
  assign n38289 = n38288 ^ n38267;
  assign n38290 = ~n38268 & n38289;
  assign n38291 = n38290 ^ n38266;
  assign n38258 = n36654 ^ n35992;
  assign n38259 = n37334 ^ n36654;
  assign n38260 = n38258 & n38259;
  assign n38261 = n38260 ^ n35992;
  assign n38373 = n38291 ^ n38261;
  assign n38257 = n37846 ^ n37803;
  assign n38374 = n38373 ^ n38257;
  assign n38375 = n38374 ^ n34947;
  assign n38445 = n38393 ^ n38375;
  assign n38542 = n38452 ^ n38445;
  assign n38561 = n38560 ^ n38542;
  assign n38562 = n36337 ^ n27724;
  assign n38563 = n38562 ^ n1324;
  assign n38564 = n38563 ^ n26606;
  assign n38565 = n38564 ^ n38542;
  assign n38566 = ~n38561 & n38565;
  assign n38567 = n38566 ^ n38564;
  assign n38538 = n3146 ^ n1409;
  assign n38539 = n38538 ^ n32386;
  assign n38540 = n38539 ^ n26511;
  assign n38453 = ~n38445 & n38452;
  assign n38394 = n38393 ^ n38374;
  assign n38395 = ~n38375 & ~n38394;
  assign n38396 = n38395 ^ n34947;
  assign n38262 = n38261 ^ n38257;
  assign n38292 = n38291 ^ n38257;
  assign n38293 = n38262 & n38292;
  assign n38294 = n38293 ^ n38261;
  assign n38252 = n36648 ^ n35982;
  assign n38253 = n37472 ^ n36648;
  assign n38254 = n38252 & n38253;
  assign n38255 = n38254 ^ n35982;
  assign n38164 = n37853 ^ n37850;
  assign n38256 = n38255 ^ n38164;
  assign n38371 = n38294 ^ n38256;
  assign n38372 = n38371 ^ n34941;
  assign n38444 = n38396 ^ n38372;
  assign n38537 = n38453 ^ n38444;
  assign n38541 = n38540 ^ n38537;
  assign n38889 = n38567 ^ n38541;
  assign n38885 = n37499 ^ n37086;
  assign n38196 = n37887 ^ n37762;
  assign n38886 = n38196 ^ n37499;
  assign n38887 = n38885 & ~n38886;
  assign n38888 = n38887 ^ n37086;
  assign n38890 = n38889 ^ n38888;
  assign n38895 = n38564 ^ n38561;
  assign n38891 = n37298 ^ n36945;
  assign n38198 = n37884 ^ n37767;
  assign n38892 = n38198 ^ n37298;
  assign n38893 = ~n38891 & ~n38892;
  assign n38894 = n38893 ^ n36945;
  assign n38896 = n38895 ^ n38894;
  assign n38901 = n38557 ^ n38544;
  assign n38897 = n37304 ^ n36887;
  assign n38204 = n37881 ^ n37772;
  assign n38898 = n38204 ^ n37304;
  assign n38899 = n38897 & ~n38898;
  assign n38900 = n38899 ^ n36887;
  assign n38902 = n38901 ^ n38900;
  assign n38907 = n38554 ^ n1168;
  assign n38903 = n37310 ^ n36790;
  assign n38210 = n37878 ^ n37777;
  assign n38904 = n38210 ^ n37310;
  assign n38905 = n38903 & n38904;
  assign n38906 = n38905 ^ n36790;
  assign n38908 = n38907 ^ n38906;
  assign n38913 = n38550 ^ n38547;
  assign n38909 = n37316 ^ n36645;
  assign n38220 = n37875 ^ n37782;
  assign n38910 = n38220 ^ n37316;
  assign n38911 = ~n38909 & ~n38910;
  assign n38912 = n38911 ^ n36645;
  assign n38914 = n38913 ^ n38912;
  assign n38915 = n37322 ^ n36648;
  assign n38226 = n37872 ^ n37787;
  assign n38916 = n38226 ^ n37322;
  assign n38917 = ~n38915 & ~n38916;
  assign n38918 = n38917 ^ n36648;
  assign n38163 = n38162 ^ n3332;
  assign n38919 = n38918 ^ n38163;
  assign n38924 = n38158 ^ n38080;
  assign n38920 = n37328 ^ n36654;
  assign n38228 = n37869 ^ n37792;
  assign n38921 = n38228 ^ n37328;
  assign n38922 = n38920 & ~n38921;
  assign n38923 = n38922 ^ n36654;
  assign n38925 = n38924 ^ n38923;
  assign n38930 = n38155 ^ n38085;
  assign n38926 = n37472 ^ n36664;
  assign n38234 = n37866 ^ n37797;
  assign n38927 = n38234 ^ n37472;
  assign n38928 = n38926 & n38927;
  assign n38929 = n38928 ^ n36664;
  assign n38931 = n38930 ^ n38929;
  assign n38936 = n38152 ^ n38090;
  assign n38932 = n37334 ^ n36670;
  assign n38240 = n37863 ^ n37860;
  assign n38933 = n38240 ^ n37334;
  assign n38934 = ~n38932 & ~n38933;
  assign n38935 = n38934 ^ n36670;
  assign n38937 = n38936 ^ n38935;
  assign n38942 = n38149 ^ n38146;
  assign n38938 = n37340 ^ n36673;
  assign n38246 = n37856 ^ n37800;
  assign n38939 = n38246 ^ n37340;
  assign n38940 = n38938 & n38939;
  assign n38941 = n38940 ^ n36673;
  assign n38943 = n38942 ^ n38941;
  assign n38948 = n38142 ^ n38096;
  assign n38944 = n37342 ^ n36679;
  assign n38945 = n38164 ^ n37342;
  assign n38946 = ~n38944 & n38945;
  assign n38947 = n38946 ^ n36679;
  assign n38949 = n38948 ^ n38947;
  assign n38954 = n38139 ^ n38101;
  assign n38950 = n37352 ^ n36686;
  assign n38951 = n38257 ^ n37352;
  assign n38952 = ~n38950 & ~n38951;
  assign n38953 = n38952 ^ n36686;
  assign n38955 = n38954 ^ n38953;
  assign n38727 = n37364 ^ n36702;
  assign n38728 = n38269 ^ n37364;
  assign n38729 = n38727 & ~n38728;
  assign n38730 = n38729 ^ n36702;
  assign n38726 = n38133 ^ n38111;
  assign n38731 = n38730 ^ n38726;
  assign n38167 = n36708 ^ n36636;
  assign n38169 = n38168 ^ n36636;
  assign n38170 = n38167 & ~n38169;
  assign n38171 = n38170 ^ n36708;
  assign n38166 = n38130 ^ n38127;
  assign n38732 = n38171 ^ n38166;
  assign n38671 = n38123 ^ n38113;
  assign n38173 = n37266 ^ n36717;
  assign n38174 = n37981 ^ n37266;
  assign n38175 = n38173 & n38174;
  assign n38176 = n38175 ^ n36717;
  assign n38172 = n38120 ^ n38119;
  assign n38177 = n38176 ^ n38172;
  assign n38179 = n37273 ^ n36724;
  assign n38180 = n37273 ^ n37256;
  assign n38181 = ~n38179 & n38180;
  assign n38182 = n38181 ^ n36724;
  assign n38178 = n38117 ^ n38116;
  assign n38183 = n38182 ^ n38178;
  assign n38624 = n37280 ^ n36730;
  assign n38625 = n37280 ^ n37263;
  assign n38626 = n38624 & n38625;
  assign n38627 = n38626 ^ n36730;
  assign n38199 = n36428 ^ n35673;
  assign n38200 = n37714 ^ n36428;
  assign n38201 = n38199 & n38200;
  assign n38202 = n38201 ^ n35673;
  assign n38203 = n38202 ^ n38198;
  assign n38205 = n36435 ^ n35680;
  assign n38206 = n37293 ^ n36435;
  assign n38207 = n38205 & n38206;
  assign n38208 = n38207 ^ n35680;
  assign n38209 = n38208 ^ n38204;
  assign n38211 = n37179 ^ n36265;
  assign n38212 = n37499 ^ n37179;
  assign n38213 = ~n38211 & n38212;
  assign n38214 = n38213 ^ n36265;
  assign n38215 = n38214 ^ n38210;
  assign n38216 = n37132 ^ n35948;
  assign n38217 = n37298 ^ n37132;
  assign n38218 = n38216 & n38217;
  assign n38219 = n38218 ^ n35948;
  assign n38221 = n38220 ^ n38219;
  assign n38222 = n37086 ^ n35950;
  assign n38223 = n37304 ^ n37086;
  assign n38224 = n38222 & ~n38223;
  assign n38225 = n38224 ^ n35950;
  assign n38227 = n38226 ^ n38225;
  assign n38229 = n36945 ^ n35960;
  assign n38230 = n37310 ^ n36945;
  assign n38231 = n38229 & ~n38230;
  assign n38232 = n38231 ^ n35960;
  assign n38233 = n38232 ^ n38228;
  assign n38235 = n36887 ^ n35966;
  assign n38236 = n37316 ^ n36887;
  assign n38237 = ~n38235 & ~n38236;
  assign n38238 = n38237 ^ n35966;
  assign n38239 = n38238 ^ n38234;
  assign n38241 = n36790 ^ n35972;
  assign n38242 = n37322 ^ n36790;
  assign n38243 = ~n38241 & n38242;
  assign n38244 = n38243 ^ n35972;
  assign n38245 = n38244 ^ n38240;
  assign n38247 = n36645 ^ n35979;
  assign n38248 = n37328 ^ n36645;
  assign n38249 = n38247 & n38248;
  assign n38250 = n38249 ^ n35979;
  assign n38251 = n38250 ^ n38246;
  assign n38295 = n38294 ^ n38164;
  assign n38296 = n38256 & n38295;
  assign n38297 = n38296 ^ n38255;
  assign n38298 = n38297 ^ n38246;
  assign n38299 = ~n38251 & n38298;
  assign n38300 = n38299 ^ n38250;
  assign n38301 = n38300 ^ n38240;
  assign n38302 = ~n38245 & ~n38301;
  assign n38303 = n38302 ^ n38244;
  assign n38304 = n38303 ^ n38234;
  assign n38305 = n38239 & n38304;
  assign n38306 = n38305 ^ n38238;
  assign n38307 = n38306 ^ n38228;
  assign n38308 = ~n38233 & n38307;
  assign n38309 = n38308 ^ n38232;
  assign n38310 = n38309 ^ n38226;
  assign n38311 = n38227 & n38310;
  assign n38312 = n38311 ^ n38225;
  assign n38313 = n38312 ^ n38220;
  assign n38314 = ~n38221 & ~n38313;
  assign n38315 = n38314 ^ n38219;
  assign n38316 = n38315 ^ n38210;
  assign n38317 = n38215 & n38316;
  assign n38318 = n38317 ^ n38214;
  assign n38319 = n38318 ^ n38204;
  assign n38320 = ~n38209 & ~n38319;
  assign n38321 = n38320 ^ n38208;
  assign n38322 = n38321 ^ n38198;
  assign n38323 = n38203 & n38322;
  assign n38324 = n38323 ^ n38202;
  assign n38192 = n36418 ^ n35667;
  assign n38193 = n37102 ^ n36418;
  assign n38194 = n38192 & n38193;
  assign n38195 = n38194 ^ n35667;
  assign n38197 = n38196 ^ n38195;
  assign n38350 = n38324 ^ n38197;
  assign n38351 = n38350 ^ n34847;
  assign n38352 = n38321 ^ n38203;
  assign n38353 = n38352 ^ n34864;
  assign n38354 = n38318 ^ n38209;
  assign n38355 = n38354 ^ n34857;
  assign n38356 = n38315 ^ n38214;
  assign n38357 = n38356 ^ n38210;
  assign n38358 = n38357 ^ n35430;
  assign n38359 = n38312 ^ n38221;
  assign n38360 = n38359 ^ n34900;
  assign n38361 = n38309 ^ n38227;
  assign n38362 = n38361 ^ n34902;
  assign n38363 = n38306 ^ n38233;
  assign n38364 = n38363 ^ n34912;
  assign n38365 = n38303 ^ n38239;
  assign n38366 = n38365 ^ n34919;
  assign n38367 = n38300 ^ n38245;
  assign n38368 = n38367 ^ n34926;
  assign n38369 = n38297 ^ n38251;
  assign n38370 = n38369 ^ n34934;
  assign n38397 = n38396 ^ n38371;
  assign n38398 = n38372 & ~n38397;
  assign n38399 = n38398 ^ n34941;
  assign n38400 = n38399 ^ n38369;
  assign n38401 = ~n38370 & ~n38400;
  assign n38402 = n38401 ^ n34934;
  assign n38403 = n38402 ^ n38367;
  assign n38404 = n38368 & n38403;
  assign n38405 = n38404 ^ n34926;
  assign n38406 = n38405 ^ n38365;
  assign n38407 = n38366 & ~n38406;
  assign n38408 = n38407 ^ n34919;
  assign n38409 = n38408 ^ n38363;
  assign n38410 = ~n38364 & ~n38409;
  assign n38411 = n38410 ^ n34912;
  assign n38412 = n38411 ^ n38361;
  assign n38413 = n38362 & ~n38412;
  assign n38414 = n38413 ^ n34902;
  assign n38415 = n38414 ^ n38359;
  assign n38416 = ~n38360 & ~n38415;
  assign n38417 = n38416 ^ n34900;
  assign n38418 = n38417 ^ n38357;
  assign n38419 = n38358 & n38418;
  assign n38420 = n38419 ^ n35430;
  assign n38421 = n38420 ^ n38354;
  assign n38422 = n38355 & ~n38421;
  assign n38423 = n38422 ^ n34857;
  assign n38424 = n38423 ^ n38352;
  assign n38425 = n38353 & ~n38424;
  assign n38426 = n38425 ^ n34864;
  assign n38427 = n38426 ^ n38350;
  assign n38428 = ~n38351 & ~n38427;
  assign n38429 = n38428 ^ n34847;
  assign n38325 = n38324 ^ n38196;
  assign n38326 = ~n38197 & ~n38325;
  assign n38327 = n38326 ^ n38195;
  assign n38190 = n37890 ^ n37760;
  assign n38186 = n36415 ^ n35660;
  assign n38187 = n37109 ^ n36415;
  assign n38188 = ~n38186 & ~n38187;
  assign n38189 = n38188 ^ n35660;
  assign n38191 = n38190 ^ n38189;
  assign n38348 = n38327 ^ n38191;
  assign n38349 = n38348 ^ n35109;
  assign n38437 = n38429 ^ n38349;
  assign n38438 = n38423 ^ n38353;
  assign n38439 = n38420 ^ n38355;
  assign n38440 = n38417 ^ n38358;
  assign n38441 = n38414 ^ n38360;
  assign n38442 = n38408 ^ n38364;
  assign n38443 = n38399 ^ n38370;
  assign n38454 = ~n38444 & n38453;
  assign n38455 = ~n38443 & ~n38454;
  assign n38456 = n38402 ^ n38368;
  assign n38457 = ~n38455 & n38456;
  assign n38458 = n38405 ^ n38366;
  assign n38459 = n38457 & ~n38458;
  assign n38460 = ~n38442 & ~n38459;
  assign n38461 = n38411 ^ n38362;
  assign n38462 = n38460 & ~n38461;
  assign n38463 = n38441 & n38462;
  assign n38464 = ~n38440 & ~n38463;
  assign n38465 = n38439 & n38464;
  assign n38466 = n38438 & n38465;
  assign n38467 = n38426 ^ n38351;
  assign n38468 = n38466 & ~n38467;
  assign n38469 = n38437 & ~n38468;
  assign n38430 = n38429 ^ n38348;
  assign n38431 = n38349 & n38430;
  assign n38432 = n38431 ^ n35109;
  assign n38470 = n38432 ^ n35103;
  assign n38332 = n36405 ^ n35654;
  assign n38333 = n37092 ^ n36405;
  assign n38334 = n38332 & ~n38333;
  assign n38335 = n38334 ^ n35654;
  assign n38328 = n38327 ^ n38190;
  assign n38329 = n38191 & ~n38328;
  assign n38330 = n38329 ^ n38189;
  assign n38185 = n37893 ^ n37758;
  assign n38331 = n38330 ^ n38185;
  assign n38346 = n38335 ^ n38331;
  assign n38471 = n38470 ^ n38346;
  assign n38472 = n38469 & ~n38471;
  assign n38347 = n38346 ^ n35103;
  assign n38433 = n38432 ^ n38346;
  assign n38434 = n38347 & n38433;
  assign n38435 = n38434 ^ n35103;
  assign n38340 = n35946 ^ n34898;
  assign n38341 = n37147 ^ n35946;
  assign n38342 = n38340 & ~n38341;
  assign n38343 = n38342 ^ n34898;
  assign n38336 = n38335 ^ n38185;
  assign n38337 = n38331 & ~n38336;
  assign n38338 = n38337 ^ n38335;
  assign n38184 = n37897 ^ n2964;
  assign n38339 = n38338 ^ n38184;
  assign n38344 = n38343 ^ n38339;
  assign n38345 = n38344 ^ n35049;
  assign n38436 = n38435 ^ n38345;
  assign n38493 = n38472 ^ n38436;
  assign n38490 = n36285 ^ n28150;
  assign n38491 = n38490 ^ n26798;
  assign n38492 = n38491 ^ n1832;
  assign n38494 = n38493 ^ n38492;
  assign n38498 = n38471 ^ n38469;
  assign n38495 = n36290 ^ n28155;
  assign n38496 = n38495 ^ n32485;
  assign n38497 = n38496 ^ n1827;
  assign n38499 = n38498 ^ n38497;
  assign n38502 = n36297 ^ n28161;
  assign n38503 = n38502 ^ n1742;
  assign n38504 = n38503 ^ n32233;
  assign n38501 = n38467 ^ n38466;
  assign n38505 = n38504 ^ n38501;
  assign n38507 = n3002 ^ n1647;
  assign n38508 = n38507 ^ n32238;
  assign n38509 = n38508 ^ n26645;
  assign n38506 = n38465 ^ n38438;
  assign n38510 = n38509 ^ n38506;
  assign n38513 = n36307 ^ n2921;
  assign n38514 = n38513 ^ n32262;
  assign n38515 = n38514 ^ n3128;
  assign n38512 = n38463 ^ n38440;
  assign n38516 = n38515 ^ n38512;
  assign n38517 = n38462 ^ n38441;
  assign n38521 = n38520 ^ n38517;
  assign n38523 = n36317 ^ n3233;
  assign n38524 = n38523 ^ n2645;
  assign n38525 = n38524 ^ n3098;
  assign n38522 = n38461 ^ n38460;
  assign n38526 = n38525 ^ n38522;
  assign n38527 = n38459 ^ n38442;
  assign n3078 = n3077 ^ n3071;
  assign n3082 = n3081 ^ n3078;
  assign n3083 = n3082 ^ n2643;
  assign n38528 = n38527 ^ n3083;
  assign n38529 = n38458 ^ n38457;
  assign n2547 = n2546 ^ n2531;
  assign n2566 = n2565 ^ n2547;
  assign n2573 = n2572 ^ n2566;
  assign n38530 = n38529 ^ n2573;
  assign n38534 = n38456 ^ n38455;
  assign n38531 = n36325 ^ n3053;
  assign n38532 = n38531 ^ n3167;
  assign n38533 = n38532 ^ n2560;
  assign n38535 = n38534 ^ n38533;
  assign n38568 = n38567 ^ n38537;
  assign n38569 = n38541 & ~n38568;
  assign n38570 = n38569 ^ n38540;
  assign n38536 = n38454 ^ n38443;
  assign n38571 = n38570 ^ n38536;
  assign n38572 = n36331 ^ n2484;
  assign n38573 = n38572 ^ n32380;
  assign n38574 = n38573 ^ n3165;
  assign n38575 = n38574 ^ n38536;
  assign n38576 = ~n38571 & n38575;
  assign n38577 = n38576 ^ n38574;
  assign n38578 = n38577 ^ n38534;
  assign n38579 = n38535 & ~n38578;
  assign n38580 = n38579 ^ n38533;
  assign n38581 = n38580 ^ n38529;
  assign n38582 = n38530 & ~n38581;
  assign n38583 = n38582 ^ n2573;
  assign n38584 = n38583 ^ n38527;
  assign n38585 = n38528 & ~n38584;
  assign n38586 = n38585 ^ n3083;
  assign n38587 = n38586 ^ n38522;
  assign n38588 = ~n38526 & n38587;
  assign n38589 = n38588 ^ n38525;
  assign n38590 = n38589 ^ n38517;
  assign n38591 = n38521 & ~n38590;
  assign n38592 = n38591 ^ n38520;
  assign n38593 = n38592 ^ n38512;
  assign n38594 = ~n38516 & n38593;
  assign n38595 = n38594 ^ n38515;
  assign n38511 = n38464 ^ n38439;
  assign n38596 = n38595 ^ n38511;
  assign n38600 = n38599 ^ n38511;
  assign n38601 = n38596 & ~n38600;
  assign n38602 = n38601 ^ n38599;
  assign n38603 = n38602 ^ n38506;
  assign n38604 = ~n38510 & n38603;
  assign n38605 = n38604 ^ n38509;
  assign n38606 = n38605 ^ n38501;
  assign n38607 = n38505 & ~n38606;
  assign n38608 = n38607 ^ n38504;
  assign n38500 = n38468 ^ n38437;
  assign n38609 = n38608 ^ n38500;
  assign n1716 = n1715 ^ n1697;
  assign n1732 = n1731 ^ n1716;
  assign n1745 = n1744 ^ n1732;
  assign n38610 = n38500 ^ n1745;
  assign n38611 = n38609 & ~n38610;
  assign n38612 = n38611 ^ n1745;
  assign n38613 = n38612 ^ n38498;
  assign n38614 = ~n38499 & n38613;
  assign n38615 = n38614 ^ n38497;
  assign n38616 = n38615 ^ n38493;
  assign n38617 = ~n38494 & n38616;
  assign n38618 = n38617 ^ n38492;
  assign n38622 = n38621 ^ n38618;
  assign n38484 = n38435 ^ n38344;
  assign n38485 = ~n38345 & n38484;
  assign n38486 = n38485 ^ n35049;
  assign n38487 = n38486 ^ n35047;
  assign n38479 = n38343 ^ n38184;
  assign n38480 = ~n38339 & n38479;
  assign n38481 = n38480 ^ n38343;
  assign n38475 = n35940 ^ n34891;
  assign n38476 = n37192 ^ n35940;
  assign n38477 = n38475 & n38476;
  assign n38478 = n38477 ^ n34891;
  assign n38482 = n38481 ^ n38478;
  assign n38474 = n37900 ^ n37755;
  assign n38483 = n38482 ^ n38474;
  assign n38488 = n38487 ^ n38483;
  assign n38473 = ~n38436 & n38472;
  assign n38489 = n38488 ^ n38473;
  assign n38623 = n38622 ^ n38489;
  assign n38628 = n38627 ^ n38623;
  assign n38630 = n37287 ^ n36623;
  assign n38631 = n37287 ^ n37270;
  assign n38632 = ~n38630 & n38631;
  assign n38633 = n38632 ^ n36623;
  assign n38629 = n38615 ^ n38494;
  assign n38634 = n38633 ^ n38629;
  assign n38636 = n37400 ^ n36515;
  assign n38637 = n37400 ^ n37277;
  assign n38638 = ~n38636 & n38637;
  assign n38639 = n38638 ^ n36515;
  assign n38635 = n38612 ^ n38499;
  assign n38640 = n38639 ^ n38635;
  assign n38642 = n37406 ^ n36464;
  assign n38643 = n37406 ^ n37284;
  assign n38644 = n38642 & ~n38643;
  assign n38645 = n38644 ^ n36464;
  assign n38641 = n38609 ^ n1745;
  assign n38646 = n38645 ^ n38641;
  assign n38647 = n38605 ^ n38505;
  assign n38648 = n37412 ^ n35934;
  assign n38649 = n37412 ^ n37291;
  assign n38650 = n38648 & ~n38649;
  assign n38651 = n38650 ^ n35934;
  assign n38652 = n38647 & ~n38651;
  assign n38653 = n38652 ^ n38641;
  assign n38654 = n38646 & ~n38653;
  assign n38655 = n38654 ^ n38652;
  assign n38656 = n38655 ^ n38635;
  assign n38657 = n38640 & n38656;
  assign n38658 = n38657 ^ n38639;
  assign n38659 = n38658 ^ n38629;
  assign n38660 = ~n38634 & ~n38659;
  assign n38661 = n38660 ^ n38633;
  assign n38662 = n38661 ^ n38623;
  assign n38663 = n38628 & ~n38662;
  assign n38664 = n38663 ^ n38627;
  assign n38665 = n38664 ^ n38178;
  assign n38666 = n38183 & n38665;
  assign n38667 = n38666 ^ n38182;
  assign n38668 = n38667 ^ n38172;
  assign n38669 = n38177 & n38668;
  assign n38670 = n38669 ^ n38176;
  assign n38672 = n38671 ^ n38670;
  assign n38673 = n37259 ^ n36715;
  assign n38674 = n38047 ^ n37259;
  assign n38675 = ~n38673 & n38674;
  assign n38676 = n38675 ^ n36715;
  assign n38677 = n38676 ^ n38671;
  assign n38678 = n38672 & n38677;
  assign n38679 = n38678 ^ n38676;
  assign n38733 = n38679 ^ n38166;
  assign n38734 = n38732 & n38733;
  assign n38735 = n38734 ^ n38171;
  assign n38832 = n38735 ^ n38730;
  assign n38833 = ~n38731 & n38832;
  assign n38834 = n38833 ^ n38726;
  assign n38830 = n38136 ^ n38106;
  assign n38956 = n38834 ^ n38830;
  assign n38826 = n37358 ^ n35927;
  assign n38827 = n38267 ^ n37358;
  assign n38828 = ~n38826 & ~n38827;
  assign n38829 = n38828 ^ n35927;
  assign n38957 = n38834 ^ n38829;
  assign n38958 = ~n38956 & n38957;
  assign n38959 = n38958 ^ n38830;
  assign n38960 = n38959 ^ n38954;
  assign n38961 = n38955 & ~n38960;
  assign n38962 = n38961 ^ n38953;
  assign n38963 = n38962 ^ n38948;
  assign n38964 = ~n38949 & n38963;
  assign n38965 = n38964 ^ n38947;
  assign n38966 = n38965 ^ n38942;
  assign n38967 = n38943 & ~n38966;
  assign n38968 = n38967 ^ n38941;
  assign n38969 = n38968 ^ n38936;
  assign n38970 = n38937 & n38969;
  assign n38971 = n38970 ^ n38935;
  assign n38972 = n38971 ^ n38930;
  assign n38973 = ~n38931 & n38972;
  assign n38974 = n38973 ^ n38929;
  assign n38975 = n38974 ^ n38924;
  assign n38976 = n38925 & ~n38975;
  assign n38977 = n38976 ^ n38923;
  assign n38978 = n38977 ^ n38163;
  assign n38979 = ~n38919 & ~n38978;
  assign n38980 = n38979 ^ n38918;
  assign n38981 = n38980 ^ n38913;
  assign n38982 = n38914 & ~n38981;
  assign n38983 = n38982 ^ n38912;
  assign n38984 = n38983 ^ n38907;
  assign n38985 = n38908 & ~n38984;
  assign n38986 = n38985 ^ n38906;
  assign n38987 = n38986 ^ n38901;
  assign n38988 = ~n38902 & ~n38987;
  assign n38989 = n38988 ^ n38900;
  assign n38990 = n38989 ^ n38895;
  assign n38991 = ~n38896 & ~n38990;
  assign n38992 = n38991 ^ n38894;
  assign n38993 = n38992 ^ n38889;
  assign n38994 = n38890 & n38993;
  assign n38995 = n38994 ^ n38888;
  assign n38883 = n38574 ^ n38571;
  assign n38879 = n37293 ^ n37132;
  assign n38880 = n38190 ^ n37293;
  assign n38881 = ~n38879 & n38880;
  assign n38882 = n38881 ^ n37132;
  assign n38884 = n38883 ^ n38882;
  assign n39044 = n38995 ^ n38884;
  assign n39045 = n39044 ^ n35948;
  assign n39046 = n38992 ^ n38890;
  assign n39047 = n39046 ^ n35950;
  assign n39048 = n38989 ^ n38896;
  assign n39049 = n39048 ^ n35960;
  assign n39050 = n38986 ^ n38902;
  assign n39051 = n39050 ^ n35966;
  assign n39052 = n38983 ^ n38908;
  assign n39053 = n39052 ^ n35972;
  assign n39054 = n38980 ^ n38914;
  assign n39055 = n39054 ^ n35979;
  assign n39056 = n38977 ^ n38919;
  assign n39057 = n39056 ^ n35982;
  assign n39058 = n38974 ^ n38925;
  assign n39059 = n39058 ^ n35992;
  assign n39060 = n38971 ^ n38931;
  assign n39061 = n39060 ^ n35998;
  assign n39062 = n38968 ^ n38935;
  assign n39063 = n39062 ^ n38936;
  assign n39064 = n39063 ^ n36000;
  assign n39065 = n38965 ^ n38941;
  assign n39066 = n39065 ^ n38942;
  assign n39067 = n39066 ^ n36002;
  assign n39068 = n38962 ^ n38947;
  assign n39069 = n39068 ^ n38948;
  assign n39070 = n39069 ^ n36008;
  assign n39071 = n38959 ^ n38953;
  assign n39072 = n39071 ^ n38954;
  assign n39073 = n39072 ^ n36019;
  assign n38680 = n38679 ^ n38171;
  assign n38681 = n38680 ^ n38166;
  assign n38682 = n38681 ^ n36055;
  assign n38683 = n38676 ^ n38672;
  assign n38684 = n38683 ^ n36034;
  assign n38685 = n38667 ^ n38176;
  assign n38686 = n38685 ^ n38172;
  assign n38687 = n38686 ^ n36040;
  assign n38688 = n38664 ^ n38183;
  assign n38689 = n38688 ^ n35917;
  assign n38690 = n38661 ^ n38628;
  assign n38691 = n38690 ^ n35816;
  assign n38692 = n38658 ^ n38633;
  assign n38693 = n38692 ^ n38629;
  assign n38694 = n38693 ^ n35800;
  assign n38695 = n38655 ^ n38640;
  assign n38696 = n38695 ^ n35770;
  assign n38697 = n38651 ^ n38647;
  assign n38698 = n34889 & ~n38697;
  assign n38699 = n38698 ^ n35716;
  assign n38700 = n38652 ^ n38645;
  assign n38701 = n38700 ^ n38641;
  assign n38702 = n38701 ^ n38698;
  assign n38703 = n38699 & n38702;
  assign n38704 = n38703 ^ n35716;
  assign n38705 = n38704 ^ n38695;
  assign n38706 = n38696 & ~n38705;
  assign n38707 = n38706 ^ n35770;
  assign n38708 = n38707 ^ n38693;
  assign n38709 = n38694 & ~n38708;
  assign n38710 = n38709 ^ n35800;
  assign n38711 = n38710 ^ n38690;
  assign n38712 = ~n38691 & ~n38711;
  assign n38713 = n38712 ^ n35816;
  assign n38714 = n38713 ^ n38688;
  assign n38715 = n38689 & n38714;
  assign n38716 = n38715 ^ n35917;
  assign n38717 = n38716 ^ n38686;
  assign n38718 = ~n38687 & n38717;
  assign n38719 = n38718 ^ n36040;
  assign n38720 = n38719 ^ n38683;
  assign n38721 = n38684 & ~n38720;
  assign n38722 = n38721 ^ n36034;
  assign n38723 = n38722 ^ n38681;
  assign n38724 = ~n38682 & n38723;
  assign n38725 = n38724 ^ n36055;
  assign n38837 = n38725 ^ n36031;
  assign n38736 = n38735 ^ n38731;
  assign n38838 = n38736 ^ n38725;
  assign n38839 = ~n38837 & n38838;
  assign n38840 = n38839 ^ n36031;
  assign n39074 = n38840 ^ n35928;
  assign n38831 = n38830 ^ n38829;
  assign n38835 = n38834 ^ n38831;
  assign n39075 = n38840 ^ n38835;
  assign n39076 = n39074 & n39075;
  assign n39077 = n39076 ^ n35928;
  assign n39078 = n39077 ^ n39072;
  assign n39079 = ~n39073 & ~n39078;
  assign n39080 = n39079 ^ n36019;
  assign n39081 = n39080 ^ n39069;
  assign n39082 = n39070 & ~n39081;
  assign n39083 = n39082 ^ n36008;
  assign n39084 = n39083 ^ n39066;
  assign n39085 = n39067 & n39084;
  assign n39086 = n39085 ^ n36002;
  assign n39087 = n39086 ^ n39063;
  assign n39088 = n39064 & ~n39087;
  assign n39089 = n39088 ^ n36000;
  assign n39090 = n39089 ^ n39060;
  assign n39091 = n39061 & ~n39090;
  assign n39092 = n39091 ^ n35998;
  assign n39093 = n39092 ^ n39058;
  assign n39094 = n39059 & n39093;
  assign n39095 = n39094 ^ n35992;
  assign n39096 = n39095 ^ n39056;
  assign n39097 = n39057 & n39096;
  assign n39098 = n39097 ^ n35982;
  assign n39099 = n39098 ^ n39054;
  assign n39100 = n39055 & ~n39099;
  assign n39101 = n39100 ^ n35979;
  assign n39102 = n39101 ^ n39052;
  assign n39103 = ~n39053 & ~n39102;
  assign n39104 = n39103 ^ n35972;
  assign n39105 = n39104 ^ n39050;
  assign n39106 = ~n39051 & ~n39105;
  assign n39107 = n39106 ^ n35966;
  assign n39108 = n39107 ^ n39048;
  assign n39109 = n39049 & ~n39108;
  assign n39110 = n39109 ^ n35960;
  assign n39111 = n39110 ^ n39046;
  assign n39112 = ~n39047 & ~n39111;
  assign n39113 = n39112 ^ n35950;
  assign n39114 = n39113 ^ n39044;
  assign n39115 = n39045 & n39114;
  assign n39116 = n39115 ^ n35948;
  assign n38996 = n38995 ^ n38883;
  assign n38997 = ~n38884 & ~n38996;
  assign n38998 = n38997 ^ n38882;
  assign n38874 = n37714 ^ n37179;
  assign n38875 = n38185 ^ n37714;
  assign n38876 = n38874 & n38875;
  assign n38877 = n38876 ^ n37179;
  assign n39041 = n38998 ^ n38877;
  assign n38873 = n38577 ^ n38535;
  assign n39042 = n39041 ^ n38873;
  assign n39043 = n39042 ^ n36265;
  assign n39167 = n39116 ^ n39043;
  assign n39139 = n39107 ^ n39049;
  assign n39140 = n39104 ^ n39051;
  assign n39141 = n39095 ^ n39057;
  assign n39142 = n39089 ^ n39061;
  assign n39143 = n39083 ^ n39067;
  assign n39144 = n39080 ^ n39070;
  assign n39145 = n39077 ^ n39073;
  assign n38737 = n38736 ^ n36031;
  assign n38738 = n38737 ^ n38725;
  assign n38739 = n38704 ^ n38696;
  assign n38740 = n38707 ^ n38694;
  assign n38741 = ~n38739 & ~n38740;
  assign n38742 = n38710 ^ n38691;
  assign n38743 = n38741 & n38742;
  assign n38744 = n38713 ^ n38689;
  assign n38745 = ~n38743 & ~n38744;
  assign n38746 = n38716 ^ n38687;
  assign n38747 = ~n38745 & n38746;
  assign n38748 = n38719 ^ n38684;
  assign n38749 = n38747 & ~n38748;
  assign n38750 = n38722 ^ n38682;
  assign n38751 = ~n38749 & ~n38750;
  assign n38825 = n38738 & n38751;
  assign n38836 = n38835 ^ n35928;
  assign n38841 = n38840 ^ n38836;
  assign n39146 = ~n38825 & ~n38841;
  assign n39147 = ~n39145 & n39146;
  assign n39148 = ~n39144 & n39147;
  assign n39149 = ~n39143 & n39148;
  assign n39150 = n39086 ^ n36000;
  assign n39151 = n39150 ^ n39063;
  assign n39152 = ~n39149 & ~n39151;
  assign n39153 = n39142 & ~n39152;
  assign n39154 = n39092 ^ n39059;
  assign n39155 = n39153 & n39154;
  assign n39156 = ~n39141 & n39155;
  assign n39157 = n39098 ^ n39055;
  assign n39158 = ~n39156 & ~n39157;
  assign n39159 = n39101 ^ n39053;
  assign n39160 = ~n39158 & ~n39159;
  assign n39161 = n39140 & n39160;
  assign n39162 = ~n39139 & ~n39161;
  assign n39163 = n39110 ^ n39047;
  assign n39164 = n39162 & n39163;
  assign n39165 = n39113 ^ n39045;
  assign n39166 = n39164 & n39165;
  assign n39220 = n39167 ^ n39166;
  assign n2820 = n2819 ^ n2762;
  assign n2827 = n2826 ^ n2820;
  assign n2828 = n2827 ^ n1592;
  assign n39221 = n39220 ^ n2828;
  assign n39222 = n39165 ^ n39164;
  assign n3115 = n3110 ^ n3105;
  assign n3116 = n3115 ^ n2737;
  assign n3117 = n3116 ^ n2824;
  assign n39223 = n39222 ^ n3117;
  assign n39224 = n39163 ^ n39162;
  assign n2704 = n2700 ^ n2673;
  assign n2723 = n2722 ^ n2704;
  assign n2730 = n2729 ^ n2723;
  assign n39225 = n39224 ^ n2730;
  assign n39226 = n39161 ^ n39139;
  assign n3192 = n3191 ^ n2623;
  assign n3202 = n3201 ^ n3192;
  assign n3203 = n3202 ^ n2717;
  assign n39227 = n39226 ^ n3203;
  assign n39232 = n39159 ^ n39158;
  assign n39229 = n36982 ^ n3177;
  assign n39230 = n39229 ^ n33183;
  assign n39231 = n39230 ^ n27111;
  assign n39233 = n39232 ^ n39231;
  assign n39236 = n37027 ^ n28588;
  assign n39237 = n39236 ^ n1485;
  assign n39238 = n39237 ^ n3023;
  assign n39235 = n39155 ^ n39141;
  assign n39239 = n39238 ^ n39235;
  assign n39240 = n39154 ^ n39153;
  assign n1470 = n1427 ^ n1361;
  assign n1471 = n1470 ^ n1467;
  assign n1475 = n1474 ^ n1471;
  assign n39241 = n39240 ^ n1475;
  assign n39242 = n39152 ^ n39142;
  assign n1443 = n1346 ^ n1263;
  assign n1453 = n1452 ^ n1443;
  assign n1460 = n1459 ^ n1453;
  assign n39243 = n39242 ^ n1460;
  assign n39248 = n39148 ^ n39143;
  assign n39245 = n37010 ^ n1230;
  assign n39246 = n39245 ^ n33213;
  assign n39247 = n39246 ^ n1013;
  assign n39249 = n39248 ^ n39247;
  assign n39253 = n39147 ^ n39144;
  assign n39250 = n36999 ^ n3337;
  assign n39251 = n39250 ^ n878;
  assign n39252 = n39251 ^ n27130;
  assign n39254 = n39253 ^ n39252;
  assign n39258 = n39146 ^ n39145;
  assign n39255 = n36616 ^ n28673;
  assign n39256 = n39255 ^ n33220;
  assign n39257 = n39256 ^ n873;
  assign n39259 = n39258 ^ n39257;
  assign n38842 = n38841 ^ n38825;
  assign n762 = n761 ^ n740;
  assign n781 = n780 ^ n762;
  assign n788 = n787 ^ n781;
  assign n38843 = n38842 ^ n788;
  assign n38753 = n36607 ^ n28604;
  assign n38754 = n38753 ^ n33227;
  assign n38755 = n38754 ^ n774;
  assign n38752 = n38751 ^ n38738;
  assign n38756 = n38755 ^ n38752;
  assign n38758 = n38748 ^ n38747;
  assign n38762 = n38761 ^ n38758;
  assign n38764 = n36557 ^ n28616;
  assign n38765 = n38764 ^ n33242;
  assign n38766 = n38765 ^ n27174;
  assign n38763 = n38746 ^ n38745;
  assign n38767 = n38766 ^ n38763;
  assign n38771 = n38744 ^ n38743;
  assign n38768 = n36561 ^ n28648;
  assign n38769 = n38768 ^ n33247;
  assign n38770 = n38769 ^ n27167;
  assign n38772 = n38771 ^ n38770;
  assign n38776 = n38742 ^ n38741;
  assign n38773 = n36588 ^ n28621;
  assign n38774 = n38773 ^ n33251;
  assign n38775 = n38774 ^ n27158;
  assign n38777 = n38776 ^ n38775;
  assign n38779 = n36571 ^ n28625;
  assign n38780 = n38779 ^ n2231;
  assign n38781 = n38780 ^ n27147;
  assign n38782 = n38781 ^ n38739;
  assign n38785 = n36574 ^ n2222;
  assign n38786 = n38785 ^ n32500;
  assign n38787 = n38786 ^ n28628;
  assign n2046 = n2045 ^ n1979;
  assign n2059 = n2058 ^ n2046;
  assign n2066 = n2065 ^ n2059;
  assign n38783 = n38697 ^ n34889;
  assign n38784 = n2066 & ~n38783;
  assign n38788 = n38787 ^ n38784;
  assign n38789 = n38701 ^ n38699;
  assign n38790 = n38789 ^ n38787;
  assign n38791 = n38788 & n38790;
  assign n38792 = n38791 ^ n38784;
  assign n38793 = n38792 ^ n38781;
  assign n38794 = ~n38782 & ~n38793;
  assign n38795 = n38794 ^ n38739;
  assign n38778 = n38740 ^ n38739;
  assign n38796 = n38795 ^ n38778;
  assign n38797 = n33256 ^ n28639;
  assign n38798 = n38797 ^ n36567;
  assign n38799 = n38798 ^ n27142;
  assign n38800 = n38799 ^ n38778;
  assign n38801 = ~n38796 & ~n38800;
  assign n38802 = n38801 ^ n38799;
  assign n38803 = n38802 ^ n38776;
  assign n38804 = ~n38777 & n38803;
  assign n38805 = n38804 ^ n38775;
  assign n38806 = n38805 ^ n38771;
  assign n38807 = n38772 & ~n38806;
  assign n38808 = n38807 ^ n38770;
  assign n38809 = n38808 ^ n38763;
  assign n38810 = n38767 & ~n38809;
  assign n38811 = n38810 ^ n38766;
  assign n38812 = n38811 ^ n38758;
  assign n38813 = n38762 & ~n38812;
  assign n38814 = n38813 ^ n38761;
  assign n38757 = n38750 ^ n38749;
  assign n38815 = n38814 ^ n38757;
  assign n38816 = n36547 ^ n605;
  assign n38817 = n38816 ^ n33232;
  assign n38818 = n38817 ^ n3293;
  assign n38819 = n38818 ^ n38757;
  assign n38820 = ~n38815 & n38819;
  assign n38821 = n38820 ^ n38818;
  assign n38822 = n38821 ^ n38752;
  assign n38823 = n38756 & ~n38822;
  assign n38824 = n38823 ^ n38755;
  assign n39260 = n38842 ^ n38824;
  assign n39261 = ~n38843 & n39260;
  assign n39262 = n39261 ^ n788;
  assign n39263 = n39262 ^ n39257;
  assign n39264 = n39259 & ~n39263;
  assign n39265 = n39264 ^ n39258;
  assign n39266 = n39265 ^ n39253;
  assign n39267 = n39254 & ~n39266;
  assign n39268 = n39267 ^ n39252;
  assign n39269 = n39268 ^ n39248;
  assign n39270 = n39249 & ~n39269;
  assign n39271 = n39270 ^ n39247;
  assign n39244 = n39151 ^ n39149;
  assign n39272 = n39271 ^ n39244;
  assign n39273 = n3348 ^ n1245;
  assign n39274 = n39273 ^ n33208;
  assign n39275 = n39274 ^ n1450;
  assign n39276 = n39275 ^ n39244;
  assign n39277 = ~n39272 & n39276;
  assign n39278 = n39277 ^ n39275;
  assign n39279 = n39278 ^ n39242;
  assign n39280 = n39243 & ~n39279;
  assign n39281 = n39280 ^ n1460;
  assign n39282 = n39281 ^ n39240;
  assign n39283 = ~n39241 & n39282;
  assign n39284 = n39283 ^ n1475;
  assign n39285 = n39284 ^ n39235;
  assign n39286 = n39239 & ~n39285;
  assign n39287 = n39286 ^ n39238;
  assign n39234 = n39157 ^ n39156;
  assign n39288 = n39287 ^ n39234;
  assign n39289 = n36986 ^ n28583;
  assign n39290 = n39289 ^ n33190;
  assign n39291 = n39290 ^ n27116;
  assign n39292 = n39291 ^ n39234;
  assign n39293 = ~n39288 & n39292;
  assign n39294 = n39293 ^ n39291;
  assign n39295 = n39294 ^ n39232;
  assign n39296 = ~n39233 & n39295;
  assign n39297 = n39296 ^ n39231;
  assign n39228 = n39160 ^ n39140;
  assign n39298 = n39297 ^ n39228;
  assign n39299 = n36977 ^ n2614;
  assign n39300 = n39299 ^ n33178;
  assign n39301 = n39300 ^ n3199;
  assign n39302 = n39301 ^ n39228;
  assign n39303 = n39298 & ~n39302;
  assign n39304 = n39303 ^ n39301;
  assign n39305 = n39304 ^ n39226;
  assign n39306 = n39227 & ~n39305;
  assign n39307 = n39306 ^ n3203;
  assign n39308 = n39307 ^ n39224;
  assign n39309 = n39225 & ~n39308;
  assign n39310 = n39309 ^ n2730;
  assign n39311 = n39310 ^ n39222;
  assign n39312 = n39223 & ~n39311;
  assign n39313 = n39312 ^ n3117;
  assign n39314 = n39313 ^ n39220;
  assign n39315 = n39221 & ~n39314;
  assign n39316 = n39315 ^ n2828;
  assign n39168 = ~n39166 & n39167;
  assign n39117 = n39116 ^ n39042;
  assign n39118 = n39043 & n39117;
  assign n39119 = n39118 ^ n36265;
  assign n39004 = n37102 ^ n36435;
  assign n39005 = n38184 ^ n37102;
  assign n39006 = ~n39004 & n39005;
  assign n39007 = n39006 ^ n36435;
  assign n39002 = n38580 ^ n38530;
  assign n38878 = n38877 ^ n38873;
  assign n38999 = n38998 ^ n38873;
  assign n39000 = ~n38878 & n38999;
  assign n39001 = n39000 ^ n38877;
  assign n39003 = n39002 ^ n39001;
  assign n39040 = n39007 ^ n39003;
  assign n39120 = n39119 ^ n39040;
  assign n39138 = n39120 ^ n35680;
  assign n39219 = n39168 ^ n39138;
  assign n39317 = n39316 ^ n39219;
  assign n39321 = n39320 ^ n39219;
  assign n39322 = n39317 & ~n39321;
  assign n39323 = n39322 ^ n39320;
  assign n39121 = n39040 ^ n35680;
  assign n39122 = ~n39120 & ~n39121;
  assign n39123 = n39122 ^ n35680;
  assign n39008 = n39007 ^ n39002;
  assign n39009 = n39003 & ~n39008;
  assign n39010 = n39009 ^ n39007;
  assign n38871 = n38583 ^ n38528;
  assign n38867 = n37109 ^ n36428;
  assign n38868 = n38474 ^ n37109;
  assign n38869 = n38867 & ~n38868;
  assign n38870 = n38869 ^ n36428;
  assign n38872 = n38871 ^ n38870;
  assign n39038 = n39010 ^ n38872;
  assign n39039 = n39038 ^ n35673;
  assign n39170 = n39123 ^ n39039;
  assign n39169 = n39138 & n39168;
  assign n39214 = n39170 ^ n39169;
  assign n39218 = n39217 ^ n39214;
  assign n39899 = n39323 ^ n39218;
  assign n39181 = n38602 ^ n38510;
  assign n41150 = n39899 ^ n39181;
  assign n39556 = n39265 ^ n39254;
  assign n39552 = n38210 ^ n37322;
  assign n39553 = n38889 ^ n38210;
  assign n39554 = n39552 & ~n39553;
  assign n39555 = n39554 ^ n37322;
  assign n39557 = n39556 ^ n39555;
  assign n39562 = n39262 ^ n39259;
  assign n39558 = n38220 ^ n37328;
  assign n39559 = n38895 ^ n38220;
  assign n39560 = n39558 & ~n39559;
  assign n39561 = n39560 ^ n37328;
  assign n39563 = n39562 ^ n39561;
  assign n39564 = n38226 ^ n37472;
  assign n39565 = n38901 ^ n38226;
  assign n39566 = n39564 & n39565;
  assign n39567 = n39566 ^ n37472;
  assign n38844 = n38843 ^ n38824;
  assign n39568 = n39567 ^ n38844;
  assign n39569 = n38228 ^ n37334;
  assign n39570 = n38907 ^ n38228;
  assign n39571 = ~n39569 & n39570;
  assign n39572 = n39571 ^ n37334;
  assign n39454 = n38821 ^ n38756;
  assign n39573 = n39572 ^ n39454;
  assign n39574 = n38234 ^ n37340;
  assign n39575 = n38913 ^ n38234;
  assign n39576 = n39574 & ~n39575;
  assign n39577 = n39576 ^ n37340;
  assign n39461 = n38818 ^ n38815;
  assign n39578 = n39577 ^ n39461;
  assign n39579 = n38240 ^ n37342;
  assign n39580 = n38240 ^ n38163;
  assign n39581 = ~n39579 & n39580;
  assign n39582 = n39581 ^ n37342;
  assign n39468 = n38811 ^ n38762;
  assign n39583 = n39582 ^ n39468;
  assign n39584 = n38246 ^ n37352;
  assign n39585 = n38924 ^ n38246;
  assign n39586 = n39584 & ~n39585;
  assign n39587 = n39586 ^ n37352;
  assign n39475 = n38808 ^ n38767;
  assign n39588 = n39587 ^ n39475;
  assign n39589 = n38164 ^ n37358;
  assign n39590 = n38930 ^ n38164;
  assign n39591 = ~n39589 & ~n39590;
  assign n39592 = n39591 ^ n37358;
  assign n39483 = n38805 ^ n38772;
  assign n39593 = n39592 ^ n39483;
  assign n39598 = n38802 ^ n38777;
  assign n39594 = n38257 ^ n37364;
  assign n39595 = n38936 ^ n38257;
  assign n39596 = ~n39594 & ~n39595;
  assign n39597 = n39596 ^ n37364;
  assign n39599 = n39598 ^ n39597;
  assign n39604 = n38799 ^ n38796;
  assign n39600 = n38267 ^ n36636;
  assign n39601 = n38942 ^ n38267;
  assign n39602 = n39600 & n39601;
  assign n39603 = n39602 ^ n36636;
  assign n39605 = n39604 ^ n39603;
  assign n39607 = n38269 ^ n37259;
  assign n39608 = n38948 ^ n38269;
  assign n39609 = ~n39607 & n39608;
  assign n39610 = n39609 ^ n37259;
  assign n39606 = n38792 ^ n38782;
  assign n39611 = n39610 ^ n39606;
  assign n39613 = n38168 ^ n37266;
  assign n39614 = n38954 ^ n38168;
  assign n39615 = n39613 & n39614;
  assign n39616 = n39615 ^ n37266;
  assign n39612 = n38789 ^ n38788;
  assign n39617 = n39616 ^ n39612;
  assign n39437 = n38783 ^ n2066;
  assign n39433 = n38047 ^ n37273;
  assign n39434 = n38830 ^ n38047;
  assign n39435 = ~n39433 & ~n39434;
  assign n39436 = n39435 ^ n37273;
  assign n39438 = n39437 ^ n39436;
  assign n39341 = n37981 ^ n37280;
  assign n39342 = n38726 ^ n37981;
  assign n39343 = ~n39341 & n39342;
  assign n39344 = n39343 ^ n37280;
  assign n38865 = n38586 ^ n38526;
  assign n38861 = n37092 ^ n36418;
  assign n38862 = n37939 ^ n37092;
  assign n38863 = n38861 & n38862;
  assign n38864 = n38863 ^ n36418;
  assign n38866 = n38865 ^ n38864;
  assign n39011 = n39010 ^ n38871;
  assign n39012 = n38872 & n39011;
  assign n39013 = n39012 ^ n38870;
  assign n39014 = n39013 ^ n38865;
  assign n39015 = n38866 & n39014;
  assign n39016 = n39015 ^ n38864;
  assign n38855 = n37147 ^ n36415;
  assign n38856 = n37946 ^ n37147;
  assign n38857 = ~n38855 & n38856;
  assign n38858 = n38857 ^ n36415;
  assign n39033 = n39016 ^ n38858;
  assign n38859 = n38589 ^ n38521;
  assign n39034 = n39033 ^ n38859;
  assign n39035 = n39034 ^ n35660;
  assign n39036 = n39013 ^ n38866;
  assign n39037 = n39036 ^ n35667;
  assign n39124 = n39123 ^ n39038;
  assign n39125 = ~n39039 & ~n39124;
  assign n39126 = n39125 ^ n35673;
  assign n39127 = n39126 ^ n39036;
  assign n39128 = ~n39037 & ~n39127;
  assign n39129 = n39128 ^ n35667;
  assign n39130 = n39129 ^ n39034;
  assign n39131 = n39035 & ~n39130;
  assign n39132 = n39131 ^ n35660;
  assign n38860 = n38859 ^ n38858;
  assign n39017 = n39016 ^ n38859;
  assign n39018 = n38860 & n39017;
  assign n39019 = n39018 ^ n38858;
  assign n38850 = n37192 ^ n36405;
  assign n38851 = n37929 ^ n37192;
  assign n38852 = n38850 & n38851;
  assign n38853 = n38852 ^ n36405;
  assign n39030 = n39019 ^ n38853;
  assign n38849 = n38592 ^ n38516;
  assign n39031 = n39030 ^ n38849;
  assign n39032 = n39031 ^ n35654;
  assign n39137 = n39132 ^ n39032;
  assign n39171 = n39169 & ~n39170;
  assign n39172 = n39126 ^ n39037;
  assign n39173 = n39171 & n39172;
  assign n39174 = n39129 ^ n39035;
  assign n39175 = ~n39173 & ~n39174;
  assign n39176 = n39137 & n39175;
  assign n39133 = n39132 ^ n39031;
  assign n39134 = ~n39032 & n39133;
  assign n39135 = n39134 ^ n35654;
  assign n39024 = n37250 ^ n35946;
  assign n39025 = n37927 ^ n37250;
  assign n39026 = n39024 & n39025;
  assign n39027 = n39026 ^ n35946;
  assign n38854 = n38853 ^ n38849;
  assign n39020 = n39019 ^ n38849;
  assign n39021 = n38854 & n39020;
  assign n39022 = n39021 ^ n38853;
  assign n38848 = n38599 ^ n38596;
  assign n39023 = n39022 ^ n38848;
  assign n39028 = n39027 ^ n39023;
  assign n39029 = n39028 ^ n34898;
  assign n39136 = n39135 ^ n39029;
  assign n39197 = n39176 ^ n39136;
  assign n1906 = n1896 ^ n1860;
  assign n1925 = n1924 ^ n1906;
  assign n1932 = n1931 ^ n1925;
  assign n39198 = n39197 ^ n1932;
  assign n39200 = n37067 ^ n1801;
  assign n39201 = n39200 ^ n33139;
  assign n39202 = n39201 ^ n1921;
  assign n39199 = n39175 ^ n39137;
  assign n39203 = n39202 ^ n39199;
  assign n39205 = n36952 ^ n1786;
  assign n39206 = n39205 ^ n33144;
  assign n39207 = n39206 ^ n27433;
  assign n39204 = n39174 ^ n39173;
  assign n39208 = n39207 ^ n39204;
  assign n39209 = n39172 ^ n39171;
  assign n39213 = n39212 ^ n39209;
  assign n39324 = n39323 ^ n39214;
  assign n39325 = n39218 & ~n39324;
  assign n39326 = n39325 ^ n39217;
  assign n39327 = n39326 ^ n39209;
  assign n39328 = ~n39213 & n39327;
  assign n39329 = n39328 ^ n39212;
  assign n39330 = n39329 ^ n39204;
  assign n39331 = n39208 & ~n39330;
  assign n39332 = n39331 ^ n39207;
  assign n39333 = n39332 ^ n39199;
  assign n39334 = n39203 & ~n39333;
  assign n39335 = n39334 ^ n39202;
  assign n39336 = n39335 ^ n39197;
  assign n39337 = ~n39198 & n39336;
  assign n39338 = n39337 ^ n1932;
  assign n39194 = n37126 ^ n28885;
  assign n39195 = n39194 ^ n1939;
  assign n39196 = n39195 ^ n2053;
  assign n39339 = n39338 ^ n39196;
  assign n39188 = n39135 ^ n39028;
  assign n39189 = n39029 & ~n39188;
  assign n39190 = n39189 ^ n34898;
  assign n39191 = n39190 ^ n34891;
  assign n39183 = n37414 ^ n35940;
  assign n39184 = n37917 ^ n37414;
  assign n39185 = n39183 & n39184;
  assign n39186 = n39185 ^ n35940;
  assign n39178 = n39027 ^ n38848;
  assign n39179 = ~n39023 & n39178;
  assign n39180 = n39179 ^ n39027;
  assign n39182 = n39181 ^ n39180;
  assign n39187 = n39186 ^ n39182;
  assign n39192 = n39191 ^ n39187;
  assign n39177 = ~n39136 & n39176;
  assign n39193 = n39192 ^ n39177;
  assign n39340 = n39339 ^ n39193;
  assign n39345 = n39344 ^ n39340;
  assign n39347 = n37287 ^ n37256;
  assign n39348 = n38166 ^ n37256;
  assign n39349 = n39347 & n39348;
  assign n39350 = n39349 ^ n37287;
  assign n39346 = n39335 ^ n39198;
  assign n39351 = n39350 ^ n39346;
  assign n39353 = n37400 ^ n37263;
  assign n39354 = n38671 ^ n37263;
  assign n39355 = ~n39353 & ~n39354;
  assign n39356 = n39355 ^ n37400;
  assign n39352 = n39332 ^ n39203;
  assign n39357 = n39356 ^ n39352;
  assign n39364 = n37406 ^ n37270;
  assign n39365 = n38172 ^ n37270;
  assign n39366 = n39364 & ~n39365;
  assign n39367 = n39366 ^ n37406;
  assign n39358 = n39326 ^ n39213;
  assign n39359 = n37412 ^ n37277;
  assign n39360 = n38178 ^ n37277;
  assign n39361 = n39359 & ~n39360;
  assign n39362 = n39361 ^ n37412;
  assign n39363 = ~n39358 & ~n39362;
  assign n39368 = n39367 ^ n39363;
  assign n39369 = n39329 ^ n39208;
  assign n39370 = n39369 ^ n39367;
  assign n39371 = n39368 & ~n39370;
  assign n39372 = n39371 ^ n39363;
  assign n39373 = n39372 ^ n39352;
  assign n39374 = n39357 & ~n39373;
  assign n39375 = n39374 ^ n39356;
  assign n39376 = n39375 ^ n39346;
  assign n39377 = n39351 & n39376;
  assign n39378 = n39377 ^ n39350;
  assign n39439 = n39378 ^ n39340;
  assign n39440 = n39345 & n39439;
  assign n39441 = n39440 ^ n39344;
  assign n39618 = n39441 ^ n39437;
  assign n39619 = ~n39438 & n39618;
  assign n39620 = n39619 ^ n39436;
  assign n39621 = n39620 ^ n39612;
  assign n39622 = ~n39617 & n39621;
  assign n39623 = n39622 ^ n39616;
  assign n39624 = n39623 ^ n39606;
  assign n39625 = ~n39611 & n39624;
  assign n39626 = n39625 ^ n39610;
  assign n39627 = n39626 ^ n39604;
  assign n39628 = n39605 & ~n39627;
  assign n39629 = n39628 ^ n39603;
  assign n39630 = n39629 ^ n39598;
  assign n39631 = n39599 & n39630;
  assign n39632 = n39631 ^ n39597;
  assign n39633 = n39632 ^ n39483;
  assign n39634 = n39593 & n39633;
  assign n39635 = n39634 ^ n39592;
  assign n39636 = n39635 ^ n39475;
  assign n39637 = n39588 & ~n39636;
  assign n39638 = n39637 ^ n39587;
  assign n39639 = n39638 ^ n39468;
  assign n39640 = n39583 & ~n39639;
  assign n39641 = n39640 ^ n39582;
  assign n39642 = n39641 ^ n39461;
  assign n39643 = ~n39578 & ~n39642;
  assign n39644 = n39643 ^ n39577;
  assign n39645 = n39644 ^ n39454;
  assign n39646 = ~n39573 & n39645;
  assign n39647 = n39646 ^ n39572;
  assign n39648 = n39647 ^ n38844;
  assign n39649 = ~n39568 & ~n39648;
  assign n39650 = n39649 ^ n39567;
  assign n39651 = n39650 ^ n39562;
  assign n39652 = n39563 & ~n39651;
  assign n39653 = n39652 ^ n39561;
  assign n39654 = n39653 ^ n39556;
  assign n39655 = n39557 & ~n39654;
  assign n39656 = n39655 ^ n39555;
  assign n39550 = n39268 ^ n39249;
  assign n39546 = n38204 ^ n37316;
  assign n39547 = n38883 ^ n38204;
  assign n39548 = n39546 & ~n39547;
  assign n39549 = n39548 ^ n37316;
  assign n39551 = n39550 ^ n39549;
  assign n39738 = n39656 ^ n39551;
  assign n39739 = n39738 ^ n36645;
  assign n39740 = n39653 ^ n39557;
  assign n39741 = n39740 ^ n36648;
  assign n39742 = n39650 ^ n39563;
  assign n39743 = n39742 ^ n36654;
  assign n39744 = n39647 ^ n39568;
  assign n39745 = n39744 ^ n36664;
  assign n39746 = n39644 ^ n39573;
  assign n39747 = n39746 ^ n36670;
  assign n39748 = n39641 ^ n39578;
  assign n39749 = n39748 ^ n36673;
  assign n39750 = n39638 ^ n39582;
  assign n39751 = n39750 ^ n39468;
  assign n39752 = n39751 ^ n36679;
  assign n39753 = n39635 ^ n39588;
  assign n39754 = n39753 ^ n36686;
  assign n39755 = n39632 ^ n39593;
  assign n39756 = n39755 ^ n35927;
  assign n39757 = n39629 ^ n39599;
  assign n39758 = n39757 ^ n36702;
  assign n39759 = n39626 ^ n39603;
  assign n39760 = n39759 ^ n39604;
  assign n39761 = n39760 ^ n36708;
  assign n39762 = n39623 ^ n39611;
  assign n39763 = n39762 ^ n36715;
  assign n39764 = n39620 ^ n39616;
  assign n39765 = n39764 ^ n39612;
  assign n39766 = n39765 ^ n36717;
  assign n39442 = n39441 ^ n39438;
  assign n39443 = n39442 ^ n36724;
  assign n39379 = n39378 ^ n39345;
  assign n39380 = n39379 ^ n36730;
  assign n39381 = n39375 ^ n39350;
  assign n39382 = n39381 ^ n39346;
  assign n39383 = n39382 ^ n36623;
  assign n39384 = n39372 ^ n39357;
  assign n39385 = n39384 ^ n36515;
  assign n39386 = n39362 ^ n39358;
  assign n39387 = ~n35934 & n39386;
  assign n39388 = n39387 ^ n36464;
  assign n39389 = n39369 ^ n39368;
  assign n39390 = n39389 ^ n39387;
  assign n39391 = n39388 & ~n39390;
  assign n39392 = n39391 ^ n36464;
  assign n39393 = n39392 ^ n39384;
  assign n39394 = ~n39385 & ~n39393;
  assign n39395 = n39394 ^ n36515;
  assign n39396 = n39395 ^ n39382;
  assign n39397 = n39383 & n39396;
  assign n39398 = n39397 ^ n36623;
  assign n39444 = n39398 ^ n39379;
  assign n39445 = ~n39380 & n39444;
  assign n39446 = n39445 ^ n36730;
  assign n39767 = n39446 ^ n39442;
  assign n39768 = n39443 & n39767;
  assign n39769 = n39768 ^ n36724;
  assign n39770 = n39769 ^ n39765;
  assign n39771 = ~n39766 & ~n39770;
  assign n39772 = n39771 ^ n36717;
  assign n39773 = n39772 ^ n39762;
  assign n39774 = n39763 & n39773;
  assign n39775 = n39774 ^ n36715;
  assign n39776 = n39775 ^ n39760;
  assign n39777 = n39761 & n39776;
  assign n39778 = n39777 ^ n36708;
  assign n39779 = n39778 ^ n39757;
  assign n39780 = ~n39758 & ~n39779;
  assign n39781 = n39780 ^ n36702;
  assign n39782 = n39781 ^ n39755;
  assign n39783 = n39756 & ~n39782;
  assign n39784 = n39783 ^ n35927;
  assign n39785 = n39784 ^ n39753;
  assign n39786 = ~n39754 & n39785;
  assign n39787 = n39786 ^ n36686;
  assign n39788 = n39787 ^ n39751;
  assign n39789 = ~n39752 & n39788;
  assign n39790 = n39789 ^ n36679;
  assign n39791 = n39790 ^ n39748;
  assign n39792 = n39749 & ~n39791;
  assign n39793 = n39792 ^ n36673;
  assign n39794 = n39793 ^ n39746;
  assign n39795 = n39747 & n39794;
  assign n39796 = n39795 ^ n36670;
  assign n39797 = n39796 ^ n39744;
  assign n39798 = n39745 & ~n39797;
  assign n39799 = n39798 ^ n36664;
  assign n39800 = n39799 ^ n39742;
  assign n39801 = n39743 & ~n39800;
  assign n39802 = n39801 ^ n36654;
  assign n39803 = n39802 ^ n39740;
  assign n39804 = ~n39741 & ~n39803;
  assign n39805 = n39804 ^ n36648;
  assign n39806 = n39805 ^ n39738;
  assign n39807 = ~n39739 & n39806;
  assign n39808 = n39807 ^ n36645;
  assign n39657 = n39656 ^ n39550;
  assign n39658 = n39551 & ~n39657;
  assign n39659 = n39658 ^ n39549;
  assign n39544 = n39275 ^ n39272;
  assign n39540 = n38198 ^ n37310;
  assign n39541 = n38873 ^ n38198;
  assign n39542 = ~n39540 & ~n39541;
  assign n39543 = n39542 ^ n37310;
  assign n39545 = n39544 ^ n39543;
  assign n39736 = n39659 ^ n39545;
  assign n39737 = n39736 ^ n36790;
  assign n39847 = n39808 ^ n39737;
  assign n39848 = n39802 ^ n39741;
  assign n39849 = n39796 ^ n39745;
  assign n39850 = n39790 ^ n39749;
  assign n39851 = n39784 ^ n39754;
  assign n39852 = n39781 ^ n39756;
  assign n39853 = n39778 ^ n39758;
  assign n39854 = n39775 ^ n39761;
  assign n39855 = n39772 ^ n39763;
  assign n39447 = n39446 ^ n39443;
  assign n39399 = n39398 ^ n39380;
  assign n39400 = n39392 ^ n39385;
  assign n39401 = n39395 ^ n39383;
  assign n39402 = n39400 & n39401;
  assign n39448 = n39399 & n39402;
  assign n39856 = n39447 & ~n39448;
  assign n39857 = n39769 ^ n39766;
  assign n39858 = ~n39856 & ~n39857;
  assign n39859 = ~n39855 & n39858;
  assign n39860 = ~n39854 & ~n39859;
  assign n39861 = ~n39853 & n39860;
  assign n39862 = n39852 & ~n39861;
  assign n39863 = ~n39851 & n39862;
  assign n39864 = n39787 ^ n39752;
  assign n39865 = n39863 & ~n39864;
  assign n39866 = n39850 & n39865;
  assign n39867 = n39793 ^ n39747;
  assign n39868 = ~n39866 & ~n39867;
  assign n39869 = ~n39849 & ~n39868;
  assign n39870 = n39799 ^ n39743;
  assign n39871 = n39869 & ~n39870;
  assign n39872 = n39848 & n39871;
  assign n39873 = n39805 ^ n39739;
  assign n39874 = ~n39872 & n39873;
  assign n39875 = n39847 & ~n39874;
  assign n39809 = n39808 ^ n39736;
  assign n39810 = n39737 & ~n39809;
  assign n39811 = n39810 ^ n36790;
  assign n39660 = n39659 ^ n39544;
  assign n39661 = ~n39545 & ~n39660;
  assign n39662 = n39661 ^ n39543;
  assign n39538 = n39278 ^ n39243;
  assign n39534 = n38196 ^ n37304;
  assign n39535 = n39002 ^ n38196;
  assign n39536 = n39534 & ~n39535;
  assign n39537 = n39536 ^ n37304;
  assign n39539 = n39538 ^ n39537;
  assign n39734 = n39662 ^ n39539;
  assign n39735 = n39734 ^ n36887;
  assign n39876 = n39811 ^ n39735;
  assign n39877 = n39875 & ~n39876;
  assign n39812 = n39811 ^ n39734;
  assign n39813 = ~n39735 & ~n39812;
  assign n39814 = n39813 ^ n36887;
  assign n39668 = n38190 ^ n37298;
  assign n39669 = n38871 ^ n38190;
  assign n39670 = ~n39668 & n39669;
  assign n39671 = n39670 ^ n37298;
  assign n39666 = n39281 ^ n39241;
  assign n39663 = n39662 ^ n39538;
  assign n39664 = n39539 & n39663;
  assign n39665 = n39664 ^ n39537;
  assign n39667 = n39666 ^ n39665;
  assign n39732 = n39671 ^ n39667;
  assign n39733 = n39732 ^ n36945;
  assign n39878 = n39814 ^ n39733;
  assign n39879 = ~n39877 & n39878;
  assign n39815 = n39814 ^ n39732;
  assign n39816 = n39733 & n39815;
  assign n39817 = n39816 ^ n36945;
  assign n39845 = n39817 ^ n37086;
  assign n39677 = n38185 ^ n37499;
  assign n39678 = n38865 ^ n38185;
  assign n39679 = n39677 & n39678;
  assign n39680 = n39679 ^ n37499;
  assign n39675 = n39284 ^ n39239;
  assign n39672 = n39671 ^ n39666;
  assign n39673 = n39667 & ~n39672;
  assign n39674 = n39673 ^ n39671;
  assign n39676 = n39675 ^ n39674;
  assign n39730 = n39680 ^ n39676;
  assign n39846 = n39845 ^ n39730;
  assign n39937 = n39879 ^ n39846;
  assign n39941 = n39940 ^ n39937;
  assign n39945 = n39878 ^ n39877;
  assign n39942 = n37770 ^ n3211;
  assign n39943 = n39942 ^ n34007;
  assign n39944 = n39943 ^ n3077;
  assign n39946 = n39945 ^ n39944;
  assign n39951 = n39874 ^ n39847;
  assign n39948 = n37780 ^ n29410;
  assign n39949 = n39948 ^ n2492;
  assign n39950 = n39949 ^ n3053;
  assign n39952 = n39951 ^ n39950;
  assign n39957 = n39871 ^ n39848;
  assign n39954 = n37790 ^ n2429;
  assign n39955 = n39954 ^ n34023;
  assign n39956 = n39955 ^ n3146;
  assign n39958 = n39957 ^ n39956;
  assign n39960 = n37796 ^ n29418;
  assign n39961 = n39960 ^ n1301;
  assign n39962 = n39961 ^ n27724;
  assign n39959 = n39870 ^ n39869;
  assign n39963 = n39962 ^ n39959;
  assign n39965 = n37863 ^ n29424;
  assign n39966 = n39965 ^ n33961;
  assign n39967 = n39966 ^ n1293;
  assign n39964 = n39868 ^ n39849;
  assign n39968 = n39967 ^ n39964;
  assign n39969 = n39867 ^ n39866;
  assign n1101 = n1100 ^ n1034;
  assign n1117 = n1116 ^ n1101;
  assign n1124 = n1123 ^ n1117;
  assign n39970 = n39969 ^ n1124;
  assign n39974 = n39865 ^ n39850;
  assign n39971 = n37853 ^ n29095;
  assign n39972 = n39971 ^ n994;
  assign n39973 = n39972 ^ n1107;
  assign n39975 = n39974 ^ n39973;
  assign n39977 = n39862 ^ n39851;
  assign n39981 = n39980 ^ n39977;
  assign n39983 = n37808 ^ n832;
  assign n39984 = n39983 ^ n33539;
  assign n39985 = n39984 ^ n3312;
  assign n39982 = n39861 ^ n39852;
  assign n39986 = n39985 ^ n39982;
  assign n39987 = n39860 ^ n39853;
  assign n39991 = n39990 ^ n39987;
  assign n39993 = n37814 ^ n29021;
  assign n39994 = n39993 ^ n33469;
  assign n39995 = n39994 ^ n27742;
  assign n39992 = n39859 ^ n39854;
  assign n39996 = n39995 ^ n39992;
  assign n40000 = n39858 ^ n39855;
  assign n39997 = n37818 ^ n29026;
  assign n39998 = n39997 ^ n33473;
  assign n39999 = n39998 ^ n27747;
  assign n40001 = n40000 ^ n39999;
  assign n40005 = n39857 ^ n39856;
  assign n40002 = n37236 ^ n29031;
  assign n40003 = n40002 ^ n33478;
  assign n40004 = n40003 ^ n708;
  assign n40006 = n40005 ^ n40004;
  assign n39449 = n39448 ^ n39447;
  assign n39430 = n37207 ^ n29035;
  assign n39431 = n39430 ^ n33483;
  assign n39432 = n39431 ^ n27753;
  assign n39450 = n39449 ^ n39432;
  assign n39404 = n37212 ^ n29039;
  assign n39405 = n39404 ^ n33489;
  assign n39406 = n39405 ^ n27759;
  assign n39403 = n39402 ^ n39399;
  assign n39407 = n39406 ^ n39403;
  assign n2335 = n2324 ^ n2247;
  assign n2345 = n2344 ^ n2335;
  assign n2352 = n2351 ^ n2345;
  assign n39409 = n39400 ^ n2352;
  assign n2183 = n2143 ^ n2092;
  assign n2184 = n2183 ^ n2182;
  assign n2185 = n2184 ^ n2170;
  assign n39410 = n39386 ^ n35934;
  assign n39411 = n2185 & ~n39410;
  assign n2195 = n2192 ^ n2158;
  assign n2196 = n2195 ^ n2110;
  assign n2203 = n2202 ^ n2196;
  assign n39412 = n39411 ^ n2203;
  assign n39413 = n39389 ^ n39388;
  assign n39414 = n39413 ^ n2203;
  assign n39415 = n39412 & ~n39414;
  assign n39416 = n39415 ^ n39411;
  assign n39417 = n39416 ^ n39400;
  assign n39418 = n39409 & ~n39417;
  assign n39419 = n39418 ^ n2352;
  assign n39408 = n39401 ^ n39400;
  assign n39420 = n39419 ^ n39408;
  assign n39421 = n37216 ^ n28809;
  assign n39422 = n39421 ^ n2362;
  assign n39423 = n39422 ^ n27763;
  assign n39424 = n39423 ^ n39408;
  assign n39425 = n39420 & ~n39424;
  assign n39426 = n39425 ^ n39423;
  assign n39427 = n39426 ^ n39403;
  assign n39428 = ~n39407 & n39427;
  assign n39429 = n39428 ^ n39406;
  assign n40007 = n39449 ^ n39429;
  assign n40008 = ~n39450 & n40007;
  assign n40009 = n40008 ^ n39432;
  assign n40010 = n40009 ^ n40005;
  assign n40011 = ~n40006 & n40010;
  assign n40012 = n40011 ^ n40004;
  assign n40013 = n40012 ^ n40000;
  assign n40014 = n40001 & ~n40013;
  assign n40015 = n40014 ^ n39999;
  assign n40016 = n40015 ^ n39992;
  assign n40017 = n39996 & ~n40016;
  assign n40018 = n40017 ^ n39995;
  assign n40019 = n40018 ^ n39987;
  assign n40020 = ~n39991 & n40019;
  assign n40021 = n40020 ^ n39990;
  assign n40022 = n40021 ^ n39982;
  assign n40023 = n39986 & ~n40022;
  assign n40024 = n40023 ^ n39985;
  assign n40025 = n40024 ^ n39977;
  assign n40026 = n39981 & ~n40025;
  assign n40027 = n40026 ^ n39980;
  assign n39976 = n39864 ^ n39863;
  assign n40028 = n40027 ^ n39976;
  assign n952 = n942 ^ n906;
  assign n977 = n976 ^ n952;
  assign n984 = n983 ^ n977;
  assign n40029 = n39976 ^ n984;
  assign n40030 = ~n40028 & n40029;
  assign n40031 = n40030 ^ n984;
  assign n40032 = n40031 ^ n39974;
  assign n40033 = ~n39975 & n40032;
  assign n40034 = n40033 ^ n39973;
  assign n40035 = n40034 ^ n39969;
  assign n40036 = n39970 & ~n40035;
  assign n40037 = n40036 ^ n1124;
  assign n40038 = n40037 ^ n39964;
  assign n40039 = ~n39968 & n40038;
  assign n40040 = n40039 ^ n39967;
  assign n40041 = n40040 ^ n39959;
  assign n40042 = n39963 & ~n40041;
  assign n40043 = n40042 ^ n39962;
  assign n40044 = n40043 ^ n39957;
  assign n40045 = ~n39958 & n40044;
  assign n40046 = n40045 ^ n39956;
  assign n39953 = n39873 ^ n39872;
  assign n40047 = n40046 ^ n39953;
  assign n40048 = n37785 ^ n3035;
  assign n40049 = n40048 ^ n34018;
  assign n40050 = n40049 ^ n2484;
  assign n40051 = n40050 ^ n39953;
  assign n40052 = n40047 & ~n40051;
  assign n40053 = n40052 ^ n40050;
  assign n40054 = n40053 ^ n39951;
  assign n40055 = n39952 & ~n40054;
  assign n40056 = n40055 ^ n39950;
  assign n39947 = n39876 ^ n39875;
  assign n40057 = n40056 ^ n39947;
  assign n40058 = n37775 ^ n29405;
  assign n40059 = n40058 ^ n3059;
  assign n40060 = n40059 ^ n2546;
  assign n40061 = n40060 ^ n39947;
  assign n40062 = ~n40057 & n40061;
  assign n40063 = n40062 ^ n40060;
  assign n40064 = n40063 ^ n39945;
  assign n40065 = ~n39946 & n40064;
  assign n40066 = n40065 ^ n39944;
  assign n40067 = n40066 ^ n39937;
  assign n40068 = ~n39941 & n40067;
  assign n40069 = n40068 ^ n39940;
  assign n39731 = n39730 ^ n37086;
  assign n39818 = n39817 ^ n39730;
  assign n39819 = n39731 & n39818;
  assign n39820 = n39819 ^ n37086;
  assign n39881 = n39820 ^ n37132;
  assign n39681 = n39680 ^ n39675;
  assign n39682 = ~n39676 & n39681;
  assign n39683 = n39682 ^ n39680;
  assign n39529 = n38184 ^ n37293;
  assign n39530 = n38859 ^ n38184;
  assign n39531 = ~n39529 & n39530;
  assign n39532 = n39531 ^ n37293;
  assign n39727 = n39683 ^ n39532;
  assign n39528 = n39291 ^ n39288;
  assign n39728 = n39727 ^ n39528;
  assign n39882 = n39881 ^ n39728;
  assign n39880 = ~n39846 & n39879;
  assign n39936 = n39882 ^ n39880;
  assign n40070 = n40069 ^ n39936;
  assign n3229 = n3225 ^ n2795;
  assign n3236 = n3235 ^ n3229;
  assign n3237 = n3236 ^ n2911;
  assign n40071 = n39936 ^ n3237;
  assign n40072 = n40070 & ~n40071;
  assign n40073 = n40072 ^ n3237;
  assign n39729 = n39728 ^ n37132;
  assign n39821 = n39820 ^ n39728;
  assign n39822 = ~n39729 & ~n39821;
  assign n39823 = n39822 ^ n37132;
  assign n39533 = n39532 ^ n39528;
  assign n39684 = n39683 ^ n39528;
  assign n39685 = n39533 & ~n39684;
  assign n39686 = n39685 ^ n39532;
  assign n39523 = n38474 ^ n37714;
  assign n39524 = n38849 ^ n38474;
  assign n39525 = ~n39523 & n39524;
  assign n39526 = n39525 ^ n37714;
  assign n39724 = n39686 ^ n39526;
  assign n39522 = n39294 ^ n39233;
  assign n39725 = n39724 ^ n39522;
  assign n39726 = n39725 ^ n37179;
  assign n39884 = n39823 ^ n39726;
  assign n39883 = n39880 & ~n39882;
  assign n39934 = n39884 ^ n39883;
  assign n2896 = n2890 ^ n2854;
  assign n2915 = n2914 ^ n2896;
  assign n2922 = n2921 ^ n2915;
  assign n39935 = n39934 ^ n2922;
  assign n40456 = n40073 ^ n39935;
  assign n41151 = n40456 ^ n39899;
  assign n41152 = ~n41150 & n41151;
  assign n41153 = n41152 ^ n39181;
  assign n40755 = n38540 ^ n3155;
  assign n40756 = n40755 ^ n34746;
  assign n40757 = n40756 ^ n28583;
  assign n40534 = n38883 ^ n38220;
  assign n40535 = n39666 ^ n38883;
  assign n40536 = n40534 & n40535;
  assign n40537 = n40536 ^ n38220;
  assign n40533 = n40024 ^ n39981;
  assign n40538 = n40537 ^ n40533;
  assign n40412 = n38889 ^ n38226;
  assign n40413 = n39538 ^ n38889;
  assign n40414 = n40412 & ~n40413;
  assign n40415 = n40414 ^ n38226;
  assign n40411 = n40021 ^ n39986;
  assign n40416 = n40415 ^ n40411;
  assign n40287 = n38895 ^ n38228;
  assign n40288 = n39544 ^ n38895;
  assign n40289 = n40287 & ~n40288;
  assign n40290 = n40289 ^ n38228;
  assign n40286 = n40018 ^ n39991;
  assign n40291 = n40290 ^ n40286;
  assign n40249 = n38901 ^ n38234;
  assign n40250 = n39550 ^ n38901;
  assign n40251 = n40249 & n40250;
  assign n40252 = n40251 ^ n38234;
  assign n40248 = n40015 ^ n39996;
  assign n40253 = n40252 ^ n40248;
  assign n40239 = n40012 ^ n40001;
  assign n40235 = n38907 ^ n38240;
  assign n40236 = n39556 ^ n38907;
  assign n40237 = n40235 & n40236;
  assign n40238 = n40237 ^ n38240;
  assign n40240 = n40239 ^ n40238;
  assign n40168 = n40009 ^ n40006;
  assign n40164 = n38913 ^ n38246;
  assign n40165 = n39562 ^ n38913;
  assign n40166 = ~n40164 & n40165;
  assign n40167 = n40166 ^ n38246;
  assign n40169 = n40168 ^ n40167;
  assign n39451 = n39450 ^ n39429;
  assign n38165 = n38164 ^ n38163;
  assign n38845 = n38844 ^ n38163;
  assign n38846 = ~n38165 & n38845;
  assign n38847 = n38846 ^ n38164;
  assign n39452 = n39451 ^ n38847;
  assign n39458 = n39426 ^ n39407;
  assign n39453 = n38924 ^ n38257;
  assign n39455 = n39454 ^ n38924;
  assign n39456 = n39453 & ~n39455;
  assign n39457 = n39456 ^ n38257;
  assign n39459 = n39458 ^ n39457;
  assign n39465 = n39423 ^ n39420;
  assign n39460 = n38930 ^ n38267;
  assign n39462 = n39461 ^ n38930;
  assign n39463 = ~n39460 & n39462;
  assign n39464 = n39463 ^ n38267;
  assign n39466 = n39465 ^ n39464;
  assign n39472 = n39416 ^ n39409;
  assign n39467 = n38936 ^ n38269;
  assign n39469 = n39468 ^ n38936;
  assign n39470 = ~n39467 & ~n39469;
  assign n39471 = n39470 ^ n38269;
  assign n39473 = n39472 ^ n39471;
  assign n39479 = n39413 ^ n39412;
  assign n39474 = n38942 ^ n38168;
  assign n39476 = n39475 ^ n38942;
  assign n39477 = ~n39474 & n39476;
  assign n39478 = n39477 ^ n38168;
  assign n39480 = n39479 ^ n39478;
  assign n39482 = n38948 ^ n38047;
  assign n39484 = n39483 ^ n38948;
  assign n39485 = ~n39482 & ~n39484;
  assign n39486 = n39485 ^ n38047;
  assign n39481 = n39410 ^ n2185;
  assign n39487 = n39486 ^ n39481;
  assign n40105 = n38954 ^ n37981;
  assign n40106 = n39598 ^ n38954;
  assign n40107 = n40105 & ~n40106;
  assign n40108 = n40107 ^ n37981;
  assign n39511 = n37946 ^ n37109;
  assign n39512 = n39181 ^ n37946;
  assign n39513 = n39511 & n39512;
  assign n39514 = n39513 ^ n37109;
  assign n39510 = n39304 ^ n39227;
  assign n39515 = n39514 ^ n39510;
  assign n39517 = n37939 ^ n37102;
  assign n39518 = n38848 ^ n37939;
  assign n39519 = n39517 & n39518;
  assign n39520 = n39519 ^ n37102;
  assign n39516 = n39301 ^ n39298;
  assign n39521 = n39520 ^ n39516;
  assign n39527 = n39526 ^ n39522;
  assign n39687 = n39686 ^ n39522;
  assign n39688 = n39527 & n39687;
  assign n39689 = n39688 ^ n39526;
  assign n39690 = n39689 ^ n39516;
  assign n39691 = ~n39521 & ~n39690;
  assign n39692 = n39691 ^ n39520;
  assign n39693 = n39692 ^ n39510;
  assign n39694 = n39515 & ~n39693;
  assign n39695 = n39694 ^ n39514;
  assign n39505 = n37929 ^ n37092;
  assign n39506 = n38647 ^ n37929;
  assign n39507 = ~n39505 & ~n39506;
  assign n39508 = n39507 ^ n37092;
  assign n39715 = n39695 ^ n39508;
  assign n39504 = n39307 ^ n39225;
  assign n39716 = n39715 ^ n39504;
  assign n39717 = n39716 ^ n36418;
  assign n39718 = n39692 ^ n39514;
  assign n39719 = n39718 ^ n39510;
  assign n39720 = n39719 ^ n36428;
  assign n39721 = n39689 ^ n39520;
  assign n39722 = n39721 ^ n39516;
  assign n39723 = n39722 ^ n36435;
  assign n39824 = n39823 ^ n39725;
  assign n39825 = ~n39726 & n39824;
  assign n39826 = n39825 ^ n37179;
  assign n39827 = n39826 ^ n39722;
  assign n39828 = ~n39723 & n39827;
  assign n39829 = n39828 ^ n36435;
  assign n39830 = n39829 ^ n39719;
  assign n39831 = n39720 & n39830;
  assign n39832 = n39831 ^ n36428;
  assign n39833 = n39832 ^ n39716;
  assign n39834 = n39717 & n39833;
  assign n39835 = n39834 ^ n36418;
  assign n39509 = n39508 ^ n39504;
  assign n39696 = n39695 ^ n39504;
  assign n39697 = ~n39509 & ~n39696;
  assign n39698 = n39697 ^ n39508;
  assign n39499 = n37927 ^ n37147;
  assign n39500 = n38641 ^ n37927;
  assign n39501 = ~n39499 & n39500;
  assign n39502 = n39501 ^ n37147;
  assign n39712 = n39698 ^ n39502;
  assign n39498 = n39310 ^ n39223;
  assign n39713 = n39712 ^ n39498;
  assign n39714 = n39713 ^ n36415;
  assign n39843 = n39835 ^ n39714;
  assign n39844 = n39829 ^ n39720;
  assign n39885 = ~n39883 & ~n39884;
  assign n39886 = n39826 ^ n39723;
  assign n39887 = n39885 & ~n39886;
  assign n39888 = n39844 & n39887;
  assign n39889 = n39832 ^ n39717;
  assign n39890 = n39888 & ~n39889;
  assign n39891 = ~n39843 & ~n39890;
  assign n39836 = n39835 ^ n39713;
  assign n39837 = n39714 & n39836;
  assign n39838 = n39837 ^ n36415;
  assign n39503 = n39502 ^ n39498;
  assign n39699 = n39698 ^ n39498;
  assign n39700 = ~n39503 & n39699;
  assign n39701 = n39700 ^ n39502;
  assign n39493 = n37917 ^ n37192;
  assign n39494 = n38635 ^ n37917;
  assign n39495 = n39493 & ~n39494;
  assign n39496 = n39495 ^ n37192;
  assign n39709 = n39701 ^ n39496;
  assign n39492 = n39313 ^ n39221;
  assign n39710 = n39709 ^ n39492;
  assign n39711 = n39710 ^ n36405;
  assign n39892 = n39838 ^ n39711;
  assign n39893 = n39891 & ~n39892;
  assign n39839 = n39838 ^ n39710;
  assign n39840 = ~n39711 & ~n39839;
  assign n39841 = n39840 ^ n36405;
  assign n39706 = n39320 ^ n39317;
  assign n39497 = n39496 ^ n39492;
  assign n39702 = n39701 ^ n39492;
  assign n39703 = ~n39497 & n39702;
  assign n39704 = n39703 ^ n39496;
  assign n39488 = n37291 ^ n37250;
  assign n39489 = n38629 ^ n37291;
  assign n39490 = n39488 & ~n39489;
  assign n39491 = n39490 ^ n37250;
  assign n39705 = n39704 ^ n39491;
  assign n39707 = n39706 ^ n39705;
  assign n39708 = n39707 ^ n35946;
  assign n39842 = n39841 ^ n39708;
  assign n39912 = n39893 ^ n39842;
  assign n39916 = n39915 ^ n39912;
  assign n39918 = n37744 ^ n29376;
  assign n39919 = n39918 ^ n33940;
  assign n39920 = n39919 ^ n28155;
  assign n39917 = n39892 ^ n39891;
  assign n39921 = n39920 ^ n39917;
  assign n39923 = n37749 ^ n29381;
  assign n39924 = n39923 ^ n33944;
  assign n39925 = n39924 ^ n1731;
  assign n39922 = n39890 ^ n39843;
  assign n39926 = n39925 ^ n39922;
  assign n39931 = n39887 ^ n39844;
  assign n39928 = n29391 ^ n2964;
  assign n39929 = n39928 ^ n33951;
  assign n39930 = n39929 ^ n1647;
  assign n39932 = n39931 ^ n39930;
  assign n40074 = n40073 ^ n39934;
  assign n40075 = ~n39935 & n40074;
  assign n40076 = n40075 ^ n2922;
  assign n39933 = n39886 ^ n39885;
  assign n40077 = n40076 ^ n39933;
  assign n2933 = n2869 ^ n1601;
  assign n2934 = n2933 ^ n2930;
  assign n2938 = n2937 ^ n2934;
  assign n40078 = n39933 ^ n2938;
  assign n40079 = ~n40077 & n40078;
  assign n40080 = n40079 ^ n2938;
  assign n40081 = n40080 ^ n39931;
  assign n40082 = ~n39932 & n40081;
  assign n40083 = n40082 ^ n39930;
  assign n39927 = n39889 ^ n39888;
  assign n40084 = n40083 ^ n39927;
  assign n40085 = n37754 ^ n29386;
  assign n40086 = n40085 ^ n1655;
  assign n40087 = n40086 ^ n28161;
  assign n40088 = n40087 ^ n39927;
  assign n40089 = ~n40084 & n40088;
  assign n40090 = n40089 ^ n40087;
  assign n40091 = n40090 ^ n39922;
  assign n40092 = n39926 & ~n40091;
  assign n40093 = n40092 ^ n39925;
  assign n40094 = n40093 ^ n39917;
  assign n40095 = ~n39921 & n40094;
  assign n40096 = n40095 ^ n39920;
  assign n40097 = n40096 ^ n39912;
  assign n40098 = ~n39916 & n40097;
  assign n40099 = n40098 ^ n39915;
  assign n40103 = n40102 ^ n40099;
  assign n39907 = n39841 ^ n39707;
  assign n39908 = n39708 & ~n39907;
  assign n39909 = n39908 ^ n35946;
  assign n39901 = n39706 ^ n39491;
  assign n39902 = n39706 ^ n39704;
  assign n39903 = n39901 & ~n39902;
  assign n39904 = n39903 ^ n39491;
  assign n39895 = n37414 ^ n37284;
  assign n39896 = n38623 ^ n37284;
  assign n39897 = n39895 & ~n39896;
  assign n39898 = n39897 ^ n37414;
  assign n39900 = n39899 ^ n39898;
  assign n39905 = n39904 ^ n39900;
  assign n39906 = n39905 ^ n35940;
  assign n39910 = n39909 ^ n39906;
  assign n39894 = ~n39842 & n39893;
  assign n39911 = n39910 ^ n39894;
  assign n40104 = n40103 ^ n39911;
  assign n40109 = n40108 ^ n40104;
  assign n40114 = n40096 ^ n39916;
  assign n40110 = n38830 ^ n37256;
  assign n40111 = n39604 ^ n38830;
  assign n40112 = n40110 & n40111;
  assign n40113 = n40112 ^ n37256;
  assign n40115 = n40114 ^ n40113;
  assign n40117 = n38726 ^ n37263;
  assign n40118 = n39606 ^ n38726;
  assign n40119 = ~n40117 & n40118;
  assign n40120 = n40119 ^ n37263;
  assign n40116 = n40093 ^ n39921;
  assign n40121 = n40120 ^ n40116;
  assign n40123 = n38166 ^ n37270;
  assign n40124 = n39612 ^ n38166;
  assign n40125 = n40123 & n40124;
  assign n40126 = n40125 ^ n37270;
  assign n40122 = n40090 ^ n39926;
  assign n40127 = n40126 ^ n40122;
  assign n40128 = n40087 ^ n40084;
  assign n40129 = n38671 ^ n37277;
  assign n40130 = n39437 ^ n38671;
  assign n40131 = n40129 & ~n40130;
  assign n40132 = n40131 ^ n37277;
  assign n40133 = n40128 & ~n40132;
  assign n40134 = n40133 ^ n40122;
  assign n40135 = ~n40127 & n40134;
  assign n40136 = n40135 ^ n40133;
  assign n40137 = n40136 ^ n40116;
  assign n40138 = n40121 & n40137;
  assign n40139 = n40138 ^ n40120;
  assign n40140 = n40139 ^ n40114;
  assign n40141 = n40115 & ~n40140;
  assign n40142 = n40141 ^ n40113;
  assign n40143 = n40142 ^ n40104;
  assign n40144 = n40109 & ~n40143;
  assign n40145 = n40144 ^ n40108;
  assign n40146 = n40145 ^ n39481;
  assign n40147 = n39487 & ~n40146;
  assign n40148 = n40147 ^ n39486;
  assign n40149 = n40148 ^ n39479;
  assign n40150 = n39480 & n40149;
  assign n40151 = n40150 ^ n39478;
  assign n40152 = n40151 ^ n39472;
  assign n40153 = ~n39473 & ~n40152;
  assign n40154 = n40153 ^ n39471;
  assign n40155 = n40154 ^ n39465;
  assign n40156 = ~n39466 & ~n40155;
  assign n40157 = n40156 ^ n39464;
  assign n40158 = n40157 ^ n39458;
  assign n40159 = ~n39459 & n40158;
  assign n40160 = n40159 ^ n39457;
  assign n40161 = n40160 ^ n39451;
  assign n40162 = n39452 & n40161;
  assign n40163 = n40162 ^ n38847;
  assign n40232 = n40168 ^ n40163;
  assign n40233 = ~n40169 & ~n40232;
  assign n40234 = n40233 ^ n40167;
  assign n40245 = n40239 ^ n40234;
  assign n40246 = ~n40240 & ~n40245;
  assign n40247 = n40246 ^ n40238;
  assign n40283 = n40248 ^ n40247;
  assign n40284 = ~n40253 & n40283;
  assign n40285 = n40284 ^ n40252;
  assign n40408 = n40286 ^ n40285;
  assign n40409 = ~n40291 & ~n40408;
  assign n40410 = n40409 ^ n40290;
  assign n40539 = n40411 ^ n40410;
  assign n40540 = n40416 & ~n40539;
  assign n40541 = n40540 ^ n40415;
  assign n40542 = n40541 ^ n40533;
  assign n40543 = n40538 & ~n40542;
  assign n40544 = n40543 ^ n40537;
  assign n40528 = n38873 ^ n38210;
  assign n40529 = n39675 ^ n38873;
  assign n40530 = n40528 & ~n40529;
  assign n40531 = n40530 ^ n38210;
  assign n40527 = n40028 ^ n984;
  assign n40532 = n40531 ^ n40527;
  assign n40619 = n40544 ^ n40532;
  assign n40620 = n40619 ^ n37322;
  assign n40621 = n40541 ^ n40538;
  assign n40622 = n40621 ^ n37328;
  assign n40417 = n40416 ^ n40410;
  assign n40418 = n40417 ^ n37472;
  assign n40292 = n40291 ^ n40285;
  assign n40293 = n40292 ^ n37334;
  assign n40254 = n40253 ^ n40247;
  assign n40255 = n40254 ^ n37340;
  assign n40170 = n40169 ^ n40163;
  assign n40171 = n40170 ^ n37352;
  assign n40172 = n40160 ^ n39452;
  assign n40173 = n40172 ^ n37358;
  assign n40174 = n40157 ^ n39459;
  assign n40175 = n40174 ^ n37364;
  assign n40176 = n40154 ^ n39464;
  assign n40177 = n40176 ^ n39465;
  assign n40178 = n40177 ^ n36636;
  assign n40179 = n40151 ^ n39473;
  assign n40180 = n40179 ^ n37259;
  assign n40181 = n40148 ^ n39478;
  assign n40182 = n40181 ^ n39479;
  assign n40183 = n40182 ^ n37266;
  assign n40184 = n40145 ^ n39487;
  assign n40185 = n40184 ^ n37273;
  assign n40186 = n40142 ^ n40109;
  assign n40187 = n40186 ^ n37280;
  assign n40188 = n40139 ^ n40113;
  assign n40189 = n40188 ^ n40114;
  assign n40190 = n40189 ^ n37287;
  assign n40191 = n40136 ^ n40121;
  assign n40192 = n40191 ^ n37400;
  assign n40193 = n40132 ^ n40128;
  assign n40194 = ~n37412 & ~n40193;
  assign n40195 = n40194 ^ n37406;
  assign n40196 = n40133 ^ n40126;
  assign n40197 = n40196 ^ n40122;
  assign n40198 = n40197 ^ n40194;
  assign n40199 = n40195 & ~n40198;
  assign n40200 = n40199 ^ n37406;
  assign n40201 = n40200 ^ n40191;
  assign n40202 = n40192 & ~n40201;
  assign n40203 = n40202 ^ n37400;
  assign n40204 = n40203 ^ n40189;
  assign n40205 = n40190 & n40204;
  assign n40206 = n40205 ^ n37287;
  assign n40207 = n40206 ^ n40186;
  assign n40208 = ~n40187 & ~n40207;
  assign n40209 = n40208 ^ n37280;
  assign n40210 = n40209 ^ n40184;
  assign n40211 = ~n40185 & n40210;
  assign n40212 = n40211 ^ n37273;
  assign n40213 = n40212 ^ n40182;
  assign n40214 = ~n40183 & n40213;
  assign n40215 = n40214 ^ n37266;
  assign n40216 = n40215 ^ n40179;
  assign n40217 = ~n40180 & n40216;
  assign n40218 = n40217 ^ n37259;
  assign n40219 = n40218 ^ n40177;
  assign n40220 = n40178 & ~n40219;
  assign n40221 = n40220 ^ n36636;
  assign n40222 = n40221 ^ n40174;
  assign n40223 = n40175 & n40222;
  assign n40224 = n40223 ^ n37364;
  assign n40225 = n40224 ^ n40172;
  assign n40226 = n40173 & n40225;
  assign n40227 = n40226 ^ n37358;
  assign n40228 = n40227 ^ n40170;
  assign n40229 = n40171 & ~n40228;
  assign n40230 = n40229 ^ n37352;
  assign n40231 = n40230 ^ n37342;
  assign n40241 = n40240 ^ n40234;
  assign n40242 = n40241 ^ n40230;
  assign n40243 = n40231 & n40242;
  assign n40244 = n40243 ^ n37342;
  assign n40280 = n40254 ^ n40244;
  assign n40281 = ~n40255 & ~n40280;
  assign n40282 = n40281 ^ n37340;
  assign n40405 = n40292 ^ n40282;
  assign n40406 = ~n40293 & n40405;
  assign n40407 = n40406 ^ n37334;
  assign n40623 = n40417 ^ n40407;
  assign n40624 = n40418 & n40623;
  assign n40625 = n40624 ^ n37472;
  assign n40626 = n40625 ^ n40621;
  assign n40627 = n40622 & ~n40626;
  assign n40628 = n40627 ^ n37328;
  assign n40629 = n40628 ^ n40619;
  assign n40630 = n40620 & ~n40629;
  assign n40631 = n40630 ^ n37322;
  assign n40545 = n40544 ^ n40527;
  assign n40546 = n40532 & ~n40545;
  assign n40547 = n40546 ^ n40531;
  assign n40522 = n39002 ^ n38204;
  assign n40523 = n39528 ^ n39002;
  assign n40524 = n40522 & ~n40523;
  assign n40525 = n40524 ^ n38204;
  assign n40521 = n40031 ^ n39975;
  assign n40526 = n40525 ^ n40521;
  assign n40617 = n40547 ^ n40526;
  assign n40618 = n40617 ^ n37316;
  assign n40679 = n40631 ^ n40618;
  assign n40674 = n40625 ^ n40622;
  assign n40419 = n40418 ^ n40407;
  assign n40256 = n40255 ^ n40244;
  assign n40257 = n40241 ^ n37342;
  assign n40258 = n40257 ^ n40230;
  assign n40259 = n40221 ^ n40175;
  assign n40260 = n40218 ^ n40178;
  assign n40261 = n40215 ^ n40180;
  assign n40262 = n40212 ^ n40183;
  assign n40263 = n40209 ^ n40185;
  assign n40264 = n40200 ^ n40192;
  assign n40265 = n40203 ^ n40190;
  assign n40266 = ~n40264 & ~n40265;
  assign n40267 = n40206 ^ n40187;
  assign n40268 = n40266 & ~n40267;
  assign n40269 = ~n40263 & ~n40268;
  assign n40270 = n40262 & ~n40269;
  assign n40271 = n40261 & n40270;
  assign n40272 = n40260 & ~n40271;
  assign n40273 = n40259 & n40272;
  assign n40274 = n40224 ^ n40173;
  assign n40275 = ~n40273 & n40274;
  assign n40276 = n40227 ^ n40171;
  assign n40277 = n40275 & ~n40276;
  assign n40278 = n40258 & n40277;
  assign n40279 = n40256 & n40278;
  assign n40294 = n40293 ^ n40282;
  assign n40420 = ~n40279 & n40294;
  assign n40675 = n40419 & ~n40420;
  assign n40676 = ~n40674 & n40675;
  assign n40677 = n40628 ^ n40620;
  assign n40678 = n40676 & ~n40677;
  assign n40754 = n40679 ^ n40678;
  assign n40758 = n40757 ^ n40754;
  assign n40760 = n38564 ^ n30220;
  assign n40761 = n40760 ^ n1438;
  assign n40762 = n40761 ^ n28588;
  assign n40759 = n40677 ^ n40676;
  assign n40763 = n40762 ^ n40759;
  assign n40764 = n40675 ^ n40674;
  assign n1411 = n1401 ^ n1317;
  assign n1421 = n1420 ^ n1411;
  assign n1428 = n1427 ^ n1421;
  assign n40765 = n40764 ^ n1428;
  assign n40421 = n40420 ^ n40419;
  assign n1256 = n1216 ^ n1168;
  assign n1257 = n1256 ^ n1253;
  assign n1264 = n1263 ^ n1257;
  assign n40422 = n40421 ^ n1264;
  assign n40296 = n40278 ^ n40256;
  assign n3333 = n3332 ^ n1067;
  assign n3340 = n3339 ^ n3333;
  assign n3341 = n3340 ^ n1230;
  assign n40297 = n40296 ^ n3341;
  assign n40299 = n40276 ^ n40275;
  assign n40303 = n40302 ^ n40299;
  assign n40307 = n40274 ^ n40273;
  assign n40304 = n38088 ^ n30194;
  assign n40305 = n40304 ^ n34769;
  assign n40306 = n40305 ^ n761;
  assign n40308 = n40307 ^ n40306;
  assign n40312 = n40272 ^ n40259;
  assign n40309 = n38149 ^ n30175;
  assign n40310 = n40309 ^ n732;
  assign n40311 = n40310 ^ n28604;
  assign n40313 = n40312 ^ n40311;
  assign n40316 = n38099 ^ n714;
  assign n40317 = n40316 ^ n34236;
  assign n40318 = n40317 ^ n28611;
  assign n40315 = n40270 ^ n40261;
  assign n40319 = n40318 ^ n40315;
  assign n40321 = n38105 ^ n29643;
  assign n40322 = n40321 ^ n34241;
  assign n40323 = n40322 ^ n28616;
  assign n40320 = n40269 ^ n40262;
  assign n40324 = n40323 ^ n40320;
  assign n40326 = n38109 ^ n29670;
  assign n40327 = n40326 ^ n34246;
  assign n40328 = n40327 ^ n28648;
  assign n40325 = n40268 ^ n40263;
  assign n40329 = n40328 ^ n40325;
  assign n40331 = n38130 ^ n29649;
  assign n40332 = n40331 ^ n34250;
  assign n40333 = n40332 ^ n28621;
  assign n40330 = n40267 ^ n40266;
  assign n40334 = n40333 ^ n40330;
  assign n40336 = n34264 ^ n2381;
  assign n40337 = n40336 ^ n2298;
  assign n40338 = n40337 ^ n28625;
  assign n40339 = n40338 ^ n40264;
  assign n40343 = n38621 ^ n2268;
  assign n40344 = n40343 ^ n35101;
  assign n40345 = n40344 ^ n2045;
  assign n40346 = n40193 ^ n37412;
  assign n40347 = n40345 & n40346;
  assign n40340 = n38116 ^ n2280;
  assign n40341 = n40340 ^ n34259;
  assign n40342 = n40341 ^ n28628;
  assign n40348 = n40347 ^ n40342;
  assign n40349 = n40197 ^ n40195;
  assign n40350 = n40349 ^ n40342;
  assign n40351 = n40348 & ~n40350;
  assign n40352 = n40351 ^ n40347;
  assign n40353 = n40352 ^ n40264;
  assign n40354 = ~n40339 & n40353;
  assign n40355 = n40354 ^ n40338;
  assign n40335 = n40265 ^ n40264;
  assign n40356 = n40355 ^ n40335;
  assign n40357 = n29660 ^ n2396;
  assign n40358 = n40357 ^ n34255;
  assign n40359 = n40358 ^ n28639;
  assign n40360 = n40359 ^ n40335;
  assign n40361 = n40356 & ~n40360;
  assign n40362 = n40361 ^ n40359;
  assign n40363 = n40362 ^ n40330;
  assign n40364 = n40334 & ~n40363;
  assign n40365 = n40364 ^ n40333;
  assign n40366 = n40365 ^ n40325;
  assign n40367 = n40329 & ~n40366;
  assign n40368 = n40367 ^ n40328;
  assign n40369 = n40368 ^ n40320;
  assign n40370 = n40324 & ~n40369;
  assign n40371 = n40370 ^ n40323;
  assign n40372 = n40371 ^ n40315;
  assign n40373 = ~n40319 & n40372;
  assign n40374 = n40373 ^ n40318;
  assign n40314 = n40271 ^ n40260;
  assign n40375 = n40374 ^ n40314;
  assign n40376 = n38094 ^ n30180;
  assign n40377 = n40376 ^ n34287;
  assign n40378 = n40377 ^ n605;
  assign n40379 = n40378 ^ n40314;
  assign n40380 = n40375 & ~n40379;
  assign n40381 = n40380 ^ n40378;
  assign n40382 = n40381 ^ n40312;
  assign n40383 = n40313 & ~n40382;
  assign n40384 = n40383 ^ n40311;
  assign n40385 = n40384 ^ n40307;
  assign n40386 = n40308 & ~n40385;
  assign n40387 = n40386 ^ n40306;
  assign n40388 = n40387 ^ n40299;
  assign n40389 = n40303 & ~n40388;
  assign n40390 = n40389 ^ n40302;
  assign n40298 = n40277 ^ n40258;
  assign n40391 = n40390 ^ n40298;
  assign n40395 = n40394 ^ n40298;
  assign n40396 = n40391 & ~n40395;
  assign n40397 = n40396 ^ n40394;
  assign n40398 = n40397 ^ n40296;
  assign n40399 = ~n40297 & n40398;
  assign n40400 = n40399 ^ n3341;
  assign n40295 = n40294 ^ n40279;
  assign n40401 = n40400 ^ n40295;
  assign n1220 = n1201 ^ n1150;
  assign n1239 = n1238 ^ n1220;
  assign n1246 = n1245 ^ n1239;
  assign n40402 = n40295 ^ n1246;
  assign n40403 = n40401 & ~n40402;
  assign n40404 = n40403 ^ n1246;
  assign n40766 = n40421 ^ n40404;
  assign n40767 = n40422 & ~n40766;
  assign n40768 = n40767 ^ n1264;
  assign n40769 = n40768 ^ n40764;
  assign n40770 = n40765 & ~n40769;
  assign n40771 = n40770 ^ n1428;
  assign n40772 = n40771 ^ n40759;
  assign n40773 = n40763 & ~n40772;
  assign n40774 = n40773 ^ n40762;
  assign n40775 = n40774 ^ n40754;
  assign n40776 = n40758 & ~n40775;
  assign n40777 = n40776 ^ n40757;
  assign n40750 = n38574 ^ n2523;
  assign n40751 = n40750 ^ n34741;
  assign n40752 = n40751 ^ n3177;
  assign n40680 = ~n40678 & ~n40679;
  assign n40632 = n40631 ^ n40617;
  assign n40633 = ~n40618 & n40632;
  assign n40634 = n40633 ^ n37316;
  assign n40548 = n40547 ^ n40521;
  assign n40549 = ~n40526 & n40548;
  assign n40550 = n40549 ^ n40525;
  assign n40516 = n38871 ^ n38198;
  assign n40517 = n39522 ^ n38871;
  assign n40518 = n40516 & n40517;
  assign n40519 = n40518 ^ n38198;
  assign n40515 = n40034 ^ n39970;
  assign n40520 = n40519 ^ n40515;
  assign n40615 = n40550 ^ n40520;
  assign n40616 = n40615 ^ n37310;
  assign n40673 = n40634 ^ n40616;
  assign n40749 = n40680 ^ n40673;
  assign n40753 = n40752 ^ n40749;
  assign n41149 = n40777 ^ n40753;
  assign n41154 = n41153 ^ n41149;
  assign n41156 = n39706 ^ n38848;
  assign n40466 = n40070 ^ n3237;
  assign n41157 = n40466 ^ n39706;
  assign n41158 = n41156 & ~n41157;
  assign n41159 = n41158 ^ n38848;
  assign n41155 = n40774 ^ n40758;
  assign n41160 = n41159 ^ n41155;
  assign n41162 = n39492 ^ n38849;
  assign n40472 = n40066 ^ n39941;
  assign n41163 = n40472 ^ n39492;
  assign n41164 = ~n41162 & n41163;
  assign n41165 = n41164 ^ n38849;
  assign n41161 = n40771 ^ n40763;
  assign n41166 = n41165 ^ n41161;
  assign n41169 = n39498 ^ n38859;
  assign n40478 = n40063 ^ n39946;
  assign n41170 = n40478 ^ n39498;
  assign n41171 = n41169 & n41170;
  assign n41172 = n41171 ^ n38859;
  assign n41167 = n40768 ^ n1428;
  assign n41168 = n41167 ^ n40764;
  assign n41173 = n41172 ^ n41168;
  assign n41174 = n39504 ^ n38865;
  assign n40484 = n40060 ^ n40057;
  assign n41175 = n40484 ^ n39504;
  assign n41176 = ~n41174 & ~n41175;
  assign n41177 = n41176 ^ n38865;
  assign n40423 = n40422 ^ n40404;
  assign n41178 = n41177 ^ n40423;
  assign n41183 = n40401 ^ n1246;
  assign n41179 = n39510 ^ n38871;
  assign n40490 = n40053 ^ n39952;
  assign n41180 = n40490 ^ n39510;
  assign n41181 = n41179 & ~n41180;
  assign n41182 = n41181 ^ n38871;
  assign n41184 = n41183 ^ n41182;
  assign n41189 = n40397 ^ n40297;
  assign n41185 = n39516 ^ n39002;
  assign n40496 = n40050 ^ n40047;
  assign n41186 = n40496 ^ n39516;
  assign n41187 = ~n41185 & ~n41186;
  assign n41188 = n41187 ^ n39002;
  assign n41190 = n41189 ^ n41188;
  assign n41195 = n40394 ^ n40391;
  assign n41191 = n39522 ^ n38873;
  assign n40498 = n40043 ^ n39958;
  assign n41192 = n40498 ^ n39522;
  assign n41193 = ~n41191 & ~n41192;
  assign n41194 = n41193 ^ n38873;
  assign n41196 = n41195 ^ n41194;
  assign n41201 = n40387 ^ n40303;
  assign n41197 = n39528 ^ n38883;
  assign n40504 = n40040 ^ n39963;
  assign n41198 = n40504 ^ n39528;
  assign n41199 = n41197 & ~n41198;
  assign n41200 = n41199 ^ n38883;
  assign n41202 = n41201 ^ n41200;
  assign n41207 = n40384 ^ n40308;
  assign n41203 = n39675 ^ n38889;
  assign n40424 = n40037 ^ n39968;
  assign n41204 = n40424 ^ n39675;
  assign n41205 = n41203 & n41204;
  assign n41206 = n41205 ^ n38889;
  assign n41208 = n41207 ^ n41206;
  assign n41213 = n40381 ^ n40313;
  assign n41209 = n39666 ^ n38895;
  assign n41210 = n40515 ^ n39666;
  assign n41211 = ~n41209 & n41210;
  assign n41212 = n41211 ^ n38895;
  assign n41214 = n41213 ^ n41212;
  assign n41109 = n40378 ^ n40375;
  assign n41104 = n39538 ^ n38901;
  assign n41105 = n40521 ^ n39538;
  assign n41106 = ~n41104 & n41105;
  assign n41107 = n41106 ^ n38901;
  assign n41215 = n41109 ^ n41107;
  assign n40972 = n39544 ^ n38907;
  assign n40973 = n40527 ^ n39544;
  assign n40974 = ~n40972 & ~n40973;
  assign n40975 = n40974 ^ n38907;
  assign n40971 = n40371 ^ n40319;
  assign n40976 = n40975 ^ n40971;
  assign n40901 = n40368 ^ n40324;
  assign n40896 = n39550 ^ n38913;
  assign n40897 = n40533 ^ n39550;
  assign n40898 = ~n40896 & ~n40897;
  assign n40899 = n40898 ^ n38913;
  assign n40967 = n40901 ^ n40899;
  assign n40427 = n39556 ^ n38163;
  assign n40428 = n40411 ^ n39556;
  assign n40429 = n40427 & ~n40428;
  assign n40430 = n40429 ^ n38163;
  assign n40426 = n40365 ^ n40329;
  assign n40431 = n40430 ^ n40426;
  assign n40433 = n39562 ^ n38924;
  assign n40434 = n40286 ^ n39562;
  assign n40435 = n40433 & n40434;
  assign n40436 = n40435 ^ n38924;
  assign n40432 = n40362 ^ n40334;
  assign n40437 = n40436 ^ n40432;
  assign n40439 = n38930 ^ n38844;
  assign n40440 = n40248 ^ n38844;
  assign n40441 = n40439 & n40440;
  assign n40442 = n40441 ^ n38930;
  assign n40438 = n40359 ^ n40356;
  assign n40443 = n40442 ^ n40438;
  assign n40878 = n40352 ^ n40339;
  assign n40448 = n40349 ^ n40348;
  assign n40444 = n39461 ^ n38942;
  assign n40445 = n40168 ^ n39461;
  assign n40446 = ~n40444 & n40445;
  assign n40447 = n40446 ^ n38942;
  assign n40449 = n40448 ^ n40447;
  assign n40454 = n40346 ^ n40345;
  assign n40450 = n39468 ^ n38948;
  assign n40451 = n39468 ^ n39451;
  assign n40452 = n40450 & n40451;
  assign n40453 = n40452 ^ n38948;
  assign n40455 = n40454 ^ n40453;
  assign n40831 = n39475 ^ n38954;
  assign n40832 = n39475 ^ n39458;
  assign n40833 = ~n40831 & n40832;
  assign n40834 = n40833 ^ n38954;
  assign n40826 = n38492 ^ n30125;
  assign n40827 = n40826 ^ n1904;
  assign n40828 = n40827 ^ n28885;
  assign n40480 = n38647 ^ n37939;
  assign n40481 = n39706 ^ n38647;
  assign n40482 = n40480 & n40481;
  assign n40483 = n40482 ^ n37939;
  assign n40485 = n40484 ^ n40483;
  assign n40486 = n39181 ^ n38474;
  assign n40487 = n39492 ^ n39181;
  assign n40488 = ~n40486 & n40487;
  assign n40489 = n40488 ^ n38474;
  assign n40491 = n40490 ^ n40489;
  assign n40492 = n38848 ^ n38184;
  assign n40493 = n39498 ^ n38848;
  assign n40494 = n40492 & n40493;
  assign n40495 = n40494 ^ n38184;
  assign n40497 = n40496 ^ n40495;
  assign n40499 = n38849 ^ n38185;
  assign n40500 = n39504 ^ n38849;
  assign n40501 = ~n40499 & n40500;
  assign n40502 = n40501 ^ n38185;
  assign n40503 = n40502 ^ n40498;
  assign n40505 = n38859 ^ n38190;
  assign n40506 = n39510 ^ n38859;
  assign n40507 = ~n40505 & ~n40506;
  assign n40508 = n40507 ^ n38190;
  assign n40509 = n40508 ^ n40504;
  assign n40510 = n38865 ^ n38196;
  assign n40511 = n39516 ^ n38865;
  assign n40512 = ~n40510 & ~n40511;
  assign n40513 = n40512 ^ n38196;
  assign n40514 = n40513 ^ n40424;
  assign n40551 = n40550 ^ n40515;
  assign n40552 = n40520 & ~n40551;
  assign n40553 = n40552 ^ n40519;
  assign n40554 = n40553 ^ n40424;
  assign n40555 = ~n40514 & n40554;
  assign n40556 = n40555 ^ n40513;
  assign n40557 = n40556 ^ n40504;
  assign n40558 = ~n40509 & ~n40557;
  assign n40559 = n40558 ^ n40508;
  assign n40560 = n40559 ^ n40498;
  assign n40561 = ~n40503 & ~n40560;
  assign n40562 = n40561 ^ n40502;
  assign n40563 = n40562 ^ n40496;
  assign n40564 = n40497 & n40563;
  assign n40565 = n40564 ^ n40495;
  assign n40566 = n40565 ^ n40490;
  assign n40567 = n40491 & n40566;
  assign n40568 = n40567 ^ n40489;
  assign n40569 = n40568 ^ n40484;
  assign n40570 = n40485 & ~n40569;
  assign n40571 = n40570 ^ n40483;
  assign n40474 = n38641 ^ n37946;
  assign n40475 = n39899 ^ n38641;
  assign n40476 = ~n40474 & n40475;
  assign n40477 = n40476 ^ n37946;
  assign n40479 = n40478 ^ n40477;
  assign n40600 = n40571 ^ n40479;
  assign n40601 = n40600 ^ n37109;
  assign n40602 = n40568 ^ n40485;
  assign n40603 = n40602 ^ n37102;
  assign n40604 = n40565 ^ n40489;
  assign n40605 = n40604 ^ n40490;
  assign n40606 = n40605 ^ n37714;
  assign n40607 = n40562 ^ n40497;
  assign n40608 = n40607 ^ n37293;
  assign n40609 = n40559 ^ n40503;
  assign n40610 = n40609 ^ n37499;
  assign n40611 = n40556 ^ n40509;
  assign n40612 = n40611 ^ n37298;
  assign n40613 = n40553 ^ n40514;
  assign n40614 = n40613 ^ n37304;
  assign n40635 = n40634 ^ n40615;
  assign n40636 = ~n40616 & ~n40635;
  assign n40637 = n40636 ^ n37310;
  assign n40638 = n40637 ^ n40613;
  assign n40639 = ~n40614 & ~n40638;
  assign n40640 = n40639 ^ n37304;
  assign n40641 = n40640 ^ n40611;
  assign n40642 = ~n40612 & n40641;
  assign n40643 = n40642 ^ n37298;
  assign n40644 = n40643 ^ n40609;
  assign n40645 = n40610 & ~n40644;
  assign n40646 = n40645 ^ n37499;
  assign n40647 = n40646 ^ n40607;
  assign n40648 = n40608 & ~n40647;
  assign n40649 = n40648 ^ n37293;
  assign n40650 = n40649 ^ n40605;
  assign n40651 = n40606 & n40650;
  assign n40652 = n40651 ^ n37714;
  assign n40653 = n40652 ^ n40602;
  assign n40654 = n40603 & n40653;
  assign n40655 = n40654 ^ n37102;
  assign n40656 = n40655 ^ n40600;
  assign n40657 = ~n40601 & n40656;
  assign n40658 = n40657 ^ n37109;
  assign n40572 = n40571 ^ n40478;
  assign n40573 = ~n40479 & n40572;
  assign n40574 = n40573 ^ n40477;
  assign n40468 = n38635 ^ n37929;
  assign n40469 = n39358 ^ n38635;
  assign n40470 = ~n40468 & ~n40469;
  assign n40471 = n40470 ^ n37929;
  assign n40473 = n40472 ^ n40471;
  assign n40598 = n40574 ^ n40473;
  assign n40599 = n40598 ^ n37092;
  assign n40669 = n40658 ^ n40599;
  assign n40670 = n40652 ^ n40603;
  assign n40671 = n40646 ^ n40608;
  assign n40672 = n40643 ^ n40610;
  assign n40681 = n40673 & ~n40680;
  assign n40682 = n40637 ^ n40614;
  assign n40683 = n40681 & ~n40682;
  assign n40684 = n40640 ^ n40612;
  assign n40685 = ~n40683 & ~n40684;
  assign n40686 = n40672 & n40685;
  assign n40687 = n40671 & n40686;
  assign n40688 = n40649 ^ n40606;
  assign n40689 = ~n40687 & ~n40688;
  assign n40690 = n40670 & n40689;
  assign n40691 = n40655 ^ n40601;
  assign n40692 = n40690 & n40691;
  assign n40693 = ~n40669 & n40692;
  assign n40659 = n40658 ^ n40598;
  assign n40660 = n40599 & n40659;
  assign n40661 = n40660 ^ n37092;
  assign n40575 = n40574 ^ n40472;
  assign n40576 = ~n40473 & n40575;
  assign n40577 = n40576 ^ n40471;
  assign n40462 = n38629 ^ n37927;
  assign n40463 = n39369 ^ n38629;
  assign n40464 = ~n40462 & n40463;
  assign n40465 = n40464 ^ n37927;
  assign n40595 = n40577 ^ n40465;
  assign n40596 = n40595 ^ n40466;
  assign n40597 = n40596 ^ n37147;
  assign n40694 = n40661 ^ n40597;
  assign n40695 = ~n40693 & ~n40694;
  assign n40662 = n40661 ^ n40596;
  assign n40663 = n40597 & ~n40662;
  assign n40664 = n40663 ^ n37147;
  assign n40467 = n40466 ^ n40465;
  assign n40578 = n40577 ^ n40466;
  assign n40579 = ~n40467 & n40578;
  assign n40580 = n40579 ^ n40465;
  assign n40457 = n38623 ^ n37917;
  assign n40458 = n39352 ^ n38623;
  assign n40459 = ~n40457 & ~n40458;
  assign n40460 = n40459 ^ n37917;
  assign n40592 = n40580 ^ n40460;
  assign n40593 = n40592 ^ n40456;
  assign n40594 = n40593 ^ n37192;
  assign n40696 = n40664 ^ n40594;
  assign n40697 = n40695 & n40696;
  assign n40665 = n40664 ^ n40593;
  assign n40666 = ~n40594 & n40665;
  assign n40667 = n40666 ^ n37192;
  assign n40586 = n38178 ^ n37291;
  assign n40587 = n39346 ^ n38178;
  assign n40588 = n40586 & ~n40587;
  assign n40589 = n40588 ^ n37291;
  assign n40584 = n40077 ^ n2938;
  assign n40461 = n40460 ^ n40456;
  assign n40581 = n40580 ^ n40456;
  assign n40582 = n40461 & n40581;
  assign n40583 = n40582 ^ n40460;
  assign n40585 = n40584 ^ n40583;
  assign n40590 = n40589 ^ n40585;
  assign n40591 = n40590 ^ n37250;
  assign n40668 = n40667 ^ n40591;
  assign n40718 = n40697 ^ n40668;
  assign n40715 = n38497 ^ n30130;
  assign n40716 = n40715 ^ n34709;
  assign n40717 = n40716 ^ n1896;
  assign n40719 = n40718 ^ n40717;
  assign n40720 = n40696 ^ n40695;
  assign n1767 = n1766 ^ n1745;
  assign n1795 = n1794 ^ n1767;
  assign n1802 = n1801 ^ n1795;
  assign n40721 = n40720 ^ n1802;
  assign n40724 = n38509 ^ n1689;
  assign n40725 = n40724 ^ n34716;
  assign n40726 = n40725 ^ n28556;
  assign n40723 = n40692 ^ n40669;
  assign n40727 = n40726 ^ n40723;
  assign n40728 = n40691 ^ n40690;
  assign n40732 = n40731 ^ n40728;
  assign n40734 = n40688 ^ n40687;
  assign n40738 = n40737 ^ n40734;
  assign n40740 = n38525 ^ n30149;
  assign n40741 = n40740 ^ n2702;
  assign n40742 = n40741 ^ n3110;
  assign n40739 = n40686 ^ n40671;
  assign n40743 = n40742 ^ n40739;
  assign n40744 = n40685 ^ n40672;
  assign n3090 = n3089 ^ n3083;
  assign n3094 = n3093 ^ n3090;
  assign n3095 = n3094 ^ n2700;
  assign n40745 = n40744 ^ n3095;
  assign n40746 = n40684 ^ n40683;
  assign n2589 = n2588 ^ n2573;
  assign n2617 = n2616 ^ n2589;
  assign n2624 = n2623 ^ n2617;
  assign n40747 = n40746 ^ n2624;
  assign n40778 = n40777 ^ n40749;
  assign n40779 = n40753 & ~n40778;
  assign n40780 = n40779 ^ n40752;
  assign n40748 = n40682 ^ n40681;
  assign n40781 = n40780 ^ n40748;
  assign n40782 = n38533 ^ n3069;
  assign n40783 = n40782 ^ n3179;
  assign n40784 = n40783 ^ n2614;
  assign n40785 = n40784 ^ n40748;
  assign n40786 = ~n40781 & n40785;
  assign n40787 = n40786 ^ n40784;
  assign n40788 = n40787 ^ n40746;
  assign n40789 = n40747 & ~n40788;
  assign n40790 = n40789 ^ n2624;
  assign n40791 = n40790 ^ n40744;
  assign n40792 = n40745 & ~n40791;
  assign n40793 = n40792 ^ n3095;
  assign n40794 = n40793 ^ n40739;
  assign n40795 = n40743 & ~n40794;
  assign n40796 = n40795 ^ n40742;
  assign n40797 = n40796 ^ n40734;
  assign n40798 = ~n40738 & n40797;
  assign n40799 = n40798 ^ n40737;
  assign n40733 = n40689 ^ n40670;
  assign n40800 = n40799 ^ n40733;
  assign n40801 = n38515 ^ n2994;
  assign n40802 = n40801 ^ n34726;
  assign n40803 = n40802 ^ n28566;
  assign n40804 = n40803 ^ n40733;
  assign n40805 = n40800 & ~n40804;
  assign n40806 = n40805 ^ n40803;
  assign n40807 = n40806 ^ n40728;
  assign n40808 = ~n40732 & n40807;
  assign n40809 = n40808 ^ n40731;
  assign n40810 = n40809 ^ n40723;
  assign n40811 = n40727 & ~n40810;
  assign n40812 = n40811 ^ n40726;
  assign n40722 = n40694 ^ n40693;
  assign n40813 = n40812 ^ n40722;
  assign n40814 = n38504 ^ n30136;
  assign n40815 = n40814 ^ n34839;
  assign n40816 = n40815 ^ n1786;
  assign n40817 = n40816 ^ n40722;
  assign n40818 = ~n40813 & n40817;
  assign n40819 = n40818 ^ n40816;
  assign n40820 = n40819 ^ n40720;
  assign n40821 = n40721 & ~n40820;
  assign n40822 = n40821 ^ n1802;
  assign n40823 = n40822 ^ n40718;
  assign n40824 = n40719 & ~n40823;
  assign n40825 = n40824 ^ n40717;
  assign n40829 = n40828 ^ n40825;
  assign n40709 = n40667 ^ n40590;
  assign n40710 = ~n40591 & n40709;
  assign n40711 = n40710 ^ n37250;
  assign n40712 = n40711 ^ n37414;
  assign n40707 = n40080 ^ n39932;
  assign n40703 = n40589 ^ n40584;
  assign n40704 = n40585 & ~n40703;
  assign n40705 = n40704 ^ n40589;
  assign n40699 = n38172 ^ n37284;
  assign n40700 = n39340 ^ n38172;
  assign n40701 = n40699 & ~n40700;
  assign n40702 = n40701 ^ n37284;
  assign n40706 = n40705 ^ n40702;
  assign n40708 = n40707 ^ n40706;
  assign n40713 = n40712 ^ n40708;
  assign n40698 = n40668 & n40697;
  assign n40714 = n40713 ^ n40698;
  assign n40830 = n40829 ^ n40714;
  assign n40835 = n40834 ^ n40830;
  assign n40837 = n39483 ^ n38830;
  assign n40838 = n39483 ^ n39465;
  assign n40839 = ~n40837 & n40838;
  assign n40840 = n40839 ^ n38830;
  assign n40836 = n40822 ^ n40719;
  assign n40841 = n40840 ^ n40836;
  assign n40843 = n39598 ^ n38726;
  assign n40844 = n39598 ^ n39472;
  assign n40845 = ~n40843 & n40844;
  assign n40846 = n40845 ^ n38726;
  assign n40842 = n40819 ^ n40721;
  assign n40847 = n40846 ^ n40842;
  assign n40849 = n39604 ^ n38166;
  assign n40850 = n39604 ^ n39479;
  assign n40851 = n40849 & ~n40850;
  assign n40852 = n40851 ^ n38166;
  assign n40848 = n40816 ^ n40813;
  assign n40853 = n40852 ^ n40848;
  assign n40854 = n39606 ^ n38671;
  assign n40855 = n39606 ^ n39481;
  assign n40856 = n40854 & ~n40855;
  assign n40857 = n40856 ^ n38671;
  assign n40858 = n40809 ^ n40727;
  assign n40859 = ~n40857 & n40858;
  assign n40860 = n40859 ^ n40848;
  assign n40861 = ~n40853 & n40860;
  assign n40862 = n40861 ^ n40859;
  assign n40863 = n40862 ^ n40842;
  assign n40864 = n40847 & ~n40863;
  assign n40865 = n40864 ^ n40846;
  assign n40866 = n40865 ^ n40836;
  assign n40867 = ~n40841 & ~n40866;
  assign n40868 = n40867 ^ n40840;
  assign n40869 = n40868 ^ n40830;
  assign n40870 = ~n40835 & n40869;
  assign n40871 = n40870 ^ n40834;
  assign n40872 = n40871 ^ n40454;
  assign n40873 = n40455 & n40872;
  assign n40874 = n40873 ^ n40453;
  assign n40875 = n40874 ^ n40448;
  assign n40876 = ~n40449 & ~n40875;
  assign n40877 = n40876 ^ n40447;
  assign n40879 = n40878 ^ n40877;
  assign n40880 = n39454 ^ n38936;
  assign n40881 = n40239 ^ n39454;
  assign n40882 = n40880 & ~n40881;
  assign n40883 = n40882 ^ n38936;
  assign n40884 = n40883 ^ n40877;
  assign n40885 = n40879 & n40884;
  assign n40886 = n40885 ^ n40878;
  assign n40887 = n40886 ^ n40438;
  assign n40888 = n40443 & ~n40887;
  assign n40889 = n40888 ^ n40442;
  assign n40890 = n40889 ^ n40432;
  assign n40891 = n40437 & n40890;
  assign n40892 = n40891 ^ n40436;
  assign n40893 = n40892 ^ n40426;
  assign n40894 = n40431 & ~n40893;
  assign n40895 = n40894 ^ n40430;
  assign n40968 = n40901 ^ n40895;
  assign n40969 = ~n40967 & ~n40968;
  assign n40970 = n40969 ^ n40899;
  assign n41101 = n40971 ^ n40970;
  assign n41102 = n40976 & ~n41101;
  assign n41103 = n41102 ^ n40975;
  assign n41216 = n41109 ^ n41103;
  assign n41217 = n41215 & ~n41216;
  assign n41218 = n41217 ^ n41107;
  assign n41219 = n41218 ^ n41213;
  assign n41220 = n41214 & n41219;
  assign n41221 = n41220 ^ n41212;
  assign n41222 = n41221 ^ n41207;
  assign n41223 = n41208 & ~n41222;
  assign n41224 = n41223 ^ n41206;
  assign n41225 = n41224 ^ n41201;
  assign n41226 = n41202 & ~n41225;
  assign n41227 = n41226 ^ n41200;
  assign n41228 = n41227 ^ n41195;
  assign n41229 = ~n41196 & n41228;
  assign n41230 = n41229 ^ n41194;
  assign n41231 = n41230 ^ n41189;
  assign n41232 = ~n41190 & n41231;
  assign n41233 = n41232 ^ n41188;
  assign n41234 = n41233 ^ n41183;
  assign n41235 = ~n41184 & n41234;
  assign n41236 = n41235 ^ n41182;
  assign n41237 = n41236 ^ n40423;
  assign n41238 = ~n41178 & ~n41237;
  assign n41239 = n41238 ^ n41177;
  assign n41240 = n41239 ^ n41168;
  assign n41241 = n41173 & n41240;
  assign n41242 = n41241 ^ n41172;
  assign n41243 = n41242 ^ n41161;
  assign n41244 = ~n41166 & ~n41243;
  assign n41245 = n41244 ^ n41165;
  assign n41246 = n41245 ^ n41155;
  assign n41247 = ~n41160 & n41246;
  assign n41248 = n41247 ^ n41159;
  assign n41249 = n41248 ^ n41149;
  assign n41250 = ~n41154 & n41249;
  assign n41251 = n41250 ^ n41153;
  assign n41144 = n39358 ^ n38647;
  assign n41145 = n40584 ^ n39358;
  assign n41146 = ~n41144 & n41145;
  assign n41147 = n41146 ^ n38647;
  assign n41143 = n40784 ^ n40781;
  assign n41148 = n41147 ^ n41143;
  assign n41268 = n41251 ^ n41148;
  assign n41269 = n41268 ^ n37939;
  assign n41270 = n41248 ^ n41153;
  assign n41271 = n41270 ^ n41149;
  assign n41272 = n41271 ^ n38474;
  assign n41273 = n41245 ^ n41160;
  assign n41274 = n41273 ^ n38184;
  assign n41275 = n41242 ^ n41166;
  assign n41276 = n41275 ^ n38185;
  assign n41277 = n41239 ^ n41173;
  assign n41278 = n41277 ^ n38190;
  assign n41279 = n41236 ^ n41178;
  assign n41280 = n41279 ^ n38196;
  assign n41281 = n41233 ^ n41184;
  assign n41282 = n41281 ^ n38198;
  assign n41283 = n41230 ^ n41190;
  assign n41284 = n41283 ^ n38204;
  assign n41285 = n41227 ^ n41196;
  assign n41286 = n41285 ^ n38210;
  assign n41287 = n41224 ^ n41200;
  assign n41288 = n41287 ^ n41201;
  assign n41289 = n41288 ^ n38220;
  assign n41290 = n41221 ^ n41208;
  assign n41291 = n41290 ^ n38226;
  assign n41292 = n41218 ^ n41212;
  assign n41293 = n41292 ^ n41213;
  assign n41294 = n41293 ^ n38228;
  assign n41108 = n41107 ^ n41103;
  assign n41110 = n41109 ^ n41108;
  assign n41111 = n41110 ^ n38234;
  assign n40977 = n40976 ^ n40970;
  assign n40978 = n40977 ^ n38240;
  assign n40900 = n40899 ^ n40895;
  assign n40902 = n40901 ^ n40900;
  assign n40903 = n40902 ^ n38246;
  assign n40904 = n40892 ^ n40430;
  assign n40905 = n40904 ^ n40426;
  assign n40906 = n40905 ^ n38164;
  assign n40907 = n40889 ^ n40436;
  assign n40908 = n40907 ^ n40432;
  assign n40909 = n40908 ^ n38257;
  assign n40910 = n40886 ^ n40442;
  assign n40911 = n40910 ^ n40438;
  assign n40912 = n40911 ^ n38267;
  assign n40913 = n40874 ^ n40447;
  assign n40914 = n40913 ^ n40448;
  assign n40915 = n40914 ^ n38168;
  assign n40917 = n40868 ^ n40835;
  assign n40918 = n40917 ^ n37981;
  assign n40919 = n40865 ^ n40840;
  assign n40920 = n40919 ^ n40836;
  assign n40921 = n40920 ^ n37256;
  assign n40922 = n40862 ^ n40846;
  assign n40923 = n40922 ^ n40842;
  assign n40924 = n40923 ^ n37263;
  assign n40925 = n40858 ^ n40857;
  assign n40926 = ~n37277 & ~n40925;
  assign n40927 = n40926 ^ n37270;
  assign n40928 = n40859 ^ n40852;
  assign n40929 = n40928 ^ n40848;
  assign n40930 = n40929 ^ n40926;
  assign n40931 = n40927 & ~n40930;
  assign n40932 = n40931 ^ n37270;
  assign n40933 = n40932 ^ n40923;
  assign n40934 = ~n40924 & ~n40933;
  assign n40935 = n40934 ^ n37263;
  assign n40936 = n40935 ^ n40920;
  assign n40937 = n40921 & ~n40936;
  assign n40938 = n40937 ^ n37256;
  assign n40939 = n40938 ^ n40917;
  assign n40940 = ~n40918 & n40939;
  assign n40941 = n40940 ^ n37981;
  assign n40916 = n40871 ^ n40455;
  assign n40942 = n40941 ^ n40916;
  assign n40943 = n40916 ^ n38047;
  assign n40944 = ~n40942 & n40943;
  assign n40945 = n40944 ^ n38047;
  assign n40946 = n40945 ^ n40914;
  assign n40947 = ~n40915 & ~n40946;
  assign n40948 = n40947 ^ n38168;
  assign n40949 = n40948 ^ n38269;
  assign n40950 = n40883 ^ n40878;
  assign n40951 = n40950 ^ n40877;
  assign n40952 = n40951 ^ n40948;
  assign n40953 = ~n40949 & ~n40952;
  assign n40954 = n40953 ^ n38269;
  assign n40955 = n40954 ^ n40911;
  assign n40956 = ~n40912 & ~n40955;
  assign n40957 = n40956 ^ n38267;
  assign n40958 = n40957 ^ n40908;
  assign n40959 = ~n40909 & n40958;
  assign n40960 = n40959 ^ n38257;
  assign n40961 = n40960 ^ n40905;
  assign n40962 = ~n40906 & ~n40961;
  assign n40963 = n40962 ^ n38164;
  assign n40964 = n40963 ^ n40902;
  assign n40965 = ~n40903 & ~n40964;
  assign n40966 = n40965 ^ n38246;
  assign n41098 = n40977 ^ n40966;
  assign n41099 = n40978 & n41098;
  assign n41100 = n41099 ^ n38240;
  assign n41295 = n41110 ^ n41100;
  assign n41296 = n41111 & ~n41295;
  assign n41297 = n41296 ^ n38234;
  assign n41298 = n41297 ^ n41293;
  assign n41299 = ~n41294 & ~n41298;
  assign n41300 = n41299 ^ n38228;
  assign n41301 = n41300 ^ n41290;
  assign n41302 = n41291 & ~n41301;
  assign n41303 = n41302 ^ n38226;
  assign n41304 = n41303 ^ n41288;
  assign n41305 = n41289 & ~n41304;
  assign n41306 = n41305 ^ n38220;
  assign n41307 = n41306 ^ n41285;
  assign n41308 = ~n41286 & n41307;
  assign n41309 = n41308 ^ n38210;
  assign n41310 = n41309 ^ n41283;
  assign n41311 = ~n41284 & n41310;
  assign n41312 = n41311 ^ n38204;
  assign n41313 = n41312 ^ n41281;
  assign n41314 = ~n41282 & n41313;
  assign n41315 = n41314 ^ n38198;
  assign n41316 = n41315 ^ n41279;
  assign n41317 = ~n41280 & n41316;
  assign n41318 = n41317 ^ n38196;
  assign n41319 = n41318 ^ n41277;
  assign n41320 = n41278 & n41319;
  assign n41321 = n41320 ^ n38190;
  assign n41322 = n41321 ^ n41275;
  assign n41323 = ~n41276 & ~n41322;
  assign n41324 = n41323 ^ n38185;
  assign n41325 = n41324 ^ n41273;
  assign n41326 = ~n41274 & ~n41325;
  assign n41327 = n41326 ^ n38184;
  assign n41328 = n41327 ^ n41271;
  assign n41329 = n41272 & n41328;
  assign n41330 = n41329 ^ n38474;
  assign n41331 = n41330 ^ n41268;
  assign n41332 = ~n41269 & n41331;
  assign n41333 = n41332 ^ n37939;
  assign n41252 = n41251 ^ n41143;
  assign n41253 = n41148 & n41252;
  assign n41254 = n41253 ^ n41147;
  assign n41138 = n39369 ^ n38641;
  assign n41139 = n40707 ^ n39369;
  assign n41140 = ~n41138 & n41139;
  assign n41141 = n41140 ^ n38641;
  assign n41137 = n40787 ^ n40747;
  assign n41142 = n41141 ^ n41137;
  assign n41266 = n41254 ^ n41142;
  assign n41267 = n41266 ^ n37946;
  assign n41368 = n41333 ^ n41267;
  assign n41342 = n41330 ^ n41269;
  assign n41343 = n41312 ^ n41282;
  assign n41344 = n41306 ^ n41286;
  assign n41345 = n41303 ^ n41289;
  assign n41346 = n41300 ^ n41291;
  assign n40979 = n40978 ^ n40966;
  assign n40980 = n40963 ^ n40903;
  assign n40981 = n40957 ^ n40909;
  assign n40982 = n40951 ^ n38269;
  assign n40983 = n40982 ^ n40948;
  assign n40984 = n40945 ^ n40915;
  assign n40985 = n40942 ^ n38047;
  assign n40986 = n40938 ^ n40918;
  assign n40987 = n40932 ^ n40924;
  assign n40988 = n40935 ^ n40921;
  assign n40989 = n40987 & n40988;
  assign n40990 = ~n40986 & n40989;
  assign n40991 = ~n40985 & ~n40990;
  assign n40992 = ~n40984 & ~n40991;
  assign n40993 = n40983 & n40992;
  assign n40994 = n40954 ^ n40912;
  assign n40995 = ~n40993 & n40994;
  assign n40996 = ~n40981 & n40995;
  assign n40997 = n40960 ^ n40906;
  assign n40998 = ~n40996 & n40997;
  assign n40999 = ~n40980 & n40998;
  assign n41097 = ~n40979 & n40999;
  assign n41112 = n41111 ^ n41100;
  assign n41347 = n41097 & n41112;
  assign n41348 = n41297 ^ n38228;
  assign n41349 = n41348 ^ n41293;
  assign n41350 = ~n41347 & n41349;
  assign n41351 = ~n41346 & ~n41350;
  assign n41352 = ~n41345 & n41351;
  assign n41353 = n41344 & n41352;
  assign n41354 = n41309 ^ n41284;
  assign n41355 = ~n41353 & ~n41354;
  assign n41356 = n41343 & ~n41355;
  assign n41357 = n41315 ^ n41280;
  assign n41358 = n41356 & n41357;
  assign n41359 = n41318 ^ n41278;
  assign n41360 = ~n41358 & n41359;
  assign n41361 = n41321 ^ n41276;
  assign n41362 = n41360 & n41361;
  assign n41363 = n41324 ^ n41274;
  assign n41364 = n41362 & ~n41363;
  assign n41365 = n41327 ^ n41272;
  assign n41366 = ~n41364 & n41365;
  assign n41367 = n41342 & n41366;
  assign n41441 = n41368 ^ n41367;
  assign n41445 = n41444 ^ n41441;
  assign n41447 = n41365 ^ n41364;
  assign n3133 = n3125 ^ n3117;
  assign n3134 = n3133 ^ n2803;
  assign n3135 = n3134 ^ n2890;
  assign n41448 = n41447 ^ n3135;
  assign n41449 = n41363 ^ n41362;
  assign n2764 = n2760 ^ n2730;
  assign n2789 = n2788 ^ n2764;
  assign n2796 = n2795 ^ n2789;
  assign n41450 = n41449 ^ n2796;
  assign n41451 = n41361 ^ n41360;
  assign n3204 = n3203 ^ n2680;
  assign n3214 = n3213 ^ n3204;
  assign n3215 = n3214 ^ n2780;
  assign n41452 = n41451 ^ n3215;
  assign n41456 = n41359 ^ n41358;
  assign n41453 = n39301 ^ n2665;
  assign n41454 = n41453 ^ n35485;
  assign n41455 = n41454 ^ n3211;
  assign n41457 = n41456 ^ n41455;
  assign n41461 = n41357 ^ n41356;
  assign n41458 = n39231 ^ n3189;
  assign n41459 = n41458 ^ n35489;
  assign n41460 = n41459 ^ n29405;
  assign n41462 = n41461 ^ n41460;
  assign n41465 = n39238 ^ n31006;
  assign n41466 = n41465 ^ n35499;
  assign n41467 = n41466 ^ n3035;
  assign n41464 = n41354 ^ n41353;
  assign n41468 = n41467 ^ n41464;
  assign n41472 = n41352 ^ n41344;
  assign n41469 = n31001 ^ n1475;
  assign n41470 = n41469 ^ n35504;
  assign n41471 = n41470 ^ n2429;
  assign n41473 = n41472 ^ n41471;
  assign n41476 = n39275 ^ n1353;
  assign n41477 = n41476 ^ n35515;
  assign n41478 = n41477 ^ n29424;
  assign n41475 = n41350 ^ n41346;
  assign n41479 = n41478 ^ n41475;
  assign n41113 = n41112 ^ n41097;
  assign n41094 = n39252 ^ n3347;
  assign n41095 = n41094 ^ n950;
  assign n41096 = n41095 ^ n29095;
  assign n41114 = n41113 ^ n41096;
  assign n41003 = n38755 ^ n30469;
  assign n41004 = n41003 ^ n35534;
  assign n41005 = n41004 ^ n832;
  assign n41002 = n40997 ^ n40996;
  assign n41006 = n41005 ^ n41002;
  assign n41008 = n38818 ^ n632;
  assign n41009 = n41008 ^ n35539;
  assign n41010 = n41009 ^ n3296;
  assign n41007 = n40995 ^ n40981;
  assign n41011 = n41010 ^ n41007;
  assign n41014 = n38766 ^ n30501;
  assign n41015 = n41014 ^ n35549;
  assign n41016 = n41015 ^ n29026;
  assign n41013 = n40992 ^ n40983;
  assign n41017 = n41016 ^ n41013;
  assign n41021 = n40991 ^ n40984;
  assign n41018 = n38770 ^ n30506;
  assign n41019 = n41018 ^ n35553;
  assign n41020 = n41019 ^ n29031;
  assign n41022 = n41021 ^ n41020;
  assign n41026 = n40990 ^ n40985;
  assign n41023 = n38775 ^ n30511;
  assign n41024 = n41023 ^ n35558;
  assign n41025 = n41024 ^ n29035;
  assign n41027 = n41026 ^ n41025;
  assign n41029 = n38799 ^ n30534;
  assign n41030 = n41029 ^ n35564;
  assign n41031 = n41030 ^ n29039;
  assign n41028 = n40989 ^ n40986;
  assign n41032 = n41031 ^ n41028;
  assign n41034 = n38781 ^ n30526;
  assign n41035 = n41034 ^ n2333;
  assign n41036 = n41035 ^ n28809;
  assign n41033 = n40988 ^ n40987;
  assign n41037 = n41036 ^ n41033;
  assign n41038 = n38787 ^ n30518;
  assign n41039 = n41038 ^ n34883;
  assign n41040 = n41039 ^ n2324;
  assign n41041 = n41040 ^ n40987;
  assign n41042 = n39196 ^ n30971;
  assign n41043 = n41042 ^ n2023;
  assign n41044 = n41043 ^ n2143;
  assign n41045 = n40925 ^ n37277;
  assign n41046 = n41044 & n41045;
  assign n2136 = n2135 ^ n2066;
  assign n2152 = n2151 ^ n2136;
  assign n2159 = n2158 ^ n2152;
  assign n41047 = n41046 ^ n2159;
  assign n41048 = n40929 ^ n40927;
  assign n41049 = n41048 ^ n2159;
  assign n41050 = n41047 & ~n41049;
  assign n41051 = n41050 ^ n41046;
  assign n41052 = n41051 ^ n40987;
  assign n41053 = n41041 & ~n41052;
  assign n41054 = n41053 ^ n41040;
  assign n41055 = n41054 ^ n41033;
  assign n41056 = ~n41037 & n41055;
  assign n41057 = n41056 ^ n41036;
  assign n41058 = n41057 ^ n41028;
  assign n41059 = n41032 & ~n41058;
  assign n41060 = n41059 ^ n41031;
  assign n41061 = n41060 ^ n41026;
  assign n41062 = n41027 & ~n41061;
  assign n41063 = n41062 ^ n41025;
  assign n41064 = n41063 ^ n41021;
  assign n41065 = ~n41022 & n41064;
  assign n41066 = n41065 ^ n41020;
  assign n41067 = n41066 ^ n41013;
  assign n41068 = ~n41017 & n41067;
  assign n41069 = n41068 ^ n41016;
  assign n41012 = n40994 ^ n40993;
  assign n41070 = n41069 ^ n41012;
  assign n41074 = n41073 ^ n41012;
  assign n41075 = n41070 & ~n41074;
  assign n41076 = n41075 ^ n41073;
  assign n41077 = n41076 ^ n41007;
  assign n41078 = ~n41011 & n41077;
  assign n41079 = n41078 ^ n41010;
  assign n41080 = n41079 ^ n41002;
  assign n41081 = n41006 & ~n41080;
  assign n41082 = n41081 ^ n41005;
  assign n41001 = n40998 ^ n40980;
  assign n41083 = n41082 ^ n41001;
  assign n813 = n812 ^ n788;
  assign n841 = n840 ^ n813;
  assign n848 = n847 ^ n841;
  assign n41084 = n41001 ^ n848;
  assign n41085 = ~n41083 & n41084;
  assign n41086 = n41085 ^ n848;
  assign n41000 = n40999 ^ n40979;
  assign n41087 = n41086 ^ n41000;
  assign n41088 = n39257 ^ n30484;
  assign n41089 = n41088 ^ n35527;
  assign n41090 = n41089 ^ n942;
  assign n41091 = n41090 ^ n41000;
  assign n41092 = ~n41087 & n41091;
  assign n41093 = n41092 ^ n41090;
  assign n41481 = n41113 ^ n41093;
  assign n41482 = ~n41114 & n41481;
  assign n41483 = n41482 ^ n41096;
  assign n41480 = n41349 ^ n41347;
  assign n41484 = n41483 ^ n41480;
  assign n41485 = n39247 ^ n1338;
  assign n41486 = n41485 ^ n35520;
  assign n41487 = n41486 ^ n1100;
  assign n41488 = n41487 ^ n41480;
  assign n41489 = n41484 & ~n41488;
  assign n41490 = n41489 ^ n41487;
  assign n41491 = n41490 ^ n41475;
  assign n41492 = ~n41479 & n41491;
  assign n41493 = n41492 ^ n41478;
  assign n41474 = n41351 ^ n41345;
  assign n41494 = n41493 ^ n41474;
  assign n41495 = n1460 ^ n1371;
  assign n41496 = n41495 ^ n35509;
  assign n41497 = n41496 ^ n29418;
  assign n41498 = n41497 ^ n41474;
  assign n41499 = ~n41494 & n41498;
  assign n41500 = n41499 ^ n41497;
  assign n41501 = n41500 ^ n41472;
  assign n41502 = ~n41473 & n41501;
  assign n41503 = n41502 ^ n41471;
  assign n41504 = n41503 ^ n41464;
  assign n41505 = n41468 & ~n41504;
  assign n41506 = n41505 ^ n41467;
  assign n41463 = n41355 ^ n41343;
  assign n41507 = n41506 ^ n41463;
  assign n41508 = n39291 ^ n30996;
  assign n41509 = n41508 ^ n35494;
  assign n41510 = n41509 ^ n29410;
  assign n41511 = n41510 ^ n41463;
  assign n41512 = ~n41507 & n41511;
  assign n41513 = n41512 ^ n41510;
  assign n41514 = n41513 ^ n41461;
  assign n41515 = ~n41462 & n41514;
  assign n41516 = n41515 ^ n41460;
  assign n41517 = n41516 ^ n41456;
  assign n41518 = ~n41457 & n41517;
  assign n41519 = n41518 ^ n41455;
  assign n41520 = n41519 ^ n41451;
  assign n41521 = n41452 & ~n41520;
  assign n41522 = n41521 ^ n3215;
  assign n41523 = n41522 ^ n41449;
  assign n41524 = ~n41450 & n41523;
  assign n41525 = n41524 ^ n2796;
  assign n41526 = n41525 ^ n41447;
  assign n41527 = n41448 & ~n41526;
  assign n41528 = n41527 ^ n3135;
  assign n41446 = n41366 ^ n41342;
  assign n41529 = n41528 ^ n41446;
  assign n2886 = n2885 ^ n2828;
  assign n2893 = n2892 ^ n2886;
  assign n2894 = n2893 ^ n1601;
  assign n41530 = n41446 ^ n2894;
  assign n41531 = n41529 & ~n41530;
  assign n41532 = n41531 ^ n2894;
  assign n41533 = n41532 ^ n41441;
  assign n41534 = ~n41445 & n41533;
  assign n41535 = n41534 ^ n41444;
  assign n41369 = n41367 & n41368;
  assign n41334 = n41333 ^ n41266;
  assign n41335 = ~n41267 & n41334;
  assign n41336 = n41335 ^ n37946;
  assign n41255 = n41254 ^ n41137;
  assign n41256 = ~n41142 & ~n41255;
  assign n41257 = n41256 ^ n41141;
  assign n41135 = n40790 ^ n40745;
  assign n41131 = n39352 ^ n38635;
  assign n41132 = n40128 ^ n39352;
  assign n41133 = ~n41131 & ~n41132;
  assign n41134 = n41133 ^ n38635;
  assign n41136 = n41135 ^ n41134;
  assign n41264 = n41257 ^ n41136;
  assign n41265 = n41264 ^ n37929;
  assign n41341 = n41336 ^ n41265;
  assign n41436 = n41369 ^ n41341;
  assign n41440 = n41439 ^ n41436;
  assign n41577 = n41535 ^ n41440;
  assign n41573 = n39606 ^ n39472;
  assign n41574 = n40454 ^ n39472;
  assign n41575 = ~n41573 & ~n41574;
  assign n41576 = n41575 ^ n39606;
  assign n41600 = n41577 ^ n41576;
  assign n41699 = n41600 ^ n38671;
  assign n41700 = n41698 & n41699;
  assign n2258 = n2246 ^ n2185;
  assign n2274 = n2273 ^ n2258;
  assign n2281 = n2280 ^ n2274;
  assign n41701 = n41700 ^ n2281;
  assign n41578 = ~n41576 & n41577;
  assign n41568 = n39604 ^ n39465;
  assign n41569 = n40448 ^ n39465;
  assign n41570 = ~n41568 & n41569;
  assign n41571 = n41570 ^ n39604;
  assign n41603 = n41578 ^ n41571;
  assign n41536 = n41535 ^ n41436;
  assign n41537 = n41440 & ~n41536;
  assign n41538 = n41537 ^ n41439;
  assign n41370 = ~n41341 & n41369;
  assign n41337 = n41336 ^ n41264;
  assign n41338 = n41265 & ~n41337;
  assign n41339 = n41338 ^ n37929;
  assign n41258 = n41257 ^ n41135;
  assign n41259 = ~n41136 & n41258;
  assign n41260 = n41259 ^ n41134;
  assign n41127 = n39346 ^ n38629;
  assign n41128 = n40122 ^ n39346;
  assign n41129 = n41127 & n41128;
  assign n41130 = n41129 ^ n38629;
  assign n41261 = n41260 ^ n41130;
  assign n41126 = n40793 ^ n40743;
  assign n41262 = n41261 ^ n41126;
  assign n41263 = n41262 ^ n37927;
  assign n41340 = n41339 ^ n41263;
  assign n41434 = n41370 ^ n41340;
  assign n41431 = n39212 ^ n31061;
  assign n41432 = n41431 ^ n35462;
  assign n41433 = n41432 ^ n29381;
  assign n41435 = n41434 ^ n41433;
  assign n41567 = n41538 ^ n41435;
  assign n41604 = n41603 ^ n41567;
  assign n41601 = ~n38671 & ~n41600;
  assign n41602 = n41601 ^ n38166;
  assign n41702 = n41604 ^ n41602;
  assign n41703 = n41702 ^ n2281;
  assign n41704 = n41701 & n41703;
  assign n41705 = n41704 ^ n41700;
  assign n41605 = n41604 ^ n41601;
  assign n41606 = n41602 & n41605;
  assign n41607 = n41606 ^ n38166;
  assign n41572 = n41571 ^ n41567;
  assign n41579 = n41578 ^ n41567;
  assign n41580 = n41572 & ~n41579;
  assign n41581 = n41580 ^ n41578;
  assign n41562 = n39598 ^ n39458;
  assign n41563 = n40878 ^ n39458;
  assign n41564 = n41562 & ~n41563;
  assign n41565 = n41564 ^ n39598;
  assign n41539 = n41538 ^ n41434;
  assign n41540 = ~n41435 & n41539;
  assign n41541 = n41540 ^ n41433;
  assign n41427 = n39207 ^ n1852;
  assign n41428 = n41427 ^ n35457;
  assign n41429 = n41428 ^ n29376;
  assign n41384 = n41339 ^ n41262;
  assign n41385 = n41263 & ~n41384;
  assign n41386 = n41385 ^ n37927;
  assign n41378 = n39340 ^ n38623;
  assign n41379 = n40116 ^ n39340;
  assign n41380 = n41378 & n41379;
  assign n41381 = n41380 ^ n38623;
  assign n41373 = n41130 ^ n41126;
  assign n41374 = n41260 ^ n41126;
  assign n41375 = ~n41373 & n41374;
  assign n41376 = n41375 ^ n41130;
  assign n41372 = n40796 ^ n40738;
  assign n41377 = n41376 ^ n41372;
  assign n41382 = n41381 ^ n41377;
  assign n41383 = n41382 ^ n37917;
  assign n41387 = n41386 ^ n41383;
  assign n41371 = n41340 & ~n41370;
  assign n41426 = n41387 ^ n41371;
  assign n41430 = n41429 ^ n41426;
  assign n41561 = n41541 ^ n41430;
  assign n41566 = n41565 ^ n41561;
  assign n41598 = n41581 ^ n41566;
  assign n41599 = n41598 ^ n38726;
  assign n41619 = n41607 ^ n41599;
  assign n2291 = n2254 ^ n2203;
  assign n2292 = n2291 ^ n2288;
  assign n2299 = n2298 ^ n2292;
  assign n41695 = n41619 ^ n2299;
  assign n41751 = n41705 ^ n41695;
  assign n41644 = n41051 ^ n41041;
  assign n43667 = n41751 ^ n41644;
  assign n42527 = n40828 ^ n32743;
  assign n42528 = n42527 ^ n1979;
  assign n42529 = n42528 ^ n30971;
  assign n42291 = n39930 ^ n31788;
  assign n42292 = n42291 ^ n36297;
  assign n42293 = n42292 ^ n1689;
  assign n41797 = n40707 ^ n39899;
  assign n41798 = n41372 ^ n40707;
  assign n41799 = ~n41797 & ~n41798;
  assign n41800 = n41799 ^ n39899;
  assign n41796 = n41510 ^ n41507;
  assign n41801 = n41800 ^ n41796;
  assign n41803 = n40584 ^ n39706;
  assign n41804 = n41126 ^ n40584;
  assign n41805 = ~n41803 & ~n41804;
  assign n41806 = n41805 ^ n39706;
  assign n41802 = n41503 ^ n41468;
  assign n41807 = n41806 ^ n41802;
  assign n41921 = n41500 ^ n41473;
  assign n41812 = n41497 ^ n41494;
  assign n41808 = n40466 ^ n39498;
  assign n41809 = n41137 ^ n40466;
  assign n41810 = ~n41808 & n41809;
  assign n41811 = n41810 ^ n39498;
  assign n41813 = n41812 ^ n41811;
  assign n41815 = n40472 ^ n39504;
  assign n41816 = n41143 ^ n40472;
  assign n41817 = ~n41815 & n41816;
  assign n41818 = n41817 ^ n39504;
  assign n41814 = n41490 ^ n41479;
  assign n41819 = n41818 ^ n41814;
  assign n41824 = n41487 ^ n41484;
  assign n41820 = n40478 ^ n39510;
  assign n41821 = n41149 ^ n40478;
  assign n41822 = ~n41820 & n41821;
  assign n41823 = n41822 ^ n39510;
  assign n41825 = n41824 ^ n41823;
  assign n41826 = n40484 ^ n39516;
  assign n41827 = n41155 ^ n40484;
  assign n41828 = ~n41826 & ~n41827;
  assign n41829 = n41828 ^ n39516;
  assign n41115 = n41114 ^ n41093;
  assign n41830 = n41829 ^ n41115;
  assign n41831 = n40490 ^ n39522;
  assign n41832 = n41161 ^ n40490;
  assign n41833 = ~n41831 & ~n41832;
  assign n41834 = n41833 ^ n39522;
  assign n41731 = n41090 ^ n41087;
  assign n41835 = n41834 ^ n41731;
  assign n41836 = n40496 ^ n39528;
  assign n41837 = n41168 ^ n40496;
  assign n41838 = ~n41836 & n41837;
  assign n41839 = n41838 ^ n39528;
  assign n41736 = n41083 ^ n848;
  assign n41840 = n41839 ^ n41736;
  assign n41841 = n40498 ^ n39675;
  assign n41842 = n40498 ^ n40423;
  assign n41843 = ~n41841 & n41842;
  assign n41844 = n41843 ^ n39675;
  assign n41741 = n41079 ^ n41006;
  assign n41845 = n41844 ^ n41741;
  assign n41850 = n41076 ^ n41011;
  assign n41846 = n40504 ^ n39666;
  assign n41847 = n41183 ^ n40504;
  assign n41848 = ~n41846 & n41847;
  assign n41849 = n41848 ^ n39666;
  assign n41851 = n41850 ^ n41849;
  assign n41852 = n40424 ^ n39538;
  assign n41853 = n41189 ^ n40424;
  assign n41854 = ~n41852 & ~n41853;
  assign n41855 = n41854 ^ n39538;
  assign n41747 = n41073 ^ n41070;
  assign n41856 = n41855 ^ n41747;
  assign n41857 = n40515 ^ n39544;
  assign n41858 = n41195 ^ n40515;
  assign n41859 = n41857 & n41858;
  assign n41860 = n41859 ^ n39544;
  assign n41753 = n41066 ^ n41017;
  assign n41861 = n41860 ^ n41753;
  assign n41862 = n40521 ^ n39550;
  assign n41863 = n41201 ^ n40521;
  assign n41864 = ~n41862 & n41863;
  assign n41865 = n41864 ^ n39550;
  assign n41756 = n41063 ^ n41022;
  assign n41866 = n41865 ^ n41756;
  assign n41867 = n40527 ^ n39556;
  assign n41868 = n41207 ^ n40527;
  assign n41869 = n41867 & ~n41868;
  assign n41870 = n41869 ^ n39556;
  assign n41762 = n41060 ^ n41027;
  assign n41871 = n41870 ^ n41762;
  assign n41876 = n41057 ^ n41032;
  assign n41872 = n40533 ^ n39562;
  assign n41873 = n41213 ^ n40533;
  assign n41874 = n41872 & ~n41873;
  assign n41875 = n41874 ^ n39562;
  assign n41877 = n41876 ^ n41875;
  assign n41668 = n41054 ^ n41036;
  assign n41669 = n41668 ^ n41033;
  assign n41663 = n40411 ^ n38844;
  assign n41664 = n41109 ^ n40411;
  assign n41665 = ~n41663 & n41664;
  assign n41666 = n41665 ^ n38844;
  assign n41878 = n41669 ^ n41666;
  assign n41640 = n40286 ^ n39454;
  assign n41641 = n40971 ^ n40286;
  assign n41642 = ~n41640 & ~n41641;
  assign n41643 = n41642 ^ n39454;
  assign n41645 = n41644 ^ n41643;
  assign n41625 = n40248 ^ n39461;
  assign n41626 = n40901 ^ n40248;
  assign n41627 = n41625 & ~n41626;
  assign n41628 = n41627 ^ n39461;
  assign n41624 = n41048 ^ n41047;
  assign n41646 = n41628 ^ n41624;
  assign n41124 = n41045 ^ n41044;
  assign n41120 = n40239 ^ n39468;
  assign n41121 = n40426 ^ n40239;
  assign n41122 = n41120 & ~n41121;
  assign n41123 = n41122 ^ n39468;
  assign n41125 = n41124 ^ n41123;
  assign n41550 = n40168 ^ n39475;
  assign n41551 = n40432 ^ n40168;
  assign n41552 = ~n41550 & n41551;
  assign n41553 = n41552 ^ n39475;
  assign n41422 = n39202 ^ n1867;
  assign n41423 = n41422 ^ n35452;
  assign n41424 = n41423 ^ n2002;
  assign n41400 = n41386 ^ n41382;
  assign n41401 = ~n41383 & ~n41400;
  assign n41402 = n41401 ^ n37917;
  assign n41394 = n39437 ^ n38178;
  assign n41395 = n40114 ^ n39437;
  assign n41396 = n41394 & ~n41395;
  assign n41397 = n41396 ^ n38178;
  assign n41390 = n41381 ^ n41372;
  assign n41391 = ~n41377 & ~n41390;
  assign n41392 = n41391 ^ n41381;
  assign n41389 = n40803 ^ n40800;
  assign n41393 = n41392 ^ n41389;
  assign n41398 = n41397 ^ n41393;
  assign n41399 = n41398 ^ n37291;
  assign n41403 = n41402 ^ n41399;
  assign n41388 = n41371 & ~n41387;
  assign n41421 = n41403 ^ n41388;
  assign n41425 = n41424 ^ n41421;
  assign n41542 = n41541 ^ n41426;
  assign n41543 = ~n41430 & n41542;
  assign n41544 = n41543 ^ n41429;
  assign n41545 = n41544 ^ n41421;
  assign n41546 = n41425 & ~n41545;
  assign n41547 = n41546 ^ n41424;
  assign n1981 = n1978 ^ n1932;
  assign n2006 = n2005 ^ n1981;
  assign n2013 = n2012 ^ n2006;
  assign n41548 = n41547 ^ n2013;
  assign n41415 = n41402 ^ n41398;
  assign n41416 = ~n41399 & n41415;
  assign n41417 = n41416 ^ n37291;
  assign n41418 = n41417 ^ n37284;
  assign n41410 = n41397 ^ n41389;
  assign n41411 = n41393 & n41410;
  assign n41412 = n41411 ^ n41397;
  assign n41406 = n39612 ^ n38172;
  assign n41407 = n40104 ^ n39612;
  assign n41408 = ~n41406 & ~n41407;
  assign n41409 = n41408 ^ n38172;
  assign n41413 = n41412 ^ n41409;
  assign n41405 = n40806 ^ n40732;
  assign n41414 = n41413 ^ n41405;
  assign n41419 = n41418 ^ n41414;
  assign n41404 = n41388 & n41403;
  assign n41420 = n41419 ^ n41404;
  assign n41549 = n41548 ^ n41420;
  assign n41554 = n41553 ^ n41549;
  assign n41559 = n41544 ^ n41425;
  assign n41555 = n39483 ^ n39451;
  assign n41556 = n40438 ^ n39451;
  assign n41557 = ~n41555 & ~n41556;
  assign n41558 = n41557 ^ n39483;
  assign n41560 = n41559 ^ n41558;
  assign n41582 = n41581 ^ n41561;
  assign n41583 = n41566 & n41582;
  assign n41584 = n41583 ^ n41565;
  assign n41585 = n41584 ^ n41559;
  assign n41586 = n41560 & n41585;
  assign n41587 = n41586 ^ n41558;
  assign n41588 = n41587 ^ n41549;
  assign n41589 = n41554 & ~n41588;
  assign n41590 = n41589 ^ n41553;
  assign n41629 = n41590 ^ n41124;
  assign n41630 = n41125 & ~n41629;
  assign n41631 = n41630 ^ n41123;
  assign n41647 = n41631 ^ n41624;
  assign n41648 = n41646 & ~n41647;
  assign n41649 = n41648 ^ n41628;
  assign n41660 = n41649 ^ n41644;
  assign n41661 = n41645 & ~n41660;
  assign n41662 = n41661 ^ n41643;
  assign n41879 = n41669 ^ n41662;
  assign n41880 = n41878 & n41879;
  assign n41881 = n41880 ^ n41666;
  assign n41882 = n41881 ^ n41876;
  assign n41883 = n41877 & n41882;
  assign n41884 = n41883 ^ n41875;
  assign n41885 = n41884 ^ n41762;
  assign n41886 = n41871 & ~n41885;
  assign n41887 = n41886 ^ n41870;
  assign n41888 = n41887 ^ n41756;
  assign n41889 = ~n41866 & n41888;
  assign n41890 = n41889 ^ n41865;
  assign n41891 = n41890 ^ n41753;
  assign n41892 = ~n41861 & n41891;
  assign n41893 = n41892 ^ n41860;
  assign n41894 = n41893 ^ n41747;
  assign n41895 = ~n41856 & n41894;
  assign n41896 = n41895 ^ n41855;
  assign n41897 = n41896 ^ n41850;
  assign n41898 = n41851 & n41897;
  assign n41899 = n41898 ^ n41849;
  assign n41900 = n41899 ^ n41741;
  assign n41901 = n41845 & n41900;
  assign n41902 = n41901 ^ n41844;
  assign n41903 = n41902 ^ n41736;
  assign n41904 = n41840 & ~n41903;
  assign n41905 = n41904 ^ n41839;
  assign n41906 = n41905 ^ n41731;
  assign n41907 = ~n41835 & ~n41906;
  assign n41908 = n41907 ^ n41834;
  assign n41909 = n41908 ^ n41115;
  assign n41910 = n41830 & ~n41909;
  assign n41911 = n41910 ^ n41829;
  assign n41912 = n41911 ^ n41824;
  assign n41913 = ~n41825 & ~n41912;
  assign n41914 = n41913 ^ n41823;
  assign n41915 = n41914 ^ n41814;
  assign n41916 = ~n41819 & n41915;
  assign n41917 = n41916 ^ n41818;
  assign n41918 = n41917 ^ n41812;
  assign n41919 = n41813 & ~n41918;
  assign n41920 = n41919 ^ n41811;
  assign n41922 = n41921 ^ n41920;
  assign n41923 = n40456 ^ n39492;
  assign n41924 = n41135 ^ n40456;
  assign n41925 = ~n41923 & n41924;
  assign n41926 = n41925 ^ n39492;
  assign n41927 = n41926 ^ n41921;
  assign n41928 = n41922 & ~n41927;
  assign n41929 = n41928 ^ n41926;
  assign n41930 = n41929 ^ n41802;
  assign n41931 = ~n41807 & ~n41930;
  assign n41932 = n41931 ^ n41806;
  assign n41933 = n41932 ^ n41796;
  assign n41934 = n41801 & n41933;
  assign n41935 = n41934 ^ n41800;
  assign n41791 = n40128 ^ n39358;
  assign n41792 = n41389 ^ n40128;
  assign n41793 = ~n41791 & n41792;
  assign n41794 = n41793 ^ n39358;
  assign n41970 = n41935 ^ n41794;
  assign n41790 = n41513 ^ n41462;
  assign n41971 = n41970 ^ n41790;
  assign n41972 = n41971 ^ n38647;
  assign n41973 = n41932 ^ n41800;
  assign n41974 = n41973 ^ n41796;
  assign n41975 = n41974 ^ n39181;
  assign n41976 = n41929 ^ n41806;
  assign n41977 = n41976 ^ n41802;
  assign n41978 = n41977 ^ n38848;
  assign n41979 = n41926 ^ n41922;
  assign n41980 = n41979 ^ n38849;
  assign n41981 = n41917 ^ n41811;
  assign n41982 = n41981 ^ n41812;
  assign n41983 = n41982 ^ n38859;
  assign n41984 = n41914 ^ n41818;
  assign n41985 = n41984 ^ n41814;
  assign n41986 = n41985 ^ n38865;
  assign n41987 = n41911 ^ n41825;
  assign n41988 = n41987 ^ n38871;
  assign n41989 = n41908 ^ n41830;
  assign n41990 = n41989 ^ n39002;
  assign n41991 = n41905 ^ n41835;
  assign n41992 = n41991 ^ n38873;
  assign n41993 = n41902 ^ n41839;
  assign n41994 = n41993 ^ n41736;
  assign n41995 = n41994 ^ n38883;
  assign n41996 = n41899 ^ n41845;
  assign n41997 = n41996 ^ n38889;
  assign n41998 = n41896 ^ n41851;
  assign n41999 = n41998 ^ n38895;
  assign n42000 = n41893 ^ n41856;
  assign n42001 = n42000 ^ n38901;
  assign n42002 = n41890 ^ n41860;
  assign n42003 = n42002 ^ n41753;
  assign n42004 = n42003 ^ n38907;
  assign n42005 = n41887 ^ n41865;
  assign n42006 = n42005 ^ n41756;
  assign n42007 = n42006 ^ n38913;
  assign n42008 = n41884 ^ n41870;
  assign n42009 = n42008 ^ n41762;
  assign n42010 = n42009 ^ n38163;
  assign n42011 = n41881 ^ n41875;
  assign n42012 = n42011 ^ n41876;
  assign n42013 = n42012 ^ n38924;
  assign n41667 = n41666 ^ n41662;
  assign n41670 = n41669 ^ n41667;
  assign n41671 = n41670 ^ n38930;
  assign n41650 = n41649 ^ n41645;
  assign n41651 = n41650 ^ n38936;
  assign n41632 = n41631 ^ n41628;
  assign n41633 = n41632 ^ n41624;
  assign n41634 = n41633 ^ n38942;
  assign n41591 = n41590 ^ n41125;
  assign n41592 = n41591 ^ n38948;
  assign n41593 = n41587 ^ n41554;
  assign n41594 = n41593 ^ n38954;
  assign n41595 = n41584 ^ n41558;
  assign n41596 = n41595 ^ n41559;
  assign n41597 = n41596 ^ n38830;
  assign n41608 = n41607 ^ n41598;
  assign n41609 = n41599 & ~n41608;
  assign n41610 = n41609 ^ n38726;
  assign n41611 = n41610 ^ n41596;
  assign n41612 = n41597 & n41611;
  assign n41613 = n41612 ^ n38830;
  assign n41614 = n41613 ^ n41593;
  assign n41615 = ~n41594 & n41614;
  assign n41616 = n41615 ^ n38954;
  assign n41635 = n41616 ^ n41591;
  assign n41636 = n41592 & n41635;
  assign n41637 = n41636 ^ n38948;
  assign n41652 = n41637 ^ n41633;
  assign n41653 = ~n41634 & ~n41652;
  assign n41654 = n41653 ^ n38942;
  assign n41657 = n41654 ^ n41650;
  assign n41658 = n41651 & n41657;
  assign n41659 = n41658 ^ n38936;
  assign n42014 = n41670 ^ n41659;
  assign n42015 = ~n41671 & ~n42014;
  assign n42016 = n42015 ^ n38930;
  assign n42017 = n42016 ^ n42012;
  assign n42018 = ~n42013 & ~n42017;
  assign n42019 = n42018 ^ n38924;
  assign n42020 = n42019 ^ n42009;
  assign n42021 = n42010 & ~n42020;
  assign n42022 = n42021 ^ n38163;
  assign n42023 = n42022 ^ n42006;
  assign n42024 = n42007 & n42023;
  assign n42025 = n42024 ^ n38913;
  assign n42026 = n42025 ^ n42003;
  assign n42027 = n42004 & ~n42026;
  assign n42028 = n42027 ^ n38907;
  assign n42029 = n42028 ^ n42000;
  assign n42030 = n42001 & ~n42029;
  assign n42031 = n42030 ^ n38901;
  assign n42032 = n42031 ^ n41998;
  assign n42033 = n41999 & n42032;
  assign n42034 = n42033 ^ n38895;
  assign n42035 = n42034 ^ n41996;
  assign n42036 = ~n41997 & n42035;
  assign n42037 = n42036 ^ n38889;
  assign n42038 = n42037 ^ n41994;
  assign n42039 = n41995 & ~n42038;
  assign n42040 = n42039 ^ n38883;
  assign n42041 = n42040 ^ n41991;
  assign n42042 = ~n41992 & n42041;
  assign n42043 = n42042 ^ n38873;
  assign n42044 = n42043 ^ n41989;
  assign n42045 = ~n41990 & n42044;
  assign n42046 = n42045 ^ n39002;
  assign n42047 = n42046 ^ n41987;
  assign n42048 = n41988 & ~n42047;
  assign n42049 = n42048 ^ n38871;
  assign n42050 = n42049 ^ n41985;
  assign n42051 = n41986 & n42050;
  assign n42052 = n42051 ^ n38865;
  assign n42053 = n42052 ^ n41982;
  assign n42054 = n41983 & n42053;
  assign n42055 = n42054 ^ n38859;
  assign n42056 = n42055 ^ n41979;
  assign n42057 = n41980 & n42056;
  assign n42058 = n42057 ^ n38849;
  assign n42059 = n42058 ^ n41977;
  assign n42060 = n41978 & ~n42059;
  assign n42061 = n42060 ^ n38848;
  assign n42062 = n42061 ^ n41974;
  assign n42063 = n41975 & ~n42062;
  assign n42064 = n42063 ^ n39181;
  assign n42065 = n42064 ^ n41971;
  assign n42066 = n41972 & n42065;
  assign n42067 = n42066 ^ n38647;
  assign n41795 = n41794 ^ n41790;
  assign n41936 = n41935 ^ n41790;
  assign n41937 = n41795 & n41936;
  assign n41938 = n41937 ^ n41794;
  assign n41784 = n40122 ^ n39369;
  assign n41785 = n41405 ^ n40122;
  assign n41786 = n41784 & n41785;
  assign n41787 = n41786 ^ n39369;
  assign n41967 = n41938 ^ n41787;
  assign n41788 = n41516 ^ n41457;
  assign n41968 = n41967 ^ n41788;
  assign n41969 = n41968 ^ n38641;
  assign n42118 = n42067 ^ n41969;
  assign n42081 = n42064 ^ n41972;
  assign n42082 = n42061 ^ n41975;
  assign n42083 = n42058 ^ n38848;
  assign n42084 = n42083 ^ n41977;
  assign n42085 = n42055 ^ n38849;
  assign n42086 = n42085 ^ n41979;
  assign n42087 = n42052 ^ n41983;
  assign n42088 = n42049 ^ n41986;
  assign n42089 = n42046 ^ n41988;
  assign n42090 = n42040 ^ n41992;
  assign n42091 = n42037 ^ n41995;
  assign n42092 = n42025 ^ n42004;
  assign n42093 = n42019 ^ n42010;
  assign n41617 = n41616 ^ n41592;
  assign n41618 = n41613 ^ n41594;
  assign n41620 = n41610 ^ n41597;
  assign n41621 = ~n41619 & ~n41620;
  assign n41622 = ~n41618 & n41621;
  assign n41623 = ~n41617 & ~n41622;
  assign n41638 = n41637 ^ n41634;
  assign n41639 = ~n41623 & n41638;
  assign n41655 = n41654 ^ n41651;
  assign n41656 = n41639 & n41655;
  assign n41672 = n41671 ^ n41659;
  assign n42094 = ~n41656 & ~n41672;
  assign n42095 = n42016 ^ n42013;
  assign n42096 = n42094 & n42095;
  assign n42097 = ~n42093 & ~n42096;
  assign n42098 = n42022 ^ n42007;
  assign n42099 = n42097 & ~n42098;
  assign n42100 = n42092 & n42099;
  assign n42101 = n42028 ^ n42001;
  assign n42102 = n42100 & n42101;
  assign n42103 = n42031 ^ n41999;
  assign n42104 = ~n42102 & ~n42103;
  assign n42105 = n42034 ^ n41997;
  assign n42106 = ~n42104 & n42105;
  assign n42107 = ~n42091 & n42106;
  assign n42108 = n42090 & n42107;
  assign n42109 = n42043 ^ n41990;
  assign n42110 = ~n42108 & ~n42109;
  assign n42111 = ~n42089 & ~n42110;
  assign n42112 = ~n42088 & n42111;
  assign n42113 = ~n42087 & ~n42112;
  assign n42114 = n42086 & n42113;
  assign n42115 = ~n42084 & n42114;
  assign n42116 = n42082 & ~n42115;
  assign n42117 = n42081 & n42116;
  assign n42155 = n42118 ^ n42117;
  assign n3005 = n2938 ^ n1613;
  assign n3006 = n3005 ^ n3002;
  assign n3010 = n3009 ^ n3006;
  assign n42156 = n42155 ^ n3010;
  assign n42161 = n42115 ^ n42082;
  assign n42158 = n3237 ^ n2861;
  assign n42159 = n42158 ^ n36307;
  assign n42160 = n42159 ^ n2984;
  assign n42162 = n42161 ^ n42160;
  assign n42163 = n42114 ^ n42084;
  assign n42167 = n42166 ^ n42163;
  assign n42171 = n42113 ^ n42086;
  assign n42168 = n39944 ^ n3223;
  assign n42169 = n42168 ^ n36317;
  assign n42170 = n42169 ^ n3089;
  assign n42172 = n42171 ^ n42170;
  assign n42176 = n42112 ^ n42087;
  assign n42173 = n40060 ^ n31345;
  assign n42174 = n42173 ^ n3071;
  assign n42175 = n42174 ^ n2588;
  assign n42177 = n42176 ^ n42175;
  assign n42181 = n42111 ^ n42088;
  assign n42178 = n39950 ^ n31350;
  assign n42179 = n42178 ^ n2531;
  assign n42180 = n42179 ^ n3069;
  assign n42182 = n42181 ^ n42180;
  assign n42186 = n42110 ^ n42089;
  assign n42183 = n40050 ^ n3047;
  assign n42184 = n42183 ^ n36325;
  assign n42185 = n42184 ^ n2523;
  assign n42187 = n42186 ^ n42185;
  assign n42190 = n39962 ^ n31358;
  assign n42191 = n42190 ^ n1409;
  assign n42192 = n42191 ^ n30220;
  assign n42189 = n42107 ^ n42090;
  assign n42193 = n42192 ^ n42189;
  assign n42195 = n42105 ^ n42104;
  assign n1194 = n1193 ^ n1124;
  assign n1210 = n1209 ^ n1194;
  assign n1217 = n1216 ^ n1210;
  assign n42196 = n42195 ^ n1217;
  assign n42198 = n42101 ^ n42100;
  assign n1036 = n1026 ^ n984;
  assign n1061 = n1060 ^ n1036;
  assign n1068 = n1067 ^ n1061;
  assign n42199 = n42198 ^ n1068;
  assign n42202 = n39985 ^ n898;
  assign n42203 = n42202 ^ n35830;
  assign n42204 = n42203 ^ n3321;
  assign n42201 = n42098 ^ n42097;
  assign n42205 = n42204 ^ n42201;
  assign n42206 = n42096 ^ n42093;
  assign n42210 = n42209 ^ n42206;
  assign n42212 = n39995 ^ n31384;
  assign n42213 = n42212 ^ n35839;
  assign n42214 = n42213 ^ n30175;
  assign n42211 = n42095 ^ n42094;
  assign n42215 = n42214 ^ n42211;
  assign n41677 = n41655 ^ n41639;
  assign n41674 = n40004 ^ n31394;
  assign n41675 = n41674 ^ n35849;
  assign n41676 = n41675 ^ n714;
  assign n41678 = n41677 ^ n41676;
  assign n41682 = n41638 ^ n41623;
  assign n41679 = n39432 ^ n31398;
  assign n41680 = n41679 ^ n35854;
  assign n41681 = n41680 ^ n29643;
  assign n41683 = n41682 ^ n41681;
  assign n41685 = n39406 ^ n31404;
  assign n41686 = n41685 ^ n35860;
  assign n41687 = n41686 ^ n29670;
  assign n41684 = n41622 ^ n41617;
  assign n41688 = n41687 ^ n41684;
  assign n41690 = n39423 ^ n31409;
  assign n41691 = n41690 ^ n35865;
  assign n41692 = n41691 ^ n29649;
  assign n41689 = n41621 ^ n41618;
  assign n41693 = n41692 ^ n41689;
  assign n41706 = n41705 ^ n41619;
  assign n41707 = ~n41695 & n41706;
  assign n41708 = n41707 ^ n2299;
  assign n41694 = n41620 ^ n41619;
  assign n41709 = n41708 ^ n41694;
  assign n41710 = n31421 ^ n2352;
  assign n41711 = n41710 ^ n35869;
  assign n41712 = n41711 ^ n29660;
  assign n41713 = n41712 ^ n41694;
  assign n41714 = n41709 & ~n41713;
  assign n41715 = n41714 ^ n41712;
  assign n41716 = n41715 ^ n41689;
  assign n41717 = n41693 & ~n41716;
  assign n41718 = n41717 ^ n41692;
  assign n41719 = n41718 ^ n41684;
  assign n41720 = n41688 & ~n41719;
  assign n41721 = n41720 ^ n41687;
  assign n41722 = n41721 ^ n41682;
  assign n41723 = n41683 & ~n41722;
  assign n41724 = n41723 ^ n41681;
  assign n41725 = n41724 ^ n41677;
  assign n41726 = ~n41678 & n41725;
  assign n41727 = n41726 ^ n41676;
  assign n41673 = n41672 ^ n41656;
  assign n41728 = n41727 ^ n41673;
  assign n41117 = n39999 ^ n31389;
  assign n41118 = n41117 ^ n35844;
  assign n41119 = n41118 ^ n30180;
  assign n42216 = n41673 ^ n41119;
  assign n42217 = ~n41728 & n42216;
  assign n42218 = n42217 ^ n41119;
  assign n42219 = n42218 ^ n42211;
  assign n42220 = n42215 & ~n42219;
  assign n42221 = n42220 ^ n42214;
  assign n42222 = n42221 ^ n42206;
  assign n42223 = ~n42210 & n42222;
  assign n42224 = n42223 ^ n42209;
  assign n42225 = n42224 ^ n42201;
  assign n42226 = n42205 & ~n42225;
  assign n42227 = n42226 ^ n42204;
  assign n42200 = n42099 ^ n42092;
  assign n42228 = n42227 ^ n42200;
  assign n42232 = n42231 ^ n42200;
  assign n42233 = n42228 & ~n42232;
  assign n42234 = n42233 ^ n42231;
  assign n42235 = n42234 ^ n42198;
  assign n42236 = ~n42199 & n42235;
  assign n42237 = n42236 ^ n1068;
  assign n42197 = n42103 ^ n42102;
  assign n42238 = n42237 ^ n42197;
  assign n42239 = n39973 ^ n31371;
  assign n42240 = n42239 ^ n1078;
  assign n42241 = n42240 ^ n1201;
  assign n42242 = n42241 ^ n42197;
  assign n42243 = ~n42238 & n42242;
  assign n42244 = n42243 ^ n42241;
  assign n42245 = n42244 ^ n42195;
  assign n42246 = n42196 & ~n42245;
  assign n42247 = n42246 ^ n1217;
  assign n42194 = n42106 ^ n42091;
  assign n42248 = n42247 ^ n42194;
  assign n42249 = n39967 ^ n31364;
  assign n42250 = n42249 ^ n36337;
  assign n42251 = n42250 ^ n1401;
  assign n42252 = n42251 ^ n42194;
  assign n42253 = ~n42248 & n42252;
  assign n42254 = n42253 ^ n42251;
  assign n42255 = n42254 ^ n42189;
  assign n42256 = ~n42193 & n42255;
  assign n42257 = n42256 ^ n42192;
  assign n42188 = n42109 ^ n42108;
  assign n42258 = n42257 ^ n42188;
  assign n42259 = n39956 ^ n2453;
  assign n42260 = n42259 ^ n36331;
  assign n42261 = n42260 ^ n3155;
  assign n42262 = n42261 ^ n42188;
  assign n42263 = ~n42258 & n42262;
  assign n42264 = n42263 ^ n42261;
  assign n42265 = n42264 ^ n42186;
  assign n42266 = ~n42187 & n42265;
  assign n42267 = n42266 ^ n42185;
  assign n42268 = n42267 ^ n42181;
  assign n42269 = n42182 & ~n42268;
  assign n42270 = n42269 ^ n42180;
  assign n42271 = n42270 ^ n42176;
  assign n42272 = n42177 & ~n42271;
  assign n42273 = n42272 ^ n42175;
  assign n42274 = n42273 ^ n42171;
  assign n42275 = n42172 & ~n42274;
  assign n42276 = n42275 ^ n42170;
  assign n42277 = n42276 ^ n42163;
  assign n42278 = ~n42167 & n42277;
  assign n42279 = n42278 ^ n42166;
  assign n42280 = n42279 ^ n42161;
  assign n42281 = n42162 & ~n42280;
  assign n42282 = n42281 ^ n42160;
  assign n42157 = n42116 ^ n42081;
  assign n42283 = n42282 ^ n42157;
  assign n2969 = n2962 ^ n2922;
  assign n2988 = n2987 ^ n2969;
  assign n2995 = n2994 ^ n2988;
  assign n42284 = n42157 ^ n2995;
  assign n42285 = n42283 & ~n42284;
  assign n42286 = n42285 ^ n2995;
  assign n42287 = n42286 ^ n3010;
  assign n42288 = ~n42156 & ~n42287;
  assign n42289 = n42288 ^ n42155;
  assign n42068 = n42067 ^ n41968;
  assign n42069 = ~n41969 & ~n42068;
  assign n42070 = n42069 ^ n38641;
  assign n41789 = n41788 ^ n41787;
  assign n41939 = n41938 ^ n41788;
  assign n41940 = ~n41789 & ~n41939;
  assign n41941 = n41940 ^ n41787;
  assign n41778 = n40116 ^ n39352;
  assign n41779 = n40858 ^ n40116;
  assign n41780 = ~n41778 & n41779;
  assign n41781 = n41780 ^ n39352;
  assign n41964 = n41941 ^ n41781;
  assign n41782 = n41519 ^ n41452;
  assign n41965 = n41964 ^ n41782;
  assign n41966 = n41965 ^ n38635;
  assign n42120 = n42070 ^ n41966;
  assign n42119 = n42117 & n42118;
  assign n42154 = n42120 ^ n42119;
  assign n42290 = n42289 ^ n42154;
  assign n42322 = n42293 ^ n42290;
  assign n42320 = n40878 ^ n39472;
  assign n42321 = n42320 ^ n41124;
  assign n42397 = n42322 ^ n42321;
  assign n42526 = n42397 ^ n39606;
  assign n42637 = n42529 ^ n42526;
  assign n43668 = n43667 ^ n42637;
  assign n43481 = n33156 ^ n3135;
  assign n43482 = n43481 ^ n2869;
  assign n43483 = n43482 ^ n2962;
  assign n42446 = n42218 ^ n42215;
  assign n42444 = n41168 ^ n40504;
  assign n42445 = n42444 ^ n41824;
  assign n42447 = n42446 ^ n42445;
  assign n41733 = n41724 ^ n41678;
  assign n41730 = n41183 ^ n40515;
  assign n41732 = n41731 ^ n41730;
  assign n41734 = n41733 ^ n41732;
  assign n41738 = n41721 ^ n41683;
  assign n41735 = n41189 ^ n40521;
  assign n41737 = n41736 ^ n41735;
  assign n41739 = n41738 ^ n41737;
  assign n41743 = n41718 ^ n41688;
  assign n41740 = n41195 ^ n40527;
  assign n41742 = n41741 ^ n41740;
  assign n41744 = n41743 ^ n41742;
  assign n41749 = n41712 ^ n41709;
  assign n41746 = n41207 ^ n40411;
  assign n41748 = n41747 ^ n41746;
  assign n41750 = n41749 ^ n41748;
  assign n41752 = n41213 ^ n40286;
  assign n41754 = n41753 ^ n41752;
  assign n41755 = n41754 ^ n41751;
  assign n41759 = n41702 ^ n41701;
  assign n41757 = n41756 ^ n41109;
  assign n41758 = n41757 ^ n40248;
  assign n41760 = n41759 ^ n41758;
  assign n41764 = n41699 ^ n41698;
  assign n41761 = n40971 ^ n40239;
  assign n41763 = n41762 ^ n41761;
  assign n41765 = n41764 ^ n41763;
  assign n42316 = n40426 ^ n39451;
  assign n42317 = n42316 ^ n41669;
  assign n41783 = n41782 ^ n41781;
  assign n41942 = n41941 ^ n41782;
  assign n41943 = n41783 & ~n41942;
  assign n41944 = n41943 ^ n41781;
  assign n41773 = n40114 ^ n39346;
  assign n41774 = n40848 ^ n40114;
  assign n41775 = n41773 & n41774;
  assign n41776 = n41775 ^ n39346;
  assign n41961 = n41944 ^ n41776;
  assign n41772 = n41522 ^ n41450;
  assign n41962 = n41961 ^ n41772;
  assign n41963 = n41962 ^ n38629;
  assign n42071 = n42070 ^ n41965;
  assign n42072 = ~n41966 & n42071;
  assign n42073 = n42072 ^ n38635;
  assign n42074 = n42073 ^ n41962;
  assign n42075 = ~n41963 & n42074;
  assign n42076 = n42075 ^ n38629;
  assign n41777 = n41776 ^ n41772;
  assign n41945 = n41944 ^ n41772;
  assign n41946 = n41777 & n41945;
  assign n41947 = n41946 ^ n41776;
  assign n41770 = n41525 ^ n41448;
  assign n41766 = n40104 ^ n39340;
  assign n41767 = n40842 ^ n40104;
  assign n41768 = ~n41766 & n41767;
  assign n41769 = n41768 ^ n39340;
  assign n41771 = n41770 ^ n41769;
  assign n41959 = n41947 ^ n41771;
  assign n41960 = n41959 ^ n38623;
  assign n42124 = n42076 ^ n41960;
  assign n42121 = n42119 & ~n42120;
  assign n42122 = n42073 ^ n41963;
  assign n42123 = ~n42121 & n42122;
  assign n42151 = n42124 ^ n42123;
  assign n42148 = n39925 ^ n31778;
  assign n42149 = n42148 ^ n36290;
  assign n42150 = n42149 ^ n1766;
  assign n42152 = n42151 ^ n42150;
  assign n42294 = n42293 ^ n42154;
  assign n42295 = n42290 & n42294;
  assign n42296 = n42295 ^ n42293;
  assign n42153 = n42122 ^ n42121;
  assign n42297 = n42296 ^ n42153;
  assign n42298 = n40087 ^ n31783;
  assign n42299 = n42298 ^ n1697;
  assign n42300 = n42299 ^ n30136;
  assign n42301 = n42300 ^ n42153;
  assign n42302 = n42297 & ~n42301;
  assign n42303 = n42302 ^ n42300;
  assign n42304 = n42303 ^ n42151;
  assign n42305 = n42152 & ~n42304;
  assign n42306 = n42305 ^ n42150;
  assign n42144 = n39920 ^ n31773;
  assign n42145 = n42144 ^ n36285;
  assign n42146 = n42145 ^ n30130;
  assign n42125 = n42123 & n42124;
  assign n42077 = n42076 ^ n41959;
  assign n42078 = ~n41960 & ~n42077;
  assign n42079 = n42078 ^ n38623;
  assign n41953 = n39481 ^ n39437;
  assign n41954 = n40836 ^ n39481;
  assign n41955 = n41953 & n41954;
  assign n41956 = n41955 ^ n39437;
  assign n41951 = n41529 ^ n2894;
  assign n41948 = n41947 ^ n41770;
  assign n41949 = n41771 & n41948;
  assign n41950 = n41949 ^ n41769;
  assign n41952 = n41951 ^ n41950;
  assign n41957 = n41956 ^ n41952;
  assign n41958 = n41957 ^ n38178;
  assign n42080 = n42079 ^ n41958;
  assign n42143 = n42125 ^ n42080;
  assign n42147 = n42146 ^ n42143;
  assign n42315 = n42306 ^ n42147;
  assign n42318 = n42317 ^ n42315;
  assign n42324 = n40438 ^ n39465;
  assign n42325 = n42324 ^ n41624;
  assign n42323 = ~n42321 & ~n42322;
  assign n42326 = n42325 ^ n42323;
  assign n42327 = n42300 ^ n42297;
  assign n42328 = n42327 ^ n42325;
  assign n42329 = n42326 & n42328;
  assign n42330 = n42329 ^ n42323;
  assign n42319 = n42303 ^ n42152;
  assign n42331 = n42330 ^ n42319;
  assign n42332 = n40432 ^ n39458;
  assign n42333 = n42332 ^ n41644;
  assign n42334 = n42333 ^ n42319;
  assign n42335 = ~n42331 & ~n42334;
  assign n42336 = n42335 ^ n42333;
  assign n42337 = n42336 ^ n42315;
  assign n42338 = ~n42318 & ~n42337;
  assign n42339 = n42338 ^ n42317;
  assign n42307 = n42306 ^ n42143;
  assign n42308 = ~n42147 & n42307;
  assign n42309 = n42308 ^ n42146;
  assign n42313 = n42312 ^ n42309;
  assign n42137 = n42079 ^ n41957;
  assign n42138 = ~n41958 & ~n42137;
  assign n42139 = n42138 ^ n38178;
  assign n42140 = n42139 ^ n38172;
  assign n42135 = n41532 ^ n41445;
  assign n42131 = n41956 ^ n41951;
  assign n42132 = n41952 & n42131;
  assign n42133 = n42132 ^ n41956;
  assign n42127 = n39612 ^ n39479;
  assign n42128 = n40830 ^ n39479;
  assign n42129 = ~n42127 & ~n42128;
  assign n42130 = n42129 ^ n39612;
  assign n42134 = n42133 ^ n42130;
  assign n42136 = n42135 ^ n42134;
  assign n42141 = n42140 ^ n42136;
  assign n42126 = ~n42080 & n42125;
  assign n42142 = n42141 ^ n42126;
  assign n42314 = n42313 ^ n42142;
  assign n42340 = n42339 ^ n42314;
  assign n42341 = n40901 ^ n40168;
  assign n42342 = n42341 ^ n41876;
  assign n42343 = n42342 ^ n42314;
  assign n42344 = n42340 & n42343;
  assign n42345 = n42344 ^ n42342;
  assign n42346 = n42345 ^ n41764;
  assign n42347 = ~n41765 & n42346;
  assign n42348 = n42347 ^ n41763;
  assign n42349 = n42348 ^ n41759;
  assign n42350 = ~n41760 & ~n42349;
  assign n42351 = n42350 ^ n41758;
  assign n42352 = n42351 ^ n41751;
  assign n42353 = ~n41755 & n42352;
  assign n42354 = n42353 ^ n41754;
  assign n42355 = n42354 ^ n41749;
  assign n42356 = n41750 & n42355;
  assign n42357 = n42356 ^ n41748;
  assign n41745 = n41715 ^ n41693;
  assign n42358 = n42357 ^ n41745;
  assign n42359 = n41201 ^ n40533;
  assign n42360 = n42359 ^ n41850;
  assign n42361 = n42360 ^ n41745;
  assign n42362 = n42358 & ~n42361;
  assign n42363 = n42362 ^ n42360;
  assign n42364 = n42363 ^ n41743;
  assign n42365 = ~n41744 & n42364;
  assign n42366 = n42365 ^ n41742;
  assign n42367 = n42366 ^ n41738;
  assign n42368 = n41739 & n42367;
  assign n42369 = n42368 ^ n41737;
  assign n42370 = n42369 ^ n41733;
  assign n42371 = n41734 & n42370;
  assign n42372 = n42371 ^ n41732;
  assign n41729 = n41728 ^ n41119;
  assign n42373 = n42372 ^ n41729;
  assign n40425 = n40424 ^ n40423;
  assign n41116 = n41115 ^ n40425;
  assign n42441 = n41729 ^ n41116;
  assign n42442 = n42373 & n42441;
  assign n42443 = n42442 ^ n41116;
  assign n42596 = n42446 ^ n42443;
  assign n42597 = ~n42447 & ~n42596;
  assign n42598 = n42597 ^ n42445;
  assign n42595 = n42221 ^ n42210;
  assign n42599 = n42598 ^ n42595;
  assign n42593 = n41161 ^ n40498;
  assign n42594 = n42593 ^ n41814;
  assign n42600 = n42599 ^ n42594;
  assign n42601 = n42600 ^ n39675;
  assign n42448 = n42447 ^ n42443;
  assign n42449 = n42448 ^ n39666;
  assign n42374 = n42373 ^ n41116;
  assign n42375 = n42374 ^ n39538;
  assign n42376 = n42369 ^ n41734;
  assign n42377 = n42376 ^ n39544;
  assign n42378 = n42366 ^ n41739;
  assign n42379 = n42378 ^ n39550;
  assign n42380 = n42363 ^ n41744;
  assign n42381 = n42380 ^ n39556;
  assign n42382 = n42360 ^ n42358;
  assign n42383 = n42382 ^ n39562;
  assign n42385 = n42351 ^ n41755;
  assign n42386 = n42385 ^ n39454;
  assign n42387 = n42348 ^ n41760;
  assign n42388 = n42387 ^ n39461;
  assign n42389 = n42345 ^ n41765;
  assign n42390 = n42389 ^ n39468;
  assign n42391 = n42342 ^ n42340;
  assign n42392 = n42391 ^ n39475;
  assign n42393 = n42336 ^ n42318;
  assign n42394 = n42393 ^ n39483;
  assign n42395 = n42333 ^ n42331;
  assign n42396 = n42395 ^ n39598;
  assign n42398 = ~n39606 & n42397;
  assign n42399 = n42398 ^ n39604;
  assign n42400 = n42327 ^ n42326;
  assign n42401 = n42400 ^ n42398;
  assign n42402 = n42399 & n42401;
  assign n42403 = n42402 ^ n39604;
  assign n42404 = n42403 ^ n42395;
  assign n42405 = n42396 & n42404;
  assign n42406 = n42405 ^ n39598;
  assign n42407 = n42406 ^ n42393;
  assign n42408 = n42394 & n42407;
  assign n42409 = n42408 ^ n39483;
  assign n42410 = n42409 ^ n42391;
  assign n42411 = n42392 & ~n42410;
  assign n42412 = n42411 ^ n39475;
  assign n42413 = n42412 ^ n42389;
  assign n42414 = n42390 & ~n42413;
  assign n42415 = n42414 ^ n39468;
  assign n42416 = n42415 ^ n42387;
  assign n42417 = n42388 & ~n42416;
  assign n42418 = n42417 ^ n39461;
  assign n42419 = n42418 ^ n42385;
  assign n42420 = ~n42386 & n42419;
  assign n42421 = n42420 ^ n39454;
  assign n42384 = n42354 ^ n41750;
  assign n42422 = n42421 ^ n42384;
  assign n42423 = n42384 ^ n38844;
  assign n42424 = ~n42422 & ~n42423;
  assign n42425 = n42424 ^ n38844;
  assign n42426 = n42425 ^ n42382;
  assign n42427 = n42383 & n42426;
  assign n42428 = n42427 ^ n39562;
  assign n42429 = n42428 ^ n42380;
  assign n42430 = n42381 & ~n42429;
  assign n42431 = n42430 ^ n39556;
  assign n42432 = n42431 ^ n42378;
  assign n42433 = ~n42379 & n42432;
  assign n42434 = n42433 ^ n39550;
  assign n42435 = n42434 ^ n42376;
  assign n42436 = n42377 & ~n42435;
  assign n42437 = n42436 ^ n39544;
  assign n42438 = n42437 ^ n42374;
  assign n42439 = ~n42375 & n42438;
  assign n42440 = n42439 ^ n39538;
  assign n42590 = n42448 ^ n42440;
  assign n42591 = n42449 & n42590;
  assign n42592 = n42591 ^ n39666;
  assign n42602 = n42601 ^ n42592;
  assign n42450 = n42449 ^ n42440;
  assign n42451 = n42437 ^ n42375;
  assign n42452 = n42434 ^ n42377;
  assign n42453 = n42431 ^ n42379;
  assign n42454 = n42422 ^ n38844;
  assign n42455 = n42418 ^ n42386;
  assign n42456 = n42415 ^ n42388;
  assign n42457 = n42412 ^ n42390;
  assign n42458 = n42406 ^ n42394;
  assign n42459 = n42400 ^ n42399;
  assign n42460 = n42403 ^ n42396;
  assign n42461 = n42459 & ~n42460;
  assign n42462 = ~n42458 & ~n42461;
  assign n42463 = n42409 ^ n42392;
  assign n42464 = ~n42462 & ~n42463;
  assign n42465 = n42457 & ~n42464;
  assign n42466 = ~n42456 & ~n42465;
  assign n42467 = n42455 & n42466;
  assign n42468 = n42454 & n42467;
  assign n42469 = n42425 ^ n42383;
  assign n42470 = ~n42468 & ~n42469;
  assign n42471 = n42428 ^ n42381;
  assign n42472 = n42470 & n42471;
  assign n42473 = ~n42453 & n42472;
  assign n42474 = n42452 & n42473;
  assign n42475 = ~n42451 & n42474;
  assign n42589 = ~n42450 & ~n42475;
  assign n42603 = n42602 ^ n42589;
  assign n1328 = n1309 ^ n1246;
  assign n1347 = n1346 ^ n1328;
  assign n1354 = n1353 ^ n1347;
  assign n42604 = n42603 ^ n1354;
  assign n42476 = n42475 ^ n42450;
  assign n3342 = n3341 ^ n1157;
  assign n3349 = n3348 ^ n3342;
  assign n3350 = n3349 ^ n1338;
  assign n42477 = n42476 ^ n3350;
  assign n42478 = n42474 ^ n42451;
  assign n42482 = n42481 ^ n42478;
  assign n42483 = n42473 ^ n42452;
  assign n42487 = n42486 ^ n42483;
  assign n42491 = n42472 ^ n42453;
  assign n42488 = n40306 ^ n32292;
  assign n42489 = n42488 ^ n36616;
  assign n42490 = n42489 ^ n812;
  assign n42492 = n42491 ^ n42490;
  assign n42496 = n42471 ^ n42470;
  assign n42493 = n40311 ^ n32297;
  assign n42494 = n42493 ^ n740;
  assign n42495 = n42494 ^ n30469;
  assign n42497 = n42496 ^ n42495;
  assign n42500 = n40318 ^ n723;
  assign n42501 = n42500 ^ n36547;
  assign n42502 = n42501 ^ n30496;
  assign n42499 = n42467 ^ n42454;
  assign n42503 = n42502 ^ n42499;
  assign n42506 = n40328 ^ n32313;
  assign n42507 = n42506 ^ n36557;
  assign n42508 = n42507 ^ n30506;
  assign n42505 = n42465 ^ n42456;
  assign n42509 = n42508 ^ n42505;
  assign n42514 = n42463 ^ n42462;
  assign n42511 = n40359 ^ n32324;
  assign n42512 = n42511 ^ n36588;
  assign n42513 = n42512 ^ n30534;
  assign n42515 = n42514 ^ n42513;
  assign n42519 = n42461 ^ n42458;
  assign n42516 = n40338 ^ n2406;
  assign n42517 = n42516 ^ n36567;
  assign n42518 = n42517 ^ n30526;
  assign n42520 = n42519 ^ n42518;
  assign n42524 = n42460 ^ n42459;
  assign n42521 = n40342 ^ n2388;
  assign n42522 = n42521 ^ n36571;
  assign n42523 = n42522 ^ n30518;
  assign n42525 = n42524 ^ n42523;
  assign n42531 = n40345 ^ n2380;
  assign n42532 = n42531 ^ n36574;
  assign n42533 = n42532 ^ n2135;
  assign n42530 = ~n42526 & n42529;
  assign n42534 = n42533 ^ n42530;
  assign n42535 = n42530 ^ n42459;
  assign n42536 = n42534 & ~n42535;
  assign n42537 = n42536 ^ n42533;
  assign n42538 = n42537 ^ n42524;
  assign n42539 = n42525 & ~n42538;
  assign n42540 = n42539 ^ n42523;
  assign n42541 = n42540 ^ n42519;
  assign n42542 = n42520 & ~n42541;
  assign n42543 = n42542 ^ n42518;
  assign n42544 = n42543 ^ n42514;
  assign n42545 = ~n42515 & n42544;
  assign n42546 = n42545 ^ n42513;
  assign n42510 = n42464 ^ n42457;
  assign n42547 = n42546 ^ n42510;
  assign n42548 = n40333 ^ n32319;
  assign n42549 = n42548 ^ n36561;
  assign n42550 = n42549 ^ n30511;
  assign n42551 = n42550 ^ n42510;
  assign n42552 = n42547 & ~n42551;
  assign n42553 = n42552 ^ n42550;
  assign n42554 = n42553 ^ n42505;
  assign n42555 = ~n42509 & n42554;
  assign n42556 = n42555 ^ n42508;
  assign n42504 = n42466 ^ n42455;
  assign n42557 = n42556 ^ n42504;
  assign n42558 = n40323 ^ n32308;
  assign n42559 = n42558 ^ n36552;
  assign n42560 = n42559 ^ n30501;
  assign n42561 = n42560 ^ n42504;
  assign n42562 = n42557 & ~n42561;
  assign n42563 = n42562 ^ n42560;
  assign n42564 = n42563 ^ n42499;
  assign n42565 = ~n42503 & n42564;
  assign n42566 = n42565 ^ n42502;
  assign n42498 = n42469 ^ n42468;
  assign n42567 = n42566 ^ n42498;
  assign n42568 = n40378 ^ n32301;
  assign n42569 = n42568 ^ n36607;
  assign n42570 = n42569 ^ n632;
  assign n42571 = n42570 ^ n42498;
  assign n42572 = ~n42567 & n42571;
  assign n42573 = n42572 ^ n42570;
  assign n42574 = n42573 ^ n42496;
  assign n42575 = n42497 & ~n42574;
  assign n42576 = n42575 ^ n42495;
  assign n42577 = n42576 ^ n42491;
  assign n42578 = ~n42492 & n42577;
  assign n42579 = n42578 ^ n42490;
  assign n42580 = n42579 ^ n42483;
  assign n42581 = n42487 & ~n42580;
  assign n42582 = n42581 ^ n42486;
  assign n42583 = n42582 ^ n42478;
  assign n42584 = ~n42482 & n42583;
  assign n42585 = n42584 ^ n42481;
  assign n42586 = n42585 ^ n42476;
  assign n42587 = ~n42477 & n42586;
  assign n42588 = n42587 ^ n3350;
  assign n42917 = n42603 ^ n42588;
  assign n42918 = ~n42604 & n42917;
  assign n42919 = n42918 ^ n1354;
  assign n42824 = n42589 & n42602;
  assign n42770 = n42600 ^ n42592;
  assign n42771 = n42601 & n42770;
  assign n42772 = n42771 ^ n39675;
  assign n42669 = n42595 ^ n42594;
  assign n42670 = ~n42599 & ~n42669;
  assign n42671 = n42670 ^ n42594;
  assign n42666 = n41155 ^ n40496;
  assign n42667 = n42666 ^ n41812;
  assign n42665 = n42224 ^ n42205;
  assign n42668 = n42667 ^ n42665;
  assign n42768 = n42671 ^ n42668;
  assign n42769 = n42768 ^ n39528;
  assign n42823 = n42772 ^ n42769;
  assign n42916 = n42824 ^ n42823;
  assign n42920 = n42919 ^ n42916;
  assign n1364 = n1324 ^ n1264;
  assign n1365 = n1364 ^ n1361;
  assign n1372 = n1371 ^ n1365;
  assign n43094 = n42920 ^ n1372;
  assign n43091 = n41772 ^ n41126;
  assign n42714 = n42270 ^ n42177;
  assign n43092 = n43091 ^ n42714;
  assign n43206 = n43094 ^ n43092;
  assign n42614 = n42570 ^ n42567;
  assign n42612 = n42241 ^ n42238;
  assign n42611 = n41812 ^ n41168;
  assign n42613 = n42612 ^ n42611;
  assign n42615 = n42614 ^ n42613;
  assign n42618 = n42234 ^ n42199;
  assign n42617 = n41814 ^ n40423;
  assign n42619 = n42618 ^ n42617;
  assign n42616 = n42563 ^ n42503;
  assign n42620 = n42619 ^ n42616;
  assign n42624 = n42560 ^ n42557;
  assign n42622 = n42231 ^ n42228;
  assign n42621 = n41824 ^ n41183;
  assign n42623 = n42622 ^ n42621;
  assign n42625 = n42624 ^ n42623;
  assign n43039 = n42553 ^ n42509;
  assign n43032 = n42550 ^ n42547;
  assign n42632 = n42533 ^ n42459;
  assign n42633 = n42632 ^ n42530;
  assign n42630 = n41747 ^ n41109;
  assign n42631 = n42630 ^ n41738;
  assign n42634 = n42633 ^ n42631;
  assign n42635 = n41753 ^ n40971;
  assign n42636 = n42635 ^ n41743;
  assign n42638 = n42637 ^ n42636;
  assign n42655 = n42254 ^ n42193;
  assign n42653 = n41372 ^ n40456;
  assign n42654 = n42653 ^ n41782;
  assign n42656 = n42655 ^ n42654;
  assign n42659 = n41137 ^ n40478;
  assign n42660 = n42659 ^ n41796;
  assign n42661 = n42660 ^ n42612;
  assign n42662 = n41149 ^ n40490;
  assign n42663 = n42662 ^ n41921;
  assign n42664 = n42663 ^ n42622;
  assign n42672 = n42671 ^ n42665;
  assign n42673 = ~n42668 & ~n42672;
  assign n42674 = n42673 ^ n42667;
  assign n42675 = n42674 ^ n42622;
  assign n42676 = n42664 & ~n42675;
  assign n42677 = n42676 ^ n42663;
  assign n42678 = n42677 ^ n42618;
  assign n42679 = n41143 ^ n40484;
  assign n42680 = n42679 ^ n41802;
  assign n42681 = n42680 ^ n42618;
  assign n42682 = ~n42678 & ~n42681;
  assign n42683 = n42682 ^ n42680;
  assign n42684 = n42683 ^ n42612;
  assign n42685 = ~n42661 & ~n42684;
  assign n42686 = n42685 ^ n42660;
  assign n42658 = n42244 ^ n42196;
  assign n42687 = n42686 ^ n42658;
  assign n42688 = n41135 ^ n40472;
  assign n42689 = n42688 ^ n41790;
  assign n42690 = n42689 ^ n42658;
  assign n42691 = n42687 & n42690;
  assign n42692 = n42691 ^ n42689;
  assign n42657 = n42251 ^ n42248;
  assign n42693 = n42692 ^ n42657;
  assign n42694 = n41126 ^ n40466;
  assign n42695 = n42694 ^ n41788;
  assign n42696 = n42695 ^ n42657;
  assign n42697 = ~n42693 & n42696;
  assign n42698 = n42697 ^ n42695;
  assign n42699 = n42698 ^ n42655;
  assign n42700 = ~n42656 & n42699;
  assign n42701 = n42700 ^ n42654;
  assign n42652 = n42261 ^ n42258;
  assign n42702 = n42701 ^ n42652;
  assign n42703 = n41389 ^ n40584;
  assign n42704 = n42703 ^ n41772;
  assign n42705 = n42704 ^ n42652;
  assign n42706 = ~n42702 & n42705;
  assign n42707 = n42706 ^ n42704;
  assign n42650 = n42264 ^ n42187;
  assign n42648 = n41405 ^ n40707;
  assign n42649 = n42648 ^ n41770;
  assign n42651 = n42650 ^ n42649;
  assign n42753 = n42707 ^ n42651;
  assign n42754 = n42753 ^ n39899;
  assign n42755 = n42704 ^ n42702;
  assign n42756 = n42755 ^ n39706;
  assign n42757 = n42698 ^ n42656;
  assign n42758 = n42757 ^ n39492;
  assign n42760 = n42689 ^ n42687;
  assign n42761 = n42760 ^ n39504;
  assign n42762 = n42683 ^ n42661;
  assign n42763 = n42762 ^ n39510;
  assign n42764 = n42680 ^ n42678;
  assign n42765 = n42764 ^ n39516;
  assign n42766 = n42674 ^ n42664;
  assign n42767 = n42766 ^ n39522;
  assign n42773 = n42772 ^ n42768;
  assign n42774 = ~n42769 & n42773;
  assign n42775 = n42774 ^ n39528;
  assign n42776 = n42775 ^ n42766;
  assign n42777 = n42767 & n42776;
  assign n42778 = n42777 ^ n39522;
  assign n42779 = n42778 ^ n42764;
  assign n42780 = ~n42765 & n42779;
  assign n42781 = n42780 ^ n39516;
  assign n42782 = n42781 ^ n42762;
  assign n42783 = ~n42763 & ~n42782;
  assign n42784 = n42783 ^ n39510;
  assign n42785 = n42784 ^ n42760;
  assign n42786 = ~n42761 & n42785;
  assign n42787 = n42786 ^ n39504;
  assign n42759 = n42695 ^ n42693;
  assign n42788 = n42787 ^ n42759;
  assign n42789 = n42759 ^ n39498;
  assign n42790 = ~n42788 & n42789;
  assign n42791 = n42790 ^ n39498;
  assign n42792 = n42791 ^ n42757;
  assign n42793 = ~n42758 & n42792;
  assign n42794 = n42793 ^ n39492;
  assign n42795 = n42794 ^ n42755;
  assign n42796 = ~n42756 & ~n42795;
  assign n42797 = n42796 ^ n39706;
  assign n42798 = n42797 ^ n42753;
  assign n42799 = ~n42754 & ~n42798;
  assign n42800 = n42799 ^ n39899;
  assign n42708 = n42707 ^ n42650;
  assign n42709 = ~n42651 & n42708;
  assign n42710 = n42709 ^ n42649;
  assign n42646 = n42267 ^ n42182;
  assign n42644 = n40858 ^ n40128;
  assign n42645 = n42644 ^ n41951;
  assign n42647 = n42646 ^ n42645;
  assign n42751 = n42710 ^ n42647;
  assign n42752 = n42751 ^ n39358;
  assign n42818 = n42800 ^ n42752;
  assign n42819 = n42797 ^ n42754;
  assign n42820 = n42794 ^ n42756;
  assign n42821 = n42788 ^ n39498;
  assign n42822 = n42775 ^ n42767;
  assign n42825 = ~n42823 & ~n42824;
  assign n42826 = ~n42822 & ~n42825;
  assign n42827 = n42778 ^ n42765;
  assign n42828 = ~n42826 & n42827;
  assign n42829 = n42781 ^ n42763;
  assign n42830 = n42828 & n42829;
  assign n42831 = n42784 ^ n42761;
  assign n42832 = n42830 & ~n42831;
  assign n42833 = ~n42821 & ~n42832;
  assign n42834 = n42791 ^ n42758;
  assign n42835 = n42833 & n42834;
  assign n42836 = ~n42820 & ~n42835;
  assign n42837 = n42819 & n42836;
  assign n42838 = ~n42818 & ~n42837;
  assign n42801 = n42800 ^ n42751;
  assign n42802 = n42752 & n42801;
  assign n42803 = n42802 ^ n39358;
  assign n42716 = n40848 ^ n40122;
  assign n42717 = n42716 ^ n42135;
  assign n42711 = n42710 ^ n42646;
  assign n42712 = ~n42647 & ~n42711;
  assign n42713 = n42712 ^ n42645;
  assign n42715 = n42714 ^ n42713;
  assign n42749 = n42717 ^ n42715;
  assign n42750 = n42749 ^ n39369;
  assign n42839 = n42803 ^ n42750;
  assign n42840 = ~n42838 & ~n42839;
  assign n42804 = n42803 ^ n42749;
  assign n42805 = n42750 & n42804;
  assign n42806 = n42805 ^ n39369;
  assign n42722 = n40842 ^ n40116;
  assign n42723 = n42722 ^ n41577;
  assign n42718 = n42717 ^ n42714;
  assign n42719 = n42715 & ~n42718;
  assign n42720 = n42719 ^ n42717;
  assign n42643 = n42273 ^ n42172;
  assign n42721 = n42720 ^ n42643;
  assign n42747 = n42723 ^ n42721;
  assign n42748 = n42747 ^ n39352;
  assign n42841 = n42806 ^ n42748;
  assign n42842 = ~n42840 & ~n42841;
  assign n42807 = n42806 ^ n42747;
  assign n42808 = n42748 & ~n42807;
  assign n42809 = n42808 ^ n39352;
  assign n42728 = n40836 ^ n40114;
  assign n42729 = n42728 ^ n41567;
  assign n42724 = n42723 ^ n42643;
  assign n42725 = n42721 & ~n42724;
  assign n42726 = n42725 ^ n42723;
  assign n42642 = n42276 ^ n42167;
  assign n42727 = n42726 ^ n42642;
  assign n42745 = n42729 ^ n42727;
  assign n42746 = n42745 ^ n39346;
  assign n42843 = n42809 ^ n42746;
  assign n42844 = ~n42842 & ~n42843;
  assign n42810 = n42809 ^ n42745;
  assign n42811 = ~n42746 & ~n42810;
  assign n42812 = n42811 ^ n39346;
  assign n42735 = n40830 ^ n40104;
  assign n42736 = n42735 ^ n41561;
  assign n42733 = n42279 ^ n42162;
  assign n42730 = n42729 ^ n42642;
  assign n42731 = ~n42727 & ~n42730;
  assign n42732 = n42731 ^ n42729;
  assign n42734 = n42733 ^ n42732;
  assign n42743 = n42736 ^ n42734;
  assign n42744 = n42743 ^ n39340;
  assign n42817 = n42812 ^ n42744;
  assign n42869 = n42844 ^ n42817;
  assign n42866 = n40816 ^ n32485;
  assign n42867 = n42866 ^ n37067;
  assign n42868 = n42867 ^ n1852;
  assign n42870 = n42869 ^ n42868;
  assign n42872 = n40726 ^ n1744;
  assign n42873 = n42872 ^ n36952;
  assign n42874 = n42873 ^ n31061;
  assign n42871 = n42843 ^ n42842;
  assign n42875 = n42874 ^ n42871;
  assign n42878 = n40803 ^ n32238;
  assign n42879 = n42878 ^ n36962;
  assign n42880 = n42879 ^ n31050;
  assign n42877 = n42839 ^ n42838;
  assign n42881 = n42880 ^ n42877;
  assign n42882 = n42837 ^ n42818;
  assign n42886 = n42885 ^ n42882;
  assign n42888 = n42835 ^ n42820;
  assign n3102 = n3101 ^ n3095;
  assign n3106 = n3105 ^ n3102;
  assign n3107 = n3106 ^ n2760;
  assign n42889 = n42888 ^ n3107;
  assign n42892 = n40784 ^ n3081;
  assign n42893 = n42892 ^ n3191;
  assign n42894 = n42893 ^ n2665;
  assign n42891 = n42832 ^ n42821;
  assign n42895 = n42894 ^ n42891;
  assign n42897 = n40752 ^ n2565;
  assign n42898 = n42897 ^ n36977;
  assign n42899 = n42898 ^ n3189;
  assign n42896 = n42831 ^ n42830;
  assign n42900 = n42899 ^ n42896;
  assign n42902 = n40757 ^ n3167;
  assign n42903 = n42902 ^ n36982;
  assign n42904 = n42903 ^ n30996;
  assign n42901 = n42829 ^ n42828;
  assign n42905 = n42904 ^ n42901;
  assign n42909 = n42827 ^ n42826;
  assign n42906 = n40762 ^ n32380;
  assign n42907 = n42906 ^ n36986;
  assign n42908 = n42907 ^ n31006;
  assign n42910 = n42909 ^ n42908;
  assign n42914 = n42825 ^ n42822;
  assign n42911 = n32386 ^ n1428;
  assign n42912 = n42911 ^ n37027;
  assign n42913 = n42912 ^ n31001;
  assign n42915 = n42914 ^ n42913;
  assign n42921 = n42916 ^ n1372;
  assign n42922 = ~n42920 & n42921;
  assign n42923 = n42922 ^ n1372;
  assign n42924 = n42923 ^ n42914;
  assign n42925 = ~n42915 & n42924;
  assign n42926 = n42925 ^ n42913;
  assign n42927 = n42926 ^ n42909;
  assign n42928 = ~n42910 & n42927;
  assign n42929 = n42928 ^ n42908;
  assign n42930 = n42929 ^ n42901;
  assign n42931 = n42905 & ~n42930;
  assign n42932 = n42931 ^ n42904;
  assign n42933 = n42932 ^ n42896;
  assign n42934 = ~n42900 & n42933;
  assign n42935 = n42934 ^ n42899;
  assign n42936 = n42935 ^ n42891;
  assign n42937 = ~n42895 & n42936;
  assign n42938 = n42937 ^ n42894;
  assign n42890 = n42834 ^ n42833;
  assign n42939 = n42938 ^ n42890;
  assign n2646 = n2645 ^ n2624;
  assign n2674 = n2673 ^ n2646;
  assign n2681 = n2680 ^ n2674;
  assign n42940 = n42890 ^ n2681;
  assign n42941 = n42939 & ~n42940;
  assign n42942 = n42941 ^ n2681;
  assign n42943 = n42942 ^ n42888;
  assign n42944 = n42889 & ~n42943;
  assign n42945 = n42944 ^ n3107;
  assign n42887 = n42836 ^ n42819;
  assign n42946 = n42945 ^ n42887;
  assign n42947 = n40742 ^ n32262;
  assign n42948 = n42947 ^ n2762;
  assign n42949 = n42948 ^ n3125;
  assign n42950 = n42949 ^ n42887;
  assign n42951 = ~n42946 & n42950;
  assign n42952 = n42951 ^ n42949;
  assign n42953 = n42952 ^ n42882;
  assign n42954 = ~n42886 & n42953;
  assign n42955 = n42954 ^ n42885;
  assign n42956 = n42955 ^ n42877;
  assign n42957 = n42881 & ~n42956;
  assign n42958 = n42957 ^ n42880;
  assign n42876 = n42841 ^ n42840;
  assign n42959 = n42958 ^ n42876;
  assign n42963 = n42962 ^ n42876;
  assign n42964 = n42959 & ~n42963;
  assign n42965 = n42964 ^ n42962;
  assign n42966 = n42965 ^ n42871;
  assign n42967 = n42875 & ~n42966;
  assign n42968 = n42967 ^ n42874;
  assign n42969 = n42968 ^ n42869;
  assign n42970 = ~n42870 & n42969;
  assign n42971 = n42970 ^ n42868;
  assign n42845 = ~n42817 & n42844;
  assign n42813 = n42812 ^ n42743;
  assign n42814 = n42744 & n42813;
  assign n42815 = n42814 ^ n39340;
  assign n42737 = n42736 ^ n42733;
  assign n42738 = ~n42734 & n42737;
  assign n42739 = n42738 ^ n42736;
  assign n42641 = n42283 ^ n2995;
  assign n42740 = n42739 ^ n42641;
  assign n42639 = n40454 ^ n39481;
  assign n42640 = n42639 ^ n41559;
  assign n42741 = n42740 ^ n42640;
  assign n42742 = n42741 ^ n39437;
  assign n42816 = n42815 ^ n42742;
  assign n42865 = n42845 ^ n42816;
  assign n42972 = n42971 ^ n42865;
  assign n1833 = n1832 ^ n1802;
  assign n1861 = n1860 ^ n1833;
  assign n1868 = n1867 ^ n1861;
  assign n42979 = n42972 ^ n1868;
  assign n42977 = n41762 ^ n40426;
  assign n42978 = n42977 ^ n41749;
  assign n42980 = n42979 ^ n42978;
  assign n42986 = n41669 ^ n40438;
  assign n42987 = n42986 ^ n41759;
  assign n42982 = n42962 ^ n42959;
  assign n42983 = n41644 ^ n40878;
  assign n42984 = n42983 ^ n41764;
  assign n42985 = ~n42982 & ~n42984;
  assign n42988 = n42987 ^ n42985;
  assign n42989 = n42965 ^ n42875;
  assign n42990 = n42989 ^ n42987;
  assign n42991 = ~n42988 & n42990;
  assign n42992 = n42991 ^ n42985;
  assign n42981 = n42968 ^ n42870;
  assign n42993 = n42992 ^ n42981;
  assign n42994 = n41876 ^ n40432;
  assign n42995 = n42994 ^ n41751;
  assign n42996 = n42995 ^ n42981;
  assign n42997 = n42993 & n42996;
  assign n42998 = n42997 ^ n42995;
  assign n42999 = n42998 ^ n42979;
  assign n43000 = ~n42980 & n42999;
  assign n43001 = n43000 ^ n42978;
  assign n42973 = n42865 ^ n1868;
  assign n42974 = ~n42972 & n42973;
  assign n42975 = n42974 ^ n1868;
  assign n42858 = n42815 ^ n42741;
  assign n42859 = ~n42742 & ~n42858;
  assign n42860 = n42859 ^ n39437;
  assign n42861 = n42860 ^ n39612;
  assign n42854 = n42641 ^ n42640;
  assign n42855 = n42740 & n42854;
  assign n42856 = n42855 ^ n42640;
  assign n42852 = n42286 ^ n42156;
  assign n42850 = n40448 ^ n39479;
  assign n42851 = n42850 ^ n41549;
  assign n42853 = n42852 ^ n42851;
  assign n42857 = n42856 ^ n42853;
  assign n42862 = n42861 ^ n42857;
  assign n42847 = n40717 ^ n32748;
  assign n42848 = n42847 ^ n37126;
  assign n42849 = n42848 ^ n1978;
  assign n42863 = n42862 ^ n42849;
  assign n42846 = n42816 & ~n42845;
  assign n42864 = n42863 ^ n42846;
  assign n42976 = n42975 ^ n42864;
  assign n43002 = n43001 ^ n42976;
  assign n43003 = n41756 ^ n40901;
  assign n43004 = n43003 ^ n41745;
  assign n43005 = n43004 ^ n42976;
  assign n43006 = n43002 & ~n43005;
  assign n43007 = n43006 ^ n43004;
  assign n43008 = n43007 ^ n42637;
  assign n43009 = ~n42638 & ~n43008;
  assign n43010 = n43009 ^ n42636;
  assign n43011 = n43010 ^ n42633;
  assign n43012 = n42634 & ~n43011;
  assign n43013 = n43012 ^ n42631;
  assign n42628 = n42537 ^ n42523;
  assign n42629 = n42628 ^ n42524;
  assign n43014 = n43013 ^ n42629;
  assign n43015 = n41850 ^ n41213;
  assign n43016 = n43015 ^ n41733;
  assign n43017 = n43016 ^ n42629;
  assign n43018 = ~n43014 & n43017;
  assign n43019 = n43018 ^ n43016;
  assign n42627 = n42540 ^ n42520;
  assign n43020 = n43019 ^ n42627;
  assign n43021 = n41741 ^ n41207;
  assign n43022 = n43021 ^ n41729;
  assign n43023 = n43022 ^ n42627;
  assign n43024 = ~n43020 & n43023;
  assign n43025 = n43024 ^ n43022;
  assign n42626 = n42543 ^ n42515;
  assign n43026 = n43025 ^ n42626;
  assign n43027 = n41736 ^ n41201;
  assign n43028 = n43027 ^ n42446;
  assign n43029 = n43028 ^ n42626;
  assign n43030 = n43026 & ~n43029;
  assign n43031 = n43030 ^ n43028;
  assign n43033 = n43032 ^ n43031;
  assign n43034 = n41731 ^ n41195;
  assign n43035 = n43034 ^ n42595;
  assign n43036 = n43035 ^ n43032;
  assign n43037 = n43033 & ~n43036;
  assign n43038 = n43037 ^ n43035;
  assign n43040 = n43039 ^ n43038;
  assign n43041 = n41189 ^ n41115;
  assign n43042 = n43041 ^ n42665;
  assign n43043 = n43042 ^ n43039;
  assign n43044 = n43040 & ~n43043;
  assign n43045 = n43044 ^ n43042;
  assign n43046 = n43045 ^ n42624;
  assign n43047 = n42625 & n43046;
  assign n43048 = n43047 ^ n42623;
  assign n43049 = n43048 ^ n42616;
  assign n43050 = ~n42620 & ~n43049;
  assign n43051 = n43050 ^ n42619;
  assign n43052 = n43051 ^ n42614;
  assign n43053 = n42615 & ~n43052;
  assign n43054 = n43053 ^ n42613;
  assign n42610 = n42573 ^ n42497;
  assign n43055 = n43054 ^ n42610;
  assign n43056 = n41921 ^ n41161;
  assign n43057 = n43056 ^ n42658;
  assign n43058 = n43057 ^ n42610;
  assign n43059 = ~n43055 & ~n43058;
  assign n43060 = n43059 ^ n43057;
  assign n42609 = n42576 ^ n42492;
  assign n43061 = n43060 ^ n42609;
  assign n43062 = n41802 ^ n41155;
  assign n43063 = n43062 ^ n42657;
  assign n43064 = n43063 ^ n42609;
  assign n43065 = ~n43061 & ~n43064;
  assign n43066 = n43065 ^ n43063;
  assign n42608 = n42579 ^ n42487;
  assign n43067 = n43066 ^ n42608;
  assign n43068 = n41796 ^ n41149;
  assign n43069 = n43068 ^ n42655;
  assign n43070 = n43069 ^ n42608;
  assign n43071 = ~n43067 & ~n43070;
  assign n43072 = n43071 ^ n43069;
  assign n42607 = n42582 ^ n42482;
  assign n43073 = n43072 ^ n42607;
  assign n43074 = n41790 ^ n41143;
  assign n43075 = n43074 ^ n42652;
  assign n43076 = n43075 ^ n42607;
  assign n43077 = ~n43073 & n43076;
  assign n43078 = n43077 ^ n43075;
  assign n42606 = n42585 ^ n42477;
  assign n43079 = n43078 ^ n42606;
  assign n43080 = n41788 ^ n41137;
  assign n43081 = n43080 ^ n42650;
  assign n43082 = n43081 ^ n42606;
  assign n43083 = ~n43079 & ~n43082;
  assign n43084 = n43083 ^ n43081;
  assign n42605 = n42604 ^ n42588;
  assign n43085 = n43084 ^ n42605;
  assign n43086 = n41782 ^ n41135;
  assign n43087 = n43086 ^ n42646;
  assign n43088 = n43087 ^ n42605;
  assign n43089 = n43085 & ~n43088;
  assign n43090 = n43089 ^ n43087;
  assign n43207 = n43094 ^ n43090;
  assign n43208 = ~n43206 & ~n43207;
  assign n43209 = n43208 ^ n43092;
  assign n43205 = n42923 ^ n42915;
  assign n43210 = n43209 ^ n43205;
  assign n43203 = n41770 ^ n41372;
  assign n43204 = n43203 ^ n42643;
  assign n43211 = n43210 ^ n43204;
  assign n43093 = n43092 ^ n43090;
  assign n43095 = n43094 ^ n43093;
  assign n43096 = n43095 ^ n40466;
  assign n43097 = n43087 ^ n43085;
  assign n43098 = n43097 ^ n40472;
  assign n43099 = n43081 ^ n43079;
  assign n43100 = n43099 ^ n40478;
  assign n43101 = n43075 ^ n43073;
  assign n43102 = n43101 ^ n40484;
  assign n43103 = n43069 ^ n43067;
  assign n43104 = n43103 ^ n40490;
  assign n43105 = n43063 ^ n43061;
  assign n43106 = n43105 ^ n40496;
  assign n43107 = n43057 ^ n43055;
  assign n43108 = n43107 ^ n40498;
  assign n43109 = n43051 ^ n42615;
  assign n43110 = n43109 ^ n40504;
  assign n43111 = n43048 ^ n42620;
  assign n43112 = n43111 ^ n40424;
  assign n43113 = n43045 ^ n42625;
  assign n43114 = n43113 ^ n40515;
  assign n43116 = n43035 ^ n43033;
  assign n43117 = n43116 ^ n40527;
  assign n43119 = n43022 ^ n43020;
  assign n43120 = n43119 ^ n40411;
  assign n43121 = n43016 ^ n43014;
  assign n43122 = n43121 ^ n40286;
  assign n43123 = n43010 ^ n42634;
  assign n43124 = n43123 ^ n40248;
  assign n43126 = n43004 ^ n43002;
  assign n43127 = n43126 ^ n40168;
  assign n43128 = n42998 ^ n42980;
  assign n43129 = n43128 ^ n39451;
  assign n43130 = n42995 ^ n42993;
  assign n43131 = n43130 ^ n39458;
  assign n43132 = n42984 ^ n42982;
  assign n43133 = n39472 & n43132;
  assign n43134 = n43133 ^ n39465;
  assign n43135 = n42989 ^ n42988;
  assign n43136 = n43135 ^ n43133;
  assign n43137 = ~n43134 & n43136;
  assign n43138 = n43137 ^ n39465;
  assign n43139 = n43138 ^ n43130;
  assign n43140 = ~n43131 & n43139;
  assign n43141 = n43140 ^ n39458;
  assign n43142 = n43141 ^ n43128;
  assign n43143 = ~n43129 & n43142;
  assign n43144 = n43143 ^ n39451;
  assign n43145 = n43144 ^ n43126;
  assign n43146 = ~n43127 & n43145;
  assign n43147 = n43146 ^ n40168;
  assign n43125 = n43007 ^ n42638;
  assign n43148 = n43147 ^ n43125;
  assign n43149 = n43125 ^ n40239;
  assign n43150 = n43148 & n43149;
  assign n43151 = n43150 ^ n40239;
  assign n43152 = n43151 ^ n43123;
  assign n43153 = n43124 & ~n43152;
  assign n43154 = n43153 ^ n40248;
  assign n43155 = n43154 ^ n43121;
  assign n43156 = ~n43122 & ~n43155;
  assign n43157 = n43156 ^ n40286;
  assign n43158 = n43157 ^ n43119;
  assign n43159 = n43120 & n43158;
  assign n43160 = n43159 ^ n40411;
  assign n43118 = n43028 ^ n43026;
  assign n43161 = n43160 ^ n43118;
  assign n43162 = n43118 ^ n40533;
  assign n43163 = n43161 & ~n43162;
  assign n43164 = n43163 ^ n40533;
  assign n43165 = n43164 ^ n43116;
  assign n43166 = ~n43117 & n43165;
  assign n43167 = n43166 ^ n40527;
  assign n43115 = n43042 ^ n43040;
  assign n43168 = n43167 ^ n43115;
  assign n43169 = n43115 ^ n40521;
  assign n43170 = n43168 & n43169;
  assign n43171 = n43170 ^ n40521;
  assign n43172 = n43171 ^ n43113;
  assign n43173 = n43114 & n43172;
  assign n43174 = n43173 ^ n40515;
  assign n43175 = n43174 ^ n43111;
  assign n43176 = ~n43112 & ~n43175;
  assign n43177 = n43176 ^ n40424;
  assign n43178 = n43177 ^ n43109;
  assign n43179 = n43110 & n43178;
  assign n43180 = n43179 ^ n40504;
  assign n43181 = n43180 ^ n43107;
  assign n43182 = n43108 & n43181;
  assign n43183 = n43182 ^ n40498;
  assign n43184 = n43183 ^ n43105;
  assign n43185 = ~n43106 & n43184;
  assign n43186 = n43185 ^ n40496;
  assign n43187 = n43186 ^ n43103;
  assign n43188 = ~n43104 & ~n43187;
  assign n43189 = n43188 ^ n40490;
  assign n43190 = n43189 ^ n43101;
  assign n43191 = ~n43102 & n43190;
  assign n43192 = n43191 ^ n40484;
  assign n43193 = n43192 ^ n43099;
  assign n43194 = ~n43100 & ~n43193;
  assign n43195 = n43194 ^ n40478;
  assign n43196 = n43195 ^ n43097;
  assign n43197 = n43098 & ~n43196;
  assign n43198 = n43197 ^ n40472;
  assign n43199 = n43198 ^ n43095;
  assign n43200 = n43096 & ~n43199;
  assign n43201 = n43200 ^ n40466;
  assign n43202 = n43201 ^ n40456;
  assign n43212 = n43211 ^ n43202;
  assign n43213 = n43192 ^ n43100;
  assign n43214 = n43189 ^ n43102;
  assign n43215 = n43180 ^ n43108;
  assign n43216 = n43177 ^ n43110;
  assign n43217 = n43174 ^ n43112;
  assign n43218 = n43171 ^ n43114;
  assign n43219 = n43164 ^ n43117;
  assign n43220 = n43161 ^ n40533;
  assign n43221 = n43157 ^ n43120;
  assign n43222 = n43154 ^ n43122;
  assign n43223 = n43135 ^ n43134;
  assign n43224 = n43138 ^ n43131;
  assign n43225 = ~n43223 & ~n43224;
  assign n43226 = n43141 ^ n39451;
  assign n43227 = n43226 ^ n43128;
  assign n43228 = ~n43225 & n43227;
  assign n43229 = n43144 ^ n43127;
  assign n43230 = ~n43228 & ~n43229;
  assign n43231 = n43148 ^ n40239;
  assign n43232 = ~n43230 & ~n43231;
  assign n43233 = n43151 ^ n43124;
  assign n43234 = ~n43232 & ~n43233;
  assign n43235 = n43222 & n43234;
  assign n43236 = n43221 & n43235;
  assign n43237 = ~n43220 & ~n43236;
  assign n43238 = ~n43219 & n43237;
  assign n43239 = n43168 ^ n40521;
  assign n43240 = n43238 & n43239;
  assign n43241 = ~n43218 & n43240;
  assign n43242 = ~n43217 & n43241;
  assign n43243 = n43216 & ~n43242;
  assign n43244 = ~n43215 & n43243;
  assign n43245 = n43183 ^ n43106;
  assign n43246 = ~n43244 & n43245;
  assign n43247 = n43186 ^ n43104;
  assign n43248 = ~n43246 & ~n43247;
  assign n43249 = ~n43214 & ~n43248;
  assign n43250 = ~n43213 & n43249;
  assign n43251 = n43195 ^ n43098;
  assign n43252 = n43250 & ~n43251;
  assign n43253 = n43198 ^ n43096;
  assign n43254 = ~n43252 & n43253;
  assign n43255 = n43212 & n43254;
  assign n43266 = n41951 ^ n41389;
  assign n43267 = n43266 ^ n42642;
  assign n43262 = n43205 ^ n43204;
  assign n43263 = ~n43210 & n43262;
  assign n43264 = n43263 ^ n43204;
  assign n43261 = n42926 ^ n42910;
  assign n43265 = n43264 ^ n43261;
  assign n43268 = n43267 ^ n43265;
  assign n43256 = n43211 ^ n40456;
  assign n43257 = n43211 ^ n43201;
  assign n43258 = n43256 & ~n43257;
  assign n43259 = n43258 ^ n40456;
  assign n43260 = n43259 ^ n40584;
  assign n43269 = n43268 ^ n43260;
  assign n43270 = ~n43255 & n43269;
  assign n43280 = n43268 ^ n40584;
  assign n43281 = n43268 ^ n43259;
  assign n43282 = ~n43280 & ~n43281;
  assign n43283 = n43282 ^ n40584;
  assign n43276 = n42135 ^ n41405;
  assign n43277 = n43276 ^ n42733;
  assign n43272 = n43267 ^ n43261;
  assign n43273 = ~n43265 & n43272;
  assign n43274 = n43273 ^ n43267;
  assign n43271 = n42929 ^ n42905;
  assign n43275 = n43274 ^ n43271;
  assign n43278 = n43277 ^ n43275;
  assign n43279 = n43278 ^ n40707;
  assign n43284 = n43283 ^ n43279;
  assign n43479 = n43270 & n43284;
  assign n43475 = n43283 ^ n43278;
  assign n43476 = n43279 & n43475;
  assign n43477 = n43476 ^ n40707;
  assign n43471 = n41577 ^ n40858;
  assign n43472 = n43471 ^ n42641;
  assign n43469 = n42932 ^ n42900;
  assign n43466 = n43277 ^ n43271;
  assign n43467 = n43275 & n43466;
  assign n43468 = n43467 ^ n43277;
  assign n43470 = n43469 ^ n43468;
  assign n43473 = n43472 ^ n43470;
  assign n43474 = n43473 ^ n40128;
  assign n43478 = n43477 ^ n43474;
  assign n43480 = n43479 ^ n43478;
  assign n43484 = n43483 ^ n43480;
  assign n43285 = n43284 ^ n43270;
  assign n2830 = n2826 ^ n2796;
  assign n2855 = n2854 ^ n2830;
  assign n2862 = n2861 ^ n2855;
  assign n43286 = n43285 ^ n2862;
  assign n43287 = n43269 ^ n43255;
  assign n3216 = n3215 ^ n2737;
  assign n3226 = n3225 ^ n3216;
  assign n3227 = n3226 ^ n2846;
  assign n43288 = n43287 ^ n3227;
  assign n43293 = n43253 ^ n43252;
  assign n43290 = n41460 ^ n3201;
  assign n43291 = n43290 ^ n37770;
  assign n43292 = n43291 ^ n31345;
  assign n43294 = n43293 ^ n43292;
  assign n43298 = n43251 ^ n43250;
  assign n43295 = n41510 ^ n33178;
  assign n43296 = n43295 ^ n37775;
  assign n43297 = n43296 ^ n31350;
  assign n43299 = n43298 ^ n43297;
  assign n43301 = n41467 ^ n33183;
  assign n43302 = n43301 ^ n37780;
  assign n43303 = n43302 ^ n3047;
  assign n43300 = n43249 ^ n43213;
  assign n43304 = n43303 ^ n43300;
  assign n43308 = n43248 ^ n43214;
  assign n43305 = n41471 ^ n33190;
  assign n43306 = n43305 ^ n37785;
  assign n43307 = n43306 ^ n2453;
  assign n43309 = n43308 ^ n43307;
  assign n43315 = n43243 ^ n43215;
  assign n43312 = n41487 ^ n1452;
  assign n43313 = n43312 ^ n37863;
  assign n43314 = n43313 ^ n1193;
  assign n43316 = n43315 ^ n43314;
  assign n43320 = n43242 ^ n43216;
  assign n43317 = n41096 ^ n33208;
  assign n43318 = n43317 ^ n1034;
  assign n43319 = n43318 ^ n31371;
  assign n43321 = n43320 ^ n43319;
  assign n43325 = n43241 ^ n43217;
  assign n43322 = n41090 ^ n33213;
  assign n43323 = n43322 ^ n37853;
  assign n43324 = n43323 ^ n1026;
  assign n43326 = n43325 ^ n43324;
  assign n43327 = n43240 ^ n43218;
  assign n879 = n878 ^ n848;
  assign n907 = n906 ^ n879;
  assign n914 = n913 ^ n907;
  assign n43328 = n43327 ^ n914;
  assign n43330 = n41005 ^ n33220;
  assign n43331 = n43330 ^ n37843;
  assign n43332 = n43331 ^ n898;
  assign n43329 = n43239 ^ n43238;
  assign n43333 = n43332 ^ n43329;
  assign n43337 = n37814 ^ n33232;
  assign n43338 = n43337 ^ n41016;
  assign n43339 = n43338 ^ n31389;
  assign n43336 = n43235 ^ n43221;
  assign n43340 = n43339 ^ n43336;
  assign n43345 = n43233 ^ n43232;
  assign n43342 = n41025 ^ n33242;
  assign n43343 = n43342 ^ n37236;
  assign n43344 = n43343 ^ n31398;
  assign n43346 = n43345 ^ n43344;
  assign n43349 = n41036 ^ n33251;
  assign n43350 = n43349 ^ n37212;
  assign n43351 = n43350 ^ n31409;
  assign n43348 = n43229 ^ n43228;
  assign n43352 = n43351 ^ n43348;
  assign n43354 = n41040 ^ n33256;
  assign n43355 = n43354 ^ n37216;
  assign n43356 = n43355 ^ n31421;
  assign n43353 = n43227 ^ n43225;
  assign n43357 = n43356 ^ n43353;
  assign n43358 = n43224 ^ n43223;
  assign n2232 = n2231 ^ n2159;
  assign n2248 = n2247 ^ n2232;
  assign n2255 = n2254 ^ n2248;
  assign n43359 = n43358 ^ n2255;
  assign n2068 = n2058 ^ n2013;
  assign n2093 = n2092 ^ n2068;
  assign n2100 = n2099 ^ n2093;
  assign n43363 = n43132 ^ n39472;
  assign n43364 = n2100 & n43363;
  assign n43360 = n41044 ^ n32500;
  assign n43361 = n43360 ^ n2110;
  assign n43362 = n43361 ^ n2246;
  assign n43365 = n43364 ^ n43362;
  assign n43366 = n43364 ^ n43223;
  assign n43367 = n43365 & n43366;
  assign n43368 = n43367 ^ n43362;
  assign n43369 = n43368 ^ n43358;
  assign n43370 = ~n43359 & n43369;
  assign n43371 = n43370 ^ n2255;
  assign n43372 = n43371 ^ n43353;
  assign n43373 = ~n43357 & n43372;
  assign n43374 = n43373 ^ n43356;
  assign n43375 = n43374 ^ n43348;
  assign n43376 = ~n43352 & n43375;
  assign n43377 = n43376 ^ n43351;
  assign n43347 = n43231 ^ n43230;
  assign n43378 = n43377 ^ n43347;
  assign n43379 = n41031 ^ n33247;
  assign n43380 = n43379 ^ n37207;
  assign n43381 = n43380 ^ n31404;
  assign n43382 = n43381 ^ n43347;
  assign n43383 = ~n43378 & n43382;
  assign n43384 = n43383 ^ n43381;
  assign n43385 = n43384 ^ n43345;
  assign n43386 = ~n43346 & n43385;
  assign n43387 = n43386 ^ n43344;
  assign n43341 = n43234 ^ n43222;
  assign n43388 = n43387 ^ n43341;
  assign n43389 = n41020 ^ n33237;
  assign n43390 = n43389 ^ n37818;
  assign n43391 = n43390 ^ n31394;
  assign n43392 = n43391 ^ n43387;
  assign n43393 = n43388 & n43392;
  assign n43394 = n43393 ^ n43391;
  assign n43395 = n43394 ^ n43336;
  assign n43396 = ~n43340 & n43395;
  assign n43397 = n43396 ^ n43339;
  assign n43335 = n43236 ^ n43220;
  assign n43398 = n43397 ^ n43335;
  assign n43402 = n43401 ^ n43335;
  assign n43403 = ~n43398 & n43402;
  assign n43404 = n43403 ^ n43401;
  assign n43334 = n43237 ^ n43219;
  assign n43405 = n43404 ^ n43334;
  assign n43406 = n41010 ^ n780;
  assign n43407 = n43406 ^ n37808;
  assign n43408 = n43407 ^ n3305;
  assign n43409 = n43408 ^ n43334;
  assign n43410 = n43405 & ~n43409;
  assign n43411 = n43410 ^ n43408;
  assign n43412 = n43411 ^ n43329;
  assign n43413 = n43333 & ~n43412;
  assign n43414 = n43413 ^ n43332;
  assign n43415 = n43414 ^ n43327;
  assign n43416 = ~n43328 & n43415;
  assign n43417 = n43416 ^ n914;
  assign n43418 = n43417 ^ n43325;
  assign n43419 = ~n43326 & n43418;
  assign n43420 = n43419 ^ n43324;
  assign n43421 = n43420 ^ n43320;
  assign n43422 = n43321 & ~n43421;
  assign n43423 = n43422 ^ n43319;
  assign n43424 = n43423 ^ n43315;
  assign n43425 = n43316 & ~n43424;
  assign n43426 = n43425 ^ n43314;
  assign n43311 = n43245 ^ n43244;
  assign n43427 = n43426 ^ n43311;
  assign n43428 = n41478 ^ n1467;
  assign n43429 = n43428 ^ n37796;
  assign n43430 = n43429 ^ n31364;
  assign n43431 = n43430 ^ n43311;
  assign n43432 = n43427 & ~n43431;
  assign n43433 = n43432 ^ n43430;
  assign n43310 = n43247 ^ n43246;
  assign n43434 = n43433 ^ n43310;
  assign n43435 = n41497 ^ n1485;
  assign n43436 = n43435 ^ n37790;
  assign n43437 = n43436 ^ n31358;
  assign n43438 = n43437 ^ n43310;
  assign n43439 = n43434 & ~n43438;
  assign n43440 = n43439 ^ n43437;
  assign n43441 = n43440 ^ n43308;
  assign n43442 = n43309 & ~n43441;
  assign n43443 = n43442 ^ n43307;
  assign n43444 = n43443 ^ n43300;
  assign n43445 = ~n43304 & n43444;
  assign n43446 = n43445 ^ n43303;
  assign n43447 = n43446 ^ n43298;
  assign n43448 = ~n43299 & n43447;
  assign n43449 = n43448 ^ n43297;
  assign n43450 = n43449 ^ n43293;
  assign n43451 = n43294 & ~n43450;
  assign n43452 = n43451 ^ n43292;
  assign n43289 = n43254 ^ n43212;
  assign n43453 = n43452 ^ n43289;
  assign n43454 = n41455 ^ n2722;
  assign n43455 = n43454 ^ n37766;
  assign n43456 = n43455 ^ n3223;
  assign n43457 = n43456 ^ n43289;
  assign n43458 = n43453 & ~n43457;
  assign n43459 = n43458 ^ n43456;
  assign n43460 = n43459 ^ n43287;
  assign n43461 = ~n43288 & n43460;
  assign n43462 = n43461 ^ n3227;
  assign n43463 = n43462 ^ n43285;
  assign n43464 = n43286 & ~n43463;
  assign n43465 = n43464 ^ n2862;
  assign n43641 = n43480 ^ n43465;
  assign n43642 = n43484 & ~n43641;
  assign n43643 = n43642 ^ n43483;
  assign n43587 = n43478 & ~n43479;
  assign n43572 = n43477 ^ n43473;
  assign n43573 = n43474 & n43572;
  assign n43574 = n43573 ^ n40128;
  assign n43544 = n41567 ^ n40848;
  assign n43545 = n43544 ^ n42852;
  assign n43540 = n43472 ^ n43469;
  assign n43541 = n43470 & n43540;
  assign n43542 = n43541 ^ n43472;
  assign n43539 = n42935 ^ n42895;
  assign n43543 = n43542 ^ n43539;
  assign n43570 = n43545 ^ n43543;
  assign n43571 = n43570 ^ n40122;
  assign n43586 = n43574 ^ n43571;
  assign n43640 = n43587 ^ n43586;
  assign n43644 = n43643 ^ n43640;
  assign n2958 = n2957 ^ n2894;
  assign n2965 = n2964 ^ n2958;
  assign n2966 = n2965 ^ n1613;
  assign n43645 = n43640 ^ n2966;
  assign n43646 = n43644 & ~n43645;
  assign n43647 = n43646 ^ n2966;
  assign n43588 = n43586 & ~n43587;
  assign n43575 = n43574 ^ n43570;
  assign n43576 = n43571 & ~n43575;
  assign n43577 = n43576 ^ n40122;
  assign n43550 = n41561 ^ n40842;
  assign n43551 = n43550 ^ n42322;
  assign n43546 = n43545 ^ n43539;
  assign n43547 = ~n43543 & ~n43546;
  assign n43548 = n43547 ^ n43545;
  assign n43538 = n42939 ^ n2681;
  assign n43549 = n43548 ^ n43538;
  assign n43568 = n43551 ^ n43549;
  assign n43569 = n43568 ^ n40116;
  assign n43585 = n43577 ^ n43569;
  assign n43639 = n43588 ^ n43585;
  assign n43648 = n43647 ^ n43639;
  assign n43666 = n43651 ^ n43648;
  assign n43815 = n43668 ^ n43666;
  assign n44004 = n43815 ^ n40878;
  assign n44005 = n44003 & n44004;
  assign n43998 = n41698 ^ n2192;
  assign n43999 = n43998 ^ n38116;
  assign n44000 = n43999 ^ n2380;
  assign n44006 = n44005 ^ n44000;
  assign n43652 = n43651 ^ n43639;
  assign n43653 = n43648 & ~n43652;
  assign n43654 = n43653 ^ n43651;
  assign n43578 = n43577 ^ n43568;
  assign n43579 = n43569 & n43578;
  assign n43580 = n43579 ^ n40116;
  assign n43556 = n41559 ^ n40836;
  assign n43557 = n43556 ^ n42327;
  assign n43552 = n43551 ^ n43538;
  assign n43553 = n43549 & ~n43552;
  assign n43554 = n43553 ^ n43551;
  assign n43537 = n42942 ^ n42889;
  assign n43555 = n43554 ^ n43537;
  assign n43566 = n43557 ^ n43555;
  assign n43567 = n43566 ^ n40114;
  assign n43590 = n43580 ^ n43567;
  assign n43589 = ~n43585 & ~n43588;
  assign n43634 = n43590 ^ n43589;
  assign n43638 = n43637 ^ n43634;
  assign n43673 = n43654 ^ n43638;
  assign n43670 = n41749 ^ n41669;
  assign n43671 = n43670 ^ n42633;
  assign n43669 = ~n43666 & n43668;
  assign n43672 = n43671 ^ n43669;
  assign n43818 = n43673 ^ n43672;
  assign n43816 = ~n40878 & ~n43815;
  assign n43817 = n43816 ^ n40438;
  assign n43894 = n43818 ^ n43817;
  assign n44007 = n44005 ^ n43894;
  assign n44008 = n44006 & ~n44007;
  assign n44009 = n44008 ^ n44000;
  assign n43819 = n43818 ^ n43816;
  assign n43820 = ~n43817 & ~n43819;
  assign n43821 = n43820 ^ n40438;
  assign n43679 = n41876 ^ n41745;
  assign n43680 = n43679 ^ n42629;
  assign n43655 = n43654 ^ n43634;
  assign n43656 = n43638 & ~n43655;
  assign n43657 = n43656 ^ n43637;
  assign n43630 = n41433 ^ n33139;
  assign n43631 = n43630 ^ n37744;
  assign n43632 = n43631 ^ n31778;
  assign n43591 = ~n43589 & ~n43590;
  assign n43581 = n43580 ^ n43566;
  assign n43582 = n43567 & ~n43581;
  assign n43583 = n43582 ^ n40114;
  assign n43562 = n41549 ^ n40830;
  assign n43563 = n43562 ^ n42319;
  assign n43558 = n43557 ^ n43537;
  assign n43559 = ~n43555 & ~n43558;
  assign n43560 = n43559 ^ n43557;
  assign n43536 = n42949 ^ n42946;
  assign n43561 = n43560 ^ n43536;
  assign n43564 = n43563 ^ n43561;
  assign n43565 = n43564 ^ n40104;
  assign n43584 = n43583 ^ n43565;
  assign n43629 = n43591 ^ n43584;
  assign n43633 = n43632 ^ n43629;
  assign n43677 = n43657 ^ n43633;
  assign n43674 = n43673 ^ n43671;
  assign n43675 = n43672 & ~n43674;
  assign n43676 = n43675 ^ n43669;
  assign n43678 = n43677 ^ n43676;
  assign n43813 = n43680 ^ n43678;
  assign n43814 = n43813 ^ n40432;
  assign n43893 = n43821 ^ n43814;
  assign n43996 = n43894 ^ n43893;
  assign n2366 = n2344 ^ n2281;
  assign n2382 = n2381 ^ n2366;
  assign n2389 = n2388 ^ n2382;
  assign n43997 = n43996 ^ n2389;
  assign n44130 = n44009 ^ n43997;
  assign n44997 = n42880 ^ n34716;
  assign n44998 = n44997 ^ n39217;
  assign n44999 = n44998 ^ n33149;
  assign n43947 = n42251 ^ n34023;
  assign n43948 = n43947 ^ n38564;
  assign n43949 = n43948 ^ n32386;
  assign n43509 = n43401 ^ n43398;
  assign n43507 = n42657 ^ n41812;
  assign n43508 = n43507 ^ n42606;
  assign n43510 = n43509 ^ n43508;
  assign n43513 = n43394 ^ n43340;
  assign n43511 = n42658 ^ n41814;
  assign n43512 = n43511 ^ n42607;
  assign n43514 = n43513 ^ n43512;
  assign n43517 = n43391 ^ n43388;
  assign n43515 = n42612 ^ n41824;
  assign n43516 = n43515 ^ n42608;
  assign n43518 = n43517 ^ n43516;
  assign n43722 = n43384 ^ n43346;
  assign n43521 = n43381 ^ n43378;
  assign n43519 = n42622 ^ n41731;
  assign n43520 = n43519 ^ n42610;
  assign n43522 = n43521 ^ n43520;
  assign n43712 = n43374 ^ n43352;
  assign n43525 = n43371 ^ n43357;
  assign n43523 = n42595 ^ n41741;
  assign n43524 = n43523 ^ n42616;
  assign n43526 = n43525 ^ n43524;
  assign n43702 = n43368 ^ n43359;
  assign n43529 = n43362 ^ n43223;
  assign n43530 = n43529 ^ n43364;
  assign n43527 = n41747 ^ n41729;
  assign n43528 = n43527 ^ n43039;
  assign n43531 = n43530 ^ n43528;
  assign n43533 = n41753 ^ n41733;
  assign n43534 = n43533 ^ n43032;
  assign n43532 = n43363 ^ n2100;
  assign n43535 = n43534 ^ n43532;
  assign n43681 = n43680 ^ n43677;
  assign n43682 = n43678 & ~n43681;
  assign n43683 = n43682 ^ n43680;
  assign n43658 = n43657 ^ n43629;
  assign n43659 = ~n43633 & n43658;
  assign n43660 = n43659 ^ n43632;
  assign n43625 = n41429 ^ n1924;
  assign n43626 = n43625 ^ n37739;
  assign n43627 = n43626 ^ n31773;
  assign n43600 = n43583 ^ n43564;
  assign n43601 = n43565 & ~n43600;
  assign n43602 = n43601 ^ n40104;
  assign n43595 = n43563 ^ n43536;
  assign n43596 = n43561 & n43595;
  assign n43597 = n43596 ^ n43563;
  assign n43486 = n42952 ^ n42886;
  assign n43598 = n43597 ^ n43486;
  assign n43593 = n41124 ^ n40454;
  assign n43594 = n43593 ^ n42315;
  assign n43599 = n43598 ^ n43594;
  assign n43603 = n43602 ^ n43599;
  assign n43604 = n43603 ^ n39481;
  assign n43592 = ~n43584 & n43591;
  assign n43624 = n43604 ^ n43592;
  assign n43628 = n43627 ^ n43624;
  assign n43665 = n43660 ^ n43628;
  assign n43684 = n43683 ^ n43665;
  assign n43685 = n41762 ^ n41743;
  assign n43686 = n43685 ^ n42627;
  assign n43687 = n43686 ^ n43665;
  assign n43688 = n43684 & ~n43687;
  assign n43689 = n43688 ^ n43686;
  assign n43661 = n43660 ^ n43624;
  assign n43662 = ~n43628 & n43661;
  assign n43663 = n43662 ^ n43627;
  assign n43620 = n41424 ^ n1939;
  assign n43621 = n43620 ^ n37734;
  assign n43622 = n43621 ^ n2083;
  assign n43614 = n43599 ^ n39481;
  assign n43615 = n43603 & ~n43614;
  assign n43616 = n43615 ^ n39481;
  assign n43617 = n43616 ^ n39479;
  assign n43612 = n42955 ^ n42881;
  assign n43608 = n43594 ^ n43486;
  assign n43609 = n43598 & n43608;
  assign n43610 = n43609 ^ n43594;
  assign n43606 = n41624 ^ n40448;
  assign n43607 = n43606 ^ n42314;
  assign n43611 = n43610 ^ n43607;
  assign n43613 = n43612 ^ n43611;
  assign n43618 = n43617 ^ n43613;
  assign n43605 = ~n43592 & ~n43604;
  assign n43619 = n43618 ^ n43605;
  assign n43623 = n43622 ^ n43619;
  assign n43664 = n43663 ^ n43623;
  assign n43690 = n43689 ^ n43664;
  assign n43691 = n41756 ^ n41738;
  assign n43692 = n43691 ^ n42626;
  assign n43693 = n43692 ^ n43664;
  assign n43694 = n43690 & ~n43693;
  assign n43695 = n43694 ^ n43692;
  assign n43696 = n43695 ^ n43532;
  assign n43697 = ~n43535 & ~n43696;
  assign n43698 = n43697 ^ n43534;
  assign n43699 = n43698 ^ n43530;
  assign n43700 = ~n43531 & ~n43699;
  assign n43701 = n43700 ^ n43528;
  assign n43703 = n43702 ^ n43701;
  assign n43704 = n42446 ^ n41850;
  assign n43705 = n43704 ^ n42624;
  assign n43706 = n43705 ^ n43702;
  assign n43707 = n43703 & ~n43706;
  assign n43708 = n43707 ^ n43705;
  assign n43709 = n43708 ^ n43525;
  assign n43710 = ~n43526 & n43709;
  assign n43711 = n43710 ^ n43524;
  assign n43713 = n43712 ^ n43711;
  assign n43714 = n42665 ^ n41736;
  assign n43715 = n43714 ^ n42614;
  assign n43716 = n43715 ^ n43712;
  assign n43717 = n43713 & ~n43716;
  assign n43718 = n43717 ^ n43715;
  assign n43719 = n43718 ^ n43521;
  assign n43720 = ~n43522 & ~n43719;
  assign n43721 = n43720 ^ n43520;
  assign n43723 = n43722 ^ n43721;
  assign n43724 = n42618 ^ n41115;
  assign n43725 = n43724 ^ n42609;
  assign n43726 = n43725 ^ n43722;
  assign n43727 = ~n43723 & n43726;
  assign n43728 = n43727 ^ n43725;
  assign n43729 = n43728 ^ n43517;
  assign n43730 = n43518 & ~n43729;
  assign n43731 = n43730 ^ n43516;
  assign n43732 = n43731 ^ n43513;
  assign n43733 = ~n43514 & ~n43732;
  assign n43734 = n43733 ^ n43512;
  assign n43735 = n43734 ^ n43509;
  assign n43736 = ~n43510 & ~n43735;
  assign n43737 = n43736 ^ n43508;
  assign n43506 = n43408 ^ n43405;
  assign n43738 = n43737 ^ n43506;
  assign n43739 = n42655 ^ n41921;
  assign n43740 = n43739 ^ n42605;
  assign n43741 = n43740 ^ n43506;
  assign n43742 = ~n43738 & n43741;
  assign n43743 = n43742 ^ n43740;
  assign n43504 = n43411 ^ n43333;
  assign n43502 = n43094 ^ n41802;
  assign n43503 = n43502 ^ n42652;
  assign n43505 = n43504 ^ n43503;
  assign n43787 = n43743 ^ n43505;
  assign n43788 = n43787 ^ n41155;
  assign n43789 = n43740 ^ n43738;
  assign n43790 = n43789 ^ n41161;
  assign n43791 = n43734 ^ n43510;
  assign n43792 = n43791 ^ n41168;
  assign n43793 = n43728 ^ n43518;
  assign n43794 = n43793 ^ n41183;
  assign n43795 = n43725 ^ n43723;
  assign n43796 = n43795 ^ n41189;
  assign n43797 = n43718 ^ n43522;
  assign n43798 = n43797 ^ n41195;
  assign n43799 = n43715 ^ n43713;
  assign n43800 = n43799 ^ n41201;
  assign n43801 = n43708 ^ n43526;
  assign n43802 = n43801 ^ n41207;
  assign n43804 = n43698 ^ n43531;
  assign n43805 = n43804 ^ n41109;
  assign n43806 = n43695 ^ n43534;
  assign n43807 = n43806 ^ n43532;
  assign n43808 = n43807 ^ n40971;
  assign n43809 = n43692 ^ n43690;
  assign n43810 = n43809 ^ n40901;
  assign n43811 = n43686 ^ n43684;
  assign n43812 = n43811 ^ n40426;
  assign n43822 = n43821 ^ n43813;
  assign n43823 = ~n43814 & ~n43822;
  assign n43824 = n43823 ^ n40432;
  assign n43825 = n43824 ^ n43811;
  assign n43826 = ~n43812 & n43825;
  assign n43827 = n43826 ^ n40426;
  assign n43828 = n43827 ^ n43809;
  assign n43829 = ~n43810 & n43828;
  assign n43830 = n43829 ^ n40901;
  assign n43831 = n43830 ^ n43807;
  assign n43832 = n43808 & n43831;
  assign n43833 = n43832 ^ n40971;
  assign n43834 = n43833 ^ n43804;
  assign n43835 = ~n43805 & n43834;
  assign n43836 = n43835 ^ n41109;
  assign n43803 = n43705 ^ n43703;
  assign n43837 = n43836 ^ n43803;
  assign n43838 = n43803 ^ n41213;
  assign n43839 = ~n43837 & ~n43838;
  assign n43840 = n43839 ^ n41213;
  assign n43841 = n43840 ^ n43801;
  assign n43842 = ~n43802 & n43841;
  assign n43843 = n43842 ^ n41207;
  assign n43844 = n43843 ^ n43799;
  assign n43845 = ~n43800 & n43844;
  assign n43846 = n43845 ^ n41201;
  assign n43847 = n43846 ^ n43797;
  assign n43848 = n43798 & n43847;
  assign n43849 = n43848 ^ n41195;
  assign n43850 = n43849 ^ n43795;
  assign n43851 = n43796 & ~n43850;
  assign n43852 = n43851 ^ n41189;
  assign n43853 = n43852 ^ n43793;
  assign n43854 = n43794 & ~n43853;
  assign n43855 = n43854 ^ n41183;
  assign n43856 = n43855 ^ n40423;
  assign n43857 = n43731 ^ n43514;
  assign n43858 = n43857 ^ n43855;
  assign n43859 = ~n43856 & n43858;
  assign n43860 = n43859 ^ n40423;
  assign n43861 = n43860 ^ n43791;
  assign n43862 = ~n43792 & n43861;
  assign n43863 = n43862 ^ n41168;
  assign n43864 = n43863 ^ n43789;
  assign n43865 = ~n43790 & n43864;
  assign n43866 = n43865 ^ n41161;
  assign n43867 = n43866 ^ n43787;
  assign n43868 = ~n43788 & n43867;
  assign n43869 = n43868 ^ n41155;
  assign n43744 = n43743 ^ n43504;
  assign n43745 = n43505 & n43744;
  assign n43746 = n43745 ^ n43503;
  assign n43500 = n43414 ^ n43328;
  assign n43498 = n42650 ^ n41796;
  assign n43499 = n43498 ^ n43205;
  assign n43501 = n43500 ^ n43499;
  assign n43785 = n43746 ^ n43501;
  assign n43786 = n43785 ^ n41149;
  assign n43920 = n43869 ^ n43786;
  assign n43888 = n43860 ^ n43792;
  assign n43889 = n43849 ^ n43796;
  assign n43890 = n43846 ^ n43798;
  assign n43891 = n43843 ^ n43800;
  assign n43892 = n43840 ^ n43802;
  assign n43895 = ~n43893 & n43894;
  assign n43896 = n43824 ^ n43812;
  assign n43897 = ~n43895 & ~n43896;
  assign n43898 = n43827 ^ n43810;
  assign n43899 = ~n43897 & n43898;
  assign n43900 = n43830 ^ n43808;
  assign n43901 = ~n43899 & n43900;
  assign n43902 = n43833 ^ n43805;
  assign n43903 = ~n43901 & ~n43902;
  assign n43904 = n43837 ^ n41213;
  assign n43905 = n43903 & ~n43904;
  assign n43906 = n43892 & n43905;
  assign n43907 = ~n43891 & ~n43906;
  assign n43908 = n43890 & n43907;
  assign n43909 = ~n43889 & n43908;
  assign n43910 = n43852 ^ n43794;
  assign n43911 = n43909 & ~n43910;
  assign n43912 = n43857 ^ n40423;
  assign n43913 = n43912 ^ n43855;
  assign n43914 = n43911 & ~n43913;
  assign n43915 = n43888 & ~n43914;
  assign n43916 = n43863 ^ n43790;
  assign n43917 = n43915 & n43916;
  assign n43918 = n43866 ^ n43788;
  assign n43919 = ~n43917 & ~n43918;
  assign n43946 = n43920 ^ n43919;
  assign n43950 = n43949 ^ n43946;
  assign n43951 = n43918 ^ n43917;
  assign n1302 = n1301 ^ n1217;
  assign n1318 = n1317 ^ n1302;
  assign n1325 = n1324 ^ n1318;
  assign n43952 = n43951 ^ n1325;
  assign n43956 = n43916 ^ n43915;
  assign n43953 = n42241 ^ n33961;
  assign n43954 = n43953 ^ n1168;
  assign n43955 = n43954 ^ n1309;
  assign n43957 = n43956 ^ n43955;
  assign n43958 = n43914 ^ n43888;
  assign n1126 = n1116 ^ n1068;
  assign n1151 = n1150 ^ n1126;
  assign n1158 = n1157 ^ n1151;
  assign n43959 = n43958 ^ n1158;
  assign n43960 = n43913 ^ n43911;
  assign n43964 = n43963 ^ n43960;
  assign n43968 = n43910 ^ n43909;
  assign n43965 = n42204 ^ n976;
  assign n43966 = n43965 ^ n38079;
  assign n43967 = n43966 ^ n3330;
  assign n43969 = n43968 ^ n43967;
  assign n43970 = n43908 ^ n43889;
  assign n43974 = n43973 ^ n43970;
  assign n43978 = n43907 ^ n43890;
  assign n43975 = n42214 ^ n33539;
  assign n43976 = n43975 ^ n38088;
  assign n43977 = n43976 ^ n32297;
  assign n43979 = n43978 ^ n43977;
  assign n43984 = n41687 ^ n33478;
  assign n43985 = n43984 ^ n38105;
  assign n43986 = n43985 ^ n32313;
  assign n43983 = n43902 ^ n43901;
  assign n43987 = n43986 ^ n43983;
  assign n43992 = n43898 ^ n43897;
  assign n43989 = n41712 ^ n33489;
  assign n43990 = n43989 ^ n38130;
  assign n43991 = n43990 ^ n32324;
  assign n43993 = n43992 ^ n43991;
  assign n43994 = n43896 ^ n43895;
  assign n2399 = n2362 ^ n2299;
  assign n2400 = n2399 ^ n2396;
  assign n2407 = n2406 ^ n2400;
  assign n43995 = n43994 ^ n2407;
  assign n44010 = n44009 ^ n43996;
  assign n44011 = n43997 & ~n44010;
  assign n44012 = n44011 ^ n2389;
  assign n44013 = n44012 ^ n43994;
  assign n44014 = n43995 & ~n44013;
  assign n44015 = n44014 ^ n2407;
  assign n44016 = n44015 ^ n43992;
  assign n44017 = n43993 & ~n44016;
  assign n44018 = n44017 ^ n43991;
  assign n43988 = n43900 ^ n43899;
  assign n44019 = n44018 ^ n43988;
  assign n44020 = n41692 ^ n33483;
  assign n44021 = n44020 ^ n38109;
  assign n44022 = n44021 ^ n32319;
  assign n44023 = n44022 ^ n43988;
  assign n44024 = n44019 & ~n44023;
  assign n44025 = n44024 ^ n44022;
  assign n44026 = n44025 ^ n43983;
  assign n44027 = ~n43987 & n44026;
  assign n44028 = n44027 ^ n43986;
  assign n43982 = n43904 ^ n43903;
  assign n44029 = n44028 ^ n43982;
  assign n44030 = n41681 ^ n33473;
  assign n44031 = n44030 ^ n38099;
  assign n44032 = n44031 ^ n32308;
  assign n44033 = n44032 ^ n43982;
  assign n44034 = ~n44029 & n44033;
  assign n44035 = n44034 ^ n44032;
  assign n43981 = n43905 ^ n43892;
  assign n44036 = n44035 ^ n43981;
  assign n44037 = n41676 ^ n33469;
  assign n44038 = n44037 ^ n38094;
  assign n44039 = n44038 ^ n723;
  assign n44040 = n44039 ^ n43981;
  assign n44041 = n44036 & ~n44040;
  assign n44042 = n44041 ^ n44039;
  assign n43980 = n43906 ^ n43891;
  assign n44043 = n44042 ^ n43980;
  assign n44044 = n41119 ^ n33464;
  assign n44045 = n44044 ^ n38149;
  assign n44046 = n44045 ^ n32301;
  assign n44047 = n44046 ^ n43980;
  assign n44048 = ~n44043 & n44047;
  assign n44049 = n44048 ^ n44046;
  assign n44050 = n44049 ^ n43978;
  assign n44051 = n43979 & ~n44050;
  assign n44052 = n44051 ^ n43977;
  assign n44053 = n44052 ^ n43970;
  assign n44054 = ~n43974 & n44053;
  assign n44055 = n44054 ^ n43973;
  assign n44056 = n44055 ^ n43968;
  assign n44057 = ~n43969 & n44056;
  assign n44058 = n44057 ^ n43967;
  assign n44059 = n44058 ^ n43960;
  assign n44060 = ~n43964 & n44059;
  assign n44061 = n44060 ^ n43963;
  assign n44062 = n44061 ^ n43958;
  assign n44063 = n43959 & ~n44062;
  assign n44064 = n44063 ^ n1158;
  assign n44065 = n44064 ^ n43956;
  assign n44066 = ~n43957 & n44065;
  assign n44067 = n44066 ^ n43955;
  assign n44068 = n44067 ^ n43951;
  assign n44069 = n43952 & ~n44068;
  assign n44070 = n44069 ^ n1325;
  assign n44071 = n44070 ^ n43949;
  assign n44072 = n43950 & ~n44071;
  assign n44073 = n44072 ^ n43946;
  assign n43942 = n42192 ^ n34018;
  assign n43943 = n43942 ^ n38540;
  assign n43944 = n43943 ^ n32380;
  assign n43921 = ~n43919 & n43920;
  assign n43870 = n43869 ^ n43785;
  assign n43871 = ~n43786 & n43870;
  assign n43872 = n43871 ^ n41149;
  assign n43751 = n42646 ^ n41790;
  assign n43752 = n43751 ^ n43261;
  assign n43747 = n43746 ^ n43500;
  assign n43748 = ~n43501 & n43747;
  assign n43749 = n43748 ^ n43499;
  assign n43497 = n43417 ^ n43326;
  assign n43750 = n43749 ^ n43497;
  assign n43783 = n43752 ^ n43750;
  assign n43784 = n43783 ^ n41143;
  assign n43887 = n43872 ^ n43784;
  assign n43941 = n43921 ^ n43887;
  assign n43945 = n43944 ^ n43941;
  assign n44782 = n44073 ^ n43945;
  assign n44755 = n43536 ^ n42733;
  assign n44172 = n43456 ^ n43453;
  assign n44756 = n44755 ^ n44172;
  assign n44696 = n44070 ^ n43950;
  assign n44757 = n44756 ^ n44696;
  assign n44758 = n43537 ^ n42642;
  assign n44165 = n43449 ^ n43294;
  assign n44759 = n44758 ^ n44165;
  assign n44701 = n44067 ^ n43952;
  assign n44760 = n44759 ^ n44701;
  assign n44761 = n43539 ^ n42714;
  assign n44154 = n43443 ^ n43304;
  assign n44762 = n44761 ^ n44154;
  assign n44711 = n44061 ^ n43959;
  assign n44763 = n44762 ^ n44711;
  assign n44412 = n44055 ^ n43969;
  assign n44405 = n44052 ^ n43974;
  assign n44392 = n44046 ^ n44043;
  assign n44385 = n44039 ^ n44036;
  assign n44378 = n44032 ^ n44029;
  assign n44371 = n44025 ^ n43987;
  assign n44123 = n44022 ^ n44019;
  assign n44121 = n42622 ^ n42608;
  assign n44122 = n44121 ^ n43506;
  assign n44124 = n44123 ^ n44122;
  assign n44128 = n44012 ^ n43995;
  assign n44126 = n42610 ^ n42595;
  assign n44127 = n44126 ^ n43513;
  assign n44129 = n44128 ^ n44127;
  assign n44133 = n44000 ^ n43894;
  assign n44134 = n44133 ^ n44005;
  assign n44131 = n42616 ^ n41729;
  assign n44132 = n44131 ^ n43722;
  assign n44135 = n44134 ^ n44132;
  assign n44138 = n44004 ^ n44003;
  assign n44136 = n42624 ^ n41733;
  assign n44137 = n44136 ^ n43521;
  assign n44139 = n44138 ^ n44137;
  assign n44308 = n42150 ^ n33935;
  assign n44309 = n44308 ^ n38497;
  assign n44310 = n44309 ^ n1832;
  assign n44150 = n43446 ^ n43299;
  assign n44148 = n42322 ^ n41577;
  assign n44149 = n44148 ^ n43486;
  assign n44151 = n44150 ^ n44149;
  assign n44152 = n42852 ^ n42135;
  assign n44153 = n44152 ^ n43536;
  assign n44155 = n44154 ^ n44153;
  assign n44105 = n43440 ^ n43309;
  assign n43772 = n42733 ^ n41770;
  assign n43773 = n43772 ^ n43538;
  assign n43771 = n43437 ^ n43434;
  assign n43774 = n43773 ^ n43771;
  assign n43495 = n43420 ^ n43321;
  assign n43493 = n42714 ^ n41788;
  assign n43494 = n43493 ^ n43271;
  assign n43496 = n43495 ^ n43494;
  assign n43753 = n43752 ^ n43497;
  assign n43754 = n43750 & ~n43753;
  assign n43755 = n43754 ^ n43752;
  assign n43756 = n43755 ^ n43495;
  assign n43757 = ~n43496 & ~n43756;
  assign n43758 = n43757 ^ n43494;
  assign n43492 = n43423 ^ n43316;
  assign n43759 = n43758 ^ n43492;
  assign n43760 = n43469 ^ n41782;
  assign n43761 = n43760 ^ n42643;
  assign n43762 = n43761 ^ n43492;
  assign n43763 = n43759 & ~n43762;
  assign n43764 = n43763 ^ n43761;
  assign n43491 = n43430 ^ n43427;
  assign n43765 = n43764 ^ n43491;
  assign n43766 = n42642 ^ n41772;
  assign n43767 = n43766 ^ n43539;
  assign n43768 = n43767 ^ n43491;
  assign n43769 = ~n43765 & n43768;
  assign n43770 = n43769 ^ n43767;
  assign n44102 = n43773 ^ n43770;
  assign n44103 = n43774 & ~n44102;
  assign n44104 = n44103 ^ n43771;
  assign n44106 = n44105 ^ n44104;
  assign n44100 = n42641 ^ n41951;
  assign n44101 = n44100 ^ n43537;
  assign n44156 = n44105 ^ n44101;
  assign n44157 = n44106 & n44156;
  assign n44158 = n44157 ^ n44101;
  assign n44159 = n44158 ^ n44154;
  assign n44160 = ~n44155 & n44159;
  assign n44161 = n44160 ^ n44153;
  assign n44162 = n44161 ^ n44150;
  assign n44163 = ~n44151 & n44162;
  assign n44164 = n44163 ^ n44149;
  assign n44166 = n44165 ^ n44164;
  assign n44167 = n43612 ^ n41567;
  assign n44168 = n44167 ^ n42327;
  assign n44169 = n44168 ^ n44165;
  assign n44170 = ~n44166 & n44169;
  assign n44171 = n44170 ^ n44168;
  assign n44173 = n44172 ^ n44171;
  assign n44174 = n42982 ^ n42319;
  assign n44175 = n44174 ^ n41561;
  assign n44176 = n44175 ^ n44172;
  assign n44177 = n44173 & ~n44176;
  assign n44178 = n44177 ^ n44175;
  assign n44145 = n42315 ^ n41559;
  assign n44146 = n44145 ^ n42989;
  assign n44144 = n43459 ^ n43288;
  assign n44147 = n44146 ^ n44144;
  assign n44214 = n44178 ^ n44147;
  assign n44215 = n44214 ^ n40836;
  assign n44191 = n44175 ^ n44173;
  assign n44192 = n44191 ^ n40842;
  assign n44193 = n44168 ^ n44166;
  assign n44194 = n44193 ^ n40848;
  assign n44195 = n44161 ^ n44151;
  assign n44196 = n44195 ^ n40858;
  assign n44197 = n44158 ^ n44155;
  assign n44198 = n44197 ^ n41405;
  assign n44107 = n44106 ^ n44101;
  assign n44108 = n44107 ^ n41389;
  assign n43777 = n43767 ^ n43765;
  assign n43778 = n43777 ^ n41126;
  assign n43779 = n43761 ^ n43759;
  assign n43780 = n43779 ^ n41135;
  assign n43781 = n43755 ^ n43496;
  assign n43782 = n43781 ^ n41137;
  assign n43873 = n43872 ^ n43783;
  assign n43874 = ~n43784 & n43873;
  assign n43875 = n43874 ^ n41143;
  assign n43876 = n43875 ^ n43781;
  assign n43877 = ~n43782 & n43876;
  assign n43878 = n43877 ^ n41137;
  assign n43879 = n43878 ^ n43779;
  assign n43880 = n43780 & ~n43879;
  assign n43881 = n43880 ^ n41135;
  assign n43882 = n43881 ^ n43777;
  assign n43883 = ~n43778 & n43882;
  assign n43884 = n43883 ^ n41126;
  assign n44096 = n43884 ^ n41372;
  assign n43775 = n43774 ^ n43770;
  assign n44097 = n43884 ^ n43775;
  assign n44098 = ~n44096 & n44097;
  assign n44099 = n44098 ^ n41372;
  assign n44199 = n44107 ^ n44099;
  assign n44200 = n44108 & ~n44199;
  assign n44201 = n44200 ^ n41389;
  assign n44202 = n44201 ^ n44197;
  assign n44203 = n44198 & ~n44202;
  assign n44204 = n44203 ^ n41405;
  assign n44205 = n44204 ^ n44195;
  assign n44206 = ~n44196 & ~n44205;
  assign n44207 = n44206 ^ n40858;
  assign n44208 = n44207 ^ n44193;
  assign n44209 = n44194 & ~n44208;
  assign n44210 = n44209 ^ n40848;
  assign n44211 = n44210 ^ n44191;
  assign n44212 = ~n44192 & n44211;
  assign n44213 = n44212 ^ n40842;
  assign n44229 = n44214 ^ n44213;
  assign n44230 = n44215 & ~n44229;
  assign n44231 = n44230 ^ n40836;
  assign n44183 = n42314 ^ n41549;
  assign n44184 = n44183 ^ n42981;
  assign n44179 = n44178 ^ n44144;
  assign n44180 = n44147 & n44179;
  assign n44181 = n44180 ^ n44146;
  assign n44143 = n43462 ^ n43286;
  assign n44182 = n44181 ^ n44143;
  assign n44227 = n44184 ^ n44182;
  assign n44228 = n44227 ^ n40830;
  assign n44232 = n44231 ^ n44228;
  assign n44216 = n44215 ^ n44213;
  assign n44217 = n44201 ^ n44198;
  assign n44109 = n44108 ^ n44099;
  assign n43776 = n43775 ^ n41372;
  assign n43885 = n43884 ^ n43776;
  assign n43886 = n43878 ^ n43780;
  assign n43922 = ~n43887 & ~n43921;
  assign n43923 = n43875 ^ n43782;
  assign n43924 = n43922 & ~n43923;
  assign n43925 = n43886 & n43924;
  assign n43926 = n43881 ^ n43778;
  assign n43927 = ~n43925 & n43926;
  assign n44110 = ~n43885 & n43927;
  assign n44218 = ~n44109 & ~n44110;
  assign n44219 = ~n44217 & n44218;
  assign n44220 = n44204 ^ n44196;
  assign n44221 = ~n44219 & ~n44220;
  assign n44222 = n44207 ^ n44194;
  assign n44223 = ~n44221 & n44222;
  assign n44224 = n44210 ^ n44192;
  assign n44225 = ~n44223 & n44224;
  assign n44226 = n44216 & ~n44225;
  assign n44259 = n44232 ^ n44226;
  assign n44256 = n42300 ^ n33940;
  assign n44257 = n44256 ^ n1745;
  assign n44258 = n44257 ^ n32485;
  assign n44260 = n44259 ^ n44258;
  assign n44264 = n44225 ^ n44216;
  assign n44261 = n42293 ^ n33944;
  assign n44262 = n44261 ^ n38504;
  assign n44263 = n44262 ^ n1744;
  assign n44265 = n44264 ^ n44263;
  assign n44267 = n3010 ^ n1655;
  assign n44268 = n44267 ^ n38509;
  assign n44269 = n44268 ^ n32233;
  assign n44266 = n44224 ^ n44223;
  assign n44270 = n44269 ^ n44266;
  assign n44275 = n44218 ^ n44217;
  assign n44279 = n44278 ^ n44275;
  assign n44111 = n44110 ^ n44109;
  assign n44093 = n38525 ^ n3235;
  assign n44094 = n44093 ^ n42170;
  assign n44095 = n44094 ^ n3101;
  assign n44112 = n44111 ^ n44095;
  assign n43928 = n43927 ^ n43885;
  assign n43488 = n42175 ^ n34002;
  assign n43489 = n43488 ^ n3083;
  assign n43490 = n43489 ^ n2645;
  assign n43929 = n43928 ^ n43490;
  assign n43933 = n43926 ^ n43925;
  assign n43930 = n42180 ^ n34007;
  assign n43931 = n43930 ^ n2573;
  assign n43932 = n43931 ^ n3081;
  assign n43934 = n43933 ^ n43932;
  assign n43938 = n43924 ^ n43886;
  assign n43935 = n42185 ^ n3059;
  assign n43936 = n43935 ^ n38533;
  assign n43937 = n43936 ^ n2565;
  assign n43939 = n43938 ^ n43937;
  assign n44074 = n44073 ^ n43941;
  assign n44075 = n43945 & ~n44074;
  assign n44076 = n44075 ^ n43944;
  assign n43940 = n43923 ^ n43922;
  assign n44077 = n44076 ^ n43940;
  assign n44078 = n42261 ^ n2492;
  assign n44079 = n44078 ^ n38574;
  assign n44080 = n44079 ^ n3167;
  assign n44081 = n44080 ^ n43940;
  assign n44082 = n44077 & ~n44081;
  assign n44083 = n44082 ^ n44080;
  assign n44084 = n44083 ^ n43938;
  assign n44085 = n43939 & ~n44084;
  assign n44086 = n44085 ^ n43937;
  assign n44087 = n44086 ^ n43933;
  assign n44088 = n43934 & ~n44087;
  assign n44089 = n44088 ^ n43932;
  assign n44090 = n44089 ^ n43928;
  assign n44091 = n43929 & ~n44090;
  assign n44092 = n44091 ^ n43490;
  assign n44280 = n44111 ^ n44092;
  assign n44281 = n44112 & ~n44280;
  assign n44282 = n44281 ^ n44095;
  assign n44283 = n44282 ^ n44278;
  assign n44284 = ~n44279 & ~n44283;
  assign n44285 = n44284 ^ n44275;
  assign n44274 = n44220 ^ n44219;
  assign n44286 = n44285 ^ n44274;
  assign n44287 = n42160 ^ n2930;
  assign n44288 = n44287 ^ n38515;
  assign n44289 = n44288 ^ n32242;
  assign n44290 = n44289 ^ n44274;
  assign n44291 = ~n44286 & ~n44290;
  assign n44292 = n44291 ^ n44289;
  assign n44271 = n33951 ^ n2995;
  assign n44272 = n44271 ^ n38599;
  assign n44273 = n44272 ^ n32238;
  assign n44293 = n44292 ^ n44273;
  assign n44294 = n44222 ^ n44221;
  assign n44295 = n44294 ^ n44292;
  assign n44296 = n44293 & n44295;
  assign n44297 = n44296 ^ n44273;
  assign n44298 = n44297 ^ n44266;
  assign n44299 = n44270 & ~n44298;
  assign n44300 = n44299 ^ n44269;
  assign n44301 = n44300 ^ n44264;
  assign n44302 = ~n44265 & n44301;
  assign n44303 = n44302 ^ n44263;
  assign n44304 = n44303 ^ n44259;
  assign n44305 = ~n44260 & n44304;
  assign n44306 = n44305 ^ n44258;
  assign n44236 = n44231 ^ n44227;
  assign n44237 = ~n44228 & n44236;
  assign n44238 = n44237 ^ n40830;
  assign n44185 = n44184 ^ n44143;
  assign n44186 = n44182 & n44185;
  assign n44187 = n44186 ^ n44184;
  assign n44140 = n41764 ^ n41124;
  assign n44141 = n44140 ^ n42979;
  assign n43485 = n43484 ^ n43465;
  assign n44142 = n44141 ^ n43485;
  assign n44234 = n44187 ^ n44142;
  assign n44235 = n44234 ^ n40454;
  assign n44239 = n44238 ^ n44235;
  assign n44233 = n44226 & ~n44232;
  assign n44255 = n44239 ^ n44233;
  assign n44307 = n44306 ^ n44255;
  assign n44317 = n44310 ^ n44307;
  assign n44315 = n43032 ^ n41743;
  assign n44316 = n44315 ^ n43525;
  assign n44318 = n44317 ^ n44316;
  assign n44321 = n44303 ^ n44258;
  assign n44322 = n44321 ^ n44259;
  assign n44319 = n43702 ^ n42626;
  assign n44320 = n44319 ^ n41745;
  assign n44323 = n44322 ^ n44320;
  assign n44328 = n42627 ^ n41749;
  assign n44329 = n44328 ^ n43530;
  assign n44324 = n44297 ^ n44270;
  assign n44325 = n42629 ^ n41751;
  assign n44326 = n44325 ^ n43532;
  assign n44327 = n44324 & ~n44326;
  assign n44330 = n44329 ^ n44327;
  assign n44331 = n44300 ^ n44265;
  assign n44332 = n44331 ^ n44329;
  assign n44333 = n44330 & n44332;
  assign n44334 = n44333 ^ n44327;
  assign n44335 = n44334 ^ n44322;
  assign n44336 = ~n44323 & n44335;
  assign n44337 = n44336 ^ n44320;
  assign n44338 = n44337 ^ n44317;
  assign n44339 = ~n44318 & n44338;
  assign n44340 = n44339 ^ n44316;
  assign n44311 = n44310 ^ n44255;
  assign n44312 = n44307 & ~n44311;
  assign n44313 = n44312 ^ n44310;
  assign n44250 = n44238 ^ n44234;
  assign n44251 = n44235 & ~n44250;
  assign n44252 = n44251 ^ n40454;
  assign n44246 = n43644 ^ n2966;
  assign n44241 = n42146 ^ n34106;
  assign n44242 = n44241 ^ n38492;
  assign n44243 = n44242 ^ n32748;
  assign n44240 = ~n44233 & ~n44239;
  assign n44244 = n44243 ^ n44240;
  assign n44245 = n44244 ^ n43606;
  assign n44247 = n44246 ^ n44245;
  assign n44248 = n44247 ^ n41759;
  assign n44188 = n44187 ^ n43485;
  assign n44189 = n44142 & ~n44188;
  assign n44190 = n44189 ^ n44141;
  assign n44249 = n44248 ^ n44190;
  assign n44253 = n44252 ^ n44249;
  assign n44254 = n44253 ^ n42976;
  assign n44314 = n44313 ^ n44254;
  assign n44341 = n44340 ^ n44314;
  assign n44342 = n43039 ^ n41738;
  assign n44343 = n44342 ^ n43712;
  assign n44344 = n44343 ^ n44314;
  assign n44345 = ~n44341 & n44344;
  assign n44346 = n44345 ^ n44343;
  assign n44347 = n44346 ^ n44138;
  assign n44348 = n44139 & ~n44347;
  assign n44349 = n44348 ^ n44137;
  assign n44350 = n44349 ^ n44134;
  assign n44351 = n44135 & ~n44350;
  assign n44352 = n44351 ^ n44132;
  assign n44353 = n44352 ^ n44130;
  assign n44354 = n42614 ^ n42446;
  assign n44355 = n44354 ^ n43517;
  assign n44356 = n44355 ^ n44130;
  assign n44357 = ~n44353 & ~n44356;
  assign n44358 = n44357 ^ n44355;
  assign n44359 = n44358 ^ n44128;
  assign n44360 = n44129 & n44359;
  assign n44361 = n44360 ^ n44127;
  assign n44125 = n44015 ^ n43993;
  assign n44362 = n44361 ^ n44125;
  assign n44363 = n42665 ^ n42609;
  assign n44364 = n44363 ^ n43509;
  assign n44365 = n44364 ^ n44125;
  assign n44366 = ~n44362 & ~n44365;
  assign n44367 = n44366 ^ n44364;
  assign n44368 = n44367 ^ n44123;
  assign n44369 = ~n44124 & ~n44368;
  assign n44370 = n44369 ^ n44122;
  assign n44372 = n44371 ^ n44370;
  assign n44373 = n42618 ^ n42607;
  assign n44374 = n44373 ^ n43504;
  assign n44375 = n44374 ^ n44371;
  assign n44376 = n44372 & ~n44375;
  assign n44377 = n44376 ^ n44374;
  assign n44379 = n44378 ^ n44377;
  assign n44380 = n42612 ^ n42606;
  assign n44381 = n44380 ^ n43500;
  assign n44382 = n44381 ^ n44378;
  assign n44383 = ~n44379 & n44382;
  assign n44384 = n44383 ^ n44381;
  assign n44386 = n44385 ^ n44384;
  assign n44387 = n42658 ^ n42605;
  assign n44388 = n44387 ^ n43497;
  assign n44389 = n44388 ^ n44385;
  assign n44390 = n44386 & ~n44389;
  assign n44391 = n44390 ^ n44388;
  assign n44393 = n44392 ^ n44391;
  assign n44394 = n43094 ^ n42657;
  assign n44395 = n44394 ^ n43495;
  assign n44396 = n44395 ^ n44392;
  assign n44397 = ~n44393 & n44396;
  assign n44398 = n44397 ^ n44395;
  assign n44120 = n44049 ^ n43979;
  assign n44399 = n44398 ^ n44120;
  assign n44400 = n43205 ^ n42655;
  assign n44401 = n44400 ^ n43492;
  assign n44402 = n44401 ^ n44120;
  assign n44403 = ~n44399 & n44402;
  assign n44404 = n44403 ^ n44401;
  assign n44406 = n44405 ^ n44404;
  assign n44407 = n43261 ^ n42652;
  assign n44408 = n44407 ^ n43491;
  assign n44409 = n44408 ^ n44405;
  assign n44410 = n44406 & ~n44409;
  assign n44411 = n44410 ^ n44408;
  assign n44413 = n44412 ^ n44411;
  assign n44118 = n43271 ^ n42650;
  assign n44119 = n44118 ^ n43771;
  assign n44504 = n44412 ^ n44119;
  assign n44505 = n44413 & ~n44504;
  assign n44506 = n44505 ^ n44119;
  assign n44503 = n44058 ^ n43964;
  assign n44507 = n44506 ^ n44503;
  assign n44501 = n43469 ^ n42646;
  assign n44502 = n44501 ^ n44105;
  assign n44764 = n44503 ^ n44502;
  assign n44765 = n44507 & n44764;
  assign n44766 = n44765 ^ n44502;
  assign n44767 = n44766 ^ n44711;
  assign n44768 = n44763 & n44767;
  assign n44769 = n44768 ^ n44762;
  assign n44706 = n44064 ^ n43957;
  assign n44770 = n44769 ^ n44706;
  assign n44771 = n43538 ^ n42643;
  assign n44772 = n44771 ^ n44150;
  assign n44773 = n44772 ^ n44706;
  assign n44774 = n44770 & ~n44773;
  assign n44775 = n44774 ^ n44772;
  assign n44776 = n44775 ^ n44701;
  assign n44777 = ~n44760 & ~n44776;
  assign n44778 = n44777 ^ n44759;
  assign n44779 = n44778 ^ n44696;
  assign n44780 = ~n44757 & n44779;
  assign n44781 = n44780 ^ n44756;
  assign n44783 = n44782 ^ n44781;
  assign n44784 = n43486 ^ n42641;
  assign n44785 = n44784 ^ n44144;
  assign n44786 = n44785 ^ n44782;
  assign n44787 = n44783 & ~n44786;
  assign n44788 = n44787 ^ n44785;
  assign n44753 = n44080 ^ n44077;
  assign n44751 = n43612 ^ n42852;
  assign n44752 = n44751 ^ n44143;
  assign n44754 = n44753 ^ n44752;
  assign n44834 = n44788 ^ n44754;
  assign n44835 = n44834 ^ n42135;
  assign n44836 = n44785 ^ n44783;
  assign n44837 = n44836 ^ n41951;
  assign n44838 = n44778 ^ n44757;
  assign n44839 = n44838 ^ n41770;
  assign n44840 = n44775 ^ n44760;
  assign n44841 = n44840 ^ n41772;
  assign n44842 = n44772 ^ n44770;
  assign n44843 = n44842 ^ n41782;
  assign n44844 = n44766 ^ n44763;
  assign n44845 = n44844 ^ n41788;
  assign n44508 = n44507 ^ n44502;
  assign n44509 = n44508 ^ n41790;
  assign n44414 = n44413 ^ n44119;
  assign n44415 = n44414 ^ n41796;
  assign n44416 = n44408 ^ n44406;
  assign n44417 = n44416 ^ n41802;
  assign n44418 = n44401 ^ n44399;
  assign n44419 = n44418 ^ n41921;
  assign n44420 = n44395 ^ n44393;
  assign n44421 = n44420 ^ n41812;
  assign n44422 = n44388 ^ n44386;
  assign n44423 = n44422 ^ n41814;
  assign n44424 = n44381 ^ n44379;
  assign n44425 = n44424 ^ n41824;
  assign n44426 = n44374 ^ n44372;
  assign n44427 = n44426 ^ n41115;
  assign n44428 = n44367 ^ n44124;
  assign n44429 = n44428 ^ n41731;
  assign n44430 = n44364 ^ n44362;
  assign n44431 = n44430 ^ n41736;
  assign n44432 = n44358 ^ n44129;
  assign n44433 = n44432 ^ n41741;
  assign n44434 = n44355 ^ n44353;
  assign n44435 = n44434 ^ n41850;
  assign n44436 = n44349 ^ n44135;
  assign n44437 = n44436 ^ n41747;
  assign n44438 = n44346 ^ n44139;
  assign n44439 = n44438 ^ n41753;
  assign n44440 = n44343 ^ n44341;
  assign n44441 = n44440 ^ n41756;
  assign n44442 = n44337 ^ n44318;
  assign n44443 = n44442 ^ n41762;
  assign n44444 = n44334 ^ n44323;
  assign n44445 = n44444 ^ n41876;
  assign n44446 = n44326 ^ n44324;
  assign n44447 = n41644 & ~n44446;
  assign n44448 = n44447 ^ n41669;
  assign n44449 = n44331 ^ n44330;
  assign n44450 = n44449 ^ n44447;
  assign n44451 = ~n44448 & n44450;
  assign n44452 = n44451 ^ n41669;
  assign n44453 = n44452 ^ n44444;
  assign n44454 = ~n44445 & ~n44453;
  assign n44455 = n44454 ^ n41876;
  assign n44456 = n44455 ^ n44442;
  assign n44457 = ~n44443 & n44456;
  assign n44458 = n44457 ^ n41762;
  assign n44459 = n44458 ^ n44440;
  assign n44460 = ~n44441 & ~n44459;
  assign n44461 = n44460 ^ n41756;
  assign n44462 = n44461 ^ n44438;
  assign n44463 = ~n44439 & n44462;
  assign n44464 = n44463 ^ n41753;
  assign n44465 = n44464 ^ n44436;
  assign n44466 = ~n44437 & n44465;
  assign n44467 = n44466 ^ n41747;
  assign n44468 = n44467 ^ n44434;
  assign n44469 = n44435 & ~n44468;
  assign n44470 = n44469 ^ n41850;
  assign n44471 = n44470 ^ n44432;
  assign n44472 = ~n44433 & ~n44471;
  assign n44473 = n44472 ^ n41741;
  assign n44474 = n44473 ^ n44430;
  assign n44475 = ~n44431 & n44474;
  assign n44476 = n44475 ^ n41736;
  assign n44477 = n44476 ^ n44428;
  assign n44478 = n44429 & ~n44477;
  assign n44479 = n44478 ^ n41731;
  assign n44480 = n44479 ^ n44426;
  assign n44481 = n44427 & n44480;
  assign n44482 = n44481 ^ n41115;
  assign n44483 = n44482 ^ n44424;
  assign n44484 = ~n44425 & n44483;
  assign n44485 = n44484 ^ n41824;
  assign n44486 = n44485 ^ n44422;
  assign n44487 = n44423 & ~n44486;
  assign n44488 = n44487 ^ n41814;
  assign n44489 = n44488 ^ n44420;
  assign n44490 = n44421 & n44489;
  assign n44491 = n44490 ^ n41812;
  assign n44492 = n44491 ^ n44418;
  assign n44493 = ~n44419 & ~n44492;
  assign n44494 = n44493 ^ n41921;
  assign n44495 = n44494 ^ n44416;
  assign n44496 = ~n44417 & ~n44495;
  assign n44497 = n44496 ^ n41802;
  assign n44498 = n44497 ^ n44414;
  assign n44499 = ~n44415 & n44498;
  assign n44500 = n44499 ^ n41796;
  assign n44846 = n44508 ^ n44500;
  assign n44847 = ~n44509 & ~n44846;
  assign n44848 = n44847 ^ n41790;
  assign n44849 = n44848 ^ n44844;
  assign n44850 = n44845 & ~n44849;
  assign n44851 = n44850 ^ n41788;
  assign n44852 = n44851 ^ n44842;
  assign n44853 = ~n44843 & ~n44852;
  assign n44854 = n44853 ^ n41782;
  assign n44855 = n44854 ^ n44840;
  assign n44856 = n44841 & n44855;
  assign n44857 = n44856 ^ n41772;
  assign n44858 = n44857 ^ n44838;
  assign n44859 = n44839 & n44858;
  assign n44860 = n44859 ^ n41770;
  assign n44861 = n44860 ^ n44836;
  assign n44862 = ~n44837 & ~n44861;
  assign n44863 = n44862 ^ n41951;
  assign n44864 = n44863 ^ n44834;
  assign n44865 = n44835 & ~n44864;
  assign n44866 = n44865 ^ n42135;
  assign n44789 = n44788 ^ n44753;
  assign n44790 = n44754 & ~n44789;
  assign n44791 = n44790 ^ n44752;
  assign n44749 = n44083 ^ n43939;
  assign n44747 = n42982 ^ n42322;
  assign n44748 = n44747 ^ n43485;
  assign n44750 = n44749 ^ n44748;
  assign n44832 = n44791 ^ n44750;
  assign n44833 = n44832 ^ n41577;
  assign n44886 = n44866 ^ n44833;
  assign n44887 = n44860 ^ n44837;
  assign n44888 = n44857 ^ n44839;
  assign n44889 = n44848 ^ n44845;
  assign n44510 = n44509 ^ n44500;
  assign n44511 = n44497 ^ n44415;
  assign n44512 = n44479 ^ n44427;
  assign n44513 = n44467 ^ n44435;
  assign n44514 = n44461 ^ n44439;
  assign n44515 = n44458 ^ n44441;
  assign n44516 = n44455 ^ n44443;
  assign n44517 = n44449 ^ n44448;
  assign n44518 = n44452 ^ n44445;
  assign n44519 = ~n44517 & ~n44518;
  assign n44520 = ~n44516 & ~n44519;
  assign n44521 = n44515 & ~n44520;
  assign n44522 = n44514 & ~n44521;
  assign n44523 = n44464 ^ n44437;
  assign n44524 = ~n44522 & ~n44523;
  assign n44525 = n44513 & n44524;
  assign n44526 = n44470 ^ n44433;
  assign n44527 = n44525 & ~n44526;
  assign n44528 = n44473 ^ n44431;
  assign n44529 = ~n44527 & ~n44528;
  assign n44530 = n44476 ^ n44429;
  assign n44531 = n44529 & n44530;
  assign n44532 = n44512 & n44531;
  assign n44533 = n44482 ^ n44425;
  assign n44534 = n44532 & n44533;
  assign n44535 = n44485 ^ n44423;
  assign n44536 = n44534 & ~n44535;
  assign n44537 = n44488 ^ n41812;
  assign n44538 = n44537 ^ n44420;
  assign n44539 = ~n44536 & n44538;
  assign n44540 = n44491 ^ n41921;
  assign n44541 = n44540 ^ n44418;
  assign n44542 = n44539 & n44541;
  assign n44543 = n44494 ^ n44417;
  assign n44544 = ~n44542 & n44543;
  assign n44545 = n44511 & ~n44544;
  assign n44890 = ~n44510 & ~n44545;
  assign n44891 = ~n44889 & n44890;
  assign n44892 = n44851 ^ n44843;
  assign n44893 = n44891 & n44892;
  assign n44894 = n44854 ^ n44841;
  assign n44895 = ~n44893 & ~n44894;
  assign n44896 = n44888 & n44895;
  assign n44897 = ~n44887 & ~n44896;
  assign n44898 = n44863 ^ n44835;
  assign n44899 = n44897 & ~n44898;
  assign n44900 = ~n44886 & ~n44899;
  assign n44867 = n44866 ^ n44832;
  assign n44868 = ~n44833 & ~n44867;
  assign n44869 = n44868 ^ n41577;
  assign n44796 = n42989 ^ n42327;
  assign n44797 = n44796 ^ n44246;
  assign n44792 = n44791 ^ n44749;
  assign n44793 = n44750 & n44792;
  assign n44794 = n44793 ^ n44748;
  assign n44692 = n44086 ^ n43934;
  assign n44795 = n44794 ^ n44692;
  assign n44830 = n44797 ^ n44795;
  assign n44831 = n44830 ^ n41567;
  assign n44885 = n44869 ^ n44831;
  assign n44935 = n44900 ^ n44885;
  assign n44939 = n44938 ^ n44935;
  assign n44941 = n42949 ^ n34726;
  assign n44942 = n44941 ^ n2828;
  assign n44943 = n44942 ^ n33156;
  assign n44940 = n44899 ^ n44886;
  assign n44944 = n44943 ^ n44940;
  assign n44946 = n44896 ^ n44887;
  assign n2703 = n2702 ^ n2681;
  assign n2731 = n2730 ^ n2703;
  assign n2738 = n2737 ^ n2731;
  assign n44947 = n44946 ^ n2738;
  assign n44952 = n44894 ^ n44893;
  assign n44949 = n42899 ^ n2616;
  assign n44950 = n44949 ^ n39301;
  assign n44951 = n44950 ^ n3201;
  assign n44953 = n44952 ^ n44951;
  assign n44957 = n44892 ^ n44891;
  assign n44954 = n42904 ^ n3179;
  assign n44955 = n44954 ^ n39231;
  assign n44956 = n44955 ^ n33178;
  assign n44958 = n44957 ^ n44956;
  assign n44548 = n44543 ^ n44542;
  assign n1442 = n1420 ^ n1354;
  assign n1461 = n1460 ^ n1442;
  assign n1468 = n1467 ^ n1461;
  assign n44549 = n44548 ^ n1468;
  assign n44553 = n44541 ^ n44539;
  assign n44550 = n3350 ^ n1253;
  assign n44551 = n44550 ^ n39275;
  assign n44552 = n44551 ^ n1452;
  assign n44554 = n44553 ^ n44552;
  assign n44558 = n44538 ^ n44536;
  assign n44555 = n42481 ^ n1238;
  assign n44556 = n44555 ^ n39247;
  assign n44557 = n44556 ^ n33208;
  assign n44559 = n44558 ^ n44557;
  assign n44563 = n44535 ^ n44534;
  assign n44560 = n42486 ^ n3339;
  assign n44561 = n44560 ^ n39252;
  assign n44562 = n44561 ^ n33213;
  assign n44564 = n44563 ^ n44562;
  assign n44568 = n44533 ^ n44532;
  assign n44565 = n42490 ^ n34760;
  assign n44566 = n44565 ^ n39257;
  assign n44567 = n44566 ^ n878;
  assign n44569 = n44568 ^ n44567;
  assign n44573 = n44531 ^ n44512;
  assign n44570 = n42495 ^ n34765;
  assign n44571 = n44570 ^ n788;
  assign n44572 = n44571 ^ n33220;
  assign n44574 = n44573 ^ n44572;
  assign n44578 = n44530 ^ n44529;
  assign n44575 = n42570 ^ n34769;
  assign n44576 = n44575 ^ n38755;
  assign n44577 = n44576 ^ n780;
  assign n44579 = n44578 ^ n44577;
  assign n44582 = n42560 ^ n34287;
  assign n44583 = n44582 ^ n38761;
  assign n44584 = n44583 ^ n33232;
  assign n44581 = n44526 ^ n44525;
  assign n44585 = n44584 ^ n44581;
  assign n44588 = n42550 ^ n34241;
  assign n44589 = n44588 ^ n38770;
  assign n44590 = n44589 ^ n33242;
  assign n44587 = n44523 ^ n44522;
  assign n44591 = n44590 ^ n44587;
  assign n44596 = n44520 ^ n44515;
  assign n44593 = n42518 ^ n34250;
  assign n44594 = n44593 ^ n38799;
  assign n44595 = n44594 ^ n33251;
  assign n44597 = n44596 ^ n44595;
  assign n44601 = n44519 ^ n44516;
  assign n44598 = n42523 ^ n34255;
  assign n44599 = n44598 ^ n38781;
  assign n44600 = n44599 ^ n33256;
  assign n44602 = n44601 ^ n44600;
  assign n44604 = n42533 ^ n34264;
  assign n44605 = n44604 ^ n38787;
  assign n44606 = n44605 ^ n2231;
  assign n44603 = n44518 ^ n44517;
  assign n44607 = n44606 ^ n44603;
  assign n44611 = n42849 ^ n35101;
  assign n44612 = n44611 ^ n39196;
  assign n44613 = n44612 ^ n2058;
  assign n44614 = n44446 ^ n41644;
  assign n44615 = n44613 & ~n44614;
  assign n44608 = n42529 ^ n34259;
  assign n44609 = n44608 ^ n2066;
  assign n44610 = n44609 ^ n32500;
  assign n44616 = n44615 ^ n44610;
  assign n44617 = n44615 ^ n44517;
  assign n44618 = n44616 & n44617;
  assign n44619 = n44618 ^ n44610;
  assign n44620 = n44619 ^ n44603;
  assign n44621 = ~n44607 & n44620;
  assign n44622 = n44621 ^ n44606;
  assign n44623 = n44622 ^ n44601;
  assign n44624 = n44602 & ~n44623;
  assign n44625 = n44624 ^ n44600;
  assign n44626 = n44625 ^ n44596;
  assign n44627 = n44597 & ~n44626;
  assign n44628 = n44627 ^ n44595;
  assign n44592 = n44521 ^ n44514;
  assign n44629 = n44628 ^ n44592;
  assign n44630 = n42513 ^ n34246;
  assign n44631 = n44630 ^ n38775;
  assign n44632 = n44631 ^ n33247;
  assign n44633 = n44632 ^ n44592;
  assign n44634 = n44629 & ~n44633;
  assign n44635 = n44634 ^ n44632;
  assign n44636 = n44635 ^ n44587;
  assign n44637 = ~n44591 & n44636;
  assign n44638 = n44637 ^ n44590;
  assign n44586 = n44524 ^ n44513;
  assign n44639 = n44638 ^ n44586;
  assign n44640 = n42508 ^ n34236;
  assign n44641 = n44640 ^ n38766;
  assign n44642 = n44641 ^ n33237;
  assign n44643 = n44642 ^ n44586;
  assign n44644 = n44639 & ~n44643;
  assign n44645 = n44644 ^ n44642;
  assign n44646 = n44645 ^ n44581;
  assign n44647 = n44585 & ~n44646;
  assign n44648 = n44647 ^ n44584;
  assign n44580 = n44528 ^ n44527;
  assign n44649 = n44648 ^ n44580;
  assign n44650 = n42502 ^ n732;
  assign n44651 = n44650 ^ n38818;
  assign n44652 = n44651 ^ n33227;
  assign n44653 = n44652 ^ n44580;
  assign n44654 = ~n44649 & n44653;
  assign n44655 = n44654 ^ n44652;
  assign n44656 = n44655 ^ n44578;
  assign n44657 = n44579 & ~n44656;
  assign n44658 = n44657 ^ n44577;
  assign n44659 = n44658 ^ n44573;
  assign n44660 = n44574 & ~n44659;
  assign n44661 = n44660 ^ n44572;
  assign n44662 = n44661 ^ n44568;
  assign n44663 = n44569 & ~n44662;
  assign n44664 = n44663 ^ n44567;
  assign n44665 = n44664 ^ n44563;
  assign n44666 = ~n44564 & n44665;
  assign n44667 = n44666 ^ n44562;
  assign n44668 = n44667 ^ n44558;
  assign n44669 = n44559 & ~n44668;
  assign n44670 = n44669 ^ n44557;
  assign n44671 = n44670 ^ n44553;
  assign n44672 = ~n44554 & n44671;
  assign n44673 = n44672 ^ n44552;
  assign n44674 = n44673 ^ n44548;
  assign n44675 = ~n44549 & n44674;
  assign n44676 = n44675 ^ n1468;
  assign n44547 = n44544 ^ n44511;
  assign n44677 = n44676 ^ n44547;
  assign n1478 = n1438 ^ n1372;
  assign n1479 = n1478 ^ n1475;
  assign n1486 = n1485 ^ n1479;
  assign n44678 = n44547 ^ n1486;
  assign n44679 = ~n44677 & n44678;
  assign n44680 = n44679 ^ n1486;
  assign n44546 = n44545 ^ n44510;
  assign n44681 = n44680 ^ n44546;
  assign n44115 = n42913 ^ n34746;
  assign n44116 = n44115 ^ n39238;
  assign n44117 = n44116 ^ n33190;
  assign n44960 = n44546 ^ n44117;
  assign n44961 = ~n44681 & n44960;
  assign n44962 = n44961 ^ n44117;
  assign n44959 = n44890 ^ n44889;
  assign n44963 = n44962 ^ n44959;
  assign n44964 = n42908 ^ n34741;
  assign n44965 = n44964 ^ n39291;
  assign n44966 = n44965 ^ n33183;
  assign n44967 = n44966 ^ n44959;
  assign n44968 = n44963 & ~n44967;
  assign n44969 = n44968 ^ n44966;
  assign n44970 = n44969 ^ n44957;
  assign n44971 = n44958 & ~n44970;
  assign n44972 = n44971 ^ n44956;
  assign n44973 = n44972 ^ n44952;
  assign n44974 = ~n44953 & n44973;
  assign n44975 = n44974 ^ n44951;
  assign n44948 = n44895 ^ n44888;
  assign n44976 = n44975 ^ n44948;
  assign n44977 = n42894 ^ n3093;
  assign n44978 = n44977 ^ n3203;
  assign n44979 = n44978 ^ n2722;
  assign n44980 = n44979 ^ n44948;
  assign n44981 = n44976 & ~n44980;
  assign n44982 = n44981 ^ n44979;
  assign n44983 = n44982 ^ n44946;
  assign n44984 = n44947 & ~n44983;
  assign n44985 = n44984 ^ n2738;
  assign n44945 = n44898 ^ n44897;
  assign n44986 = n44985 ^ n44945;
  assign n3114 = n3113 ^ n3107;
  assign n3118 = n3117 ^ n3114;
  assign n3119 = n3118 ^ n2826;
  assign n44987 = n44945 ^ n3119;
  assign n44988 = n44986 & ~n44987;
  assign n44989 = n44988 ^ n3119;
  assign n44990 = n44989 ^ n44940;
  assign n44991 = ~n44944 & n44990;
  assign n44992 = n44991 ^ n44943;
  assign n44993 = n44992 ^ n44935;
  assign n44994 = n44939 & ~n44993;
  assign n44995 = n44994 ^ n44938;
  assign n44870 = n44869 ^ n44830;
  assign n44871 = ~n44831 & ~n44870;
  assign n44872 = n44871 ^ n41567;
  assign n44802 = n42981 ^ n42319;
  assign n44803 = n44802 ^ n43666;
  assign n44798 = n44797 ^ n44692;
  assign n44799 = ~n44795 & n44798;
  assign n44800 = n44799 ^ n44797;
  assign n44685 = n44089 ^ n43929;
  assign n44801 = n44800 ^ n44685;
  assign n44828 = n44803 ^ n44801;
  assign n44829 = n44828 ^ n41561;
  assign n44902 = n44872 ^ n44829;
  assign n44901 = ~n44885 & ~n44900;
  assign n44934 = n44902 ^ n44901;
  assign n44996 = n44995 ^ n44934;
  assign n45024 = n44999 ^ n44996;
  assign n45022 = n43702 ^ n42629;
  assign n45023 = n45022 ^ n44138;
  assign n45160 = n45024 ^ n45023;
  assign n45161 = ~n41751 & n45160;
  assign n45162 = n45161 ^ n41749;
  assign n45000 = n44999 ^ n44934;
  assign n45001 = n44996 & ~n45000;
  assign n45002 = n45001 ^ n44999;
  assign n44903 = ~n44901 & ~n44902;
  assign n44873 = n44872 ^ n44828;
  assign n44874 = ~n44829 & n44873;
  assign n44875 = n44874 ^ n41561;
  assign n44808 = n42979 ^ n42315;
  assign n44809 = n44808 ^ n43673;
  assign n44804 = n44803 ^ n44685;
  assign n44805 = ~n44801 & n44804;
  assign n44806 = n44805 ^ n44803;
  assign n44113 = n44112 ^ n44092;
  assign n44807 = n44806 ^ n44113;
  assign n44826 = n44809 ^ n44807;
  assign n44827 = n44826 ^ n41559;
  assign n44884 = n44875 ^ n44827;
  assign n44929 = n44903 ^ n44884;
  assign n44933 = n44932 ^ n44929;
  assign n45029 = n45002 ^ n44933;
  assign n45026 = n43525 ^ n42627;
  assign n45027 = n45026 ^ n44134;
  assign n45025 = ~n45023 & ~n45024;
  assign n45028 = n45027 ^ n45025;
  assign n45163 = n45029 ^ n45028;
  assign n45164 = n45163 ^ n45161;
  assign n45165 = ~n45162 & ~n45164;
  assign n45166 = n45165 ^ n41749;
  assign n45034 = n43712 ^ n42626;
  assign n45035 = n45034 ^ n44130;
  assign n45030 = n45029 ^ n45027;
  assign n45031 = ~n45028 & ~n45030;
  assign n45032 = n45031 ^ n45025;
  assign n45003 = n45002 ^ n44929;
  assign n45004 = ~n44933 & n45003;
  assign n45005 = n45004 ^ n44932;
  assign n44925 = n42874 ^ n1794;
  assign n44926 = n44925 ^ n39207;
  assign n44927 = n44926 ^ n33139;
  assign n44904 = n44884 & ~n44903;
  assign n44876 = n44875 ^ n44826;
  assign n44877 = ~n44827 & ~n44876;
  assign n44878 = n44877 ^ n41559;
  assign n44815 = n42976 ^ n42314;
  assign n44816 = n44815 ^ n43677;
  assign n44813 = n44282 ^ n44279;
  assign n44810 = n44809 ^ n44113;
  assign n44811 = ~n44807 & ~n44810;
  assign n44812 = n44811 ^ n44809;
  assign n44814 = n44813 ^ n44812;
  assign n44824 = n44816 ^ n44814;
  assign n44825 = n44824 ^ n41549;
  assign n44883 = n44878 ^ n44825;
  assign n44924 = n44904 ^ n44883;
  assign n44928 = n44927 ^ n44924;
  assign n45021 = n45005 ^ n44928;
  assign n45033 = n45032 ^ n45021;
  assign n45159 = n45035 ^ n45033;
  assign n45167 = n45166 ^ n45159;
  assign n45260 = n45167 ^ n41745;
  assign n45259 = n45163 ^ n45162;
  assign n45389 = n45260 ^ n45259;
  assign n45376 = n43362 ^ n34883;
  assign n45377 = n45376 ^ n2203;
  assign n45378 = n45377 ^ n2344;
  assign n45542 = n45389 ^ n45378;
  assign n45379 = n43622 ^ n2023;
  assign n45380 = n45379 ^ n40102;
  assign n45381 = n45380 ^ n2182;
  assign n45382 = n45160 ^ n41751;
  assign n45383 = n45381 & ~n45382;
  assign n2161 = n2151 ^ n2100;
  assign n2186 = n2185 ^ n2161;
  assign n2193 = n2192 ^ n2186;
  assign n45384 = n45383 ^ n2193;
  assign n45385 = n45383 ^ n45259;
  assign n45386 = n45384 & ~n45385;
  assign n45387 = n45386 ^ n2193;
  assign n45543 = n45542 ^ n45387;
  assign n45054 = n44619 ^ n44607;
  assign n47105 = n45543 ^ n45054;
  assign n45998 = n44243 ^ n36403;
  assign n45999 = n45998 ^ n40828;
  assign n46000 = n45999 ^ n35101;
  assign n45694 = n44130 ^ n43702;
  assign n44741 = n44614 ^ n44613;
  assign n45695 = n45694 ^ n44741;
  assign n45663 = n43483 ^ n35472;
  assign n45664 = n45663 ^ n2938;
  assign n45665 = n45664 ^ n33951;
  assign n45110 = n44749 ^ n44172;
  assign n45111 = n45110 ^ n43538;
  assign n45108 = n44670 ^ n44554;
  assign n45101 = n44667 ^ n44559;
  assign n45094 = n44664 ^ n44564;
  assign n44698 = n44661 ^ n44569;
  assign n44695 = n44154 ^ n43271;
  assign n44697 = n44696 ^ n44695;
  assign n44699 = n44698 ^ n44697;
  assign n44703 = n44658 ^ n44574;
  assign n44700 = n44105 ^ n43261;
  assign n44702 = n44701 ^ n44700;
  assign n44704 = n44703 ^ n44702;
  assign n44708 = n44655 ^ n44579;
  assign n44705 = n43771 ^ n43205;
  assign n44707 = n44706 ^ n44705;
  assign n44709 = n44708 ^ n44707;
  assign n44713 = n44652 ^ n44649;
  assign n44710 = n43491 ^ n43094;
  assign n44712 = n44711 ^ n44710;
  assign n44714 = n44713 ^ n44712;
  assign n44717 = n44645 ^ n44585;
  assign n44715 = n43492 ^ n42605;
  assign n44716 = n44715 ^ n44503;
  assign n44718 = n44717 ^ n44716;
  assign n44721 = n44642 ^ n44639;
  assign n44719 = n44412 ^ n42606;
  assign n44720 = n44719 ^ n43495;
  assign n44722 = n44721 ^ n44720;
  assign n44725 = n44635 ^ n44591;
  assign n44723 = n43497 ^ n42607;
  assign n44724 = n44723 ^ n44405;
  assign n44726 = n44725 ^ n44724;
  assign n44729 = n43504 ^ n42609;
  assign n44730 = n44729 ^ n44392;
  assign n44728 = n44625 ^ n44597;
  assign n44731 = n44730 ^ n44728;
  assign n44734 = n44622 ^ n44602;
  assign n44732 = n43506 ^ n42610;
  assign n44733 = n44732 ^ n44385;
  assign n44735 = n44734 ^ n44733;
  assign n44738 = n44610 ^ n44517;
  assign n44739 = n44738 ^ n44615;
  assign n44736 = n43513 ^ n42616;
  assign n44737 = n44736 ^ n44371;
  assign n44740 = n44739 ^ n44737;
  assign n44742 = n43517 ^ n42624;
  assign n44743 = n44742 ^ n44123;
  assign n44744 = n44743 ^ n44741;
  assign n45010 = n42868 ^ n34709;
  assign n45011 = n45010 ^ n39202;
  assign n45012 = n45011 ^ n1924;
  assign n45006 = n45005 ^ n44924;
  assign n45007 = n44928 & ~n45006;
  assign n45008 = n45007 ^ n44927;
  assign n44905 = n44883 & n44904;
  assign n44879 = n44878 ^ n44824;
  assign n44880 = n44825 & ~n44879;
  assign n44881 = n44880 ^ n41549;
  assign n44820 = n44289 ^ n44286;
  assign n44817 = n44816 ^ n44813;
  assign n44818 = ~n44814 & ~n44817;
  assign n44819 = n44818 ^ n44816;
  assign n44821 = n44820 ^ n44819;
  assign n44745 = n42637 ^ n41764;
  assign n44746 = n44745 ^ n43665;
  assign n44822 = n44821 ^ n44746;
  assign n44823 = n44822 ^ n41124;
  assign n44882 = n44881 ^ n44823;
  assign n44923 = n44905 ^ n44882;
  assign n45009 = n45008 ^ n44923;
  assign n45019 = n45012 ^ n45009;
  assign n45017 = n43521 ^ n43032;
  assign n45018 = n45017 ^ n44128;
  assign n45020 = n45019 ^ n45018;
  assign n45036 = n45035 ^ n45021;
  assign n45037 = ~n45033 & n45036;
  assign n45038 = n45037 ^ n45035;
  assign n45039 = n45038 ^ n45019;
  assign n45040 = n45020 & n45039;
  assign n45041 = n45040 ^ n45018;
  assign n45013 = n45012 ^ n44923;
  assign n45014 = n45009 & ~n45013;
  assign n45015 = n45014 ^ n45012;
  assign n44916 = n44881 ^ n44822;
  assign n44917 = n44823 & ~n44916;
  assign n44918 = n44917 ^ n41124;
  assign n44919 = n44918 ^ n41624;
  assign n44911 = n44820 ^ n44746;
  assign n44912 = ~n44821 & n44911;
  assign n44913 = n44912 ^ n44746;
  assign n44909 = n42633 ^ n41759;
  assign n44910 = n44909 ^ n43664;
  assign n44914 = n44913 ^ n44910;
  assign n44907 = n44294 ^ n44273;
  assign n44908 = n44907 ^ n44292;
  assign n44915 = n44914 ^ n44908;
  assign n44920 = n44919 ^ n44915;
  assign n44906 = ~n44882 & ~n44905;
  assign n44921 = n44920 ^ n44906;
  assign n1905 = n1904 ^ n1868;
  assign n1933 = n1932 ^ n1905;
  assign n1940 = n1939 ^ n1933;
  assign n44922 = n44921 ^ n1940;
  assign n45016 = n45015 ^ n44922;
  assign n45042 = n45041 ^ n45016;
  assign n45043 = n43722 ^ n43039;
  assign n45044 = n45043 ^ n44125;
  assign n45045 = n45044 ^ n45016;
  assign n45046 = ~n45042 & ~n45045;
  assign n45047 = n45046 ^ n45044;
  assign n45048 = n45047 ^ n44741;
  assign n45049 = n44744 & n45048;
  assign n45050 = n45049 ^ n44743;
  assign n45051 = n45050 ^ n44739;
  assign n45052 = n44740 & ~n45051;
  assign n45053 = n45052 ^ n44737;
  assign n45055 = n45054 ^ n45053;
  assign n45056 = n43509 ^ n42614;
  assign n45057 = n45056 ^ n44378;
  assign n45058 = n45057 ^ n45054;
  assign n45059 = ~n45055 & ~n45058;
  assign n45060 = n45059 ^ n45057;
  assign n45061 = n45060 ^ n44734;
  assign n45062 = n44735 & ~n45061;
  assign n45063 = n45062 ^ n44733;
  assign n45064 = n45063 ^ n44730;
  assign n45065 = ~n44731 & n45064;
  assign n45066 = n45065 ^ n44728;
  assign n44727 = n44632 ^ n44629;
  assign n45067 = n45066 ^ n44727;
  assign n45068 = n43500 ^ n42608;
  assign n45069 = n45068 ^ n44120;
  assign n45070 = n45069 ^ n44727;
  assign n45071 = n45067 & n45070;
  assign n45072 = n45071 ^ n45069;
  assign n45073 = n45072 ^ n44725;
  assign n45074 = n44726 & ~n45073;
  assign n45075 = n45074 ^ n44724;
  assign n45076 = n45075 ^ n44721;
  assign n45077 = ~n44722 & ~n45076;
  assign n45078 = n45077 ^ n44720;
  assign n45079 = n45078 ^ n44717;
  assign n45080 = n44718 & ~n45079;
  assign n45081 = n45080 ^ n44716;
  assign n45082 = n45081 ^ n44712;
  assign n45083 = ~n44714 & n45082;
  assign n45084 = n45083 ^ n44713;
  assign n45085 = n45084 ^ n44707;
  assign n45086 = ~n44709 & n45085;
  assign n45087 = n45086 ^ n44708;
  assign n45088 = n45087 ^ n44703;
  assign n45089 = ~n44704 & ~n45088;
  assign n45090 = n45089 ^ n44702;
  assign n45091 = n45090 ^ n44698;
  assign n45092 = ~n44699 & n45091;
  assign n45093 = n45092 ^ n44697;
  assign n45095 = n45094 ^ n45093;
  assign n45096 = n44150 ^ n43469;
  assign n45097 = n45096 ^ n44782;
  assign n45098 = n45097 ^ n45094;
  assign n45099 = ~n45095 & ~n45098;
  assign n45100 = n45099 ^ n45097;
  assign n45102 = n45101 ^ n45100;
  assign n45103 = n44165 ^ n43539;
  assign n45104 = n45103 ^ n44753;
  assign n45105 = n45104 ^ n45101;
  assign n45106 = ~n45102 & n45105;
  assign n45107 = n45106 ^ n45104;
  assign n45109 = n45108 ^ n45107;
  assign n45132 = n45111 ^ n45109;
  assign n45133 = n45132 ^ n42643;
  assign n45134 = n45104 ^ n45102;
  assign n45135 = n45134 ^ n42714;
  assign n45136 = n45097 ^ n45095;
  assign n45137 = n45136 ^ n42646;
  assign n45138 = n45090 ^ n44699;
  assign n45139 = n45138 ^ n42650;
  assign n45141 = n45084 ^ n44709;
  assign n45142 = n45141 ^ n42655;
  assign n45143 = n45078 ^ n44718;
  assign n45144 = n45143 ^ n42658;
  assign n45190 = n45063 ^ n44731;
  assign n45149 = n45057 ^ n45055;
  assign n45150 = n45149 ^ n42446;
  assign n45151 = n45050 ^ n44740;
  assign n45152 = n45151 ^ n41729;
  assign n45153 = n45047 ^ n44744;
  assign n45154 = n45153 ^ n41733;
  assign n45155 = n45044 ^ n45042;
  assign n45156 = n45155 ^ n41738;
  assign n45157 = n45038 ^ n45020;
  assign n45158 = n45157 ^ n41743;
  assign n45168 = n45159 ^ n41745;
  assign n45169 = n45167 & n45168;
  assign n45170 = n45169 ^ n41745;
  assign n45171 = n45170 ^ n45157;
  assign n45172 = n45158 & ~n45171;
  assign n45173 = n45172 ^ n41743;
  assign n45174 = n45173 ^ n45155;
  assign n45175 = n45156 & ~n45174;
  assign n45176 = n45175 ^ n41738;
  assign n45177 = n45176 ^ n45153;
  assign n45178 = ~n45154 & ~n45177;
  assign n45179 = n45178 ^ n41733;
  assign n45180 = n45179 ^ n45151;
  assign n45181 = ~n45152 & ~n45180;
  assign n45182 = n45181 ^ n41729;
  assign n45183 = n45182 ^ n45149;
  assign n45184 = n45150 & ~n45183;
  assign n45185 = n45184 ^ n42446;
  assign n45148 = n45060 ^ n44735;
  assign n45186 = n45185 ^ n45148;
  assign n45187 = n45148 ^ n42595;
  assign n45188 = ~n45186 & ~n45187;
  assign n45189 = n45188 ^ n42595;
  assign n45191 = n45190 ^ n45189;
  assign n45192 = n45189 ^ n42665;
  assign n45193 = ~n45191 & ~n45192;
  assign n45194 = n45193 ^ n42665;
  assign n45147 = n45069 ^ n45067;
  assign n45195 = n45194 ^ n45147;
  assign n45196 = n45147 ^ n42622;
  assign n45197 = ~n45195 & ~n45196;
  assign n45198 = n45197 ^ n42622;
  assign n45146 = n45072 ^ n44726;
  assign n45199 = n45198 ^ n45146;
  assign n45200 = n45146 ^ n42618;
  assign n45201 = ~n45199 & n45200;
  assign n45202 = n45201 ^ n42618;
  assign n45145 = n45075 ^ n44722;
  assign n45203 = n45202 ^ n45145;
  assign n45204 = n45145 ^ n42612;
  assign n45205 = n45203 & n45204;
  assign n45206 = n45205 ^ n42612;
  assign n45207 = n45206 ^ n45143;
  assign n45208 = n45144 & ~n45207;
  assign n45209 = n45208 ^ n42658;
  assign n45210 = n45209 ^ n42657;
  assign n45211 = n45081 ^ n44714;
  assign n45212 = n45211 ^ n45209;
  assign n45213 = n45210 & n45212;
  assign n45214 = n45213 ^ n42657;
  assign n45215 = n45214 ^ n45141;
  assign n45216 = n45142 & n45215;
  assign n45217 = n45216 ^ n42655;
  assign n45140 = n45087 ^ n44704;
  assign n45218 = n45217 ^ n45140;
  assign n45219 = n45140 ^ n42652;
  assign n45220 = ~n45218 & ~n45219;
  assign n45221 = n45220 ^ n42652;
  assign n45222 = n45221 ^ n45138;
  assign n45223 = ~n45139 & ~n45222;
  assign n45224 = n45223 ^ n42650;
  assign n45225 = n45224 ^ n45136;
  assign n45226 = n45137 & n45225;
  assign n45227 = n45226 ^ n42646;
  assign n45228 = n45227 ^ n45134;
  assign n45229 = n45135 & ~n45228;
  assign n45230 = n45229 ^ n42714;
  assign n45231 = n45230 ^ n45132;
  assign n45232 = ~n45133 & n45231;
  assign n45233 = n45232 ^ n42643;
  assign n45112 = n45111 ^ n45108;
  assign n45113 = n45109 & ~n45112;
  assign n45114 = n45113 ^ n45111;
  assign n44691 = n44144 ^ n43537;
  assign n44693 = n44692 ^ n44691;
  assign n44689 = n44673 ^ n1468;
  assign n44690 = n44689 ^ n44548;
  assign n44694 = n44693 ^ n44690;
  assign n45131 = n45114 ^ n44694;
  assign n45234 = n45233 ^ n45131;
  assign n45235 = n45131 ^ n42642;
  assign n45236 = ~n45234 & ~n45235;
  assign n45237 = n45236 ^ n42642;
  assign n45115 = n45114 ^ n44690;
  assign n45116 = n44694 & n45115;
  assign n45117 = n45116 ^ n44693;
  assign n44686 = n44685 ^ n43536;
  assign n44687 = n44686 ^ n44143;
  assign n44684 = n44677 ^ n1486;
  assign n44688 = n44687 ^ n44684;
  assign n45130 = n45117 ^ n44688;
  assign n45238 = n45237 ^ n45130;
  assign n45239 = n45130 ^ n42733;
  assign n45240 = ~n45238 & ~n45239;
  assign n45241 = n45240 ^ n42733;
  assign n45118 = n45117 ^ n44684;
  assign n45119 = n44688 & n45118;
  assign n45120 = n45119 ^ n44687;
  assign n44682 = n44681 ^ n44117;
  assign n43487 = n43486 ^ n43485;
  assign n44114 = n44113 ^ n43487;
  assign n44683 = n44682 ^ n44114;
  assign n45129 = n45120 ^ n44683;
  assign n45242 = n45241 ^ n45129;
  assign n45243 = n45129 ^ n42641;
  assign n45244 = n45242 & n45243;
  assign n45245 = n45244 ^ n42641;
  assign n45125 = n44813 ^ n44246;
  assign n45126 = n45125 ^ n43612;
  assign n45124 = n44966 ^ n44963;
  assign n45127 = n45126 ^ n45124;
  assign n45121 = n45120 ^ n44682;
  assign n45122 = ~n44683 & ~n45121;
  assign n45123 = n45122 ^ n44114;
  assign n45128 = n45127 ^ n45123;
  assign n45246 = n45245 ^ n45128;
  assign n45487 = n45128 ^ n42852;
  assign n45488 = n45246 & ~n45487;
  assign n45489 = n45488 ^ n42852;
  assign n45483 = n44820 ^ n42982;
  assign n45484 = n45483 ^ n43666;
  assign n45482 = n44969 ^ n44958;
  assign n45485 = n45484 ^ n45482;
  assign n45479 = n45126 ^ n45123;
  assign n45480 = ~n45127 & n45479;
  assign n45481 = n45480 ^ n45124;
  assign n45486 = n45485 ^ n45481;
  assign n45490 = n45489 ^ n45486;
  assign n45605 = n45486 ^ n42322;
  assign n45606 = ~n45490 & n45605;
  assign n45607 = n45606 ^ n42322;
  assign n45573 = n45482 ^ n45481;
  assign n45574 = n45485 & n45573;
  assign n45575 = n45574 ^ n45484;
  assign n45570 = n43673 ^ n42989;
  assign n45571 = n45570 ^ n44908;
  assign n45569 = n44972 ^ n44953;
  assign n45572 = n45571 ^ n45569;
  assign n45603 = n45575 ^ n45572;
  assign n45604 = n45603 ^ n42327;
  assign n45629 = n45607 ^ n45604;
  assign n45491 = n45490 ^ n42322;
  assign n45247 = n45246 ^ n42852;
  assign n45248 = n45242 ^ n42641;
  assign n45249 = n45230 ^ n45133;
  assign n45250 = n45218 ^ n42652;
  assign n45251 = n45214 ^ n45142;
  assign n45252 = n45206 ^ n45144;
  assign n45253 = n45203 ^ n42612;
  assign n45254 = n45195 ^ n42622;
  assign n45255 = n45186 ^ n42595;
  assign n45256 = n45182 ^ n45150;
  assign n45257 = n45176 ^ n45154;
  assign n45258 = n45170 ^ n45158;
  assign n45261 = n45259 & n45260;
  assign n45262 = n45258 & ~n45261;
  assign n45263 = n45173 ^ n45156;
  assign n45264 = ~n45262 & ~n45263;
  assign n45265 = ~n45257 & ~n45264;
  assign n45266 = n45179 ^ n45152;
  assign n45267 = ~n45265 & ~n45266;
  assign n45268 = ~n45256 & n45267;
  assign n45269 = n45255 & n45268;
  assign n45270 = n45191 ^ n42665;
  assign n45271 = ~n45269 & n45270;
  assign n45272 = ~n45254 & n45271;
  assign n45273 = n45199 ^ n42618;
  assign n45274 = n45272 & ~n45273;
  assign n45275 = ~n45253 & n45274;
  assign n45276 = n45252 & n45275;
  assign n45277 = n45211 ^ n45210;
  assign n45278 = ~n45276 & n45277;
  assign n45279 = ~n45251 & n45278;
  assign n45280 = n45250 & ~n45279;
  assign n45281 = n45221 ^ n42650;
  assign n45282 = n45281 ^ n45138;
  assign n45283 = ~n45280 & n45282;
  assign n45284 = n45224 ^ n42646;
  assign n45285 = n45284 ^ n45136;
  assign n45286 = ~n45283 & ~n45285;
  assign n45287 = n45227 ^ n45135;
  assign n45288 = n45286 & n45287;
  assign n45289 = ~n45249 & n45288;
  assign n45290 = n45234 ^ n42642;
  assign n45291 = ~n45289 & n45290;
  assign n45292 = n45238 ^ n42733;
  assign n45293 = n45291 & ~n45292;
  assign n45294 = n45248 & ~n45293;
  assign n45492 = n45247 & n45294;
  assign n45628 = n45491 & ~n45492;
  assign n45662 = n45629 ^ n45628;
  assign n45666 = n45665 ^ n45662;
  assign n45493 = n45492 ^ n45491;
  assign n2923 = n2922 ^ n2892;
  assign n2924 = n2923 ^ n2862;
  assign n2931 = n2930 ^ n2924;
  assign n45494 = n45493 ^ n2931;
  assign n45295 = n45294 ^ n45247;
  assign n3228 = n3227 ^ n2803;
  assign n3238 = n3237 ^ n3228;
  assign n3239 = n3238 ^ n2914;
  assign n45296 = n45295 ^ n3239;
  assign n45298 = n43456 ^ n2788;
  assign n45299 = n45298 ^ n39940;
  assign n45300 = n45299 ^ n3235;
  assign n45297 = n45293 ^ n45248;
  assign n45301 = n45300 ^ n45297;
  assign n45306 = n45290 ^ n45289;
  assign n45303 = n43297 ^ n35485;
  assign n45304 = n45303 ^ n40060;
  assign n45305 = n45304 ^ n34007;
  assign n45307 = n45306 ^ n45305;
  assign n45312 = n45287 ^ n45286;
  assign n45309 = n43307 ^ n35494;
  assign n45310 = n45309 ^ n40050;
  assign n45311 = n45310 ^ n2492;
  assign n45313 = n45312 ^ n45311;
  assign n45317 = n45285 ^ n45283;
  assign n45314 = n43437 ^ n35499;
  assign n45315 = n45314 ^ n39956;
  assign n45316 = n45315 ^ n34018;
  assign n45318 = n45317 ^ n45316;
  assign n45320 = n43430 ^ n35504;
  assign n45321 = n45320 ^ n39962;
  assign n45322 = n45321 ^ n34023;
  assign n45319 = n45282 ^ n45280;
  assign n45323 = n45322 ^ n45319;
  assign n45327 = n45279 ^ n45250;
  assign n45324 = n43314 ^ n35509;
  assign n45325 = n45324 ^ n39967;
  assign n45326 = n45325 ^ n1301;
  assign n45328 = n45327 ^ n45326;
  assign n45335 = n45277 ^ n45276;
  assign n45332 = n43324 ^ n35520;
  assign n45333 = n45332 ^ n39973;
  assign n45334 = n45333 ^ n1116;
  assign n45336 = n45335 ^ n45334;
  assign n45340 = n45274 ^ n45253;
  assign n45337 = n43332 ^ n35527;
  assign n45338 = n45337 ^ n39980;
  assign n45339 = n45338 ^ n976;
  assign n45341 = n45340 ^ n45339;
  assign n45343 = n43408 ^ n840;
  assign n45344 = n45343 ^ n39985;
  assign n45345 = n45344 ^ n3314;
  assign n45342 = n45273 ^ n45272;
  assign n45346 = n45345 ^ n45342;
  assign n45349 = n43339 ^ n35539;
  assign n45350 = n45349 ^ n39995;
  assign n45351 = n45350 ^ n33464;
  assign n45348 = n45270 ^ n45269;
  assign n45352 = n45351 ^ n45348;
  assign n45356 = n45268 ^ n45255;
  assign n45353 = n43391 ^ n35544;
  assign n45354 = n45353 ^ n39999;
  assign n45355 = n45354 ^ n33469;
  assign n45357 = n45356 ^ n45355;
  assign n45361 = n45267 ^ n45256;
  assign n45358 = n43344 ^ n35549;
  assign n45359 = n45358 ^ n40004;
  assign n45360 = n45359 ^ n33473;
  assign n45362 = n45361 ^ n45360;
  assign n45366 = n45266 ^ n45265;
  assign n45363 = n43381 ^ n35553;
  assign n45364 = n45363 ^ n39432;
  assign n45365 = n45364 ^ n33478;
  assign n45367 = n45366 ^ n45365;
  assign n45370 = n43356 ^ n35564;
  assign n45371 = n45370 ^ n39423;
  assign n45372 = n45371 ^ n33489;
  assign n45369 = n45263 ^ n45262;
  assign n45373 = n45372 ^ n45369;
  assign n45374 = n45261 ^ n45258;
  assign n2334 = n2333 ^ n2255;
  assign n2353 = n2352 ^ n2334;
  assign n2363 = n2362 ^ n2353;
  assign n45375 = n45374 ^ n2363;
  assign n45388 = n45387 ^ n45378;
  assign n45390 = n45389 ^ n45387;
  assign n45391 = n45388 & n45390;
  assign n45392 = n45391 ^ n45378;
  assign n45393 = n45392 ^ n45374;
  assign n45394 = ~n45375 & n45393;
  assign n45395 = n45394 ^ n2363;
  assign n45396 = n45395 ^ n45369;
  assign n45397 = ~n45373 & n45396;
  assign n45398 = n45397 ^ n45372;
  assign n45368 = n45264 ^ n45257;
  assign n45399 = n45398 ^ n45368;
  assign n45400 = n43351 ^ n35558;
  assign n45401 = n45400 ^ n39406;
  assign n45402 = n45401 ^ n33483;
  assign n45403 = n45402 ^ n45368;
  assign n45404 = ~n45399 & n45403;
  assign n45405 = n45404 ^ n45402;
  assign n45406 = n45405 ^ n45365;
  assign n45407 = ~n45367 & ~n45406;
  assign n45408 = n45407 ^ n45366;
  assign n45409 = n45408 ^ n45360;
  assign n45410 = n45362 & n45409;
  assign n45411 = n45410 ^ n45361;
  assign n45412 = n45411 ^ n45356;
  assign n45413 = ~n45357 & n45412;
  assign n45414 = n45413 ^ n45355;
  assign n45415 = n45414 ^ n45348;
  assign n45416 = ~n45352 & n45415;
  assign n45417 = n45416 ^ n45351;
  assign n45347 = n45271 ^ n45254;
  assign n45418 = n45417 ^ n45347;
  assign n45422 = n45421 ^ n45417;
  assign n45423 = n45418 & n45422;
  assign n45424 = n45423 ^ n45421;
  assign n45425 = n45424 ^ n45345;
  assign n45426 = ~n45346 & ~n45425;
  assign n45427 = n45426 ^ n45342;
  assign n45428 = n45427 ^ n45339;
  assign n45429 = ~n45341 & n45428;
  assign n45430 = n45429 ^ n45340;
  assign n951 = n950 ^ n914;
  assign n985 = n984 ^ n951;
  assign n995 = n994 ^ n985;
  assign n45431 = n45430 ^ n995;
  assign n45432 = n45275 ^ n45252;
  assign n45433 = n45432 ^ n45430;
  assign n45434 = ~n45431 & n45433;
  assign n45435 = n45434 ^ n995;
  assign n45436 = n45435 ^ n45335;
  assign n45437 = n45336 & ~n45436;
  assign n45438 = n45437 ^ n45334;
  assign n45329 = n43319 ^ n35515;
  assign n45330 = n45329 ^ n1124;
  assign n45331 = n45330 ^ n33961;
  assign n45439 = n45438 ^ n45331;
  assign n45440 = n45278 ^ n45251;
  assign n45441 = n45440 ^ n45438;
  assign n45442 = n45439 & ~n45441;
  assign n45443 = n45442 ^ n45331;
  assign n45444 = n45443 ^ n45327;
  assign n45445 = ~n45328 & n45444;
  assign n45446 = n45445 ^ n45326;
  assign n45447 = n45446 ^ n45322;
  assign n45448 = n45323 & ~n45447;
  assign n45449 = n45448 ^ n45319;
  assign n45450 = n45449 ^ n45317;
  assign n45451 = n45318 & ~n45450;
  assign n45452 = n45451 ^ n45316;
  assign n45453 = n45452 ^ n45312;
  assign n45454 = n45313 & ~n45453;
  assign n45455 = n45454 ^ n45311;
  assign n45308 = n45288 ^ n45249;
  assign n45456 = n45455 ^ n45308;
  assign n45457 = n43303 ^ n35489;
  assign n45458 = n45457 ^ n39950;
  assign n45459 = n45458 ^ n3059;
  assign n45460 = n45459 ^ n45308;
  assign n45461 = n45456 & ~n45460;
  assign n45462 = n45461 ^ n45459;
  assign n45463 = n45462 ^ n45306;
  assign n45464 = n45307 & ~n45463;
  assign n45465 = n45464 ^ n45305;
  assign n45302 = n45292 ^ n45291;
  assign n45466 = n45465 ^ n45302;
  assign n45467 = n43292 ^ n3213;
  assign n45468 = n45467 ^ n39944;
  assign n45469 = n45468 ^ n34002;
  assign n45470 = n45469 ^ n45302;
  assign n45471 = ~n45466 & n45470;
  assign n45472 = n45471 ^ n45469;
  assign n45473 = n45472 ^ n45297;
  assign n45474 = ~n45301 & n45473;
  assign n45475 = n45474 ^ n45300;
  assign n45476 = n45475 ^ n45295;
  assign n45477 = n45296 & ~n45476;
  assign n45478 = n45477 ^ n3239;
  assign n45667 = n45493 ^ n45478;
  assign n45668 = n45494 & ~n45667;
  assign n45669 = n45668 ^ n2931;
  assign n45670 = n45669 ^ n45662;
  assign n45671 = ~n45666 & n45670;
  assign n45672 = n45671 ^ n45665;
  assign n45658 = n35467 ^ n2966;
  assign n45659 = n45658 ^ n39930;
  assign n45660 = n45659 ^ n1655;
  assign n45630 = ~n45628 & n45629;
  assign n45608 = n45607 ^ n45603;
  assign n45609 = ~n45604 & n45608;
  assign n45610 = n45609 ^ n42327;
  assign n45576 = n45575 ^ n45569;
  assign n45577 = n45572 & n45576;
  assign n45578 = n45577 ^ n45571;
  assign n45566 = n43677 ^ n42981;
  assign n45567 = n45566 ^ n44324;
  assign n45565 = n44979 ^ n44976;
  assign n45568 = n45567 ^ n45565;
  assign n45601 = n45578 ^ n45568;
  assign n45602 = n45601 ^ n42319;
  assign n45627 = n45610 ^ n45602;
  assign n45657 = n45630 ^ n45627;
  assign n45661 = n45660 ^ n45657;
  assign n45693 = n45672 ^ n45661;
  assign n45792 = n45695 ^ n45693;
  assign n45997 = n45792 ^ n42629;
  assign n46158 = n46000 ^ n45997;
  assign n47106 = n47105 ^ n46158;
  assign n46067 = n43949 ^ n36331;
  assign n46068 = n46067 ^ n40762;
  assign n46069 = n46068 ^ n34746;
  assign n45523 = n44711 ^ n43495;
  assign n45524 = n45523 ^ n44698;
  assign n45522 = n45408 ^ n45362;
  assign n45525 = n45524 ^ n45522;
  assign n45528 = n45405 ^ n45367;
  assign n45526 = n44503 ^ n43497;
  assign n45527 = n45526 ^ n44703;
  assign n45529 = n45528 ^ n45527;
  assign n45532 = n45402 ^ n45399;
  assign n45530 = n44412 ^ n43500;
  assign n45531 = n45530 ^ n44708;
  assign n45533 = n45532 ^ n45531;
  assign n45536 = n45395 ^ n45373;
  assign n45534 = n44405 ^ n43504;
  assign n45535 = n45534 ^ n44713;
  assign n45537 = n45536 ^ n45535;
  assign n45540 = n45392 ^ n45375;
  assign n45538 = n44120 ^ n43506;
  assign n45539 = n45538 ^ n44717;
  assign n45541 = n45540 ^ n45539;
  assign n45544 = n44392 ^ n43509;
  assign n45545 = n45544 ^ n44721;
  assign n45546 = n45545 ^ n45543;
  assign n45549 = n44385 ^ n43513;
  assign n45550 = n45549 ^ n44725;
  assign n45547 = n45259 ^ n2193;
  assign n45548 = n45547 ^ n45383;
  assign n45551 = n45550 ^ n45548;
  assign n45686 = n44371 ^ n43722;
  assign n45687 = n45686 ^ n44728;
  assign n45643 = n43632 ^ n35452;
  assign n45644 = n45643 ^ n39920;
  assign n45645 = n45644 ^ n33935;
  assign n45631 = n45627 & ~n45630;
  assign n45611 = n45610 ^ n45601;
  assign n45612 = n45602 & n45611;
  assign n45613 = n45612 ^ n42319;
  assign n45579 = n45578 ^ n45565;
  assign n45580 = ~n45568 & ~n45579;
  assign n45581 = n45580 ^ n45567;
  assign n45562 = n43665 ^ n42979;
  assign n45563 = n45562 ^ n44331;
  assign n45561 = n44982 ^ n44947;
  assign n45564 = n45563 ^ n45561;
  assign n45599 = n45581 ^ n45564;
  assign n45600 = n45599 ^ n42315;
  assign n45632 = n45613 ^ n45600;
  assign n45633 = ~n45631 & ~n45632;
  assign n45614 = n45613 ^ n45599;
  assign n45615 = ~n45600 & ~n45614;
  assign n45616 = n45615 ^ n42315;
  assign n45582 = n45581 ^ n45561;
  assign n45583 = n45564 & ~n45582;
  assign n45584 = n45583 ^ n45563;
  assign n45558 = n43664 ^ n42976;
  assign n45559 = n45558 ^ n44322;
  assign n45596 = n45584 ^ n45559;
  assign n45557 = n44986 ^ n3119;
  assign n45597 = n45596 ^ n45557;
  assign n45598 = n45597 ^ n42314;
  assign n45634 = n45616 ^ n45598;
  assign n45635 = n45633 & ~n45634;
  assign n45617 = n45616 ^ n45597;
  assign n45618 = n45598 & ~n45617;
  assign n45619 = n45618 ^ n42314;
  assign n45560 = n45559 ^ n45557;
  assign n45585 = n45584 ^ n45557;
  assign n45586 = ~n45560 & n45585;
  assign n45587 = n45586 ^ n45559;
  assign n45554 = n43532 ^ n42637;
  assign n45555 = n45554 ^ n44317;
  assign n45553 = n44989 ^ n44944;
  assign n45556 = n45555 ^ n45553;
  assign n45594 = n45587 ^ n45556;
  assign n45595 = n45594 ^ n41764;
  assign n45626 = n45619 ^ n45595;
  assign n45642 = n45635 ^ n45626;
  assign n45646 = n45645 ^ n45642;
  assign n45648 = n43637 ^ n35457;
  assign n45649 = n45648 ^ n39925;
  assign n45650 = n45649 ^ n33940;
  assign n45647 = n45634 ^ n45633;
  assign n45651 = n45650 ^ n45647;
  assign n45653 = n43651 ^ n35462;
  assign n45654 = n45653 ^ n40087;
  assign n45655 = n45654 ^ n33944;
  assign n45652 = n45632 ^ n45631;
  assign n45656 = n45655 ^ n45652;
  assign n45673 = n45672 ^ n45660;
  assign n45674 = n45661 & ~n45673;
  assign n45675 = n45674 ^ n45657;
  assign n45676 = n45675 ^ n45655;
  assign n45677 = n45656 & ~n45676;
  assign n45678 = n45677 ^ n45652;
  assign n45679 = n45678 ^ n45647;
  assign n45680 = ~n45651 & n45679;
  assign n45681 = n45680 ^ n45650;
  assign n45682 = n45681 ^ n45642;
  assign n45683 = ~n45646 & n45682;
  assign n45684 = n45683 ^ n45645;
  assign n45637 = n43627 ^ n2005;
  assign n45638 = n45637 ^ n39915;
  assign n45639 = n45638 ^ n34106;
  assign n45636 = ~n45626 & ~n45635;
  assign n45640 = n45639 ^ n45636;
  assign n45620 = n45619 ^ n45594;
  assign n45621 = ~n45595 & ~n45620;
  assign n45622 = n45621 ^ n41764;
  assign n45623 = n45622 ^ n44314;
  assign n45592 = n44992 ^ n44939;
  assign n45593 = n45592 ^ n44909;
  assign n45624 = n45623 ^ n45593;
  assign n45588 = n45587 ^ n45553;
  assign n45589 = ~n45556 & n45588;
  assign n45590 = n45589 ^ n45555;
  assign n45591 = n45590 ^ n43530;
  assign n45625 = n45624 ^ n45591;
  assign n45641 = n45640 ^ n45625;
  assign n45685 = n45684 ^ n45641;
  assign n45688 = n45687 ^ n45685;
  assign n45707 = n45681 ^ n45646;
  assign n45691 = n45678 ^ n45651;
  assign n45689 = n44125 ^ n43712;
  assign n45690 = n45689 ^ n45054;
  assign n45692 = n45691 ^ n45690;
  assign n45697 = n44128 ^ n43525;
  assign n45698 = n45697 ^ n44739;
  assign n45696 = n45693 & n45695;
  assign n45699 = n45698 ^ n45696;
  assign n45700 = n45675 ^ n45656;
  assign n45701 = n45700 ^ n45698;
  assign n45702 = n45699 & ~n45701;
  assign n45703 = n45702 ^ n45696;
  assign n45704 = n45703 ^ n45691;
  assign n45705 = ~n45692 & n45704;
  assign n45706 = n45705 ^ n45690;
  assign n45708 = n45707 ^ n45706;
  assign n45709 = n44123 ^ n43521;
  assign n45710 = n45709 ^ n44734;
  assign n45711 = n45710 ^ n45707;
  assign n45712 = n45708 & n45711;
  assign n45713 = n45712 ^ n45710;
  assign n45714 = n45713 ^ n45687;
  assign n45715 = n45688 & n45714;
  assign n45716 = n45715 ^ n45685;
  assign n45552 = n45382 ^ n45381;
  assign n45717 = n45716 ^ n45552;
  assign n45718 = n44378 ^ n43517;
  assign n45719 = n45718 ^ n44727;
  assign n45720 = n45719 ^ n45552;
  assign n45721 = n45717 & ~n45720;
  assign n45722 = n45721 ^ n45719;
  assign n45723 = n45722 ^ n45550;
  assign n45724 = ~n45551 & n45723;
  assign n45725 = n45724 ^ n45548;
  assign n45726 = n45725 ^ n45543;
  assign n45727 = n45546 & n45726;
  assign n45728 = n45727 ^ n45545;
  assign n45729 = n45728 ^ n45540;
  assign n45730 = n45541 & ~n45729;
  assign n45731 = n45730 ^ n45539;
  assign n45732 = n45731 ^ n45535;
  assign n45733 = n45537 & ~n45732;
  assign n45734 = n45733 ^ n45536;
  assign n45735 = n45734 ^ n45532;
  assign n45736 = n45533 & n45735;
  assign n45737 = n45736 ^ n45531;
  assign n45738 = n45737 ^ n45528;
  assign n45739 = ~n45529 & n45738;
  assign n45740 = n45739 ^ n45527;
  assign n45741 = n45740 ^ n45522;
  assign n45742 = ~n45525 & n45741;
  assign n45743 = n45742 ^ n45524;
  assign n45519 = n44706 ^ n43492;
  assign n45520 = n45519 ^ n45094;
  assign n45518 = n45411 ^ n45357;
  assign n45521 = n45520 ^ n45518;
  assign n45774 = n45743 ^ n45521;
  assign n45775 = n45774 ^ n42605;
  assign n45776 = n45737 ^ n45527;
  assign n45777 = n45776 ^ n45528;
  assign n45778 = n45777 ^ n42607;
  assign n45779 = n45734 ^ n45531;
  assign n45780 = n45779 ^ n45532;
  assign n45781 = n45780 ^ n42608;
  assign n45783 = n45728 ^ n45541;
  assign n45784 = n45783 ^ n42610;
  assign n45785 = n45725 ^ n45546;
  assign n45786 = n45785 ^ n42614;
  assign n45787 = n45719 ^ n45717;
  assign n45788 = n45787 ^ n42624;
  assign n45806 = n45713 ^ n45688;
  assign n45790 = n45703 ^ n45692;
  assign n45791 = n45790 ^ n42626;
  assign n45793 = n42629 & n45792;
  assign n45794 = n45793 ^ n42627;
  assign n45795 = n45700 ^ n45699;
  assign n45796 = n45795 ^ n45793;
  assign n45797 = n45794 & ~n45796;
  assign n45798 = n45797 ^ n42627;
  assign n45799 = n45798 ^ n45790;
  assign n45800 = n45791 & n45799;
  assign n45801 = n45800 ^ n42626;
  assign n45789 = n45710 ^ n45708;
  assign n45802 = n45801 ^ n45789;
  assign n45803 = n45789 ^ n43032;
  assign n45804 = n45802 & ~n45803;
  assign n45805 = n45804 ^ n43032;
  assign n45807 = n45806 ^ n45805;
  assign n45808 = n45805 ^ n43039;
  assign n45809 = ~n45807 & n45808;
  assign n45810 = n45809 ^ n43039;
  assign n45811 = n45810 ^ n45787;
  assign n45812 = n45788 & ~n45811;
  assign n45813 = n45812 ^ n42624;
  assign n45814 = n45813 ^ n42616;
  assign n45815 = n45722 ^ n45551;
  assign n45816 = n45815 ^ n45813;
  assign n45817 = n45814 & ~n45816;
  assign n45818 = n45817 ^ n42616;
  assign n45819 = n45818 ^ n45785;
  assign n45820 = n45786 & n45819;
  assign n45821 = n45820 ^ n42614;
  assign n45822 = n45821 ^ n45783;
  assign n45823 = ~n45784 & n45822;
  assign n45824 = n45823 ^ n42610;
  assign n45782 = n45731 ^ n45537;
  assign n45825 = n45824 ^ n45782;
  assign n45826 = n45782 ^ n42609;
  assign n45827 = n45825 & n45826;
  assign n45828 = n45827 ^ n42609;
  assign n45829 = n45828 ^ n45780;
  assign n45830 = ~n45781 & ~n45829;
  assign n45831 = n45830 ^ n42608;
  assign n45832 = n45831 ^ n45777;
  assign n45833 = n45778 & n45832;
  assign n45834 = n45833 ^ n42607;
  assign n45835 = n45834 ^ n42606;
  assign n45836 = n45740 ^ n45525;
  assign n45837 = n45836 ^ n45834;
  assign n45838 = n45835 & ~n45837;
  assign n45839 = n45838 ^ n42606;
  assign n45840 = n45839 ^ n45774;
  assign n45841 = n45775 & ~n45840;
  assign n45842 = n45841 ^ n42605;
  assign n45744 = n45743 ^ n45520;
  assign n45745 = ~n45521 & ~n45744;
  assign n45746 = n45745 ^ n45518;
  assign n45515 = n44701 ^ n43491;
  assign n45516 = n45515 ^ n45101;
  assign n45513 = n45414 ^ n45351;
  assign n45514 = n45513 ^ n45348;
  assign n45517 = n45516 ^ n45514;
  assign n45773 = n45746 ^ n45517;
  assign n45843 = n45842 ^ n45773;
  assign n45844 = n45773 ^ n43094;
  assign n45845 = ~n45843 & ~n45844;
  assign n45846 = n45845 ^ n43094;
  assign n45747 = n45746 ^ n45516;
  assign n45748 = n45517 & ~n45747;
  assign n45749 = n45748 ^ n45514;
  assign n45509 = n44696 ^ n43771;
  assign n45510 = n45509 ^ n45108;
  assign n45770 = n45749 ^ n45510;
  assign n45511 = n45421 ^ n45418;
  assign n45771 = n45770 ^ n45511;
  assign n45772 = n45771 ^ n43205;
  assign n45859 = n45846 ^ n45772;
  assign n45860 = n45839 ^ n42605;
  assign n45861 = n45860 ^ n45774;
  assign n45862 = n45836 ^ n42606;
  assign n45863 = n45862 ^ n45834;
  assign n45864 = n45828 ^ n45781;
  assign n45865 = n45821 ^ n45784;
  assign n45866 = n45818 ^ n42614;
  assign n45867 = n45866 ^ n45785;
  assign n45868 = n45815 ^ n42616;
  assign n45869 = n45868 ^ n45813;
  assign n45870 = n45807 ^ n43039;
  assign n45871 = n45802 ^ n43032;
  assign n45872 = n45798 ^ n45791;
  assign n45873 = n45795 ^ n45794;
  assign n45874 = ~n45872 & ~n45873;
  assign n45875 = n45871 & ~n45874;
  assign n45876 = n45870 & ~n45875;
  assign n45877 = n45810 ^ n45788;
  assign n45878 = ~n45876 & ~n45877;
  assign n45879 = n45869 & ~n45878;
  assign n45880 = n45867 & n45879;
  assign n45881 = n45865 & n45880;
  assign n45882 = n45825 ^ n42609;
  assign n45883 = ~n45881 & n45882;
  assign n45884 = n45864 & n45883;
  assign n45885 = n45831 ^ n45778;
  assign n45886 = n45884 & n45885;
  assign n45887 = ~n45863 & n45886;
  assign n45888 = ~n45861 & n45887;
  assign n45889 = n45843 ^ n43094;
  assign n45890 = ~n45888 & ~n45889;
  assign n45891 = n45859 & n45890;
  assign n45847 = n45846 ^ n45771;
  assign n45848 = ~n45772 & ~n45847;
  assign n45849 = n45848 ^ n43205;
  assign n45892 = n45849 ^ n43261;
  assign n45512 = n45511 ^ n45510;
  assign n45750 = n45749 ^ n45511;
  assign n45751 = ~n45512 & ~n45750;
  assign n45752 = n45751 ^ n45510;
  assign n45507 = n45424 ^ n45346;
  assign n45505 = n44782 ^ n44105;
  assign n45506 = n45505 ^ n44690;
  assign n45508 = n45507 ^ n45506;
  assign n45768 = n45752 ^ n45508;
  assign n45893 = n45892 ^ n45768;
  assign n45894 = ~n45891 & n45893;
  assign n45769 = n45768 ^ n43261;
  assign n45850 = n45849 ^ n45768;
  assign n45851 = ~n45769 & n45850;
  assign n45852 = n45851 ^ n43261;
  assign n45753 = n45752 ^ n45507;
  assign n45754 = n45508 & n45753;
  assign n45755 = n45754 ^ n45506;
  assign n45502 = n44753 ^ n44154;
  assign n45503 = n45502 ^ n44684;
  assign n45766 = n45755 ^ n45503;
  assign n45501 = n45427 ^ n45341;
  assign n45767 = n45766 ^ n45501;
  assign n45853 = n45852 ^ n45767;
  assign n45858 = n45853 ^ n43271;
  assign n45932 = n45894 ^ n45858;
  assign n1410 = n1409 ^ n1325;
  assign n1429 = n1428 ^ n1410;
  assign n1439 = n1438 ^ n1429;
  assign n45933 = n45932 ^ n1439;
  assign n45935 = n45890 ^ n45859;
  assign n1219 = n1209 ^ n1158;
  assign n1247 = n1246 ^ n1219;
  assign n1254 = n1253 ^ n1247;
  assign n45936 = n45935 ^ n1254;
  assign n45938 = n43963 ^ n1078;
  assign n45939 = n45938 ^ n3341;
  assign n45940 = n45939 ^ n1238;
  assign n45937 = n45889 ^ n45888;
  assign n45941 = n45940 ^ n45937;
  assign n45945 = n45887 ^ n45861;
  assign n45942 = n43967 ^ n1060;
  assign n45943 = n45942 ^ n40394;
  assign n45944 = n45943 ^ n3339;
  assign n45946 = n45945 ^ n45944;
  assign n45947 = n45886 ^ n45863;
  assign n45951 = n45950 ^ n45947;
  assign n45955 = n45885 ^ n45884;
  assign n45952 = n43977 ^ n35830;
  assign n45953 = n45952 ^ n40306;
  assign n45954 = n45953 ^ n34765;
  assign n45956 = n45955 ^ n45954;
  assign n45960 = n45883 ^ n45864;
  assign n45957 = n44046 ^ n35835;
  assign n45958 = n45957 ^ n40311;
  assign n45959 = n45958 ^ n34769;
  assign n45961 = n45960 ^ n45959;
  assign n45963 = n44039 ^ n35839;
  assign n45964 = n45963 ^ n40378;
  assign n45965 = n45964 ^ n732;
  assign n45962 = n45882 ^ n45881;
  assign n45966 = n45965 ^ n45962;
  assign n45968 = n44032 ^ n35844;
  assign n45969 = n45968 ^ n40318;
  assign n45970 = n45969 ^ n34287;
  assign n45967 = n45880 ^ n45865;
  assign n45971 = n45970 ^ n45967;
  assign n45973 = n43986 ^ n35849;
  assign n45974 = n45973 ^ n40323;
  assign n45975 = n45974 ^ n34236;
  assign n45972 = n45879 ^ n45867;
  assign n45976 = n45975 ^ n45972;
  assign n45980 = n45878 ^ n45869;
  assign n45977 = n44022 ^ n35854;
  assign n45978 = n45977 ^ n40328;
  assign n45979 = n45978 ^ n34241;
  assign n45981 = n45980 ^ n45979;
  assign n45983 = n43991 ^ n35860;
  assign n45984 = n45983 ^ n40333;
  assign n45985 = n45984 ^ n34246;
  assign n45982 = n45877 ^ n45876;
  assign n45986 = n45985 ^ n45982;
  assign n45992 = n45873 ^ n45872;
  assign n45989 = n44000 ^ n2288;
  assign n45990 = n45989 ^ n40342;
  assign n45991 = n45990 ^ n34264;
  assign n45993 = n45992 ^ n45991;
  assign n46001 = n45997 & n46000;
  assign n45994 = n40345 ^ n2273;
  assign n45995 = n45994 ^ n44003;
  assign n45996 = n45995 ^ n34259;
  assign n46002 = n46001 ^ n45996;
  assign n46003 = n46001 ^ n45873;
  assign n46004 = n46002 & n46003;
  assign n46005 = n46004 ^ n45996;
  assign n46006 = n46005 ^ n45992;
  assign n46007 = ~n45993 & n46006;
  assign n46008 = n46007 ^ n45991;
  assign n45988 = n45874 ^ n45871;
  assign n46009 = n46008 ^ n45988;
  assign n46010 = n35869 ^ n2389;
  assign n46011 = n46010 ^ n40338;
  assign n46012 = n46011 ^ n34255;
  assign n46013 = n46012 ^ n45988;
  assign n46014 = n46009 & ~n46013;
  assign n46015 = n46014 ^ n46012;
  assign n45987 = n45875 ^ n45870;
  assign n46016 = n46015 ^ n45987;
  assign n46017 = n35865 ^ n2407;
  assign n46018 = n46017 ^ n40359;
  assign n46019 = n46018 ^ n34250;
  assign n46020 = n46019 ^ n45987;
  assign n46021 = ~n46016 & n46020;
  assign n46022 = n46021 ^ n46019;
  assign n46023 = n46022 ^ n45982;
  assign n46024 = n45986 & ~n46023;
  assign n46025 = n46024 ^ n45985;
  assign n46026 = n46025 ^ n45980;
  assign n46027 = n45981 & ~n46026;
  assign n46028 = n46027 ^ n45979;
  assign n46029 = n46028 ^ n45975;
  assign n46030 = ~n45976 & ~n46029;
  assign n46031 = n46030 ^ n45972;
  assign n46032 = n46031 ^ n45970;
  assign n46033 = ~n45971 & n46032;
  assign n46034 = n46033 ^ n45967;
  assign n46035 = n46034 ^ n45965;
  assign n46036 = ~n45966 & n46035;
  assign n46037 = n46036 ^ n45962;
  assign n46038 = n46037 ^ n45960;
  assign n46039 = n45961 & n46038;
  assign n46040 = n46039 ^ n45959;
  assign n46041 = n46040 ^ n45955;
  assign n46042 = n45956 & ~n46041;
  assign n46043 = n46042 ^ n45954;
  assign n46044 = n46043 ^ n45950;
  assign n46045 = ~n45951 & ~n46044;
  assign n46046 = n46045 ^ n45947;
  assign n46047 = n46046 ^ n45945;
  assign n46048 = ~n45946 & ~n46047;
  assign n46049 = n46048 ^ n45944;
  assign n46050 = n46049 ^ n45940;
  assign n46051 = ~n45941 & ~n46050;
  assign n46052 = n46051 ^ n45937;
  assign n46053 = n46052 ^ n45935;
  assign n46054 = ~n45936 & ~n46053;
  assign n46055 = n46054 ^ n1254;
  assign n45934 = n45893 ^ n45891;
  assign n46056 = n46055 ^ n45934;
  assign n46057 = n43955 ^ n36337;
  assign n46058 = n46057 ^ n1264;
  assign n46059 = n46058 ^ n1420;
  assign n46060 = n46059 ^ n45934;
  assign n46061 = n46056 & ~n46060;
  assign n46062 = n46061 ^ n46059;
  assign n46063 = n46062 ^ n45932;
  assign n46064 = ~n45933 & n46063;
  assign n46065 = n46064 ^ n1439;
  assign n45895 = ~n45858 & ~n45894;
  assign n45854 = n45767 ^ n43271;
  assign n45855 = ~n45853 & ~n45854;
  assign n45856 = n45855 ^ n43271;
  assign n45762 = n44749 ^ n44150;
  assign n45763 = n45762 ^ n44682;
  assign n45759 = n45432 ^ n995;
  assign n45760 = n45759 ^ n45430;
  assign n45504 = n45503 ^ n45501;
  assign n45756 = n45755 ^ n45501;
  assign n45757 = n45504 & n45756;
  assign n45758 = n45757 ^ n45503;
  assign n45761 = n45760 ^ n45758;
  assign n45764 = n45763 ^ n45761;
  assign n45765 = n45764 ^ n43469;
  assign n45857 = n45856 ^ n45765;
  assign n45931 = n45895 ^ n45857;
  assign n46066 = n46065 ^ n45931;
  assign n46088 = n46069 ^ n46066;
  assign n46084 = n45472 ^ n45300;
  assign n46085 = n46084 ^ n45297;
  assign n46086 = n46085 ^ n45553;
  assign n46087 = n46086 ^ n44820;
  assign n46089 = n46088 ^ n46087;
  assign n46093 = n46062 ^ n45933;
  assign n46091 = n45557 ^ n44813;
  assign n46090 = n45469 ^ n45466;
  assign n46092 = n46091 ^ n46090;
  assign n46094 = n46093 ^ n46092;
  assign n46099 = n46059 ^ n46056;
  assign n46095 = n45462 ^ n45305;
  assign n46096 = n46095 ^ n45306;
  assign n46097 = n46096 ^ n45561;
  assign n46098 = n46097 ^ n44113;
  assign n46100 = n46099 ^ n46098;
  assign n46102 = n45459 ^ n45456;
  assign n46103 = n46102 ^ n45565;
  assign n46104 = n46103 ^ n44685;
  assign n46101 = n46052 ^ n45936;
  assign n46105 = n46104 ^ n46101;
  assign n46109 = n46049 ^ n45941;
  assign n46107 = n45569 ^ n44692;
  assign n46106 = n45452 ^ n45313;
  assign n46108 = n46107 ^ n46106;
  assign n46110 = n46109 ^ n46108;
  assign n46113 = n45449 ^ n45316;
  assign n46114 = n46113 ^ n45317;
  assign n46115 = n46114 ^ n44749;
  assign n46116 = n46115 ^ n45482;
  assign n46111 = n46046 ^ n45944;
  assign n46112 = n46111 ^ n45945;
  assign n46117 = n46116 ^ n46112;
  assign n46119 = n45446 ^ n45323;
  assign n46120 = n46119 ^ n44753;
  assign n46121 = n46120 ^ n45124;
  assign n46118 = n46043 ^ n45951;
  assign n46122 = n46121 ^ n46118;
  assign n46125 = n45443 ^ n45326;
  assign n46126 = n46125 ^ n45327;
  assign n46127 = n46126 ^ n44782;
  assign n46128 = n46127 ^ n44682;
  assign n46123 = n46040 ^ n45954;
  assign n46124 = n46123 ^ n45955;
  assign n46129 = n46128 ^ n46124;
  assign n46134 = n45108 ^ n44706;
  assign n46135 = n46134 ^ n45760;
  assign n46133 = n46031 ^ n45971;
  assign n46136 = n46135 ^ n46133;
  assign n46138 = n45501 ^ n45101;
  assign n46139 = n46138 ^ n44711;
  assign n46137 = n46028 ^ n45976;
  assign n46140 = n46139 ^ n46137;
  assign n46143 = n45507 ^ n45094;
  assign n46144 = n46143 ^ n44503;
  assign n46141 = n46025 ^ n45979;
  assign n46142 = n46141 ^ n45980;
  assign n46145 = n46144 ^ n46142;
  assign n46148 = n45511 ^ n44412;
  assign n46149 = n46148 ^ n44698;
  assign n46146 = n46022 ^ n45985;
  assign n46147 = n46146 ^ n45982;
  assign n46150 = n46149 ^ n46147;
  assign n46436 = n46005 ^ n45991;
  assign n46437 = n46436 ^ n45992;
  assign n46155 = n45996 ^ n45873;
  assign n46156 = n46155 ^ n46001;
  assign n46153 = n45528 ^ n44385;
  assign n46154 = n46153 ^ n44717;
  assign n46157 = n46156 ^ n46154;
  assign n46396 = n44725 ^ n44371;
  assign n46397 = n46396 ^ n45536;
  assign n46168 = n44322 ^ n43677;
  assign n46169 = n46168 ^ n45024;
  assign n46170 = n46169 ^ n46090;
  assign n46171 = n44331 ^ n43673;
  assign n46172 = n46171 ^ n45592;
  assign n46173 = n46172 ^ n46096;
  assign n46174 = n44324 ^ n43666;
  assign n46175 = n46174 ^ n45553;
  assign n46176 = n46175 ^ n46102;
  assign n46177 = n44908 ^ n44246;
  assign n46178 = n46177 ^ n45557;
  assign n46179 = n46178 ^ n46106;
  assign n46180 = n44820 ^ n43485;
  assign n46181 = n46180 ^ n45561;
  assign n46182 = n46181 ^ n46114;
  assign n46183 = n44813 ^ n44143;
  assign n46184 = n46183 ^ n45565;
  assign n46185 = n46184 ^ n46119;
  assign n46186 = n44144 ^ n44113;
  assign n46187 = n46186 ^ n45569;
  assign n46188 = n46187 ^ n46126;
  assign n45919 = n44685 ^ n44172;
  assign n45920 = n45919 ^ n45482;
  assign n45918 = n45440 ^ n45439;
  assign n45921 = n45920 ^ n45918;
  assign n45904 = n45763 ^ n45760;
  assign n45905 = n45761 & n45904;
  assign n45906 = n45905 ^ n45763;
  assign n45901 = n44692 ^ n44165;
  assign n45902 = n45901 ^ n45124;
  assign n45914 = n45906 ^ n45902;
  assign n45900 = n45435 ^ n45336;
  assign n45915 = n45906 ^ n45900;
  assign n45916 = n45914 & n45915;
  assign n45917 = n45916 ^ n45902;
  assign n46189 = n45918 ^ n45917;
  assign n46190 = ~n45921 & n46189;
  assign n46191 = n46190 ^ n45920;
  assign n46192 = n46191 ^ n46126;
  assign n46193 = ~n46188 & ~n46192;
  assign n46194 = n46193 ^ n46187;
  assign n46195 = n46194 ^ n46119;
  assign n46196 = n46185 & ~n46195;
  assign n46197 = n46196 ^ n46184;
  assign n46198 = n46197 ^ n46114;
  assign n46199 = n46182 & ~n46198;
  assign n46200 = n46199 ^ n46181;
  assign n46201 = n46200 ^ n46106;
  assign n46202 = ~n46179 & ~n46201;
  assign n46203 = n46202 ^ n46178;
  assign n46204 = n46203 ^ n46102;
  assign n46205 = ~n46176 & ~n46204;
  assign n46206 = n46205 ^ n46175;
  assign n46207 = n46206 ^ n46172;
  assign n46208 = ~n46173 & n46207;
  assign n46209 = n46208 ^ n46096;
  assign n46210 = n46209 ^ n46090;
  assign n46211 = ~n46170 & ~n46210;
  assign n46212 = n46211 ^ n46169;
  assign n46165 = n44317 ^ n43665;
  assign n46166 = n46165 ^ n45029;
  assign n46167 = n46166 ^ n46085;
  assign n46223 = n46212 ^ n46167;
  assign n46224 = n46223 ^ n42979;
  assign n46225 = n46209 ^ n46169;
  assign n46226 = n46225 ^ n46090;
  assign n46227 = n46226 ^ n42981;
  assign n46228 = n46206 ^ n46173;
  assign n46229 = n46228 ^ n42989;
  assign n46230 = n46203 ^ n46176;
  assign n46231 = n46230 ^ n42982;
  assign n46232 = n46200 ^ n46179;
  assign n46233 = n46232 ^ n43612;
  assign n46234 = n46197 ^ n46182;
  assign n46235 = n46234 ^ n43486;
  assign n46236 = n46194 ^ n46185;
  assign n46237 = n46236 ^ n43536;
  assign n46238 = n46191 ^ n46188;
  assign n46239 = n46238 ^ n43537;
  assign n45922 = n45921 ^ n45917;
  assign n45923 = n45922 ^ n43538;
  assign n45903 = n45902 ^ n45900;
  assign n45907 = n45906 ^ n45903;
  assign n45908 = n45907 ^ n43539;
  assign n45897 = n45856 ^ n45764;
  assign n45898 = ~n45765 & ~n45897;
  assign n45899 = n45898 ^ n43469;
  assign n45911 = n45907 ^ n45899;
  assign n45912 = ~n45908 & n45911;
  assign n45913 = n45912 ^ n43539;
  assign n46240 = n45922 ^ n45913;
  assign n46241 = ~n45923 & n46240;
  assign n46242 = n46241 ^ n43538;
  assign n46243 = n46242 ^ n46238;
  assign n46244 = n46239 & n46243;
  assign n46245 = n46244 ^ n43537;
  assign n46246 = n46245 ^ n46236;
  assign n46247 = n46237 & ~n46246;
  assign n46248 = n46247 ^ n43536;
  assign n46249 = n46248 ^ n46234;
  assign n46250 = ~n46235 & ~n46249;
  assign n46251 = n46250 ^ n43486;
  assign n46252 = n46251 ^ n46232;
  assign n46253 = ~n46233 & ~n46252;
  assign n46254 = n46253 ^ n43612;
  assign n46255 = n46254 ^ n46230;
  assign n46256 = ~n46231 & ~n46255;
  assign n46257 = n46256 ^ n42982;
  assign n46258 = n46257 ^ n46228;
  assign n46259 = ~n46229 & ~n46258;
  assign n46260 = n46259 ^ n42989;
  assign n46261 = n46260 ^ n46226;
  assign n46262 = n46227 & n46261;
  assign n46263 = n46262 ^ n42981;
  assign n46264 = n46263 ^ n46223;
  assign n46265 = ~n46224 & ~n46264;
  assign n46266 = n46265 ^ n42979;
  assign n46213 = n46212 ^ n46085;
  assign n46214 = n46167 & ~n46213;
  assign n46215 = n46214 ^ n46166;
  assign n46162 = n44314 ^ n43664;
  assign n46163 = n46162 ^ n45021;
  assign n46079 = n45475 ^ n45296;
  assign n46164 = n46163 ^ n46079;
  assign n46221 = n46215 ^ n46164;
  assign n46222 = n46221 ^ n42976;
  assign n46291 = n46266 ^ n46222;
  assign n46271 = n46257 ^ n42989;
  assign n46272 = n46271 ^ n46228;
  assign n46273 = n46254 ^ n46231;
  assign n46274 = n46251 ^ n46233;
  assign n46275 = n46248 ^ n43486;
  assign n46276 = n46275 ^ n46234;
  assign n45896 = ~n45857 & ~n45895;
  assign n45909 = n45908 ^ n45899;
  assign n45910 = n45896 & n45909;
  assign n45924 = n45923 ^ n45913;
  assign n46277 = n45910 & n45924;
  assign n46278 = n46242 ^ n43537;
  assign n46279 = n46278 ^ n46238;
  assign n46280 = ~n46277 & n46279;
  assign n46281 = n46245 ^ n46237;
  assign n46282 = n46280 & ~n46281;
  assign n46283 = ~n46276 & ~n46282;
  assign n46284 = n46274 & n46283;
  assign n46285 = n46273 & ~n46284;
  assign n46286 = n46272 & ~n46285;
  assign n46287 = n46260 ^ n46227;
  assign n46288 = ~n46286 & ~n46287;
  assign n46289 = n46263 ^ n46224;
  assign n46290 = ~n46288 & n46289;
  assign n46316 = n46291 ^ n46290;
  assign n46313 = n44263 ^ n36290;
  assign n46314 = n46313 ^ n40816;
  assign n46315 = n46314 ^ n1794;
  assign n46317 = n46316 ^ n46315;
  assign n46319 = n44269 ^ n1697;
  assign n46320 = n46319 ^ n40726;
  assign n46321 = n46320 ^ n34839;
  assign n46318 = n46289 ^ n46288;
  assign n46322 = n46321 ^ n46318;
  assign n46326 = n46287 ^ n46286;
  assign n46323 = n44273 ^ n36297;
  assign n46324 = n46323 ^ n40731;
  assign n46325 = n46324 ^ n34716;
  assign n46327 = n46326 ^ n46325;
  assign n46331 = n46285 ^ n46272;
  assign n46328 = n44289 ^ n3002;
  assign n46329 = n46328 ^ n40803;
  assign n46330 = n46329 ^ n34721;
  assign n46332 = n46331 ^ n46330;
  assign n46333 = n46284 ^ n46273;
  assign n46337 = n46336 ^ n46333;
  assign n46341 = n46283 ^ n46274;
  assign n46338 = n44095 ^ n36307;
  assign n46339 = n46338 ^ n40742;
  assign n46340 = n46339 ^ n3113;
  assign n46342 = n46341 ^ n46340;
  assign n46346 = n46282 ^ n46276;
  assign n46343 = n43490 ^ n36312;
  assign n46344 = n46343 ^ n3095;
  assign n46345 = n46344 ^ n2702;
  assign n46347 = n46346 ^ n46345;
  assign n46349 = n43932 ^ n36317;
  assign n46350 = n46349 ^ n2624;
  assign n46351 = n46350 ^ n3093;
  assign n46348 = n46281 ^ n46280;
  assign n46352 = n46351 ^ n46348;
  assign n46356 = n46279 ^ n46277;
  assign n46353 = n43937 ^ n3071;
  assign n46354 = n46353 ^ n40784;
  assign n46355 = n46354 ^ n2616;
  assign n46357 = n46356 ^ n46355;
  assign n45927 = n43944 ^ n36325;
  assign n45928 = n45927 ^ n40757;
  assign n45929 = n45928 ^ n34741;
  assign n45926 = n45909 ^ n45896;
  assign n45930 = n45929 ^ n45926;
  assign n46070 = n46069 ^ n45931;
  assign n46071 = ~n46066 & n46070;
  assign n46072 = n46071 ^ n46069;
  assign n46073 = n46072 ^ n45926;
  assign n46074 = n45930 & ~n46073;
  assign n46075 = n46074 ^ n45929;
  assign n45925 = n45924 ^ n45910;
  assign n46076 = n46075 ^ n45925;
  assign n45498 = n44080 ^ n2531;
  assign n45499 = n45498 ^ n40752;
  assign n45500 = n45499 ^ n3179;
  assign n46358 = n45925 ^ n45500;
  assign n46359 = ~n46076 & n46358;
  assign n46360 = n46359 ^ n45500;
  assign n46361 = n46360 ^ n46356;
  assign n46362 = n46357 & ~n46361;
  assign n46363 = n46362 ^ n46355;
  assign n46364 = n46363 ^ n46351;
  assign n46365 = n46352 & ~n46364;
  assign n46366 = n46365 ^ n46348;
  assign n46367 = n46366 ^ n46346;
  assign n46368 = n46347 & ~n46367;
  assign n46369 = n46368 ^ n46345;
  assign n46370 = n46369 ^ n46341;
  assign n46371 = n46342 & ~n46370;
  assign n46372 = n46371 ^ n46340;
  assign n46373 = n46372 ^ n46333;
  assign n46374 = n46337 & ~n46373;
  assign n46375 = n46374 ^ n46336;
  assign n46376 = n46375 ^ n46331;
  assign n46377 = ~n46332 & n46376;
  assign n46378 = n46377 ^ n46330;
  assign n46379 = n46378 ^ n46326;
  assign n46380 = ~n46327 & n46379;
  assign n46381 = n46380 ^ n46325;
  assign n46382 = n46381 ^ n46321;
  assign n46383 = ~n46322 & ~n46382;
  assign n46384 = n46383 ^ n46318;
  assign n46385 = n46384 ^ n46316;
  assign n46386 = n46317 & n46385;
  assign n46387 = n46386 ^ n46315;
  assign n46292 = n46290 & n46291;
  assign n46267 = n46266 ^ n46221;
  assign n46268 = n46222 & ~n46267;
  assign n46269 = n46268 ^ n42976;
  assign n46216 = n46215 ^ n46079;
  assign n46217 = ~n46164 & n46216;
  assign n46218 = n46217 ^ n46163;
  assign n46159 = n44138 ^ n43532;
  assign n46160 = n46159 ^ n45019;
  assign n45495 = n45494 ^ n45478;
  assign n46161 = n46160 ^ n45495;
  assign n46219 = n46218 ^ n46161;
  assign n46220 = n46219 ^ n42637;
  assign n46270 = n46269 ^ n46220;
  assign n46312 = n46292 ^ n46270;
  assign n46388 = n46387 ^ n46312;
  assign n46389 = n44258 ^ n36285;
  assign n46390 = n46389 ^ n1802;
  assign n46391 = n46390 ^ n34709;
  assign n46392 = n46391 ^ n46312;
  assign n46393 = ~n46388 & n46392;
  assign n46394 = n46393 ^ n46391;
  assign n46305 = n46269 ^ n46219;
  assign n46306 = ~n46220 & ~n46305;
  assign n46307 = n46306 ^ n42637;
  assign n46308 = n46307 ^ n42633;
  assign n46301 = n46218 ^ n45495;
  assign n46302 = ~n46161 & n46301;
  assign n46303 = n46302 ^ n46160;
  assign n46298 = n44134 ^ n43530;
  assign n46299 = n46298 ^ n45016;
  assign n46297 = n45669 ^ n45666;
  assign n46300 = n46299 ^ n46297;
  assign n46304 = n46303 ^ n46300;
  assign n46309 = n46308 ^ n46304;
  assign n46294 = n44310 ^ n36281;
  assign n46295 = n46294 ^ n40717;
  assign n46296 = n46295 ^ n1904;
  assign n46310 = n46309 ^ n46296;
  assign n46293 = n46270 & ~n46292;
  assign n46311 = n46310 ^ n46293;
  assign n46395 = n46394 ^ n46311;
  assign n46398 = n46397 ^ n46395;
  assign n46401 = n46391 ^ n46388;
  assign n46399 = n44727 ^ n44123;
  assign n46400 = n46399 ^ n45540;
  assign n46402 = n46401 ^ n46400;
  assign n46408 = n44734 ^ n44128;
  assign n46409 = n46408 ^ n45548;
  assign n46404 = n45054 ^ n44130;
  assign n46405 = n46404 ^ n45552;
  assign n46406 = n46378 ^ n46327;
  assign n46407 = n46405 & ~n46406;
  assign n46410 = n46409 ^ n46407;
  assign n46411 = n46381 ^ n46322;
  assign n46412 = n46411 ^ n46409;
  assign n46413 = n46410 & n46412;
  assign n46414 = n46413 ^ n46407;
  assign n46403 = n46384 ^ n46317;
  assign n46415 = n46414 ^ n46403;
  assign n46416 = n44728 ^ n44125;
  assign n46417 = n46416 ^ n45543;
  assign n46418 = n46417 ^ n46403;
  assign n46419 = n46415 & n46418;
  assign n46420 = n46419 ^ n46417;
  assign n46421 = n46420 ^ n46401;
  assign n46422 = ~n46402 & n46421;
  assign n46423 = n46422 ^ n46400;
  assign n46424 = n46423 ^ n46397;
  assign n46425 = n46398 & ~n46424;
  assign n46426 = n46425 ^ n46395;
  assign n46427 = n46426 ^ n46158;
  assign n46428 = n45532 ^ n44721;
  assign n46429 = n46428 ^ n44378;
  assign n46430 = n46429 ^ n46158;
  assign n46431 = n46427 & ~n46430;
  assign n46432 = n46431 ^ n46429;
  assign n46433 = n46432 ^ n46156;
  assign n46434 = ~n46157 & ~n46433;
  assign n46435 = n46434 ^ n46154;
  assign n46438 = n46437 ^ n46435;
  assign n46439 = n45522 ^ n44713;
  assign n46440 = n46439 ^ n44392;
  assign n46441 = n46440 ^ n46437;
  assign n46442 = n46438 & n46441;
  assign n46443 = n46442 ^ n46440;
  assign n46152 = n46012 ^ n46009;
  assign n46444 = n46443 ^ n46152;
  assign n46445 = n44708 ^ n44120;
  assign n46446 = n46445 ^ n45518;
  assign n46447 = n46446 ^ n46152;
  assign n46448 = ~n46444 & n46447;
  assign n46449 = n46448 ^ n46446;
  assign n46151 = n46019 ^ n46016;
  assign n46450 = n46449 ^ n46151;
  assign n46451 = n45514 ^ n44405;
  assign n46452 = n46451 ^ n44703;
  assign n46453 = n46452 ^ n46151;
  assign n46454 = n46450 & n46453;
  assign n46455 = n46454 ^ n46452;
  assign n46456 = n46455 ^ n46147;
  assign n46457 = n46150 & ~n46456;
  assign n46458 = n46457 ^ n46149;
  assign n46459 = n46458 ^ n46142;
  assign n46460 = ~n46145 & ~n46459;
  assign n46461 = n46460 ^ n46144;
  assign n46462 = n46461 ^ n46139;
  assign n46463 = ~n46140 & n46462;
  assign n46464 = n46463 ^ n46137;
  assign n46465 = n46464 ^ n46135;
  assign n46466 = ~n46136 & ~n46465;
  assign n46467 = n46466 ^ n46133;
  assign n46132 = n46034 ^ n45966;
  assign n46468 = n46467 ^ n46132;
  assign n46469 = n44701 ^ n44690;
  assign n46470 = n46469 ^ n45900;
  assign n46471 = n46470 ^ n46132;
  assign n46472 = ~n46468 & ~n46471;
  assign n46473 = n46472 ^ n46470;
  assign n46130 = n46037 ^ n45959;
  assign n46131 = n46130 ^ n45960;
  assign n46474 = n46473 ^ n46131;
  assign n46475 = n45918 ^ n44696;
  assign n46476 = n46475 ^ n44684;
  assign n46477 = n46476 ^ n46131;
  assign n46478 = ~n46474 & ~n46477;
  assign n46479 = n46478 ^ n46476;
  assign n46480 = n46479 ^ n46124;
  assign n46481 = ~n46129 & ~n46480;
  assign n46482 = n46481 ^ n46128;
  assign n46483 = n46482 ^ n46118;
  assign n46484 = ~n46122 & ~n46483;
  assign n46485 = n46484 ^ n46121;
  assign n46486 = n46485 ^ n46116;
  assign n46487 = n46117 & ~n46486;
  assign n46488 = n46487 ^ n46112;
  assign n46489 = n46488 ^ n46109;
  assign n46490 = n46110 & n46489;
  assign n46491 = n46490 ^ n46108;
  assign n46492 = n46491 ^ n46101;
  assign n46493 = n46105 & n46492;
  assign n46494 = n46493 ^ n46104;
  assign n46495 = n46494 ^ n46099;
  assign n46496 = ~n46100 & n46495;
  assign n46497 = n46496 ^ n46098;
  assign n46498 = n46497 ^ n46093;
  assign n46499 = ~n46094 & n46498;
  assign n46500 = n46499 ^ n46092;
  assign n46501 = n46500 ^ n46088;
  assign n46502 = n46089 & ~n46501;
  assign n46503 = n46502 ^ n46087;
  assign n46082 = n46072 ^ n45930;
  assign n46080 = n46079 ^ n44908;
  assign n46081 = n46080 ^ n45592;
  assign n46083 = n46082 ^ n46081;
  assign n46509 = n46503 ^ n46083;
  assign n46510 = n46509 ^ n44246;
  assign n46511 = n46500 ^ n46087;
  assign n46512 = n46511 ^ n46088;
  assign n46513 = n46512 ^ n43485;
  assign n46515 = n46494 ^ n46100;
  assign n46516 = n46515 ^ n44144;
  assign n46517 = n46491 ^ n46104;
  assign n46518 = n46517 ^ n46101;
  assign n46519 = n46518 ^ n44172;
  assign n46520 = n46488 ^ n46108;
  assign n46521 = n46520 ^ n46109;
  assign n46522 = n46521 ^ n44165;
  assign n46524 = n46482 ^ n46122;
  assign n46525 = n46524 ^ n44154;
  assign n46526 = n46479 ^ n46129;
  assign n46527 = n46526 ^ n44105;
  assign n46528 = n46476 ^ n46474;
  assign n46529 = n46528 ^ n43771;
  assign n46532 = n46458 ^ n46144;
  assign n46533 = n46532 ^ n46142;
  assign n46534 = n46533 ^ n43497;
  assign n46535 = n46455 ^ n46150;
  assign n46536 = n46535 ^ n43500;
  assign n46537 = n46452 ^ n46450;
  assign n46538 = n46537 ^ n43504;
  assign n46540 = n46440 ^ n46438;
  assign n46541 = n46540 ^ n43509;
  assign n46543 = n46429 ^ n46427;
  assign n46544 = n46543 ^ n43517;
  assign n46545 = n46420 ^ n46402;
  assign n46546 = n46545 ^ n43521;
  assign n46548 = n46406 ^ n46405;
  assign n46549 = ~n43702 & ~n46548;
  assign n46550 = n46549 ^ n43525;
  assign n46551 = n46411 ^ n46410;
  assign n46552 = n46551 ^ n46549;
  assign n46553 = ~n46550 & n46552;
  assign n46554 = n46553 ^ n43525;
  assign n46547 = n46417 ^ n46415;
  assign n46555 = n46554 ^ n46547;
  assign n46556 = n46547 ^ n43712;
  assign n46557 = n46555 & ~n46556;
  assign n46558 = n46557 ^ n43712;
  assign n46559 = n46558 ^ n46545;
  assign n46560 = n46546 & n46559;
  assign n46561 = n46560 ^ n43521;
  assign n46562 = n46561 ^ n43722;
  assign n46563 = n46423 ^ n46398;
  assign n46564 = n46563 ^ n46561;
  assign n46565 = ~n46562 & n46564;
  assign n46566 = n46565 ^ n43722;
  assign n46567 = n46566 ^ n46543;
  assign n46568 = ~n46544 & n46567;
  assign n46569 = n46568 ^ n43517;
  assign n46542 = n46432 ^ n46157;
  assign n46570 = n46569 ^ n46542;
  assign n46571 = n46542 ^ n43513;
  assign n46572 = n46570 & ~n46571;
  assign n46573 = n46572 ^ n43513;
  assign n46574 = n46573 ^ n46540;
  assign n46575 = n46541 & n46574;
  assign n46576 = n46575 ^ n43509;
  assign n46539 = n46446 ^ n46444;
  assign n46577 = n46576 ^ n46539;
  assign n46578 = n46539 ^ n43506;
  assign n46579 = n46577 & n46578;
  assign n46580 = n46579 ^ n43506;
  assign n46581 = n46580 ^ n46537;
  assign n46582 = ~n46538 & ~n46581;
  assign n46583 = n46582 ^ n43504;
  assign n46584 = n46583 ^ n46535;
  assign n46585 = ~n46536 & ~n46584;
  assign n46586 = n46585 ^ n43500;
  assign n46587 = n46586 ^ n46533;
  assign n46588 = n46534 & ~n46587;
  assign n46589 = n46588 ^ n43497;
  assign n46590 = n46589 ^ n43495;
  assign n46591 = n46461 ^ n46140;
  assign n46592 = n46591 ^ n46589;
  assign n46593 = ~n46590 & n46592;
  assign n46594 = n46593 ^ n43495;
  assign n46531 = n46464 ^ n46136;
  assign n46595 = n46594 ^ n46531;
  assign n46596 = n46531 ^ n43492;
  assign n46597 = ~n46595 & n46596;
  assign n46598 = n46597 ^ n43492;
  assign n46530 = n46470 ^ n46468;
  assign n46599 = n46598 ^ n46530;
  assign n46600 = n46530 ^ n43491;
  assign n46601 = n46599 & n46600;
  assign n46602 = n46601 ^ n43491;
  assign n46603 = n46602 ^ n46528;
  assign n46604 = ~n46529 & n46603;
  assign n46605 = n46604 ^ n43771;
  assign n46606 = n46605 ^ n46526;
  assign n46607 = ~n46527 & ~n46606;
  assign n46608 = n46607 ^ n44105;
  assign n46609 = n46608 ^ n46524;
  assign n46610 = ~n46525 & ~n46609;
  assign n46611 = n46610 ^ n44154;
  assign n46523 = n46485 ^ n46117;
  assign n46612 = n46611 ^ n46523;
  assign n46613 = n46523 ^ n44150;
  assign n46614 = n46612 & ~n46613;
  assign n46615 = n46614 ^ n44150;
  assign n46616 = n46615 ^ n46521;
  assign n46617 = n46522 & n46616;
  assign n46618 = n46617 ^ n44165;
  assign n46619 = n46618 ^ n46518;
  assign n46620 = n46519 & n46619;
  assign n46621 = n46620 ^ n44172;
  assign n46622 = n46621 ^ n46515;
  assign n46623 = n46516 & ~n46622;
  assign n46624 = n46623 ^ n44144;
  assign n46514 = n46497 ^ n46094;
  assign n46625 = n46624 ^ n46514;
  assign n46626 = n46514 ^ n44143;
  assign n46627 = ~n46625 & ~n46626;
  assign n46628 = n46627 ^ n44143;
  assign n46629 = n46628 ^ n46512;
  assign n46630 = n46513 & ~n46629;
  assign n46631 = n46630 ^ n43485;
  assign n46632 = n46631 ^ n46509;
  assign n46633 = n46510 & n46632;
  assign n46634 = n46633 ^ n44246;
  assign n46504 = n46503 ^ n46082;
  assign n46505 = ~n46083 & ~n46504;
  assign n46506 = n46505 ^ n46081;
  assign n46077 = n46076 ^ n45500;
  assign n45496 = n45495 ^ n44324;
  assign n45497 = n45496 ^ n45024;
  assign n46078 = n46077 ^ n45497;
  assign n46507 = n46506 ^ n46078;
  assign n46508 = n46507 ^ n43666;
  assign n46635 = n46634 ^ n46508;
  assign n46636 = n46631 ^ n46510;
  assign n46637 = n46621 ^ n46516;
  assign n46638 = n46618 ^ n46519;
  assign n46639 = n46608 ^ n44154;
  assign n46640 = n46639 ^ n46524;
  assign n46641 = n46602 ^ n46529;
  assign n46642 = n46599 ^ n43491;
  assign n46643 = n46595 ^ n43492;
  assign n46644 = n46586 ^ n46534;
  assign n46645 = n46580 ^ n46538;
  assign n46646 = n46570 ^ n43513;
  assign n46647 = n46566 ^ n46544;
  assign n46648 = n46558 ^ n46546;
  assign n46649 = n46555 ^ n43712;
  assign n46650 = n46551 ^ n46550;
  assign n46651 = ~n46649 & ~n46650;
  assign n46652 = ~n46648 & ~n46651;
  assign n46653 = n46563 ^ n46562;
  assign n46654 = ~n46652 & ~n46653;
  assign n46655 = n46647 & ~n46654;
  assign n46656 = ~n46646 & ~n46655;
  assign n46657 = n46573 ^ n46541;
  assign n46658 = n46656 & n46657;
  assign n46659 = n46577 ^ n43506;
  assign n46660 = n46658 & ~n46659;
  assign n46661 = n46645 & ~n46660;
  assign n46662 = n46583 ^ n43500;
  assign n46663 = n46662 ^ n46535;
  assign n46664 = n46661 & ~n46663;
  assign n46665 = ~n46644 & n46664;
  assign n46666 = n46591 ^ n43495;
  assign n46667 = n46666 ^ n46589;
  assign n46668 = n46665 & ~n46667;
  assign n46669 = n46643 & n46668;
  assign n46670 = ~n46642 & ~n46669;
  assign n46671 = ~n46641 & n46670;
  assign n46672 = n46605 ^ n46527;
  assign n46673 = ~n46671 & n46672;
  assign n46674 = n46640 & ~n46673;
  assign n46675 = n46612 ^ n44150;
  assign n46676 = ~n46674 & n46675;
  assign n46677 = n46615 ^ n46522;
  assign n46678 = n46676 & ~n46677;
  assign n46679 = n46638 & n46678;
  assign n46680 = n46637 & ~n46679;
  assign n46681 = n46625 ^ n44143;
  assign n46682 = n46680 & ~n46681;
  assign n46683 = n46628 ^ n46513;
  assign n46684 = ~n46682 & n46683;
  assign n46685 = n46636 & n46684;
  assign n46885 = ~n46635 & ~n46685;
  assign n46896 = n46634 ^ n46507;
  assign n46897 = n46634 ^ n43666;
  assign n46898 = n46896 & n46897;
  assign n46899 = n46898 ^ n43666;
  assign n46891 = n46506 ^ n45497;
  assign n46892 = ~n46078 & ~n46891;
  assign n46893 = n46892 ^ n46077;
  assign n46888 = n46360 ^ n46355;
  assign n46889 = n46888 ^ n46356;
  assign n46886 = n45029 ^ n44331;
  assign n46887 = n46886 ^ n46297;
  assign n46890 = n46889 ^ n46887;
  assign n46894 = n46893 ^ n46890;
  assign n46895 = n46894 ^ n43673;
  assign n46900 = n46899 ^ n46895;
  assign n47008 = ~n46885 & n46900;
  assign n46987 = n46363 ^ n46352;
  assign n46984 = n45693 ^ n45021;
  assign n46985 = n46984 ^ n44322;
  assign n47000 = n46987 ^ n46985;
  assign n46981 = n46893 ^ n46889;
  assign n46982 = ~n46890 & ~n46981;
  assign n46983 = n46982 ^ n46887;
  assign n47001 = n47000 ^ n46983;
  assign n47006 = n47001 ^ n43677;
  assign n46996 = n46899 ^ n46894;
  assign n46997 = ~n46895 & ~n46996;
  assign n46998 = n46997 ^ n43673;
  assign n47007 = n47006 ^ n46998;
  assign n47079 = n47008 ^ n47007;
  assign n47103 = n47079 ^ n47077;
  assign n46901 = n46900 ^ n46885;
  assign n46881 = n44943 ^ n36962;
  assign n46882 = n46881 ^ n2894;
  assign n46883 = n46882 ^ n35472;
  assign n47071 = n46901 ^ n46883;
  assign n46686 = n46685 ^ n46635;
  assign n3132 = n3131 ^ n3119;
  assign n3136 = n3135 ^ n3132;
  assign n3137 = n3136 ^ n2892;
  assign n46687 = n46686 ^ n3137;
  assign n46688 = n46684 ^ n46636;
  assign n2763 = n2762 ^ n2738;
  assign n2797 = n2796 ^ n2763;
  assign n2804 = n2803 ^ n2797;
  assign n46689 = n46688 ^ n2804;
  assign n46693 = n46683 ^ n46682;
  assign n46690 = n44979 ^ n3105;
  assign n46691 = n46690 ^ n3215;
  assign n46692 = n46691 ^ n2788;
  assign n46694 = n46693 ^ n46692;
  assign n46698 = n46681 ^ n46680;
  assign n46695 = n44951 ^ n2673;
  assign n46696 = n46695 ^ n41455;
  assign n46697 = n46696 ^ n3213;
  assign n46699 = n46698 ^ n46697;
  assign n46703 = n46679 ^ n46637;
  assign n46700 = n44956 ^ n3191;
  assign n46701 = n46700 ^ n41460;
  assign n46702 = n46701 ^ n35485;
  assign n46704 = n46703 ^ n46702;
  assign n46708 = n46678 ^ n46638;
  assign n46705 = n44966 ^ n36977;
  assign n46706 = n46705 ^ n41510;
  assign n46707 = n46706 ^ n35489;
  assign n46709 = n46708 ^ n46707;
  assign n46713 = n46677 ^ n46676;
  assign n46710 = n44117 ^ n36982;
  assign n46711 = n46710 ^ n41467;
  assign n46712 = n46711 ^ n35494;
  assign n46714 = n46713 ^ n46712;
  assign n46716 = n36986 ^ n1486;
  assign n46717 = n46716 ^ n41471;
  assign n46718 = n46717 ^ n35499;
  assign n46715 = n46675 ^ n46674;
  assign n46719 = n46718 ^ n46715;
  assign n46723 = n46673 ^ n46640;
  assign n46720 = n37027 ^ n1468;
  assign n46721 = n46720 ^ n41497;
  assign n46722 = n46721 ^ n35504;
  assign n46724 = n46723 ^ n46722;
  assign n46727 = n44557 ^ n1346;
  assign n46728 = n46727 ^ n41487;
  assign n46729 = n46728 ^ n35515;
  assign n46726 = n46670 ^ n46641;
  assign n46730 = n46729 ^ n46726;
  assign n46734 = n46669 ^ n46642;
  assign n46731 = n44562 ^ n3348;
  assign n46732 = n46731 ^ n41096;
  assign n46733 = n46732 ^ n35520;
  assign n46735 = n46734 ^ n46733;
  assign n46739 = n46668 ^ n46643;
  assign n46736 = n44567 ^ n37010;
  assign n46737 = n46736 ^ n41090;
  assign n46738 = n46737 ^ n950;
  assign n46740 = n46739 ^ n46738;
  assign n46744 = n46667 ^ n46665;
  assign n46741 = n44572 ^ n36999;
  assign n46742 = n46741 ^ n848;
  assign n46743 = n46742 ^ n35527;
  assign n46745 = n46744 ^ n46743;
  assign n46749 = n44584 ^ n36607;
  assign n46750 = n46749 ^ n41073;
  assign n46751 = n46750 ^ n35539;
  assign n46748 = n46660 ^ n46645;
  assign n46752 = n46751 ^ n46748;
  assign n46754 = n44642 ^ n36547;
  assign n46755 = n46754 ^ n41016;
  assign n46756 = n46755 ^ n35544;
  assign n46753 = n46659 ^ n46658;
  assign n46757 = n46756 ^ n46753;
  assign n46759 = n44590 ^ n36552;
  assign n46760 = n46759 ^ n41020;
  assign n46761 = n46760 ^ n35549;
  assign n46758 = n46657 ^ n46656;
  assign n46762 = n46761 ^ n46758;
  assign n46766 = n46655 ^ n46646;
  assign n46763 = n44632 ^ n36557;
  assign n46764 = n46763 ^ n41025;
  assign n46765 = n46764 ^ n35553;
  assign n46767 = n46766 ^ n46765;
  assign n46771 = n46654 ^ n46647;
  assign n46768 = n44595 ^ n36561;
  assign n46769 = n46768 ^ n41031;
  assign n46770 = n46769 ^ n35558;
  assign n46772 = n46771 ^ n46770;
  assign n46791 = n46651 ^ n46648;
  assign n1980 = n1979 ^ n1940;
  assign n2014 = n2013 ^ n1980;
  assign n2024 = n2023 ^ n2014;
  assign n46778 = n46548 ^ n43702;
  assign n46779 = n2024 & n46778;
  assign n46775 = n44613 ^ n36574;
  assign n46776 = n46775 ^ n41044;
  assign n46777 = n46776 ^ n2151;
  assign n46780 = n46779 ^ n46777;
  assign n46781 = n46779 ^ n46650;
  assign n46782 = n46780 & n46781;
  assign n46783 = n46782 ^ n46777;
  assign n46774 = n46650 ^ n46649;
  assign n46784 = n46783 ^ n46774;
  assign n46785 = n44610 ^ n36571;
  assign n46786 = n46785 ^ n2159;
  assign n46787 = n46786 ^ n34883;
  assign n46788 = n46787 ^ n46783;
  assign n46789 = n46784 & n46788;
  assign n46790 = n46789 ^ n46787;
  assign n46792 = n46791 ^ n46790;
  assign n46793 = n44606 ^ n36567;
  assign n46794 = n46793 ^ n41040;
  assign n46795 = n46794 ^ n2333;
  assign n46796 = n46795 ^ n46791;
  assign n46797 = ~n46792 & n46796;
  assign n46798 = n46797 ^ n46795;
  assign n46773 = n46653 ^ n46652;
  assign n46799 = n46798 ^ n46773;
  assign n46800 = n44600 ^ n36588;
  assign n46801 = n46800 ^ n41036;
  assign n46802 = n46801 ^ n35564;
  assign n46803 = n46802 ^ n46773;
  assign n46804 = n46799 & ~n46803;
  assign n46805 = n46804 ^ n46802;
  assign n46806 = n46805 ^ n46771;
  assign n46807 = ~n46772 & n46806;
  assign n46808 = n46807 ^ n46770;
  assign n46809 = n46808 ^ n46766;
  assign n46810 = ~n46767 & n46809;
  assign n46811 = n46810 ^ n46765;
  assign n46812 = n46811 ^ n46758;
  assign n46813 = ~n46762 & n46812;
  assign n46814 = n46813 ^ n46761;
  assign n46815 = n46814 ^ n46753;
  assign n46816 = n46757 & ~n46815;
  assign n46817 = n46816 ^ n46756;
  assign n46818 = n46817 ^ n46751;
  assign n46819 = ~n46752 & ~n46818;
  assign n46820 = n46819 ^ n46748;
  assign n46747 = n46663 ^ n46661;
  assign n46821 = n46820 ^ n46747;
  assign n46822 = n44652 ^ n740;
  assign n46823 = n46822 ^ n41010;
  assign n46824 = n46823 ^ n35534;
  assign n46825 = n46824 ^ n46747;
  assign n46826 = ~n46821 & ~n46825;
  assign n46827 = n46826 ^ n46824;
  assign n46746 = n46664 ^ n46644;
  assign n46828 = n46827 ^ n46746;
  assign n46829 = n44577 ^ n36616;
  assign n46830 = n46829 ^ n41005;
  assign n46831 = n46830 ^ n840;
  assign n46832 = n46831 ^ n46827;
  assign n46833 = n46828 & n46832;
  assign n46834 = n46833 ^ n46831;
  assign n46835 = n46834 ^ n46744;
  assign n46836 = ~n46745 & n46835;
  assign n46837 = n46836 ^ n46743;
  assign n46838 = n46837 ^ n46739;
  assign n46839 = n46740 & ~n46838;
  assign n46840 = n46839 ^ n46738;
  assign n46841 = n46840 ^ n46734;
  assign n46842 = ~n46735 & n46841;
  assign n46843 = n46842 ^ n46733;
  assign n46844 = n46843 ^ n46726;
  assign n46845 = n46730 & ~n46844;
  assign n46846 = n46845 ^ n46729;
  assign n46725 = n46672 ^ n46671;
  assign n46847 = n46846 ^ n46725;
  assign n46848 = n44552 ^ n1361;
  assign n46849 = n46848 ^ n41478;
  assign n46850 = n46849 ^ n35509;
  assign n46851 = n46850 ^ n46725;
  assign n46852 = n46847 & ~n46851;
  assign n46853 = n46852 ^ n46850;
  assign n46854 = n46853 ^ n46723;
  assign n46855 = n46724 & ~n46854;
  assign n46856 = n46855 ^ n46722;
  assign n46857 = n46856 ^ n46715;
  assign n46858 = ~n46719 & n46857;
  assign n46859 = n46858 ^ n46718;
  assign n46860 = n46859 ^ n46713;
  assign n46861 = ~n46714 & n46860;
  assign n46862 = n46861 ^ n46712;
  assign n46863 = n46862 ^ n46708;
  assign n46864 = n46709 & ~n46863;
  assign n46865 = n46864 ^ n46707;
  assign n46866 = n46865 ^ n46703;
  assign n46867 = n46704 & ~n46866;
  assign n46868 = n46867 ^ n46702;
  assign n46869 = n46868 ^ n46698;
  assign n46870 = n46699 & ~n46869;
  assign n46871 = n46870 ^ n46697;
  assign n46872 = n46871 ^ n46693;
  assign n46873 = ~n46694 & n46872;
  assign n46874 = n46873 ^ n46692;
  assign n46875 = n46874 ^ n46688;
  assign n46876 = n46689 & ~n46875;
  assign n46877 = n46876 ^ n2804;
  assign n46878 = n46877 ^ n46686;
  assign n46879 = ~n46687 & n46878;
  assign n46880 = n46879 ^ n3137;
  assign n47072 = n46901 ^ n46880;
  assign n47073 = ~n47071 & n47072;
  assign n47074 = n47073 ^ n46883;
  assign n47104 = n47103 ^ n47074;
  assign n47255 = n47106 ^ n47104;
  assign n47256 = n44130 & n47255;
  assign n47257 = n47256 ^ n44128;
  assign n47078 = n47077 ^ n47074;
  assign n47080 = n47079 ^ n47074;
  assign n47081 = n47078 & ~n47080;
  assign n47082 = n47081 ^ n47077;
  assign n47067 = n44999 ^ n36952;
  assign n47068 = n47067 ^ n41439;
  assign n47069 = n47068 ^ n35462;
  assign n47009 = n47007 & ~n47008;
  assign n46999 = n46998 ^ n43677;
  assign n47002 = n47001 ^ n46998;
  assign n47003 = ~n46999 & ~n47002;
  assign n47004 = n47003 ^ n43677;
  assign n46992 = n45019 ^ n44317;
  assign n46993 = n46992 ^ n45700;
  assign n46986 = n46985 ^ n46983;
  assign n46988 = n46987 ^ n46983;
  assign n46989 = n46986 & n46988;
  assign n46990 = n46989 ^ n46985;
  assign n46911 = n46366 ^ n46347;
  assign n46991 = n46990 ^ n46911;
  assign n46994 = n46993 ^ n46991;
  assign n46995 = n46994 ^ n43665;
  assign n47005 = n47004 ^ n46995;
  assign n47066 = n47009 ^ n47005;
  assign n47070 = n47069 ^ n47066;
  assign n47111 = n47082 ^ n47070;
  assign n47108 = n45540 ^ n44734;
  assign n47109 = n47108 ^ n46156;
  assign n47107 = n47104 & n47106;
  assign n47110 = n47109 ^ n47107;
  assign n47258 = n47111 ^ n47110;
  assign n47259 = n47258 ^ n47256;
  assign n47260 = n47257 & ~n47259;
  assign n47261 = n47260 ^ n44128;
  assign n47112 = n47111 ^ n47109;
  assign n47113 = n47110 & ~n47112;
  assign n47114 = n47113 ^ n47107;
  assign n47098 = n46437 ^ n44728;
  assign n47099 = n47098 ^ n45536;
  assign n47252 = n47114 ^ n47099;
  assign n47083 = n47082 ^ n47066;
  assign n47084 = n47070 & ~n47083;
  assign n47085 = n47084 ^ n47069;
  assign n47061 = n44932 ^ n37067;
  assign n47062 = n47061 ^ n41433;
  assign n47063 = n47062 ^ n35457;
  assign n47100 = n47085 ^ n47063;
  assign n47020 = n47004 ^ n46994;
  assign n47021 = n46995 & ~n47020;
  assign n47022 = n47021 ^ n43665;
  assign n47016 = n45016 ^ n44314;
  assign n47017 = n47016 ^ n45691;
  assign n47014 = n46369 ^ n46342;
  assign n47011 = n46993 ^ n46911;
  assign n47012 = n46991 & n47011;
  assign n47013 = n47012 ^ n46993;
  assign n47015 = n47014 ^ n47013;
  assign n47018 = n47017 ^ n47015;
  assign n47019 = n47018 ^ n43664;
  assign n47023 = n47022 ^ n47019;
  assign n47010 = ~n47005 & ~n47009;
  assign n47064 = n47023 ^ n47010;
  assign n47101 = n47100 ^ n47064;
  assign n47253 = n47252 ^ n47101;
  assign n47254 = n47253 ^ n44125;
  assign n47356 = n47261 ^ n47254;
  assign n47355 = n47258 ^ n47257;
  assign n47487 = n47356 ^ n47355;
  assign n2257 = n2247 ^ n2193;
  assign n2282 = n2281 ^ n2257;
  assign n2289 = n2288 ^ n2282;
  assign n47815 = n47487 ^ n2289;
  assign n47479 = n45381 ^ n2110;
  assign n47480 = n47479 ^ n41698;
  assign n47481 = n47480 ^ n2273;
  assign n47474 = n45639 ^ n2092;
  assign n47475 = n47474 ^ n42312;
  assign n47476 = n47475 ^ n36403;
  assign n47477 = n47255 ^ n44130;
  assign n47478 = n47476 & n47477;
  assign n47482 = n47481 ^ n47478;
  assign n47483 = n47478 ^ n47355;
  assign n47484 = n47482 & n47483;
  assign n47485 = n47484 ^ n47481;
  assign n47816 = n47815 ^ n47485;
  assign n47735 = n45645 ^ n37734;
  assign n47736 = n47735 ^ n42146;
  assign n47737 = n47736 ^ n36281;
  assign n49598 = n47737 ^ n40102;
  assign n49599 = n49598 ^ n44243;
  assign n49600 = n49599 ^ n38621;
  assign n46968 = n46787 ^ n46784;
  assign n49179 = n47816 ^ n46968;
  assign n48147 = n46296 ^ n38621;
  assign n48148 = n48147 ^ n42849;
  assign n48149 = n48148 ^ n1979;
  assign n47786 = n46437 ^ n45543;
  assign n46975 = n46778 ^ n2024;
  assign n47787 = n47786 ^ n46975;
  assign n47756 = n45665 ^ n37754;
  assign n47757 = n47756 ^ n3010;
  assign n47758 = n47757 ^ n36297;
  assign n47198 = n47014 ^ n45592;
  assign n47199 = n47198 ^ n46297;
  assign n46914 = n46856 ^ n46718;
  assign n46915 = n46914 ^ n46715;
  assign n46912 = n46911 ^ n45495;
  assign n46913 = n46912 ^ n45553;
  assign n46916 = n46915 ^ n46913;
  assign n47187 = n46853 ^ n46724;
  assign n46918 = n46889 ^ n45561;
  assign n46919 = n46918 ^ n46085;
  assign n46917 = n46850 ^ n46847;
  assign n46920 = n46919 ^ n46917;
  assign n46923 = n46090 ^ n46077;
  assign n46924 = n46923 ^ n45565;
  assign n46921 = n46843 ^ n46729;
  assign n46922 = n46921 ^ n46726;
  assign n46925 = n46924 ^ n46922;
  assign n46927 = n46096 ^ n46082;
  assign n46928 = n46927 ^ n45569;
  assign n46926 = n46840 ^ n46735;
  assign n46929 = n46928 ^ n46926;
  assign n46931 = n46102 ^ n45482;
  assign n46932 = n46931 ^ n46088;
  assign n46930 = n46837 ^ n46740;
  assign n46933 = n46932 ^ n46930;
  assign n46937 = n46114 ^ n44682;
  assign n46938 = n46937 ^ n46099;
  assign n46936 = n46831 ^ n46828;
  assign n46939 = n46938 ^ n46936;
  assign n46942 = n46109 ^ n44690;
  assign n46943 = n46942 ^ n46126;
  assign n46941 = n46817 ^ n46752;
  assign n46944 = n46943 ^ n46941;
  assign n46946 = n46112 ^ n45918;
  assign n46947 = n46946 ^ n45108;
  assign n46945 = n46814 ^ n46757;
  assign n46948 = n46947 ^ n46945;
  assign n46951 = n45900 ^ n45101;
  assign n46952 = n46951 ^ n46118;
  assign n46949 = n46811 ^ n46761;
  assign n46950 = n46949 ^ n46758;
  assign n46953 = n46952 ^ n46950;
  assign n46958 = n46132 ^ n45507;
  assign n46959 = n46958 ^ n44703;
  assign n46957 = n46802 ^ n46799;
  assign n46960 = n46959 ^ n46957;
  assign n46963 = n46133 ^ n44708;
  assign n46964 = n46963 ^ n45511;
  assign n46961 = n46795 ^ n46790;
  assign n46962 = n46961 ^ n46791;
  assign n46965 = n46964 ^ n46962;
  assign n46966 = n46137 ^ n44713;
  assign n46967 = n46966 ^ n45514;
  assign n46969 = n46968 ^ n46967;
  assign n46972 = n46777 ^ n46650;
  assign n46973 = n46972 ^ n46779;
  assign n46970 = n45518 ^ n44717;
  assign n46971 = n46970 ^ n46142;
  assign n46974 = n46973 ^ n46971;
  assign n46976 = n46147 ^ n45522;
  assign n46977 = n46976 ^ n44721;
  assign n46978 = n46977 ^ n46975;
  assign n47057 = n44927 ^ n1860;
  assign n47058 = n47057 ^ n41429;
  assign n47059 = n47058 ^ n35452;
  assign n47032 = n47022 ^ n47018;
  assign n47033 = ~n47019 & n47032;
  assign n47034 = n47033 ^ n43664;
  assign n47035 = n47034 ^ n43532;
  assign n47027 = n47017 ^ n47014;
  assign n47028 = ~n47015 & n47027;
  assign n47029 = n47028 ^ n47017;
  assign n46903 = n46372 ^ n46336;
  assign n46904 = n46903 ^ n46333;
  assign n47030 = n47029 ^ n46904;
  assign n47025 = n45707 ^ n44138;
  assign n47026 = n47025 ^ n44741;
  assign n47031 = n47030 ^ n47026;
  assign n47036 = n47035 ^ n47031;
  assign n47024 = n47010 & n47023;
  assign n47056 = n47036 ^ n47024;
  assign n47060 = n47059 ^ n47056;
  assign n47065 = n47064 ^ n47063;
  assign n47086 = n47085 ^ n47064;
  assign n47087 = n47065 & ~n47086;
  assign n47088 = n47087 ^ n47063;
  assign n47089 = n47088 ^ n47056;
  assign n47090 = n47060 & ~n47089;
  assign n47091 = n47090 ^ n47059;
  assign n47050 = n47026 ^ n46904;
  assign n47051 = ~n47030 & n47050;
  assign n47052 = n47051 ^ n47026;
  assign n47045 = n47031 ^ n43532;
  assign n47046 = n47034 ^ n47031;
  assign n47047 = n47045 & n47046;
  assign n47048 = n47047 ^ n43532;
  assign n47039 = n45012 ^ n37126;
  assign n47040 = n47039 ^ n41424;
  assign n47041 = n47040 ^ n2005;
  assign n47042 = n47041 ^ n44739;
  assign n47043 = n47042 ^ n46298;
  assign n47038 = n46375 ^ n46332;
  assign n47044 = n47043 ^ n47038;
  assign n47049 = n47048 ^ n47044;
  assign n47053 = n47052 ^ n47049;
  assign n47054 = n47053 ^ n45685;
  assign n47037 = ~n47024 & n47036;
  assign n47055 = n47054 ^ n47037;
  assign n47092 = n47091 ^ n47055;
  assign n46979 = n45528 ^ n44725;
  assign n46980 = n46979 ^ n46151;
  assign n47093 = n47092 ^ n46980;
  assign n47096 = n47088 ^ n47060;
  assign n47094 = n46152 ^ n44727;
  assign n47095 = n47094 ^ n45532;
  assign n47097 = n47096 ^ n47095;
  assign n47102 = n47101 ^ n47099;
  assign n47115 = n47114 ^ n47101;
  assign n47116 = n47102 & ~n47115;
  assign n47117 = n47116 ^ n47099;
  assign n47118 = n47117 ^ n47096;
  assign n47119 = n47097 & ~n47118;
  assign n47120 = n47119 ^ n47095;
  assign n47121 = n47120 ^ n47092;
  assign n47122 = ~n47093 & n47121;
  assign n47123 = n47122 ^ n46980;
  assign n47124 = n47123 ^ n46975;
  assign n47125 = n46978 & ~n47124;
  assign n47126 = n47125 ^ n46977;
  assign n47127 = n47126 ^ n46973;
  assign n47128 = n46974 & n47127;
  assign n47129 = n47128 ^ n46971;
  assign n47130 = n47129 ^ n46967;
  assign n47131 = ~n46969 & n47130;
  assign n47132 = n47131 ^ n46968;
  assign n47133 = n47132 ^ n46962;
  assign n47134 = ~n46965 & n47133;
  assign n47135 = n47134 ^ n46964;
  assign n47136 = n47135 ^ n46957;
  assign n47137 = n46960 & ~n47136;
  assign n47138 = n47137 ^ n46959;
  assign n46956 = n46805 ^ n46772;
  assign n47139 = n47138 ^ n46956;
  assign n47140 = n45501 ^ n44698;
  assign n47141 = n47140 ^ n46131;
  assign n47142 = n47141 ^ n46956;
  assign n47143 = ~n47139 & n47142;
  assign n47144 = n47143 ^ n47141;
  assign n46954 = n46808 ^ n46765;
  assign n46955 = n46954 ^ n46766;
  assign n47145 = n47144 ^ n46955;
  assign n47146 = n45760 ^ n45094;
  assign n47147 = n47146 ^ n46124;
  assign n47148 = n47147 ^ n46955;
  assign n47149 = ~n47145 & ~n47148;
  assign n47150 = n47149 ^ n47147;
  assign n47151 = n47150 ^ n46952;
  assign n47152 = n46953 & n47151;
  assign n47153 = n47152 ^ n46950;
  assign n47154 = n47153 ^ n46945;
  assign n47155 = ~n46948 & n47154;
  assign n47156 = n47155 ^ n46947;
  assign n47157 = n47156 ^ n46941;
  assign n47158 = n46944 & ~n47157;
  assign n47159 = n47158 ^ n46943;
  assign n46940 = n46824 ^ n46821;
  assign n47160 = n47159 ^ n46940;
  assign n47161 = n46119 ^ n44684;
  assign n47162 = n47161 ^ n46101;
  assign n47163 = n47162 ^ n46940;
  assign n47164 = n47160 & n47163;
  assign n47165 = n47164 ^ n47162;
  assign n47166 = n47165 ^ n46936;
  assign n47167 = n46939 & n47166;
  assign n47168 = n47167 ^ n46938;
  assign n46934 = n46834 ^ n46743;
  assign n46935 = n46934 ^ n46744;
  assign n47169 = n47168 ^ n46935;
  assign n47170 = n46093 ^ n45124;
  assign n47171 = n47170 ^ n46106;
  assign n47172 = n47171 ^ n46935;
  assign n47173 = ~n47169 & ~n47172;
  assign n47174 = n47173 ^ n47171;
  assign n47175 = n47174 ^ n46930;
  assign n47176 = ~n46933 & ~n47175;
  assign n47177 = n47176 ^ n46932;
  assign n47178 = n47177 ^ n46928;
  assign n47179 = n46929 & ~n47178;
  assign n47180 = n47179 ^ n46926;
  assign n47181 = n47180 ^ n46922;
  assign n47182 = ~n46925 & n47181;
  assign n47183 = n47182 ^ n46924;
  assign n47184 = n47183 ^ n46917;
  assign n47185 = n46920 & ~n47184;
  assign n47186 = n47185 ^ n46919;
  assign n47188 = n47187 ^ n47186;
  assign n47189 = n46079 ^ n45557;
  assign n47190 = n47189 ^ n46987;
  assign n47191 = n47190 ^ n47187;
  assign n47192 = n47188 & ~n47191;
  assign n47193 = n47192 ^ n47190;
  assign n47194 = n47193 ^ n46915;
  assign n47195 = n46916 & ~n47194;
  assign n47196 = n47195 ^ n46913;
  assign n46909 = n46859 ^ n46712;
  assign n46910 = n46909 ^ n46713;
  assign n47197 = n47196 ^ n46910;
  assign n47213 = n47199 ^ n47197;
  assign n47214 = n47213 ^ n44908;
  assign n47217 = n47183 ^ n46920;
  assign n47218 = n47217 ^ n44113;
  assign n47219 = n47180 ^ n46924;
  assign n47220 = n47219 ^ n46922;
  assign n47221 = n47220 ^ n44685;
  assign n47222 = n47177 ^ n46929;
  assign n47223 = n47222 ^ n44692;
  assign n47224 = n47174 ^ n46933;
  assign n47225 = n47224 ^ n44749;
  assign n47226 = n47171 ^ n47169;
  assign n47227 = n47226 ^ n44753;
  assign n47228 = n47165 ^ n46939;
  assign n47229 = n47228 ^ n44782;
  assign n47230 = n47162 ^ n47160;
  assign n47231 = n47230 ^ n44696;
  assign n47232 = n47156 ^ n46944;
  assign n47233 = n47232 ^ n44701;
  assign n47234 = n47153 ^ n46948;
  assign n47235 = n47234 ^ n44706;
  assign n47236 = n47150 ^ n46953;
  assign n47237 = n47236 ^ n44711;
  assign n47238 = n47147 ^ n47145;
  assign n47239 = n47238 ^ n44503;
  assign n47240 = n47141 ^ n47139;
  assign n47241 = n47240 ^ n44412;
  assign n47242 = n47135 ^ n46960;
  assign n47243 = n47242 ^ n44405;
  assign n47244 = n47132 ^ n46965;
  assign n47245 = n47244 ^ n44120;
  assign n47249 = n47117 ^ n47095;
  assign n47250 = n47249 ^ n47096;
  assign n47251 = n47250 ^ n44123;
  assign n47262 = n47261 ^ n47253;
  assign n47263 = n47254 & ~n47262;
  assign n47264 = n47263 ^ n44125;
  assign n47265 = n47264 ^ n47250;
  assign n47266 = ~n47251 & ~n47265;
  assign n47267 = n47266 ^ n44123;
  assign n47248 = n47120 ^ n47093;
  assign n47268 = n47267 ^ n47248;
  assign n47269 = n47248 ^ n44371;
  assign n47270 = ~n47268 & n47269;
  assign n47271 = n47270 ^ n44371;
  assign n47247 = n47123 ^ n46978;
  assign n47272 = n47271 ^ n47247;
  assign n47273 = n47247 ^ n44378;
  assign n47274 = n47272 & n47273;
  assign n47275 = n47274 ^ n44378;
  assign n47246 = n47126 ^ n46974;
  assign n47276 = n47275 ^ n47246;
  assign n47277 = n47246 ^ n44385;
  assign n47278 = ~n47276 & ~n47277;
  assign n47279 = n47278 ^ n44385;
  assign n47280 = n47279 ^ n44392;
  assign n47281 = n47129 ^ n46969;
  assign n47282 = n47281 ^ n47279;
  assign n47283 = ~n47280 & n47282;
  assign n47284 = n47283 ^ n44392;
  assign n47285 = n47284 ^ n47244;
  assign n47286 = n47245 & ~n47285;
  assign n47287 = n47286 ^ n44120;
  assign n47288 = n47287 ^ n47242;
  assign n47289 = n47243 & n47288;
  assign n47290 = n47289 ^ n44405;
  assign n47291 = n47290 ^ n47240;
  assign n47292 = n47241 & ~n47291;
  assign n47293 = n47292 ^ n44412;
  assign n47294 = n47293 ^ n47238;
  assign n47295 = ~n47239 & n47294;
  assign n47296 = n47295 ^ n44503;
  assign n47297 = n47296 ^ n47236;
  assign n47298 = n47237 & n47297;
  assign n47299 = n47298 ^ n44711;
  assign n47300 = n47299 ^ n47234;
  assign n47301 = ~n47235 & ~n47300;
  assign n47302 = n47301 ^ n44706;
  assign n47303 = n47302 ^ n47232;
  assign n47304 = ~n47233 & ~n47303;
  assign n47305 = n47304 ^ n44701;
  assign n47306 = n47305 ^ n47230;
  assign n47307 = ~n47231 & n47306;
  assign n47308 = n47307 ^ n44696;
  assign n47309 = n47308 ^ n47228;
  assign n47310 = n47229 & ~n47309;
  assign n47311 = n47310 ^ n44782;
  assign n47312 = n47311 ^ n47226;
  assign n47313 = ~n47227 & ~n47312;
  assign n47314 = n47313 ^ n44753;
  assign n47315 = n47314 ^ n47224;
  assign n47316 = ~n47225 & ~n47315;
  assign n47317 = n47316 ^ n44749;
  assign n47318 = n47317 ^ n47222;
  assign n47319 = ~n47223 & n47318;
  assign n47320 = n47319 ^ n44692;
  assign n47321 = n47320 ^ n47220;
  assign n47322 = n47221 & ~n47321;
  assign n47323 = n47322 ^ n44685;
  assign n47324 = n47323 ^ n47217;
  assign n47325 = ~n47218 & n47324;
  assign n47326 = n47325 ^ n44113;
  assign n47216 = n47190 ^ n47188;
  assign n47327 = n47326 ^ n47216;
  assign n47328 = n47216 ^ n44813;
  assign n47329 = ~n47327 & ~n47328;
  assign n47330 = n47329 ^ n44813;
  assign n47215 = n47193 ^ n46916;
  assign n47331 = n47330 ^ n47215;
  assign n47332 = n47215 ^ n44820;
  assign n47333 = ~n47331 & ~n47332;
  assign n47334 = n47333 ^ n44820;
  assign n47335 = n47334 ^ n47213;
  assign n47336 = n47214 & n47335;
  assign n47337 = n47336 ^ n44908;
  assign n47343 = n47337 ^ n44324;
  assign n47200 = n47199 ^ n46910;
  assign n47201 = ~n47197 & n47200;
  assign n47202 = n47201 ^ n47199;
  assign n46907 = n46862 ^ n46709;
  assign n46905 = n46904 ^ n45693;
  assign n46906 = n46905 ^ n45024;
  assign n46908 = n46907 ^ n46906;
  assign n47211 = n47202 ^ n46908;
  assign n47344 = n47343 ^ n47211;
  assign n47345 = n47334 ^ n44908;
  assign n47346 = n47345 ^ n47213;
  assign n47347 = n47331 ^ n44820;
  assign n47348 = n47320 ^ n47221;
  assign n47349 = n47314 ^ n47225;
  assign n47350 = n47302 ^ n47233;
  assign n47351 = n47299 ^ n47235;
  assign n47352 = n47296 ^ n47237;
  assign n47353 = n47290 ^ n47241;
  assign n47354 = n47276 ^ n44385;
  assign n47357 = ~n47355 & ~n47356;
  assign n47358 = n47264 ^ n44123;
  assign n47359 = n47358 ^ n47250;
  assign n47360 = ~n47357 & ~n47359;
  assign n47361 = n47268 ^ n44371;
  assign n47362 = ~n47360 & n47361;
  assign n47363 = n47272 ^ n44378;
  assign n47364 = ~n47362 & ~n47363;
  assign n47365 = n47354 & ~n47364;
  assign n47366 = n47281 ^ n44392;
  assign n47367 = n47366 ^ n47279;
  assign n47368 = n47365 & n47367;
  assign n47369 = n47284 ^ n47245;
  assign n47370 = n47368 & ~n47369;
  assign n47371 = n47287 ^ n44405;
  assign n47372 = n47371 ^ n47242;
  assign n47373 = ~n47370 & n47372;
  assign n47374 = ~n47353 & n47373;
  assign n47375 = n47293 ^ n47239;
  assign n47376 = n47374 & n47375;
  assign n47377 = ~n47352 & n47376;
  assign n47378 = ~n47351 & n47377;
  assign n47379 = ~n47350 & ~n47378;
  assign n47380 = n47305 ^ n47231;
  assign n47381 = n47379 & n47380;
  assign n47382 = n47308 ^ n47229;
  assign n47383 = ~n47381 & n47382;
  assign n47384 = n47311 ^ n47227;
  assign n47385 = ~n47383 & n47384;
  assign n47386 = n47349 & ~n47385;
  assign n47387 = n47317 ^ n44692;
  assign n47388 = n47387 ^ n47222;
  assign n47389 = n47386 & ~n47388;
  assign n47390 = n47348 & n47389;
  assign n47391 = n47323 ^ n47218;
  assign n47392 = ~n47390 & n47391;
  assign n47393 = n47327 ^ n44813;
  assign n47394 = n47392 & n47393;
  assign n47395 = n47347 & ~n47394;
  assign n47396 = n47346 & n47395;
  assign n47397 = n47344 & ~n47396;
  assign n47212 = n47211 ^ n44324;
  assign n47338 = n47337 ^ n47211;
  assign n47339 = n47212 & n47338;
  assign n47340 = n47339 ^ n44324;
  assign n47341 = n47340 ^ n44331;
  assign n47208 = n45700 ^ n45029;
  assign n47209 = n47208 ^ n47038;
  assign n47206 = n46865 ^ n46704;
  assign n47203 = n47202 ^ n46907;
  assign n47204 = ~n46908 & n47203;
  assign n47205 = n47204 ^ n46906;
  assign n47207 = n47206 ^ n47205;
  assign n47210 = n47209 ^ n47207;
  assign n47342 = n47341 ^ n47210;
  assign n47398 = n47397 ^ n47342;
  assign n2968 = n2964 ^ n2931;
  assign n2996 = n2995 ^ n2968;
  assign n3003 = n3002 ^ n2996;
  assign n47751 = n47398 ^ n3003;
  assign n47402 = n47396 ^ n47344;
  assign n47399 = n3239 ^ n2869;
  assign n47400 = n47399 ^ n42160;
  assign n47401 = n47400 ^ n2987;
  assign n47403 = n47402 ^ n47401;
  assign n47405 = n45300 ^ n2854;
  assign n47406 = n47405 ^ n42166;
  assign n47407 = n47406 ^ n36307;
  assign n47404 = n47395 ^ n47346;
  assign n47408 = n47407 ^ n47404;
  assign n47411 = n45305 ^ n37766;
  assign n47412 = n47411 ^ n42175;
  assign n47413 = n47412 ^ n36317;
  assign n47410 = n47393 ^ n47392;
  assign n47414 = n47413 ^ n47410;
  assign n47418 = n47391 ^ n47390;
  assign n47415 = n45459 ^ n37770;
  assign n47416 = n47415 ^ n42180;
  assign n47417 = n47416 ^ n3071;
  assign n47419 = n47418 ^ n47417;
  assign n47428 = n47380 ^ n47379;
  assign n47425 = n45334 ^ n37863;
  assign n47426 = n47425 ^ n42241;
  assign n47427 = n47426 ^ n1209;
  assign n47429 = n47428 ^ n47427;
  assign n47430 = n47378 ^ n47350;
  assign n1035 = n1034 ^ n995;
  assign n1069 = n1068 ^ n1035;
  assign n1079 = n1078 ^ n1069;
  assign n47431 = n47430 ^ n1079;
  assign n47435 = n47377 ^ n47351;
  assign n47432 = n45339 ^ n37853;
  assign n47433 = n47432 ^ n42231;
  assign n47434 = n47433 ^ n1060;
  assign n47436 = n47435 ^ n47434;
  assign n47439 = n45351 ^ n37808;
  assign n47440 = n47439 ^ n42214;
  assign n47441 = n47440 ^ n35835;
  assign n47438 = n47373 ^ n47353;
  assign n47442 = n47441 ^ n47438;
  assign n47446 = n47372 ^ n47370;
  assign n47443 = n45355 ^ n37833;
  assign n47444 = n47443 ^ n41119;
  assign n47445 = n47444 ^ n35839;
  assign n47447 = n47446 ^ n47445;
  assign n47451 = n47369 ^ n47368;
  assign n47448 = n45360 ^ n37814;
  assign n47449 = n47448 ^ n41676;
  assign n47450 = n47449 ^ n35844;
  assign n47452 = n47451 ^ n47450;
  assign n47456 = n47367 ^ n47365;
  assign n47453 = n45365 ^ n37818;
  assign n47454 = n47453 ^ n41681;
  assign n47455 = n47454 ^ n35849;
  assign n47457 = n47456 ^ n47455;
  assign n47459 = n45402 ^ n37236;
  assign n47460 = n47459 ^ n41687;
  assign n47461 = n47460 ^ n35854;
  assign n47458 = n47364 ^ n47354;
  assign n47462 = n47461 ^ n47458;
  assign n47464 = n45372 ^ n37207;
  assign n47465 = n47464 ^ n41692;
  assign n47466 = n47465 ^ n35860;
  assign n47463 = n47363 ^ n47362;
  assign n47467 = n47466 ^ n47463;
  assign n47472 = n47359 ^ n47357;
  assign n47469 = n45378 ^ n37216;
  assign n47470 = n47469 ^ n2299;
  assign n47471 = n47470 ^ n35869;
  assign n47473 = n47472 ^ n47471;
  assign n47486 = n47485 ^ n2289;
  assign n47488 = n47487 ^ n47485;
  assign n47489 = n47486 & n47488;
  assign n47490 = n47489 ^ n2289;
  assign n47491 = n47490 ^ n47472;
  assign n47492 = n47473 & ~n47491;
  assign n47493 = n47492 ^ n47471;
  assign n47468 = n47361 ^ n47360;
  assign n47494 = n47493 ^ n47468;
  assign n47495 = n37212 ^ n2363;
  assign n47496 = n47495 ^ n41712;
  assign n47497 = n47496 ^ n35865;
  assign n47498 = n47497 ^ n47468;
  assign n47499 = ~n47494 & n47498;
  assign n47500 = n47499 ^ n47497;
  assign n47501 = n47500 ^ n47463;
  assign n47502 = n47467 & ~n47501;
  assign n47503 = n47502 ^ n47466;
  assign n47504 = n47503 ^ n47458;
  assign n47505 = n47462 & ~n47504;
  assign n47506 = n47505 ^ n47461;
  assign n47507 = n47506 ^ n47456;
  assign n47508 = ~n47457 & n47507;
  assign n47509 = n47508 ^ n47455;
  assign n47510 = n47509 ^ n47451;
  assign n47511 = n47452 & ~n47510;
  assign n47512 = n47511 ^ n47450;
  assign n47513 = n47512 ^ n47446;
  assign n47514 = ~n47447 & n47513;
  assign n47515 = n47514 ^ n47445;
  assign n47516 = n47515 ^ n47438;
  assign n47517 = ~n47442 & n47516;
  assign n47518 = n47517 ^ n47441;
  assign n47522 = n47521 ^ n47518;
  assign n47523 = n47375 ^ n47374;
  assign n47524 = n47523 ^ n47518;
  assign n47525 = n47522 & ~n47524;
  assign n47526 = n47525 ^ n47521;
  assign n47437 = n47376 ^ n47352;
  assign n47527 = n47526 ^ n47437;
  assign n47528 = n45345 ^ n906;
  assign n47529 = n47528 ^ n42204;
  assign n47530 = n47529 ^ n3323;
  assign n47531 = n47530 ^ n47437;
  assign n47532 = n47527 & ~n47531;
  assign n47533 = n47532 ^ n47530;
  assign n47534 = n47533 ^ n47435;
  assign n47535 = ~n47436 & n47534;
  assign n47536 = n47535 ^ n47434;
  assign n47537 = n47536 ^ n47430;
  assign n47538 = ~n47431 & n47537;
  assign n47539 = n47538 ^ n1079;
  assign n47540 = n47539 ^ n47428;
  assign n47541 = ~n47429 & n47540;
  assign n47542 = n47541 ^ n47427;
  assign n47424 = n47382 ^ n47381;
  assign n47543 = n47542 ^ n47424;
  assign n47544 = n45331 ^ n37796;
  assign n47545 = n47544 ^ n1217;
  assign n47546 = n47545 ^ n36337;
  assign n47547 = n47546 ^ n47424;
  assign n47548 = n47543 & ~n47547;
  assign n47549 = n47548 ^ n47546;
  assign n47423 = n47384 ^ n47383;
  assign n47550 = n47549 ^ n47423;
  assign n47551 = n45326 ^ n37790;
  assign n47552 = n47551 ^ n42251;
  assign n47553 = n47552 ^ n1409;
  assign n47554 = n47553 ^ n47423;
  assign n47555 = ~n47550 & n47554;
  assign n47556 = n47555 ^ n47553;
  assign n47422 = n47385 ^ n47349;
  assign n47557 = n47556 ^ n47422;
  assign n47558 = n45322 ^ n37785;
  assign n47559 = n47558 ^ n42192;
  assign n47560 = n47559 ^ n36331;
  assign n47561 = n47560 ^ n47422;
  assign n47562 = n47557 & ~n47561;
  assign n47563 = n47562 ^ n47560;
  assign n47421 = n47388 ^ n47386;
  assign n47564 = n47563 ^ n47421;
  assign n47565 = n45316 ^ n37780;
  assign n47566 = n47565 ^ n42261;
  assign n47567 = n47566 ^ n36325;
  assign n47568 = n47567 ^ n47421;
  assign n47569 = n47564 & ~n47568;
  assign n47570 = n47569 ^ n47567;
  assign n47420 = n47389 ^ n47348;
  assign n47571 = n47570 ^ n47420;
  assign n47572 = n45311 ^ n37775;
  assign n47573 = n47572 ^ n42185;
  assign n47574 = n47573 ^ n2531;
  assign n47575 = n47574 ^ n47420;
  assign n47576 = ~n47571 & n47575;
  assign n47577 = n47576 ^ n47574;
  assign n47578 = n47577 ^ n47418;
  assign n47579 = n47419 & ~n47578;
  assign n47580 = n47579 ^ n47417;
  assign n47581 = n47580 ^ n47410;
  assign n47582 = ~n47414 & n47581;
  assign n47583 = n47582 ^ n47413;
  assign n47409 = n47394 ^ n47347;
  assign n47584 = n47583 ^ n47409;
  assign n47585 = n45469 ^ n3225;
  assign n47586 = n47585 ^ n42170;
  assign n47587 = n47586 ^ n36312;
  assign n47588 = n47587 ^ n47409;
  assign n47589 = n47584 & ~n47588;
  assign n47590 = n47589 ^ n47587;
  assign n47591 = n47590 ^ n47404;
  assign n47592 = n47408 & ~n47591;
  assign n47593 = n47592 ^ n47407;
  assign n47594 = n47593 ^ n47402;
  assign n47595 = n47403 & ~n47594;
  assign n47596 = n47595 ^ n47401;
  assign n47752 = n47596 ^ n47398;
  assign n47753 = ~n47751 & n47752;
  assign n47754 = n47753 ^ n3003;
  assign n47675 = n47342 & ~n47397;
  assign n47669 = n47210 ^ n44331;
  assign n47670 = n47340 ^ n47210;
  assign n47671 = n47669 & n47670;
  assign n47672 = n47671 ^ n44331;
  assign n47673 = n47672 ^ n44322;
  assign n47666 = n45691 ^ n45021;
  assign n47667 = n47666 ^ n46406;
  assign n47663 = n46868 ^ n46697;
  assign n47664 = n47663 ^ n46698;
  assign n47660 = n47209 ^ n47206;
  assign n47661 = n47207 & n47660;
  assign n47662 = n47661 ^ n47209;
  assign n47665 = n47664 ^ n47662;
  assign n47668 = n47667 ^ n47665;
  assign n47674 = n47673 ^ n47668;
  assign n47750 = n47675 ^ n47674;
  assign n47755 = n47754 ^ n47750;
  assign n47785 = n47758 ^ n47755;
  assign n47913 = n47787 ^ n47785;
  assign n48146 = n47913 ^ n45054;
  assign n48467 = n48149 ^ n48146;
  assign n49180 = n49179 ^ n48467;
  assign n48239 = n47567 ^ n47564;
  assign n48822 = n48239 ^ n46889;
  assign n48823 = n48822 ^ n47206;
  assign n47645 = n47497 ^ n47494;
  assign n47643 = n46124 ^ n45507;
  assign n47644 = n47643 ^ n46941;
  assign n47646 = n47645 ^ n47644;
  assign n47649 = n46131 ^ n45511;
  assign n47650 = n47649 ^ n46945;
  assign n47647 = n47490 ^ n47471;
  assign n47648 = n47647 ^ n47472;
  assign n47651 = n47650 ^ n47648;
  assign n47654 = n47481 ^ n47355;
  assign n47655 = n47654 ^ n47478;
  assign n47652 = n46955 ^ n45518;
  assign n47653 = n47652 ^ n46133;
  assign n47656 = n47655 ^ n47653;
  assign n47682 = n45707 ^ n45019;
  assign n47683 = n47682 ^ n46411;
  assign n47680 = n46871 ^ n46694;
  assign n47677 = n47667 ^ n47664;
  assign n47678 = ~n47665 & n47677;
  assign n47679 = n47678 ^ n47667;
  assign n47681 = n47680 ^ n47679;
  assign n47684 = n47683 ^ n47681;
  assign n47700 = n47684 ^ n44317;
  assign n47685 = n47668 ^ n44322;
  assign n47686 = n47672 ^ n47668;
  assign n47687 = ~n47685 & n47686;
  assign n47688 = n47687 ^ n44322;
  assign n47701 = n47688 ^ n47684;
  assign n47702 = ~n47700 & n47701;
  assign n47703 = n47702 ^ n44317;
  assign n47696 = n47683 ^ n47680;
  assign n47697 = n47681 & n47696;
  assign n47698 = n47697 ^ n47683;
  assign n47694 = n46874 ^ n46689;
  assign n47692 = n45685 ^ n45016;
  assign n47693 = n47692 ^ n46403;
  assign n47695 = n47694 ^ n47693;
  assign n47699 = n47698 ^ n47695;
  assign n47704 = n47703 ^ n47699;
  assign n47717 = n47699 ^ n44314;
  assign n47718 = ~n47704 & ~n47717;
  assign n47719 = n47718 ^ n44314;
  assign n47712 = n46877 ^ n3137;
  assign n47713 = n47712 ^ n46686;
  assign n47709 = n47698 ^ n47694;
  assign n47710 = n47695 & n47709;
  assign n47711 = n47710 ^ n47693;
  assign n47714 = n47713 ^ n47711;
  assign n47707 = n45552 ^ n44741;
  assign n47708 = n47707 ^ n46401;
  assign n47715 = n47714 ^ n47708;
  assign n47716 = n47715 ^ n44138;
  assign n47720 = n47719 ^ n47716;
  assign n47676 = ~n47674 & ~n47675;
  assign n47689 = n47688 ^ n44317;
  assign n47690 = n47689 ^ n47684;
  assign n47691 = ~n47676 & n47690;
  assign n47705 = n47704 ^ n44314;
  assign n47706 = n47691 & n47705;
  assign n47742 = n47720 ^ n47706;
  assign n47739 = n45650 ^ n37739;
  assign n47740 = n47739 ^ n42150;
  assign n47741 = n47740 ^ n36285;
  assign n47743 = n47742 ^ n47741;
  assign n47748 = n47690 ^ n47676;
  assign n47745 = n45660 ^ n37749;
  assign n47746 = n47745 ^ n42293;
  assign n47747 = n47746 ^ n1697;
  assign n47749 = n47748 ^ n47747;
  assign n47759 = n47758 ^ n47750;
  assign n47760 = n47755 & ~n47759;
  assign n47761 = n47760 ^ n47758;
  assign n47762 = n47761 ^ n47748;
  assign n47763 = ~n47749 & n47762;
  assign n47764 = n47763 ^ n47747;
  assign n47744 = n47705 ^ n47691;
  assign n47765 = n47764 ^ n47744;
  assign n47766 = n45655 ^ n37744;
  assign n47767 = n47766 ^ n42300;
  assign n47768 = n47767 ^ n36290;
  assign n47769 = n47768 ^ n47744;
  assign n47770 = ~n47765 & n47769;
  assign n47771 = n47770 ^ n47768;
  assign n47772 = n47771 ^ n47742;
  assign n47773 = n47743 & ~n47772;
  assign n47774 = n47773 ^ n47741;
  assign n47730 = n47719 ^ n47715;
  assign n47731 = ~n47716 & n47730;
  assign n47732 = n47731 ^ n44138;
  assign n47724 = n47713 ^ n47708;
  assign n47725 = n47714 & ~n47724;
  assign n47726 = n47725 ^ n47708;
  assign n47722 = n46395 ^ n44739;
  assign n47723 = n47722 ^ n45548;
  assign n47727 = n47726 ^ n47723;
  assign n46884 = n46883 ^ n46880;
  assign n46902 = n46901 ^ n46884;
  assign n47728 = n47727 ^ n46902;
  assign n47729 = n47728 ^ n44134;
  assign n47733 = n47732 ^ n47729;
  assign n47721 = ~n47706 & n47720;
  assign n47734 = n47733 ^ n47721;
  assign n47738 = n47737 ^ n47734;
  assign n47775 = n47774 ^ n47738;
  assign n47658 = n46957 ^ n45528;
  assign n47659 = n47658 ^ n46142;
  assign n47776 = n47775 ^ n47659;
  assign n47779 = n47771 ^ n47743;
  assign n47777 = n46147 ^ n45532;
  assign n47778 = n47777 ^ n46962;
  assign n47780 = n47779 ^ n47778;
  assign n47782 = n46968 ^ n45536;
  assign n47783 = n47782 ^ n46151;
  assign n47781 = n47768 ^ n47765;
  assign n47784 = n47783 ^ n47781;
  assign n47789 = n46152 ^ n45540;
  assign n47790 = n47789 ^ n46973;
  assign n47788 = ~n47785 & n47787;
  assign n47791 = n47790 ^ n47788;
  assign n47792 = n47761 ^ n47747;
  assign n47793 = n47792 ^ n47748;
  assign n47794 = n47793 ^ n47790;
  assign n47795 = ~n47791 & ~n47794;
  assign n47796 = n47795 ^ n47788;
  assign n47797 = n47796 ^ n47783;
  assign n47798 = n47784 & ~n47797;
  assign n47799 = n47798 ^ n47781;
  assign n47800 = n47799 ^ n47779;
  assign n47801 = n47780 & ~n47800;
  assign n47802 = n47801 ^ n47778;
  assign n47803 = n47802 ^ n47775;
  assign n47804 = ~n47776 & n47803;
  assign n47805 = n47804 ^ n47659;
  assign n47657 = n47477 ^ n47476;
  assign n47806 = n47805 ^ n47657;
  assign n47807 = n46137 ^ n45522;
  assign n47808 = n47807 ^ n46956;
  assign n47809 = n47808 ^ n47657;
  assign n47810 = ~n47806 & ~n47809;
  assign n47811 = n47810 ^ n47808;
  assign n47812 = n47811 ^ n47655;
  assign n47813 = ~n47656 & ~n47812;
  assign n47814 = n47813 ^ n47653;
  assign n47817 = n47816 ^ n47814;
  assign n47818 = n46950 ^ n46132;
  assign n47819 = n47818 ^ n45514;
  assign n47820 = n47819 ^ n47816;
  assign n47821 = n47817 & ~n47820;
  assign n47822 = n47821 ^ n47819;
  assign n47823 = n47822 ^ n47648;
  assign n47824 = n47651 & ~n47823;
  assign n47825 = n47824 ^ n47650;
  assign n47826 = n47825 ^ n47644;
  assign n47827 = n47646 & ~n47826;
  assign n47828 = n47827 ^ n47645;
  assign n47640 = n47500 ^ n47466;
  assign n47641 = n47640 ^ n47463;
  assign n47638 = n46118 ^ n45501;
  assign n47639 = n47638 ^ n46940;
  assign n47642 = n47641 ^ n47639;
  assign n47902 = n47828 ^ n47642;
  assign n47903 = n47902 ^ n44698;
  assign n47905 = n47822 ^ n47651;
  assign n47906 = n47905 ^ n44708;
  assign n47911 = n47799 ^ n47780;
  assign n47912 = n47911 ^ n44727;
  assign n47914 = ~n45054 & ~n47913;
  assign n47915 = n47914 ^ n44734;
  assign n47916 = n47793 ^ n47791;
  assign n47917 = n47916 ^ n47914;
  assign n47918 = n47915 & ~n47917;
  assign n47919 = n47918 ^ n44734;
  assign n47920 = n47919 ^ n44728;
  assign n47921 = n47796 ^ n47784;
  assign n47922 = n47921 ^ n47919;
  assign n47923 = n47920 & ~n47922;
  assign n47924 = n47923 ^ n44728;
  assign n47925 = n47924 ^ n47911;
  assign n47926 = ~n47912 & ~n47925;
  assign n47927 = n47926 ^ n44727;
  assign n47910 = n47802 ^ n47776;
  assign n47928 = n47927 ^ n47910;
  assign n47929 = n47910 ^ n44725;
  assign n47930 = ~n47928 & n47929;
  assign n47931 = n47930 ^ n44725;
  assign n47909 = n47808 ^ n47806;
  assign n47932 = n47931 ^ n47909;
  assign n47933 = n47909 ^ n44721;
  assign n47934 = ~n47932 & n47933;
  assign n47935 = n47934 ^ n44721;
  assign n47908 = n47811 ^ n47656;
  assign n47936 = n47935 ^ n47908;
  assign n47937 = n47908 ^ n44717;
  assign n47938 = n47936 & n47937;
  assign n47939 = n47938 ^ n44717;
  assign n47907 = n47819 ^ n47817;
  assign n47940 = n47939 ^ n47907;
  assign n47941 = n47907 ^ n44713;
  assign n47942 = n47940 & ~n47941;
  assign n47943 = n47942 ^ n44713;
  assign n47944 = n47943 ^ n47905;
  assign n47945 = n47906 & ~n47944;
  assign n47946 = n47945 ^ n44708;
  assign n47904 = n47825 ^ n47646;
  assign n47947 = n47946 ^ n47904;
  assign n47948 = n47904 ^ n44703;
  assign n47949 = ~n47947 & n47948;
  assign n47950 = n47949 ^ n44703;
  assign n47951 = n47950 ^ n47902;
  assign n47952 = ~n47903 & n47951;
  assign n47953 = n47952 ^ n44698;
  assign n47835 = n46936 ^ n46112;
  assign n47836 = n47835 ^ n45760;
  assign n47832 = n47503 ^ n47461;
  assign n47833 = n47832 ^ n47458;
  assign n47829 = n47828 ^ n47641;
  assign n47830 = ~n47642 & ~n47829;
  assign n47831 = n47830 ^ n47639;
  assign n47834 = n47833 ^ n47831;
  assign n47900 = n47836 ^ n47834;
  assign n47901 = n47900 ^ n45094;
  assign n48010 = n47953 ^ n47901;
  assign n48011 = n47947 ^ n44703;
  assign n48012 = n47940 ^ n44713;
  assign n48013 = n47932 ^ n44721;
  assign n48014 = n47928 ^ n44725;
  assign n48015 = n47924 ^ n44727;
  assign n48016 = n48015 ^ n47911;
  assign n48017 = n47916 ^ n47915;
  assign n48018 = n47921 ^ n47920;
  assign n48019 = ~n48017 & ~n48018;
  assign n48020 = ~n48016 & ~n48019;
  assign n48021 = n48014 & ~n48020;
  assign n48022 = ~n48013 & ~n48021;
  assign n48023 = n47936 ^ n44717;
  assign n48024 = ~n48022 & n48023;
  assign n48025 = n48012 & n48024;
  assign n48026 = n47943 ^ n47906;
  assign n48027 = n48025 & ~n48026;
  assign n48028 = n48011 & ~n48027;
  assign n48029 = n47950 ^ n47903;
  assign n48030 = n48028 & ~n48029;
  assign n48031 = n48010 & n48030;
  assign n47954 = n47953 ^ n47900;
  assign n47955 = n47901 & n47954;
  assign n47956 = n47955 ^ n45094;
  assign n47837 = n47836 ^ n47833;
  assign n47838 = n47834 & n47837;
  assign n47839 = n47838 ^ n47836;
  assign n47635 = n46109 ^ n45900;
  assign n47636 = n47635 ^ n46935;
  assign n47634 = n47506 ^ n47457;
  assign n47637 = n47636 ^ n47634;
  assign n47899 = n47839 ^ n47637;
  assign n47957 = n47956 ^ n47899;
  assign n48032 = n47957 ^ n45101;
  assign n48033 = n48031 & n48032;
  assign n47958 = n47899 ^ n45101;
  assign n47959 = ~n47957 & ~n47958;
  assign n47960 = n47959 ^ n45101;
  assign n47840 = n47839 ^ n47636;
  assign n47841 = ~n47637 & ~n47840;
  assign n47842 = n47841 ^ n47634;
  assign n47632 = n47509 ^ n47452;
  assign n47630 = n46930 ^ n45918;
  assign n47631 = n47630 ^ n46101;
  assign n47633 = n47632 ^ n47631;
  assign n47897 = n47842 ^ n47633;
  assign n47898 = n47897 ^ n45108;
  assign n48009 = n47960 ^ n47898;
  assign n48088 = n48033 ^ n48009;
  assign n48092 = n48091 ^ n48088;
  assign n48096 = n48032 ^ n48031;
  assign n48093 = n45954 ^ n38079;
  assign n48094 = n48093 ^ n42490;
  assign n48095 = n48094 ^ n36999;
  assign n48097 = n48096 ^ n48095;
  assign n48101 = n48030 ^ n48010;
  assign n48098 = n45959 ^ n38084;
  assign n48099 = n48098 ^ n42495;
  assign n48100 = n48099 ^ n36616;
  assign n48102 = n48101 ^ n48100;
  assign n48106 = n48029 ^ n48028;
  assign n48103 = n45965 ^ n38088;
  assign n48104 = n48103 ^ n42570;
  assign n48105 = n48104 ^ n740;
  assign n48107 = n48106 ^ n48105;
  assign n48111 = n48027 ^ n48011;
  assign n48108 = n45970 ^ n38149;
  assign n48109 = n48108 ^ n42502;
  assign n48110 = n48109 ^ n36607;
  assign n48112 = n48111 ^ n48110;
  assign n48114 = n45975 ^ n38094;
  assign n48115 = n48114 ^ n42560;
  assign n48116 = n48115 ^ n36547;
  assign n48113 = n48026 ^ n48025;
  assign n48117 = n48116 ^ n48113;
  assign n48121 = n48024 ^ n48012;
  assign n48118 = n45979 ^ n38099;
  assign n48119 = n48118 ^ n42508;
  assign n48120 = n48119 ^ n36552;
  assign n48122 = n48121 ^ n48120;
  assign n48126 = n48023 ^ n48022;
  assign n48123 = n45985 ^ n38105;
  assign n48124 = n48123 ^ n42550;
  assign n48125 = n48124 ^ n36557;
  assign n48127 = n48126 ^ n48125;
  assign n48131 = n48021 ^ n48013;
  assign n48128 = n46019 ^ n38109;
  assign n48129 = n48128 ^ n42513;
  assign n48130 = n48129 ^ n36561;
  assign n48132 = n48131 ^ n48130;
  assign n48136 = n48020 ^ n48014;
  assign n48133 = n46012 ^ n38130;
  assign n48134 = n48133 ^ n42518;
  assign n48135 = n48134 ^ n36588;
  assign n48137 = n48136 ^ n48135;
  assign n48141 = n48019 ^ n48016;
  assign n48138 = n45991 ^ n2396;
  assign n48139 = n48138 ^ n42523;
  assign n48140 = n48139 ^ n36567;
  assign n48142 = n48141 ^ n48140;
  assign n48151 = n46000 ^ n38116;
  assign n48152 = n48151 ^ n42529;
  assign n48153 = n48152 ^ n36574;
  assign n48150 = n48146 & n48149;
  assign n48154 = n48153 ^ n48150;
  assign n48155 = n48150 ^ n48017;
  assign n48156 = n48154 & n48155;
  assign n48157 = n48156 ^ n48153;
  assign n48143 = n45996 ^ n2381;
  assign n48144 = n48143 ^ n42533;
  assign n48145 = n48144 ^ n36571;
  assign n48158 = n48157 ^ n48145;
  assign n48159 = n48018 ^ n48017;
  assign n48160 = n48159 ^ n48157;
  assign n48161 = n48158 & n48160;
  assign n48162 = n48161 ^ n48145;
  assign n48163 = n48162 ^ n48141;
  assign n48164 = n48142 & ~n48163;
  assign n48165 = n48164 ^ n48140;
  assign n48166 = n48165 ^ n48136;
  assign n48167 = n48137 & ~n48166;
  assign n48168 = n48167 ^ n48135;
  assign n48169 = n48168 ^ n48131;
  assign n48170 = n48132 & ~n48169;
  assign n48171 = n48170 ^ n48130;
  assign n48172 = n48171 ^ n48126;
  assign n48173 = n48127 & ~n48172;
  assign n48174 = n48173 ^ n48125;
  assign n48175 = n48174 ^ n48121;
  assign n48176 = ~n48122 & n48175;
  assign n48177 = n48176 ^ n48120;
  assign n48178 = n48177 ^ n48113;
  assign n48179 = n48117 & ~n48178;
  assign n48180 = n48179 ^ n48116;
  assign n48181 = n48180 ^ n48111;
  assign n48182 = ~n48112 & n48181;
  assign n48183 = n48182 ^ n48110;
  assign n48184 = n48183 ^ n48106;
  assign n48185 = ~n48107 & n48184;
  assign n48186 = n48185 ^ n48105;
  assign n48187 = n48186 ^ n48101;
  assign n48188 = n48102 & ~n48187;
  assign n48189 = n48188 ^ n48100;
  assign n48190 = n48189 ^ n48096;
  assign n48191 = n48097 & ~n48190;
  assign n48192 = n48191 ^ n48095;
  assign n48193 = n48192 ^ n48088;
  assign n48194 = n48092 & ~n48193;
  assign n48195 = n48194 ^ n48091;
  assign n48034 = n48009 & n48033;
  assign n47961 = n47960 ^ n47897;
  assign n47962 = n47898 & n47961;
  assign n47963 = n47962 ^ n45108;
  assign n47843 = n47842 ^ n47632;
  assign n47844 = n47633 & n47843;
  assign n47845 = n47844 ^ n47631;
  assign n47627 = n46926 ^ n46099;
  assign n47628 = n47627 ^ n46126;
  assign n47894 = n47845 ^ n47628;
  assign n47625 = n47512 ^ n47445;
  assign n47626 = n47625 ^ n47446;
  assign n47895 = n47894 ^ n47626;
  assign n47896 = n47895 ^ n44690;
  assign n48008 = n47963 ^ n47896;
  assign n48086 = n48034 ^ n48008;
  assign n48083 = n45944 ^ n1150;
  assign n48084 = n48083 ^ n42481;
  assign n48085 = n48084 ^ n3348;
  assign n48087 = n48086 ^ n48085;
  assign n48821 = n48195 ^ n48087;
  assign n48824 = n48823 ^ n48821;
  assign n48664 = n48192 ^ n48092;
  assign n47999 = n47560 ^ n47557;
  assign n48661 = n47999 ^ n46077;
  assign n48662 = n48661 ^ n46907;
  assign n48817 = n48664 ^ n48662;
  assign n47603 = n47546 ^ n47543;
  assign n48602 = n47603 ^ n46915;
  assign n48603 = n48602 ^ n46088;
  assign n48601 = n48186 ^ n48102;
  assign n48604 = n48603 ^ n48601;
  assign n48518 = n48183 ^ n48107;
  assign n47607 = n47539 ^ n47429;
  assign n48515 = n47607 ^ n46093;
  assign n48516 = n48515 ^ n47187;
  assign n48597 = n48518 ^ n48516;
  assign n48258 = n48177 ^ n48117;
  assign n48256 = n46922 ^ n46101;
  assign n47609 = n47533 ^ n47436;
  assign n48257 = n48256 ^ n47609;
  assign n48259 = n48258 ^ n48257;
  assign n48262 = n48174 ^ n48122;
  assign n47613 = n47530 ^ n47527;
  assign n48260 = n47613 ^ n46926;
  assign n48261 = n48260 ^ n46109;
  assign n48263 = n48262 ^ n48261;
  assign n48496 = n48171 ^ n48127;
  assign n47621 = n47515 ^ n47442;
  assign n48265 = n47621 ^ n46935;
  assign n48266 = n48265 ^ n46118;
  assign n48264 = n48168 ^ n48132;
  assign n48267 = n48266 ^ n48264;
  assign n48486 = n48165 ^ n48137;
  assign n48271 = n46941 ^ n46132;
  assign n48272 = n48271 ^ n47634;
  assign n48270 = n48159 ^ n48158;
  assign n48273 = n48272 ^ n48270;
  assign n48276 = n47833 ^ n46133;
  assign n48277 = n48276 ^ n46945;
  assign n48274 = n48153 ^ n48017;
  assign n48275 = n48274 ^ n48150;
  assign n48278 = n48277 ^ n48275;
  assign n48436 = n47645 ^ n46142;
  assign n48437 = n48436 ^ n46955;
  assign n48385 = n46315 ^ n38497;
  assign n48386 = n48385 ^ n42868;
  assign n48387 = n48386 ^ n1860;
  assign n48293 = n47577 ^ n47419;
  assign n48291 = n46411 ^ n45700;
  assign n48292 = n48291 ^ n46902;
  assign n48294 = n48293 ^ n48292;
  assign n48297 = n47574 ^ n47571;
  assign n48295 = n47713 ^ n45693;
  assign n48296 = n48295 ^ n46406;
  assign n48298 = n48297 ^ n48296;
  assign n48237 = n47694 ^ n47038;
  assign n48238 = n48237 ^ n46297;
  assign n48240 = n48239 ^ n48238;
  assign n47996 = n47680 ^ n46904;
  assign n47997 = n47996 ^ n45495;
  assign n48233 = n47999 ^ n47997;
  assign n47877 = n47664 ^ n46079;
  assign n47878 = n47877 ^ n47014;
  assign n47876 = n47553 ^ n47550;
  assign n47879 = n47878 ^ n47876;
  assign n47604 = n46911 ^ n46085;
  assign n47605 = n47604 ^ n47206;
  assign n47606 = n47605 ^ n47603;
  assign n47610 = n46102 ^ n46077;
  assign n47611 = n47610 ^ n46915;
  assign n47612 = n47611 ^ n47609;
  assign n47614 = n47187 ^ n46082;
  assign n47615 = n47614 ^ n46106;
  assign n47616 = n47615 ^ n47613;
  assign n47618 = n46917 ^ n46114;
  assign n47619 = n47618 ^ n46088;
  assign n47617 = n47523 ^ n47522;
  assign n47620 = n47619 ^ n47617;
  assign n47622 = n46922 ^ n46119;
  assign n47623 = n47622 ^ n46093;
  assign n47624 = n47623 ^ n47621;
  assign n47629 = n47628 ^ n47626;
  assign n47846 = n47845 ^ n47626;
  assign n47847 = n47629 & n47846;
  assign n47848 = n47847 ^ n47628;
  assign n47849 = n47848 ^ n47621;
  assign n47850 = n47624 & ~n47849;
  assign n47851 = n47850 ^ n47623;
  assign n47852 = n47851 ^ n47617;
  assign n47853 = ~n47620 & n47852;
  assign n47854 = n47853 ^ n47619;
  assign n47855 = n47854 ^ n47613;
  assign n47856 = ~n47616 & ~n47855;
  assign n47857 = n47856 ^ n47615;
  assign n47858 = n47857 ^ n47609;
  assign n47859 = ~n47612 & n47858;
  assign n47860 = n47859 ^ n47611;
  assign n47608 = n47536 ^ n47431;
  assign n47861 = n47860 ^ n47608;
  assign n47862 = n46889 ^ n46096;
  assign n47863 = n47862 ^ n46910;
  assign n47864 = n47863 ^ n47608;
  assign n47865 = n47861 & n47864;
  assign n47866 = n47865 ^ n47863;
  assign n47867 = n47866 ^ n47607;
  assign n47868 = n46987 ^ n46907;
  assign n47869 = n47868 ^ n46090;
  assign n47870 = n47869 ^ n47607;
  assign n47871 = ~n47867 & ~n47870;
  assign n47872 = n47871 ^ n47869;
  assign n47873 = n47872 ^ n47603;
  assign n47874 = n47606 & n47873;
  assign n47875 = n47874 ^ n47605;
  assign n47993 = n47876 ^ n47875;
  assign n47994 = n47879 & n47993;
  assign n47995 = n47994 ^ n47878;
  assign n48234 = n47999 ^ n47995;
  assign n48235 = n48233 & n48234;
  assign n48236 = n48235 ^ n47997;
  assign n48299 = n48239 ^ n48236;
  assign n48300 = ~n48240 & ~n48299;
  assign n48301 = n48300 ^ n48238;
  assign n48302 = n48301 ^ n48297;
  assign n48303 = n48298 & ~n48302;
  assign n48304 = n48303 ^ n48296;
  assign n48305 = n48304 ^ n48293;
  assign n48306 = n48294 & ~n48305;
  assign n48307 = n48306 ^ n48292;
  assign n48288 = n47580 ^ n47413;
  assign n48289 = n48288 ^ n47410;
  assign n48286 = n47104 ^ n45691;
  assign n48287 = n48286 ^ n46403;
  assign n48290 = n48289 ^ n48287;
  assign n48333 = n48307 ^ n48290;
  assign n48334 = n48333 ^ n45021;
  assign n48335 = n48304 ^ n48294;
  assign n48336 = n48335 ^ n45029;
  assign n48337 = n48301 ^ n48296;
  assign n48338 = n48337 ^ n48297;
  assign n48339 = n48338 ^ n45024;
  assign n47998 = n47997 ^ n47995;
  assign n48000 = n47999 ^ n47998;
  assign n48001 = n48000 ^ n45553;
  assign n47880 = n47879 ^ n47875;
  assign n47881 = n47880 ^ n45557;
  assign n47882 = n47872 ^ n47606;
  assign n47883 = n47882 ^ n45561;
  assign n47884 = n47869 ^ n47867;
  assign n47885 = n47884 ^ n45565;
  assign n47887 = n47857 ^ n47612;
  assign n47888 = n47887 ^ n45482;
  assign n47889 = n47854 ^ n47616;
  assign n47890 = n47889 ^ n45124;
  assign n47891 = n47851 ^ n47620;
  assign n47892 = n47891 ^ n44682;
  assign n47964 = n47963 ^ n47895;
  assign n47965 = ~n47896 & n47964;
  assign n47966 = n47965 ^ n44690;
  assign n47893 = n47848 ^ n47624;
  assign n47967 = n47966 ^ n47893;
  assign n47968 = n47893 ^ n44684;
  assign n47969 = ~n47967 & ~n47968;
  assign n47970 = n47969 ^ n44684;
  assign n47971 = n47970 ^ n47891;
  assign n47972 = n47892 & ~n47971;
  assign n47973 = n47972 ^ n44682;
  assign n47974 = n47973 ^ n47889;
  assign n47975 = ~n47890 & ~n47974;
  assign n47976 = n47975 ^ n45124;
  assign n47977 = n47976 ^ n47887;
  assign n47978 = ~n47888 & ~n47977;
  assign n47979 = n47978 ^ n45482;
  assign n47886 = n47863 ^ n47861;
  assign n47980 = n47979 ^ n47886;
  assign n47981 = n47886 ^ n45569;
  assign n47982 = ~n47980 & ~n47981;
  assign n47983 = n47982 ^ n45569;
  assign n47984 = n47983 ^ n47884;
  assign n47985 = ~n47885 & n47984;
  assign n47986 = n47985 ^ n45565;
  assign n47987 = n47986 ^ n47882;
  assign n47988 = n47883 & n47987;
  assign n47989 = n47988 ^ n45561;
  assign n47990 = n47989 ^ n47880;
  assign n47991 = n47881 & n47990;
  assign n47992 = n47991 ^ n45557;
  assign n48242 = n48000 ^ n47992;
  assign n48243 = ~n48001 & n48242;
  assign n48244 = n48243 ^ n45553;
  assign n48241 = n48240 ^ n48236;
  assign n48245 = n48244 ^ n48241;
  assign n48340 = n48241 ^ n45592;
  assign n48341 = n48245 & n48340;
  assign n48342 = n48341 ^ n45592;
  assign n48343 = n48342 ^ n48338;
  assign n48344 = ~n48339 & ~n48343;
  assign n48345 = n48344 ^ n45024;
  assign n48346 = n48345 ^ n48335;
  assign n48347 = ~n48336 & n48346;
  assign n48348 = n48347 ^ n45029;
  assign n48349 = n48348 ^ n48333;
  assign n48350 = ~n48334 & ~n48349;
  assign n48351 = n48350 ^ n45021;
  assign n48313 = n46401 ^ n45707;
  assign n48314 = n48313 ^ n47111;
  assign n48311 = n47587 ^ n47584;
  assign n48308 = n48307 ^ n48289;
  assign n48309 = ~n48290 & n48308;
  assign n48310 = n48309 ^ n48287;
  assign n48312 = n48311 ^ n48310;
  assign n48332 = n48314 ^ n48312;
  assign n48352 = n48351 ^ n48332;
  assign n48353 = n48332 ^ n45019;
  assign n48354 = ~n48352 & ~n48353;
  assign n48355 = n48354 ^ n45019;
  assign n48320 = n47101 ^ n45685;
  assign n48321 = n48320 ^ n46395;
  assign n48318 = n47590 ^ n47408;
  assign n48315 = n48314 ^ n48311;
  assign n48316 = n48312 & n48315;
  assign n48317 = n48316 ^ n48314;
  assign n48319 = n48318 ^ n48317;
  assign n48330 = n48321 ^ n48319;
  assign n48331 = n48330 ^ n45016;
  assign n48367 = n48355 ^ n48331;
  assign n48246 = n48245 ^ n45592;
  assign n48002 = n48001 ^ n47992;
  assign n48003 = n47983 ^ n47885;
  assign n48004 = n47980 ^ n45569;
  assign n48005 = n47976 ^ n45482;
  assign n48006 = n48005 ^ n47887;
  assign n48007 = n47973 ^ n47890;
  assign n48035 = ~n48008 & ~n48034;
  assign n48036 = n47967 ^ n44684;
  assign n48037 = n48035 & ~n48036;
  assign n48038 = n47970 ^ n47892;
  assign n48039 = ~n48037 & n48038;
  assign n48040 = n48007 & ~n48039;
  assign n48041 = n48006 & ~n48040;
  assign n48042 = ~n48004 & n48041;
  assign n48043 = n48003 & n48042;
  assign n48044 = n47986 ^ n47883;
  assign n48045 = ~n48043 & n48044;
  assign n48046 = n47989 ^ n47881;
  assign n48047 = n48045 & ~n48046;
  assign n48247 = n48002 & ~n48047;
  assign n48368 = ~n48246 & n48247;
  assign n48369 = n48342 ^ n48339;
  assign n48370 = ~n48368 & n48369;
  assign n48371 = n48345 ^ n48336;
  assign n48372 = ~n48370 & n48371;
  assign n48373 = n48348 ^ n48334;
  assign n48374 = ~n48372 & ~n48373;
  assign n48375 = n48352 ^ n45019;
  assign n48376 = ~n48374 & ~n48375;
  assign n48377 = n48367 & n48376;
  assign n48322 = n48321 ^ n48318;
  assign n48323 = n48319 & ~n48322;
  assign n48324 = n48323 ^ n48321;
  assign n48284 = n47593 ^ n47403;
  assign n48282 = n46158 ^ n45552;
  assign n48283 = n48282 ^ n47096;
  assign n48285 = n48284 ^ n48283;
  assign n48360 = n48324 ^ n48285;
  assign n48365 = n48360 ^ n44741;
  assign n48356 = n48355 ^ n48330;
  assign n48357 = ~n48331 & n48356;
  assign n48358 = n48357 ^ n45016;
  assign n48366 = n48365 ^ n48358;
  assign n48384 = n48377 ^ n48366;
  assign n48388 = n48387 ^ n48384;
  assign n48393 = n48375 ^ n48374;
  assign n48390 = n46325 ^ n38504;
  assign n48391 = n48390 ^ n42962;
  assign n48392 = n48391 ^ n36952;
  assign n48394 = n48393 ^ n48392;
  assign n48396 = n46330 ^ n38509;
  assign n48397 = n48396 ^ n42880;
  assign n48398 = n48397 ^ n36957;
  assign n48395 = n48373 ^ n48372;
  assign n48399 = n48398 ^ n48395;
  assign n48400 = n48371 ^ n48370;
  assign n48404 = n48403 ^ n48400;
  assign n48408 = n48369 ^ n48368;
  assign n48405 = n46340 ^ n38515;
  assign n48406 = n48405 ^ n42949;
  assign n48407 = n48406 ^ n3131;
  assign n48409 = n48408 ^ n48407;
  assign n48248 = n48247 ^ n48246;
  assign n48230 = n46345 ^ n38520;
  assign n48231 = n48230 ^ n3107;
  assign n48232 = n48231 ^ n2762;
  assign n48249 = n48248 ^ n48232;
  assign n48048 = n48047 ^ n48002;
  assign n47600 = n46351 ^ n38525;
  assign n47601 = n47600 ^ n2681;
  assign n47602 = n47601 ^ n3105;
  assign n48049 = n48048 ^ n47602;
  assign n48051 = n46355 ^ n3083;
  assign n48052 = n48051 ^ n42894;
  assign n48053 = n48052 ^ n2673;
  assign n48050 = n48046 ^ n48045;
  assign n48054 = n48053 ^ n48050;
  assign n48056 = n45500 ^ n2573;
  assign n48057 = n48056 ^ n42899;
  assign n48058 = n48057 ^ n3191;
  assign n48055 = n48044 ^ n48043;
  assign n48059 = n48058 ^ n48055;
  assign n48061 = n45929 ^ n38533;
  assign n48062 = n48061 ^ n42904;
  assign n48063 = n48062 ^ n36977;
  assign n48060 = n48042 ^ n48003;
  assign n48064 = n48063 ^ n48060;
  assign n48068 = n48041 ^ n48004;
  assign n48065 = n46069 ^ n38574;
  assign n48066 = n48065 ^ n42908;
  assign n48067 = n48066 ^ n36982;
  assign n48069 = n48068 ^ n48067;
  assign n48074 = n48039 ^ n48007;
  assign n48071 = n46059 ^ n38564;
  assign n48072 = n48071 ^ n1372;
  assign n48073 = n48072 ^ n37027;
  assign n48075 = n48074 ^ n48073;
  assign n48076 = n48038 ^ n48037;
  assign n1327 = n1317 ^ n1254;
  assign n1355 = n1354 ^ n1327;
  assign n1362 = n1361 ^ n1355;
  assign n48077 = n48076 ^ n1362;
  assign n48081 = n48036 ^ n48035;
  assign n48078 = n45940 ^ n1168;
  assign n48079 = n48078 ^ n3350;
  assign n48080 = n48079 ^ n1346;
  assign n48082 = n48081 ^ n48080;
  assign n48196 = n48195 ^ n48086;
  assign n48197 = ~n48087 & n48196;
  assign n48198 = n48197 ^ n48085;
  assign n48199 = n48198 ^ n48081;
  assign n48200 = n48082 & ~n48199;
  assign n48201 = n48200 ^ n48080;
  assign n48202 = n48201 ^ n48076;
  assign n48203 = ~n48077 & n48202;
  assign n48204 = n48203 ^ n1362;
  assign n48205 = n48204 ^ n48074;
  assign n48206 = n48075 & ~n48205;
  assign n48207 = n48206 ^ n48073;
  assign n48070 = n48040 ^ n48006;
  assign n48208 = n48207 ^ n48070;
  assign n48209 = n38540 ^ n1439;
  assign n48210 = n48209 ^ n42913;
  assign n48211 = n48210 ^ n36986;
  assign n48212 = n48211 ^ n48070;
  assign n48213 = n48208 & ~n48212;
  assign n48214 = n48213 ^ n48211;
  assign n48215 = n48214 ^ n48067;
  assign n48216 = ~n48069 & ~n48215;
  assign n48217 = n48216 ^ n48068;
  assign n48218 = n48217 ^ n48060;
  assign n48219 = n48064 & n48218;
  assign n48220 = n48219 ^ n48063;
  assign n48221 = n48220 ^ n48055;
  assign n48222 = n48059 & ~n48221;
  assign n48223 = n48222 ^ n48058;
  assign n48224 = n48223 ^ n48053;
  assign n48225 = n48054 & ~n48224;
  assign n48226 = n48225 ^ n48050;
  assign n48227 = n48226 ^ n48048;
  assign n48228 = ~n48049 & n48227;
  assign n48229 = n48228 ^ n47602;
  assign n48410 = n48248 ^ n48229;
  assign n48411 = ~n48249 & n48410;
  assign n48412 = n48411 ^ n48232;
  assign n48413 = n48412 ^ n48408;
  assign n48414 = n48409 & ~n48413;
  assign n48415 = n48414 ^ n48407;
  assign n48416 = n48415 ^ n48400;
  assign n48417 = ~n48404 & n48416;
  assign n48418 = n48417 ^ n48403;
  assign n48419 = n48418 ^ n48398;
  assign n48420 = ~n48399 & ~n48419;
  assign n48421 = n48420 ^ n48395;
  assign n48422 = n48421 ^ n48392;
  assign n48423 = n48394 & n48422;
  assign n48424 = n48423 ^ n48393;
  assign n48389 = n48376 ^ n48367;
  assign n48425 = n48424 ^ n48389;
  assign n48426 = n46321 ^ n1745;
  assign n48427 = n48426 ^ n42874;
  assign n48428 = n48427 ^ n37067;
  assign n48429 = n48428 ^ n48389;
  assign n48430 = ~n48425 & n48429;
  assign n48431 = n48430 ^ n48428;
  assign n48432 = n48431 ^ n48387;
  assign n48433 = ~n48388 & ~n48432;
  assign n48434 = n48433 ^ n48384;
  assign n48379 = n46391 ^ n38492;
  assign n48380 = n48379 ^ n1868;
  assign n48381 = n48380 ^ n37126;
  assign n48378 = ~n48366 & ~n48377;
  assign n48382 = n48381 ^ n48378;
  assign n48359 = n48358 ^ n44741;
  assign n48361 = n48360 ^ n48358;
  assign n48362 = n48359 & n48361;
  assign n48363 = n48362 ^ n44741;
  assign n48325 = n48324 ^ n48284;
  assign n48326 = ~n48285 & n48325;
  assign n48327 = n48326 ^ n48283;
  assign n48279 = n46156 ^ n45548;
  assign n48280 = n48279 ^ n47092;
  assign n47597 = n47596 ^ n3003;
  assign n47598 = n47597 ^ n47398;
  assign n48281 = n48280 ^ n47598;
  assign n48328 = n48327 ^ n48281;
  assign n48329 = n48328 ^ n44739;
  assign n48364 = n48363 ^ n48329;
  assign n48383 = n48382 ^ n48364;
  assign n48435 = n48434 ^ n48383;
  assign n48438 = n48437 ^ n48435;
  assign n48440 = n47648 ^ n46956;
  assign n48441 = n48440 ^ n46147;
  assign n48439 = n48431 ^ n48388;
  assign n48442 = n48441 ^ n48439;
  assign n48446 = n47657 ^ n46968;
  assign n48447 = n48446 ^ n46437;
  assign n48448 = n48418 ^ n48399;
  assign n48449 = n48447 & ~n48448;
  assign n48444 = n47655 ^ n46962;
  assign n48445 = n48444 ^ n46152;
  assign n48450 = n48449 ^ n48445;
  assign n48451 = n48421 ^ n48394;
  assign n48452 = n48451 ^ n48449;
  assign n48453 = n48450 & n48452;
  assign n48454 = n48453 ^ n48445;
  assign n48443 = n48428 ^ n48425;
  assign n48455 = n48454 ^ n48443;
  assign n48456 = n46957 ^ n46151;
  assign n48457 = n48456 ^ n47816;
  assign n48458 = n48457 ^ n48443;
  assign n48459 = ~n48455 & n48458;
  assign n48460 = n48459 ^ n48457;
  assign n48461 = n48460 ^ n48441;
  assign n48462 = n48442 & n48461;
  assign n48463 = n48462 ^ n48439;
  assign n48464 = n48463 ^ n48437;
  assign n48465 = n48438 & ~n48464;
  assign n48466 = n48465 ^ n48435;
  assign n48468 = n48467 ^ n48466;
  assign n48469 = n47641 ^ n46950;
  assign n48470 = n48469 ^ n46137;
  assign n48471 = n48470 ^ n48467;
  assign n48472 = n48468 & n48471;
  assign n48473 = n48472 ^ n48470;
  assign n48474 = n48473 ^ n48275;
  assign n48475 = ~n48278 & n48474;
  assign n48476 = n48475 ^ n48277;
  assign n48477 = n48476 ^ n48270;
  assign n48478 = ~n48273 & n48477;
  assign n48479 = n48478 ^ n48272;
  assign n48268 = n48162 ^ n48140;
  assign n48269 = n48268 ^ n48141;
  assign n48480 = n48479 ^ n48269;
  assign n48481 = n47632 ^ n46940;
  assign n48482 = n48481 ^ n46131;
  assign n48483 = n48482 ^ n48269;
  assign n48484 = ~n48480 & ~n48483;
  assign n48485 = n48484 ^ n48482;
  assign n48487 = n48486 ^ n48485;
  assign n48488 = n46936 ^ n46124;
  assign n48489 = n48488 ^ n47626;
  assign n48490 = n48489 ^ n48486;
  assign n48491 = n48487 & n48490;
  assign n48492 = n48491 ^ n48489;
  assign n48493 = n48492 ^ n48264;
  assign n48494 = ~n48267 & ~n48493;
  assign n48495 = n48494 ^ n48266;
  assign n48497 = n48496 ^ n48495;
  assign n48498 = n46930 ^ n46112;
  assign n48499 = n48498 ^ n47617;
  assign n48500 = n48499 ^ n48496;
  assign n48501 = n48497 & n48500;
  assign n48502 = n48501 ^ n48499;
  assign n48503 = n48502 ^ n48261;
  assign n48504 = n48263 & n48503;
  assign n48505 = n48504 ^ n48262;
  assign n48506 = n48505 ^ n48258;
  assign n48507 = ~n48259 & n48506;
  assign n48508 = n48507 ^ n48257;
  assign n48255 = n48180 ^ n48112;
  assign n48509 = n48508 ^ n48255;
  assign n48510 = n47608 ^ n46099;
  assign n48511 = n48510 ^ n46917;
  assign n48512 = n48511 ^ n48255;
  assign n48513 = ~n48509 & n48512;
  assign n48514 = n48513 ^ n48511;
  assign n48598 = n48518 ^ n48514;
  assign n48599 = ~n48597 & ~n48598;
  assign n48600 = n48599 ^ n48516;
  assign n48646 = n48601 ^ n48600;
  assign n48647 = n48604 & ~n48646;
  assign n48648 = n48647 ^ n48603;
  assign n48644 = n48189 ^ n48095;
  assign n48645 = n48644 ^ n48096;
  assign n48649 = n48648 ^ n48645;
  assign n48642 = n47876 ^ n46910;
  assign n48643 = n48642 ^ n46082;
  assign n48658 = n48645 ^ n48643;
  assign n48659 = ~n48649 & ~n48658;
  assign n48660 = n48659 ^ n48643;
  assign n48818 = n48664 ^ n48660;
  assign n48819 = ~n48817 & n48818;
  assign n48820 = n48819 ^ n48662;
  assign n48825 = n48824 ^ n48820;
  assign n48826 = n48825 ^ n46096;
  assign n48663 = n48662 ^ n48660;
  assign n48665 = n48664 ^ n48663;
  assign n48813 = n48665 ^ n46102;
  assign n48650 = n48649 ^ n48643;
  assign n48651 = n48650 ^ n46106;
  assign n48605 = n48604 ^ n48600;
  assign n48638 = n48605 ^ n46114;
  assign n48517 = n48516 ^ n48514;
  assign n48519 = n48518 ^ n48517;
  assign n48520 = n48519 ^ n46119;
  assign n48522 = n48505 ^ n48259;
  assign n48523 = n48522 ^ n45918;
  assign n48525 = n48499 ^ n48497;
  assign n48526 = n48525 ^ n45760;
  assign n48527 = n48492 ^ n48267;
  assign n48528 = n48527 ^ n45501;
  assign n48530 = n48482 ^ n48480;
  assign n48531 = n48530 ^ n45511;
  assign n48532 = n48476 ^ n48273;
  assign n48533 = n48532 ^ n45514;
  assign n48534 = n48473 ^ n48278;
  assign n48535 = n48534 ^ n45518;
  assign n48536 = n48470 ^ n48468;
  assign n48537 = n48536 ^ n45522;
  assign n48555 = n48463 ^ n48438;
  assign n48538 = n48460 ^ n48442;
  assign n48539 = n48538 ^ n45532;
  assign n48540 = n48457 ^ n48455;
  assign n48541 = n48540 ^ n45536;
  assign n48542 = n48448 ^ n48447;
  assign n48543 = ~n45543 & ~n48542;
  assign n48544 = n48543 ^ n45540;
  assign n48545 = n48451 ^ n48450;
  assign n48546 = n48545 ^ n48543;
  assign n48547 = ~n48544 & n48546;
  assign n48548 = n48547 ^ n45540;
  assign n48549 = n48548 ^ n48540;
  assign n48550 = ~n48541 & n48549;
  assign n48551 = n48550 ^ n45536;
  assign n48552 = n48551 ^ n48538;
  assign n48553 = n48539 & n48552;
  assign n48554 = n48553 ^ n45532;
  assign n48556 = n48555 ^ n48554;
  assign n48557 = n48554 ^ n45528;
  assign n48558 = n48556 & ~n48557;
  assign n48559 = n48558 ^ n45528;
  assign n48560 = n48559 ^ n48536;
  assign n48561 = n48537 & ~n48560;
  assign n48562 = n48561 ^ n45522;
  assign n48563 = n48562 ^ n48534;
  assign n48564 = n48535 & ~n48563;
  assign n48565 = n48564 ^ n45518;
  assign n48566 = n48565 ^ n48532;
  assign n48567 = n48533 & ~n48566;
  assign n48568 = n48567 ^ n45514;
  assign n48569 = n48568 ^ n48530;
  assign n48570 = n48531 & ~n48569;
  assign n48571 = n48570 ^ n45511;
  assign n48529 = n48489 ^ n48487;
  assign n48572 = n48571 ^ n48529;
  assign n48573 = n48529 ^ n45507;
  assign n48574 = ~n48572 & n48573;
  assign n48575 = n48574 ^ n45507;
  assign n48576 = n48575 ^ n48527;
  assign n48577 = ~n48528 & ~n48576;
  assign n48578 = n48577 ^ n45501;
  assign n48579 = n48578 ^ n48525;
  assign n48580 = n48526 & n48579;
  assign n48581 = n48580 ^ n45760;
  assign n48524 = n48502 ^ n48263;
  assign n48582 = n48581 ^ n48524;
  assign n48583 = n48581 ^ n45900;
  assign n48584 = n48582 & ~n48583;
  assign n48585 = n48584 ^ n45900;
  assign n48586 = n48585 ^ n48522;
  assign n48587 = n48523 & ~n48586;
  assign n48588 = n48587 ^ n45918;
  assign n48521 = n48511 ^ n48509;
  assign n48589 = n48588 ^ n48521;
  assign n48590 = n48521 ^ n46126;
  assign n48591 = n48589 & n48590;
  assign n48592 = n48591 ^ n46126;
  assign n48593 = n48592 ^ n48519;
  assign n48594 = n48520 & n48593;
  assign n48595 = n48594 ^ n46119;
  assign n48639 = n48605 ^ n48595;
  assign n48640 = n48638 & ~n48639;
  assign n48641 = n48640 ^ n46114;
  assign n48654 = n48650 ^ n48641;
  assign n48655 = ~n48651 & n48654;
  assign n48656 = n48655 ^ n46106;
  assign n48814 = n48665 ^ n48656;
  assign n48815 = ~n48813 & ~n48814;
  assign n48816 = n48815 ^ n46102;
  assign n48827 = n48826 ^ n48816;
  assign n48596 = n48595 ^ n46114;
  assign n48606 = n48605 ^ n48596;
  assign n48607 = n48592 ^ n48520;
  assign n48608 = n48589 ^ n46126;
  assign n48609 = n48578 ^ n48526;
  assign n48610 = n48575 ^ n48528;
  assign n48611 = n48568 ^ n48531;
  assign n48612 = n48545 ^ n48544;
  assign n48613 = n48548 ^ n48541;
  assign n48614 = ~n48612 & ~n48613;
  assign n48615 = n48551 ^ n48539;
  assign n48616 = ~n48614 & ~n48615;
  assign n48617 = n48556 ^ n45528;
  assign n48618 = ~n48616 & ~n48617;
  assign n48619 = n48559 ^ n48537;
  assign n48620 = ~n48618 & ~n48619;
  assign n48621 = n48562 ^ n48535;
  assign n48622 = ~n48620 & n48621;
  assign n48623 = n48565 ^ n48533;
  assign n48624 = n48622 & n48623;
  assign n48625 = n48611 & n48624;
  assign n48626 = n48572 ^ n45507;
  assign n48627 = ~n48625 & ~n48626;
  assign n48628 = n48610 & n48627;
  assign n48629 = n48609 & n48628;
  assign n48630 = n48524 ^ n45900;
  assign n48631 = n48630 ^ n48581;
  assign n48632 = n48629 & ~n48631;
  assign n48633 = n48585 ^ n48523;
  assign n48634 = n48632 & n48633;
  assign n48635 = ~n48608 & ~n48634;
  assign n48636 = n48607 & n48635;
  assign n48637 = n48606 & ~n48636;
  assign n48652 = n48651 ^ n48641;
  assign n48653 = ~n48637 & n48652;
  assign n48657 = n48656 ^ n46102;
  assign n48666 = n48665 ^ n48657;
  assign n48828 = ~n48653 & ~n48666;
  assign n49036 = n48827 & n48828;
  assign n48994 = n48825 ^ n48816;
  assign n48995 = ~n48826 & ~n48994;
  assign n48996 = n48995 ^ n46096;
  assign n48935 = n48821 ^ n48820;
  assign n48936 = n48824 & ~n48935;
  assign n48937 = n48936 ^ n48823;
  assign n48932 = n47664 ^ n46987;
  assign n48933 = n48932 ^ n48297;
  assign n48878 = n48198 ^ n48080;
  assign n48879 = n48878 ^ n48081;
  assign n48934 = n48933 ^ n48879;
  assign n48992 = n48937 ^ n48934;
  assign n48993 = n48992 ^ n46090;
  assign n49037 = n48996 ^ n48993;
  assign n49038 = n49036 & ~n49037;
  assign n48997 = n48996 ^ n48992;
  assign n48998 = ~n48993 & n48997;
  assign n48999 = n48998 ^ n46090;
  assign n48938 = n48937 ^ n48879;
  assign n48939 = n48934 & n48938;
  assign n48940 = n48939 ^ n48933;
  assign n48929 = n47680 ^ n46911;
  assign n48930 = n48929 ^ n48293;
  assign n48872 = n48201 ^ n1362;
  assign n48873 = n48872 ^ n48076;
  assign n48931 = n48930 ^ n48873;
  assign n48990 = n48940 ^ n48931;
  assign n48991 = n48990 ^ n46085;
  assign n49039 = n48999 ^ n48991;
  assign n49040 = ~n49038 & n49039;
  assign n49000 = n48999 ^ n48990;
  assign n49001 = ~n48991 & ~n49000;
  assign n49002 = n49001 ^ n46085;
  assign n49041 = n49002 ^ n46079;
  assign n48941 = n48940 ^ n48930;
  assign n48942 = n48931 & n48941;
  assign n48943 = n48942 ^ n48873;
  assign n48926 = n47694 ^ n47014;
  assign n48927 = n48926 ^ n48289;
  assign n48869 = n48204 ^ n48075;
  assign n48928 = n48927 ^ n48869;
  assign n48988 = n48943 ^ n48928;
  assign n49042 = n49041 ^ n48988;
  assign n49043 = n49040 & n49042;
  assign n48989 = n48988 ^ n46079;
  assign n49003 = n49002 ^ n48988;
  assign n49004 = n48989 & n49003;
  assign n49005 = n49004 ^ n46079;
  assign n49044 = n49005 ^ n45495;
  assign n48944 = n48943 ^ n48869;
  assign n48945 = ~n48928 & n48944;
  assign n48946 = n48945 ^ n48927;
  assign n48923 = n47713 ^ n46904;
  assign n48924 = n48923 ^ n48311;
  assign n48862 = n48211 ^ n48208;
  assign n48925 = n48924 ^ n48862;
  assign n48986 = n48946 ^ n48925;
  assign n49045 = n49044 ^ n48986;
  assign n49046 = ~n49043 & n49045;
  assign n48987 = n48986 ^ n45495;
  assign n49006 = n49005 ^ n48986;
  assign n49007 = n48987 & ~n49006;
  assign n49008 = n49007 ^ n45495;
  assign n48947 = n48946 ^ n48862;
  assign n48948 = ~n48925 & ~n48947;
  assign n48949 = n48948 ^ n48924;
  assign n48920 = n47038 ^ n46902;
  assign n48921 = n48920 ^ n48318;
  assign n48855 = n48214 ^ n48069;
  assign n48922 = n48921 ^ n48855;
  assign n48985 = n48949 ^ n48922;
  assign n49009 = n49008 ^ n48985;
  assign n49047 = n49009 ^ n46297;
  assign n49048 = n49046 & n49047;
  assign n48950 = n48949 ^ n48855;
  assign n48951 = ~n48922 & n48950;
  assign n48952 = n48951 ^ n48921;
  assign n48917 = n47104 ^ n46406;
  assign n48918 = n48917 ^ n48284;
  assign n48848 = n48217 ^ n48063;
  assign n48849 = n48848 ^ n48060;
  assign n48919 = n48918 ^ n48849;
  assign n49014 = n48952 ^ n48919;
  assign n49010 = n48985 ^ n46297;
  assign n49011 = n49009 & n49010;
  assign n49012 = n49011 ^ n46297;
  assign n49013 = n49012 ^ n45693;
  assign n49049 = n49014 ^ n49013;
  assign n49050 = ~n49048 & n49049;
  assign n49015 = n49014 ^ n49012;
  assign n49016 = ~n49013 & n49015;
  assign n49017 = n49016 ^ n45693;
  assign n48957 = n47111 ^ n46411;
  assign n48958 = n48957 ^ n47598;
  assign n48953 = n48952 ^ n48918;
  assign n48954 = n48919 & n48953;
  assign n48955 = n48954 ^ n48849;
  assign n48842 = n48220 ^ n48058;
  assign n48843 = n48842 ^ n48055;
  assign n48956 = n48955 ^ n48843;
  assign n48983 = n48958 ^ n48956;
  assign n48984 = n48983 ^ n45700;
  assign n49035 = n49017 ^ n48984;
  assign n49097 = n49050 ^ n49035;
  assign n49094 = n39320 ^ n3137;
  assign n49095 = n49094 ^ n43483;
  assign n49096 = n49095 ^ n2964;
  assign n49098 = n49097 ^ n49096;
  assign n49099 = n49049 ^ n49048;
  assign n2829 = n2828 ^ n2804;
  assign n2863 = n2862 ^ n2829;
  assign n2870 = n2869 ^ n2863;
  assign n49100 = n49099 ^ n2870;
  assign n49104 = n49047 ^ n49046;
  assign n49101 = n46692 ^ n3117;
  assign n49102 = n49101 ^ n3227;
  assign n49103 = n49102 ^ n2854;
  assign n49105 = n49104 ^ n49103;
  assign n49109 = n49045 ^ n49043;
  assign n49106 = n46697 ^ n2730;
  assign n49107 = n49106 ^ n43456;
  assign n49108 = n49107 ^ n3225;
  assign n49110 = n49109 ^ n49108;
  assign n49114 = n49042 ^ n49040;
  assign n49111 = n46702 ^ n3203;
  assign n49112 = n49111 ^ n43292;
  assign n49113 = n49112 ^ n37766;
  assign n49115 = n49114 ^ n49113;
  assign n49119 = n49039 ^ n49038;
  assign n49116 = n46707 ^ n39301;
  assign n49117 = n49116 ^ n43297;
  assign n49118 = n49117 ^ n37770;
  assign n49120 = n49119 ^ n49118;
  assign n49122 = n46712 ^ n39231;
  assign n49123 = n49122 ^ n43303;
  assign n49124 = n49123 ^ n37775;
  assign n49121 = n49037 ^ n49036;
  assign n49125 = n49124 ^ n49121;
  assign n48829 = n48828 ^ n48827;
  assign n48809 = n46718 ^ n39291;
  assign n48810 = n48809 ^ n43307;
  assign n48811 = n48810 ^ n37780;
  assign n49126 = n48829 ^ n48811;
  assign n48667 = n48666 ^ n48653;
  assign n48252 = n46722 ^ n39238;
  assign n48253 = n48252 ^ n43437;
  assign n48254 = n48253 ^ n37785;
  assign n48668 = n48667 ^ n48254;
  assign n48672 = n48652 ^ n48637;
  assign n48669 = n46850 ^ n1475;
  assign n48670 = n48669 ^ n43430;
  assign n48671 = n48670 ^ n37790;
  assign n48673 = n48672 ^ n48671;
  assign n48677 = n48636 ^ n48606;
  assign n48674 = n46729 ^ n1460;
  assign n48675 = n48674 ^ n43314;
  assign n48676 = n48675 ^ n37796;
  assign n48678 = n48677 ^ n48676;
  assign n48682 = n48635 ^ n48607;
  assign n48679 = n46733 ^ n39275;
  assign n48680 = n48679 ^ n43319;
  assign n48681 = n48680 ^ n37863;
  assign n48683 = n48682 ^ n48681;
  assign n48687 = n48634 ^ n48608;
  assign n48684 = n46738 ^ n39247;
  assign n48685 = n48684 ^ n43324;
  assign n48686 = n48685 ^ n1034;
  assign n48688 = n48687 ^ n48686;
  assign n48692 = n48633 ^ n48632;
  assign n48689 = n46743 ^ n39252;
  assign n48690 = n48689 ^ n914;
  assign n48691 = n48690 ^ n37853;
  assign n48693 = n48692 ^ n48691;
  assign n48697 = n48631 ^ n48629;
  assign n48694 = n46831 ^ n39257;
  assign n48695 = n48694 ^ n43332;
  assign n48696 = n48695 ^ n906;
  assign n48698 = n48697 ^ n48696;
  assign n48700 = n46824 ^ n788;
  assign n48701 = n48700 ^ n43408;
  assign n48702 = n48701 ^ n37843;
  assign n48699 = n48628 ^ n48609;
  assign n48703 = n48702 ^ n48699;
  assign n48707 = n46761 ^ n38761;
  assign n48708 = n48707 ^ n43391;
  assign n48709 = n48708 ^ n37814;
  assign n48706 = n48624 ^ n48611;
  assign n48710 = n48709 ^ n48706;
  assign n48712 = n46765 ^ n38766;
  assign n48713 = n48712 ^ n43344;
  assign n48714 = n48713 ^ n37818;
  assign n48711 = n48623 ^ n48622;
  assign n48715 = n48714 ^ n48711;
  assign n48719 = n48621 ^ n48620;
  assign n48716 = n46770 ^ n38770;
  assign n48717 = n48716 ^ n43381;
  assign n48718 = n48717 ^ n37236;
  assign n48720 = n48719 ^ n48718;
  assign n48722 = n46802 ^ n38775;
  assign n48723 = n48722 ^ n43351;
  assign n48724 = n48723 ^ n37207;
  assign n48721 = n48619 ^ n48618;
  assign n48725 = n48724 ^ n48721;
  assign n48727 = n46795 ^ n38799;
  assign n48728 = n48727 ^ n43356;
  assign n48729 = n48728 ^ n37212;
  assign n48726 = n48617 ^ n48616;
  assign n48730 = n48729 ^ n48726;
  assign n48735 = n48542 ^ n45543;
  assign n48736 = n47041 ^ n39196;
  assign n48737 = n48736 ^ n43622;
  assign n48738 = n48737 ^ n2092;
  assign n48739 = n48735 & n48738;
  assign n2067 = n2066 ^ n2024;
  assign n2101 = n2100 ^ n2067;
  assign n2111 = n2110 ^ n2101;
  assign n48740 = n48739 ^ n2111;
  assign n48741 = n48739 ^ n48612;
  assign n48742 = n48740 & n48741;
  assign n48743 = n48742 ^ n2111;
  assign n48732 = n46777 ^ n38787;
  assign n48733 = n48732 ^ n43362;
  assign n48734 = n48733 ^ n2247;
  assign n48744 = n48743 ^ n48734;
  assign n48745 = n48613 ^ n48612;
  assign n48746 = n48745 ^ n48743;
  assign n48747 = n48744 & n48746;
  assign n48748 = n48747 ^ n48734;
  assign n48731 = n48615 ^ n48614;
  assign n48749 = n48748 ^ n48731;
  assign n48750 = n46787 ^ n38781;
  assign n48751 = n48750 ^ n2255;
  assign n48752 = n48751 ^ n37216;
  assign n48753 = n48752 ^ n48731;
  assign n48754 = ~n48749 & n48753;
  assign n48755 = n48754 ^ n48752;
  assign n48756 = n48755 ^ n48726;
  assign n48757 = ~n48730 & n48756;
  assign n48758 = n48757 ^ n48729;
  assign n48759 = n48758 ^ n48721;
  assign n48760 = n48725 & ~n48759;
  assign n48761 = n48760 ^ n48724;
  assign n48762 = n48761 ^ n48719;
  assign n48763 = n48720 & ~n48762;
  assign n48764 = n48763 ^ n48718;
  assign n48765 = n48764 ^ n48711;
  assign n48766 = ~n48715 & n48765;
  assign n48767 = n48766 ^ n48714;
  assign n48768 = n48767 ^ n48706;
  assign n48769 = ~n48710 & n48768;
  assign n48770 = n48769 ^ n48709;
  assign n48705 = n48626 ^ n48625;
  assign n48771 = n48770 ^ n48705;
  assign n48772 = n46756 ^ n38818;
  assign n48773 = n48772 ^ n43339;
  assign n48774 = n48773 ^ n37833;
  assign n48775 = n48774 ^ n48705;
  assign n48776 = ~n48771 & n48775;
  assign n48777 = n48776 ^ n48774;
  assign n48704 = n48627 ^ n48610;
  assign n48778 = n48777 ^ n48704;
  assign n48779 = n46751 ^ n38755;
  assign n48780 = n48779 ^ n43401;
  assign n48781 = n48780 ^ n37808;
  assign n48782 = n48781 ^ n48704;
  assign n48783 = ~n48778 & n48782;
  assign n48784 = n48783 ^ n48781;
  assign n48785 = n48784 ^ n48699;
  assign n48786 = n48703 & ~n48785;
  assign n48787 = n48786 ^ n48702;
  assign n48788 = n48787 ^ n48697;
  assign n48789 = ~n48698 & n48788;
  assign n48790 = n48789 ^ n48696;
  assign n48791 = n48790 ^ n48692;
  assign n48792 = n48693 & ~n48791;
  assign n48793 = n48792 ^ n48691;
  assign n48794 = n48793 ^ n48687;
  assign n48795 = ~n48688 & n48794;
  assign n48796 = n48795 ^ n48686;
  assign n48797 = n48796 ^ n48682;
  assign n48798 = ~n48683 & n48797;
  assign n48799 = n48798 ^ n48681;
  assign n48800 = n48799 ^ n48677;
  assign n48801 = ~n48678 & n48800;
  assign n48802 = n48801 ^ n48676;
  assign n48803 = n48802 ^ n48672;
  assign n48804 = n48673 & ~n48803;
  assign n48805 = n48804 ^ n48671;
  assign n48806 = n48805 ^ n48667;
  assign n48807 = n48668 & ~n48806;
  assign n48808 = n48807 ^ n48254;
  assign n49127 = n48829 ^ n48808;
  assign n49128 = n49126 & ~n49127;
  assign n49129 = n49128 ^ n48811;
  assign n49130 = n49129 ^ n49124;
  assign n49131 = ~n49125 & ~n49130;
  assign n49132 = n49131 ^ n49121;
  assign n49133 = n49132 ^ n49119;
  assign n49134 = n49120 & n49133;
  assign n49135 = n49134 ^ n49118;
  assign n49136 = n49135 ^ n49114;
  assign n49137 = ~n49115 & n49136;
  assign n49138 = n49137 ^ n49113;
  assign n49139 = n49138 ^ n49109;
  assign n49140 = ~n49110 & n49139;
  assign n49141 = n49140 ^ n49108;
  assign n49142 = n49141 ^ n49104;
  assign n49143 = n49105 & ~n49142;
  assign n49144 = n49143 ^ n49103;
  assign n49145 = n49144 ^ n49099;
  assign n49146 = n49100 & ~n49145;
  assign n49147 = n49146 ^ n2870;
  assign n49148 = n49147 ^ n49097;
  assign n49149 = n49098 & ~n49148;
  assign n49150 = n49149 ^ n49096;
  assign n49090 = n46883 ^ n39217;
  assign n49091 = n49090 ^ n2966;
  assign n49092 = n49091 ^ n37754;
  assign n49177 = n49150 ^ n49092;
  assign n49051 = ~n49035 & ~n49050;
  assign n49018 = n49017 ^ n48983;
  assign n49019 = ~n48984 & n49018;
  assign n49020 = n49019 ^ n45700;
  assign n48963 = n47785 ^ n47101;
  assign n48964 = n48963 ^ n46403;
  assign n48959 = n48958 ^ n48843;
  assign n48960 = n48956 & n48959;
  assign n48961 = n48960 ^ n48958;
  assign n48837 = n48223 ^ n48054;
  assign n48962 = n48961 ^ n48837;
  assign n48981 = n48964 ^ n48962;
  assign n48982 = n48981 ^ n45691;
  assign n49034 = n49020 ^ n48982;
  assign n49089 = n49051 ^ n49034;
  assign n49178 = n49177 ^ n49089;
  assign n49320 = n49180 ^ n49178;
  assign n49597 = n49320 ^ n46437;
  assign n49745 = n49600 ^ n49597;
  assign n50523 = n49745 ^ n48270;
  assign n48908 = n48745 ^ n48734;
  assign n48909 = n48908 ^ n48743;
  assign n50524 = n50523 ^ n48909;
  assign n49766 = n49144 ^ n49100;
  assign n50344 = n49766 ^ n48448;
  assign n50345 = n50344 ^ n47785;
  assign n49529 = n47560 ^ n40050;
  assign n49530 = n49529 ^ n43944;
  assign n49531 = n49530 ^ n38574;
  assign n48876 = n48784 ^ n48703;
  assign n48874 = n48873 ^ n46915;
  assign n48875 = n48874 ^ n47999;
  assign n48877 = n48876 ^ n48875;
  assign n48882 = n48781 ^ n48778;
  assign n48880 = n48879 ^ n47187;
  assign n48881 = n48880 ^ n47876;
  assign n48883 = n48882 ^ n48881;
  assign n48886 = n48774 ^ n48771;
  assign n48884 = n47603 ^ n46917;
  assign n48885 = n48884 ^ n48821;
  assign n48887 = n48886 ^ n48885;
  assign n49237 = n48767 ^ n48710;
  assign n48890 = n48764 ^ n48714;
  assign n48891 = n48890 ^ n48711;
  assign n48888 = n48645 ^ n47608;
  assign n48889 = n48888 ^ n46926;
  assign n48892 = n48891 ^ n48889;
  assign n48895 = n48761 ^ n48720;
  assign n48893 = n48601 ^ n46930;
  assign n48894 = n48893 ^ n47609;
  assign n48896 = n48895 ^ n48894;
  assign n48899 = n48758 ^ n48724;
  assign n48900 = n48899 ^ n48721;
  assign n48897 = n48518 ^ n47613;
  assign n48898 = n48897 ^ n46935;
  assign n48901 = n48900 ^ n48898;
  assign n48904 = n48755 ^ n48730;
  assign n48902 = n47617 ^ n46936;
  assign n48903 = n48902 ^ n48255;
  assign n48905 = n48904 ^ n48903;
  assign n49218 = n48752 ^ n48749;
  assign n48906 = n48262 ^ n47626;
  assign n48907 = n48906 ^ n46941;
  assign n48910 = n48909 ^ n48907;
  assign n49207 = n48612 ^ n2111;
  assign n49208 = n49207 ^ n48739;
  assign n49200 = n48738 ^ n48735;
  assign n49168 = n48486 ^ n47833;
  assign n49169 = n49168 ^ n46955;
  assign n49052 = n49034 & ~n49051;
  assign n48965 = n48964 ^ n48837;
  assign n48966 = ~n48962 & n48965;
  assign n48967 = n48966 ^ n48964;
  assign n48914 = n47096 ^ n46401;
  assign n48915 = n48914 ^ n47793;
  assign n48833 = n48226 ^ n48049;
  assign n48916 = n48915 ^ n48833;
  assign n49024 = n48967 ^ n48916;
  assign n49053 = n49024 ^ n45707;
  assign n49021 = n49020 ^ n48981;
  assign n49022 = ~n48982 & ~n49021;
  assign n49023 = n49022 ^ n45691;
  assign n49054 = n49053 ^ n49023;
  assign n49055 = ~n49052 & n49054;
  assign n49025 = n49024 ^ n49023;
  assign n49026 = n49023 ^ n45707;
  assign n49027 = n49025 & n49026;
  assign n49028 = n49027 ^ n45707;
  assign n48968 = n48967 ^ n48915;
  assign n48969 = n48916 & n48968;
  assign n48970 = n48969 ^ n48833;
  assign n48911 = n47781 ^ n47092;
  assign n48912 = n48911 ^ n46395;
  assign n48250 = n48249 ^ n48229;
  assign n48913 = n48912 ^ n48250;
  assign n48980 = n48970 ^ n48913;
  assign n49029 = n49028 ^ n48980;
  assign n49056 = n49029 ^ n45685;
  assign n49057 = n49055 & ~n49056;
  assign n49030 = n48980 ^ n45685;
  assign n49031 = n49029 & n49030;
  assign n49032 = n49031 ^ n45685;
  assign n48976 = n48412 ^ n48409;
  assign n48974 = n47779 ^ n46158;
  assign n48975 = n48974 ^ n46975;
  assign n48977 = n48976 ^ n48975;
  assign n48971 = n48970 ^ n48250;
  assign n48972 = ~n48913 & ~n48971;
  assign n48973 = n48972 ^ n48912;
  assign n48978 = n48977 ^ n48973;
  assign n48979 = n48978 ^ n45552;
  assign n49033 = n49032 ^ n48979;
  assign n49081 = n49057 ^ n49033;
  assign n49078 = n47063 ^ n39202;
  assign n49079 = n49078 ^ n43632;
  assign n49080 = n49079 ^ n37739;
  assign n49082 = n49081 ^ n49080;
  assign n49084 = n47069 ^ n39207;
  assign n49085 = n49084 ^ n43637;
  assign n49086 = n49085 ^ n37744;
  assign n49083 = n49056 ^ n49055;
  assign n49087 = n49086 ^ n49083;
  assign n49093 = n49092 ^ n49089;
  assign n49151 = n49150 ^ n49089;
  assign n49152 = n49093 & ~n49151;
  assign n49153 = n49152 ^ n49092;
  assign n49088 = n49054 ^ n49052;
  assign n49154 = n49153 ^ n49088;
  assign n49158 = n49157 ^ n49088;
  assign n49159 = n49154 & ~n49158;
  assign n49160 = n49159 ^ n49157;
  assign n49161 = n49160 ^ n49083;
  assign n49162 = ~n49087 & n49161;
  assign n49163 = n49162 ^ n49086;
  assign n49164 = n49163 ^ n49081;
  assign n49165 = n49082 & ~n49164;
  assign n49166 = n49165 ^ n49080;
  assign n49072 = n49032 ^ n48978;
  assign n49073 = ~n48979 & ~n49072;
  assign n49074 = n49073 ^ n45552;
  assign n49075 = n49074 ^ n45548;
  assign n49067 = n48975 ^ n48973;
  assign n49068 = ~n48977 & n49067;
  assign n49069 = n49068 ^ n48973;
  assign n49065 = n48415 ^ n48403;
  assign n49066 = n49065 ^ n48400;
  assign n49070 = n49069 ^ n49066;
  assign n49063 = n46973 ^ n46156;
  assign n49064 = n49063 ^ n47775;
  assign n49071 = n49070 ^ n49064;
  assign n49076 = n49075 ^ n49071;
  assign n49059 = n47059 ^ n1932;
  assign n49060 = n49059 ^ n43627;
  assign n49061 = n49060 ^ n37734;
  assign n49058 = n49033 & ~n49057;
  assign n49062 = n49061 ^ n49058;
  assign n49077 = n49076 ^ n49062;
  assign n49167 = n49166 ^ n49077;
  assign n49170 = n49169 ^ n49167;
  assign n49172 = n47641 ^ n46956;
  assign n49173 = n49172 ^ n48269;
  assign n49171 = n49163 ^ n49082;
  assign n49174 = n49173 ^ n49171;
  assign n49182 = n48275 ^ n47648;
  assign n49183 = n49182 ^ n46962;
  assign n49181 = n49178 & n49180;
  assign n49184 = n49183 ^ n49181;
  assign n49185 = n49157 ^ n49154;
  assign n49186 = n49185 ^ n49183;
  assign n49187 = ~n49184 & ~n49186;
  assign n49188 = n49187 ^ n49181;
  assign n49175 = n48270 ^ n47645;
  assign n49176 = n49175 ^ n46957;
  assign n49189 = n49188 ^ n49176;
  assign n49190 = n49160 ^ n49087;
  assign n49191 = n49190 ^ n49188;
  assign n49192 = n49189 & n49191;
  assign n49193 = n49192 ^ n49176;
  assign n49194 = n49193 ^ n49171;
  assign n49195 = ~n49174 & ~n49194;
  assign n49196 = n49195 ^ n49173;
  assign n49197 = n49196 ^ n49169;
  assign n49198 = n49170 & ~n49197;
  assign n49199 = n49198 ^ n49167;
  assign n49201 = n49200 ^ n49199;
  assign n49202 = n47634 ^ n46950;
  assign n49203 = n49202 ^ n48264;
  assign n49204 = n49203 ^ n49200;
  assign n49205 = n49201 & n49204;
  assign n49206 = n49205 ^ n49203;
  assign n49209 = n49208 ^ n49206;
  assign n49210 = n47632 ^ n46945;
  assign n49211 = n49210 ^ n48496;
  assign n49212 = n49211 ^ n49208;
  assign n49213 = n49209 & ~n49212;
  assign n49214 = n49213 ^ n49211;
  assign n49215 = n49214 ^ n48909;
  assign n49216 = n48910 & n49215;
  assign n49217 = n49216 ^ n48907;
  assign n49219 = n49218 ^ n49217;
  assign n49220 = n47621 ^ n46940;
  assign n49221 = n49220 ^ n48258;
  assign n49222 = n49221 ^ n49218;
  assign n49223 = n49219 & ~n49222;
  assign n49224 = n49223 ^ n49221;
  assign n49225 = n49224 ^ n48904;
  assign n49226 = ~n48905 & ~n49225;
  assign n49227 = n49226 ^ n48903;
  assign n49228 = n49227 ^ n48900;
  assign n49229 = ~n48901 & ~n49228;
  assign n49230 = n49229 ^ n48898;
  assign n49231 = n49230 ^ n48894;
  assign n49232 = ~n48896 & ~n49231;
  assign n49233 = n49232 ^ n48895;
  assign n49234 = n49233 ^ n48891;
  assign n49235 = ~n48892 & n49234;
  assign n49236 = n49235 ^ n48889;
  assign n49238 = n49237 ^ n49236;
  assign n49239 = n48664 ^ n46922;
  assign n49240 = n49239 ^ n47607;
  assign n49241 = n49240 ^ n49237;
  assign n49242 = n49238 & n49241;
  assign n49243 = n49242 ^ n49240;
  assign n49244 = n49243 ^ n48886;
  assign n49245 = ~n48887 & n49244;
  assign n49246 = n49245 ^ n48885;
  assign n49247 = n49246 ^ n48882;
  assign n49248 = n48883 & n49247;
  assign n49249 = n49248 ^ n48881;
  assign n49250 = n49249 ^ n48876;
  assign n49251 = ~n48877 & ~n49250;
  assign n49252 = n49251 ^ n48875;
  assign n48868 = n48239 ^ n46910;
  assign n48870 = n48869 ^ n48868;
  assign n48866 = n48787 ^ n48696;
  assign n48867 = n48866 ^ n48697;
  assign n48871 = n48870 ^ n48867;
  assign n49290 = n49252 ^ n48871;
  assign n49291 = n49290 ^ n46082;
  assign n49292 = n49249 ^ n48877;
  assign n49293 = n49292 ^ n46088;
  assign n49294 = n49246 ^ n48881;
  assign n49295 = n49294 ^ n48882;
  assign n49296 = n49295 ^ n46093;
  assign n49297 = n49243 ^ n48887;
  assign n49298 = n49297 ^ n46099;
  assign n49299 = n49240 ^ n49238;
  assign n49300 = n49299 ^ n46101;
  assign n49301 = n49233 ^ n48892;
  assign n49302 = n49301 ^ n46109;
  assign n49303 = n49230 ^ n48896;
  assign n49304 = n49303 ^ n46112;
  assign n49305 = n49227 ^ n48901;
  assign n49306 = n49305 ^ n46118;
  assign n49307 = n49224 ^ n48905;
  assign n49308 = n49307 ^ n46124;
  assign n49311 = n49211 ^ n49209;
  assign n49312 = n49311 ^ n46133;
  assign n49313 = n49203 ^ n49201;
  assign n49314 = n49313 ^ n46137;
  assign n49315 = n49196 ^ n49170;
  assign n49316 = n49315 ^ n46142;
  assign n49317 = n49193 ^ n49173;
  assign n49318 = n49317 ^ n49171;
  assign n49319 = n49318 ^ n46147;
  assign n49321 = ~n46437 & n49320;
  assign n49322 = n49321 ^ n46152;
  assign n49323 = n49185 ^ n49184;
  assign n49324 = n49323 ^ n49321;
  assign n49325 = ~n49322 & ~n49324;
  assign n49326 = n49325 ^ n46152;
  assign n49327 = n49326 ^ n46151;
  assign n49328 = n49190 ^ n49189;
  assign n49329 = n49328 ^ n49326;
  assign n49330 = ~n49327 & ~n49329;
  assign n49331 = n49330 ^ n46151;
  assign n49332 = n49331 ^ n49318;
  assign n49333 = ~n49319 & n49332;
  assign n49334 = n49333 ^ n46147;
  assign n49335 = n49334 ^ n49315;
  assign n49336 = ~n49316 & n49335;
  assign n49337 = n49336 ^ n46142;
  assign n49338 = n49337 ^ n49313;
  assign n49339 = n49314 & n49338;
  assign n49340 = n49339 ^ n46137;
  assign n49341 = n49340 ^ n49311;
  assign n49342 = ~n49312 & ~n49341;
  assign n49343 = n49342 ^ n46133;
  assign n49310 = n49214 ^ n48910;
  assign n49344 = n49343 ^ n49310;
  assign n49345 = n49310 ^ n46132;
  assign n49346 = ~n49344 & n49345;
  assign n49347 = n49346 ^ n46132;
  assign n49309 = n49221 ^ n49219;
  assign n49348 = n49347 ^ n49309;
  assign n49349 = n49309 ^ n46131;
  assign n49350 = ~n49348 & ~n49349;
  assign n49351 = n49350 ^ n46131;
  assign n49352 = n49351 ^ n49307;
  assign n49353 = n49308 & n49352;
  assign n49354 = n49353 ^ n46124;
  assign n49355 = n49354 ^ n49305;
  assign n49356 = n49306 & n49355;
  assign n49357 = n49356 ^ n46118;
  assign n49358 = n49357 ^ n49303;
  assign n49359 = n49304 & n49358;
  assign n49360 = n49359 ^ n46112;
  assign n49361 = n49360 ^ n49301;
  assign n49362 = n49302 & n49361;
  assign n49363 = n49362 ^ n46109;
  assign n49364 = n49363 ^ n49299;
  assign n49365 = n49300 & n49364;
  assign n49366 = n49365 ^ n46101;
  assign n49367 = n49366 ^ n49297;
  assign n49368 = ~n49298 & ~n49367;
  assign n49369 = n49368 ^ n46099;
  assign n49370 = n49369 ^ n49295;
  assign n49371 = n49296 & ~n49370;
  assign n49372 = n49371 ^ n46093;
  assign n49373 = n49372 ^ n49292;
  assign n49374 = ~n49293 & ~n49373;
  assign n49375 = n49374 ^ n46088;
  assign n49376 = n49375 ^ n49290;
  assign n49377 = n49291 & ~n49376;
  assign n49378 = n49377 ^ n46082;
  assign n49253 = n49252 ^ n48870;
  assign n49254 = ~n48871 & n49253;
  assign n49255 = n49254 ^ n48867;
  assign n48863 = n48862 ^ n46907;
  assign n48864 = n48863 ^ n48297;
  assign n48860 = n48790 ^ n48691;
  assign n48861 = n48860 ^ n48692;
  assign n48865 = n48864 ^ n48861;
  assign n49288 = n49255 ^ n48865;
  assign n49289 = n49288 ^ n46077;
  assign n49405 = n49378 ^ n49289;
  assign n49406 = n49372 ^ n49293;
  assign n49407 = n49363 ^ n49300;
  assign n49408 = n49360 ^ n49302;
  assign n49409 = n49357 ^ n46112;
  assign n49410 = n49409 ^ n49303;
  assign n49411 = n49348 ^ n46131;
  assign n49412 = n49344 ^ n46132;
  assign n49413 = n49340 ^ n46133;
  assign n49414 = n49413 ^ n49311;
  assign n49415 = n49334 ^ n49316;
  assign n49416 = n49323 ^ n49322;
  assign n49417 = n49328 ^ n49327;
  assign n49418 = n49416 & ~n49417;
  assign n49419 = n49331 ^ n49319;
  assign n49420 = ~n49418 & ~n49419;
  assign n49421 = n49415 & ~n49420;
  assign n49422 = n49337 ^ n49314;
  assign n49423 = ~n49421 & n49422;
  assign n49424 = ~n49414 & ~n49423;
  assign n49425 = ~n49412 & n49424;
  assign n49426 = n49411 & n49425;
  assign n49427 = n49351 ^ n49308;
  assign n49428 = ~n49426 & ~n49427;
  assign n49429 = n49354 ^ n49306;
  assign n49430 = n49428 & n49429;
  assign n49431 = ~n49410 & n49430;
  assign n49432 = n49408 & n49431;
  assign n49433 = ~n49407 & n49432;
  assign n49434 = n49366 ^ n46099;
  assign n49435 = n49434 ^ n49297;
  assign n49436 = ~n49433 & n49435;
  assign n49437 = n49369 ^ n49296;
  assign n49438 = n49436 & n49437;
  assign n49439 = n49406 & ~n49438;
  assign n49440 = n49375 ^ n49291;
  assign n49441 = ~n49439 & ~n49440;
  assign n49442 = n49405 & ~n49441;
  assign n49379 = n49378 ^ n49288;
  assign n49380 = n49289 & ~n49379;
  assign n49381 = n49380 ^ n46077;
  assign n49256 = n49255 ^ n48861;
  assign n49257 = ~n48865 & n49256;
  assign n49258 = n49257 ^ n48864;
  assign n48857 = n48793 ^ n48686;
  assign n48858 = n48857 ^ n48687;
  assign n48854 = n48293 ^ n47206;
  assign n48856 = n48855 ^ n48854;
  assign n48859 = n48858 ^ n48856;
  assign n49286 = n49258 ^ n48859;
  assign n49287 = n49286 ^ n46889;
  assign n49404 = n49381 ^ n49287;
  assign n49528 = n49442 ^ n49404;
  assign n49532 = n49531 ^ n49528;
  assign n49536 = n49441 ^ n49405;
  assign n49533 = n47553 ^ n39956;
  assign n49534 = n49533 ^ n43949;
  assign n49535 = n49534 ^ n38540;
  assign n49537 = n49536 ^ n49535;
  assign n49541 = n49440 ^ n49439;
  assign n49538 = n47546 ^ n39962;
  assign n49539 = n49538 ^ n1325;
  assign n49540 = n49539 ^ n38564;
  assign n49542 = n49541 ^ n49540;
  assign n49546 = n49438 ^ n49406;
  assign n49543 = n47427 ^ n39967;
  assign n49544 = n49543 ^ n43955;
  assign n49545 = n49544 ^ n1317;
  assign n49547 = n49546 ^ n49545;
  assign n49548 = n49437 ^ n49436;
  assign n1125 = n1124 ^ n1079;
  assign n1159 = n1158 ^ n1125;
  assign n1169 = n1168 ^ n1159;
  assign n49549 = n49548 ^ n1169;
  assign n49554 = n49432 ^ n49407;
  assign n49551 = n47530 ^ n984;
  assign n49552 = n49551 ^ n43967;
  assign n49553 = n49552 ^ n3332;
  assign n49555 = n49554 ^ n49553;
  assign n49556 = n49431 ^ n49408;
  assign n49560 = n49559 ^ n49556;
  assign n49564 = n49430 ^ n49410;
  assign n49561 = n47441 ^ n39985;
  assign n49562 = n49561 ^ n43977;
  assign n49563 = n49562 ^ n38084;
  assign n49565 = n49564 ^ n49563;
  assign n49572 = n49427 ^ n49426;
  assign n49569 = n47450 ^ n39995;
  assign n49570 = n49569 ^ n44039;
  assign n49571 = n49570 ^ n38149;
  assign n49573 = n49572 ^ n49571;
  assign n49577 = n49425 ^ n49411;
  assign n49574 = n47455 ^ n39999;
  assign n49575 = n49574 ^ n44032;
  assign n49576 = n49575 ^ n38094;
  assign n49578 = n49577 ^ n49576;
  assign n49582 = n49424 ^ n49412;
  assign n49579 = n47461 ^ n40004;
  assign n49580 = n49579 ^ n43986;
  assign n49581 = n49580 ^ n38099;
  assign n49583 = n49582 ^ n49581;
  assign n49587 = n49423 ^ n49414;
  assign n49584 = n47466 ^ n39432;
  assign n49585 = n49584 ^ n44022;
  assign n49586 = n49585 ^ n38105;
  assign n49588 = n49587 ^ n49586;
  assign n49593 = n49420 ^ n49415;
  assign n49590 = n47471 ^ n39423;
  assign n49591 = n49590 ^ n2407;
  assign n49592 = n49591 ^ n38130;
  assign n49594 = n49593 ^ n49592;
  assign n49602 = n47476 ^ n2185;
  assign n49603 = n49602 ^ n44003;
  assign n49604 = n49603 ^ n38116;
  assign n49601 = ~n49597 & n49600;
  assign n49605 = n49604 ^ n49601;
  assign n49606 = n49601 ^ n49416;
  assign n49607 = n49605 & ~n49606;
  assign n49608 = n49607 ^ n49604;
  assign n49596 = n49417 ^ n49416;
  assign n49609 = n49608 ^ n49596;
  assign n49610 = n47481 ^ n2203;
  assign n49611 = n49610 ^ n44000;
  assign n49612 = n49611 ^ n2381;
  assign n49613 = n49612 ^ n49608;
  assign n49614 = ~n49609 & n49613;
  assign n49615 = n49614 ^ n49612;
  assign n49595 = n49419 ^ n49418;
  assign n49616 = n49615 ^ n49595;
  assign n2365 = n2352 ^ n2289;
  assign n2390 = n2389 ^ n2365;
  assign n2397 = n2396 ^ n2390;
  assign n49617 = n49615 ^ n2397;
  assign n49618 = ~n49616 & n49617;
  assign n49619 = n49618 ^ n2397;
  assign n49620 = n49619 ^ n49593;
  assign n49621 = n49594 & ~n49620;
  assign n49622 = n49621 ^ n49592;
  assign n49589 = n49422 ^ n49421;
  assign n49623 = n49622 ^ n49589;
  assign n49624 = n47497 ^ n39406;
  assign n49625 = n49624 ^ n43991;
  assign n49626 = n49625 ^ n38109;
  assign n49627 = n49626 ^ n49589;
  assign n49628 = n49623 & ~n49627;
  assign n49629 = n49628 ^ n49626;
  assign n49630 = n49629 ^ n49587;
  assign n49631 = ~n49588 & n49630;
  assign n49632 = n49631 ^ n49586;
  assign n49633 = n49632 ^ n49582;
  assign n49634 = n49583 & ~n49633;
  assign n49635 = n49634 ^ n49581;
  assign n49636 = n49635 ^ n49577;
  assign n49637 = ~n49578 & n49636;
  assign n49638 = n49637 ^ n49576;
  assign n49639 = n49638 ^ n49572;
  assign n49640 = n49573 & ~n49639;
  assign n49641 = n49640 ^ n49571;
  assign n49566 = n47445 ^ n39990;
  assign n49567 = n49566 ^ n44046;
  assign n49568 = n49567 ^ n38088;
  assign n49642 = n49641 ^ n49568;
  assign n49643 = n49429 ^ n49428;
  assign n49644 = n49643 ^ n49641;
  assign n49645 = n49642 & ~n49644;
  assign n49646 = n49645 ^ n49568;
  assign n49647 = n49646 ^ n49564;
  assign n49648 = ~n49565 & n49647;
  assign n49649 = n49648 ^ n49563;
  assign n49650 = n49649 ^ n49556;
  assign n49651 = n49560 & ~n49650;
  assign n49652 = n49651 ^ n49559;
  assign n49653 = n49652 ^ n49554;
  assign n49654 = ~n49555 & n49653;
  assign n49655 = n49654 ^ n49553;
  assign n49550 = n49435 ^ n49433;
  assign n49656 = n49655 ^ n49550;
  assign n49657 = n47434 ^ n39973;
  assign n49658 = n49657 ^ n43963;
  assign n49659 = n49658 ^ n1150;
  assign n49660 = n49659 ^ n49550;
  assign n49661 = ~n49656 & n49660;
  assign n49662 = n49661 ^ n49659;
  assign n49663 = n49662 ^ n49548;
  assign n49664 = ~n49549 & n49663;
  assign n49665 = n49664 ^ n1169;
  assign n49666 = n49665 ^ n49546;
  assign n49667 = ~n49547 & n49666;
  assign n49668 = n49667 ^ n49545;
  assign n49669 = n49668 ^ n49541;
  assign n49670 = ~n49542 & n49669;
  assign n49671 = n49670 ^ n49540;
  assign n49672 = n49671 ^ n49536;
  assign n49673 = ~n49537 & n49672;
  assign n49674 = n49673 ^ n49535;
  assign n49675 = n49674 ^ n49528;
  assign n49676 = ~n49532 & n49675;
  assign n49677 = n49676 ^ n49531;
  assign n49443 = ~n49404 & n49442;
  assign n49382 = n49381 ^ n49286;
  assign n49383 = ~n49287 & n49382;
  assign n49384 = n49383 ^ n46889;
  assign n49259 = n49258 ^ n48858;
  assign n49260 = n48859 & ~n49259;
  assign n49261 = n49260 ^ n48856;
  assign n48850 = n48849 ^ n47664;
  assign n48851 = n48850 ^ n48289;
  assign n49283 = n49261 ^ n48851;
  assign n48852 = n48796 ^ n48683;
  assign n49284 = n49283 ^ n48852;
  assign n49285 = n49284 ^ n46987;
  assign n49403 = n49384 ^ n49285;
  assign n49526 = n49443 ^ n49403;
  assign n49523 = n47567 ^ n39950;
  assign n49524 = n49523 ^ n44080;
  assign n49525 = n49524 ^ n38533;
  assign n49527 = n49526 ^ n49525;
  assign n50343 = n49677 ^ n49527;
  assign n50346 = n50345 ^ n50343;
  assign n50137 = n49066 ^ n47598;
  assign n49749 = n49141 ^ n49105;
  assign n50138 = n50137 ^ n49749;
  assign n50136 = n49674 ^ n49532;
  assign n50139 = n50138 ^ n50136;
  assign n50062 = n48318 ^ n48250;
  assign n49481 = n49135 ^ n49115;
  assign n50063 = n50062 ^ n49481;
  assign n50061 = n49668 ^ n49542;
  assign n50064 = n50063 ^ n50061;
  assign n49466 = n49132 ^ n49118;
  assign n49467 = n49466 ^ n49119;
  assign n49945 = n49467 ^ n48833;
  assign n49946 = n49945 ^ n48311;
  assign n49943 = n49665 ^ n49545;
  assign n49944 = n49943 ^ n49546;
  assign n49947 = n49946 ^ n49944;
  assign n49710 = n48843 ^ n48293;
  assign n48812 = n48811 ^ n48808;
  assign n48830 = n48829 ^ n48812;
  assign n49711 = n49710 ^ n48830;
  assign n49709 = n49659 ^ n49656;
  assign n49712 = n49711 ^ n49709;
  assign n49715 = n49652 ^ n49555;
  assign n48835 = n48805 ^ n48668;
  assign n49713 = n48849 ^ n48835;
  assign n49714 = n49713 ^ n48297;
  assign n49716 = n49715 ^ n49714;
  assign n49918 = n49646 ^ n49565;
  assign n49911 = n49643 ^ n49642;
  assign n49721 = n49638 ^ n49573;
  assign n49719 = n48873 ^ n48858;
  assign n49720 = n49719 ^ n47603;
  assign n49722 = n49721 ^ n49720;
  assign n49901 = n49635 ^ n49578;
  assign n49725 = n49632 ^ n49583;
  assign n49723 = n48821 ^ n47608;
  assign n49724 = n49723 ^ n48867;
  assign n49726 = n49725 ^ n49724;
  assign n49729 = n48882 ^ n47613;
  assign n49730 = n49729 ^ n48645;
  assign n49728 = n49626 ^ n49623;
  assign n49731 = n49730 ^ n49728;
  assign n49735 = n49616 ^ n2397;
  assign n49733 = n48518 ^ n47621;
  assign n49734 = n49733 ^ n49237;
  assign n49736 = n49735 ^ n49734;
  assign n49740 = n49604 ^ n49416;
  assign n49741 = n49740 ^ n49601;
  assign n49738 = n48258 ^ n47632;
  assign n49739 = n49738 ^ n48895;
  assign n49742 = n49741 ^ n49739;
  assign n49743 = n48900 ^ n47634;
  assign n49744 = n49743 ^ n48262;
  assign n49746 = n49745 ^ n49744;
  assign n49844 = n49208 ^ n48269;
  assign n49845 = n49844 ^ n47648;
  assign n49700 = n39930 ^ n3003;
  assign n49701 = n49700 ^ n44273;
  assign n49702 = n49701 ^ n38509;
  assign n49454 = n47785 ^ n47104;
  assign n49455 = n49454 ^ n48976;
  assign n47599 = n47598 ^ n46902;
  assign n48251 = n48250 ^ n47599;
  assign n48831 = n48830 ^ n48251;
  assign n48832 = n48284 ^ n47713;
  assign n48834 = n48833 ^ n48832;
  assign n48836 = n48835 ^ n48834;
  assign n48840 = n48802 ^ n48673;
  assign n48838 = n48837 ^ n48318;
  assign n48839 = n48838 ^ n47694;
  assign n48841 = n48840 ^ n48839;
  assign n48846 = n48799 ^ n48678;
  assign n48844 = n48843 ^ n48311;
  assign n48845 = n48844 ^ n47680;
  assign n48847 = n48846 ^ n48845;
  assign n48853 = n48852 ^ n48851;
  assign n49262 = n49261 ^ n48852;
  assign n49263 = ~n48853 & ~n49262;
  assign n49264 = n49263 ^ n48851;
  assign n49265 = n49264 ^ n48846;
  assign n49266 = ~n48847 & n49265;
  assign n49267 = n49266 ^ n48845;
  assign n49268 = n49267 ^ n48840;
  assign n49269 = n48841 & ~n49268;
  assign n49270 = n49269 ^ n48839;
  assign n49271 = n49270 ^ n48835;
  assign n49272 = n48836 & ~n49271;
  assign n49273 = n49272 ^ n48834;
  assign n49450 = n49273 ^ n48251;
  assign n49451 = ~n48831 & n49450;
  assign n49452 = n49451 ^ n48830;
  assign n49449 = n49129 ^ n49125;
  assign n49453 = n49452 ^ n49449;
  assign n49456 = n49455 ^ n49453;
  assign n49473 = n49456 ^ n46406;
  assign n49275 = n49270 ^ n48836;
  assign n49276 = n49275 ^ n46904;
  assign n49277 = n49267 ^ n48839;
  assign n49278 = n49277 ^ n48840;
  assign n49279 = n49278 ^ n47014;
  assign n49280 = n49264 ^ n48845;
  assign n49281 = n49280 ^ n48846;
  assign n49282 = n49281 ^ n46911;
  assign n49385 = n49384 ^ n49284;
  assign n49386 = n49285 & ~n49385;
  assign n49387 = n49386 ^ n46987;
  assign n49388 = n49387 ^ n49281;
  assign n49389 = ~n49282 & n49388;
  assign n49390 = n49389 ^ n46911;
  assign n49391 = n49390 ^ n49278;
  assign n49392 = n49279 & ~n49391;
  assign n49393 = n49392 ^ n47014;
  assign n49394 = n49393 ^ n49275;
  assign n49395 = n49276 & ~n49394;
  assign n49396 = n49395 ^ n46904;
  assign n49274 = n49273 ^ n48831;
  assign n49397 = n49396 ^ n49274;
  assign n49457 = n49274 ^ n47038;
  assign n49458 = n49397 & n49457;
  assign n49459 = n49458 ^ n47038;
  assign n49474 = n49459 ^ n49456;
  assign n49475 = ~n49473 & n49474;
  assign n49476 = n49475 ^ n46406;
  assign n49469 = n49066 ^ n47111;
  assign n49470 = n49469 ^ n47793;
  assign n49463 = n49455 ^ n49449;
  assign n49464 = n49453 & n49463;
  assign n49465 = n49464 ^ n49455;
  assign n49468 = n49467 ^ n49465;
  assign n49471 = n49470 ^ n49468;
  assign n49472 = n49471 ^ n46411;
  assign n49477 = n49476 ^ n49472;
  assign n49398 = n49397 ^ n47038;
  assign n49399 = n49393 ^ n49276;
  assign n49400 = n49390 ^ n49279;
  assign n49401 = n49387 ^ n46911;
  assign n49402 = n49401 ^ n49281;
  assign n49444 = n49403 & n49443;
  assign n49445 = n49402 & ~n49444;
  assign n49446 = ~n49400 & n49445;
  assign n49447 = n49399 & ~n49446;
  assign n49448 = n49398 & n49447;
  assign n49460 = n49459 ^ n46406;
  assign n49461 = n49460 ^ n49456;
  assign n49462 = ~n49448 & ~n49461;
  assign n49496 = n49477 ^ n49462;
  assign n49493 = n47401 ^ n2938;
  assign n49494 = n49493 ^ n44289;
  assign n49495 = n49494 ^ n38599;
  assign n49497 = n49496 ^ n49495;
  assign n49499 = n47407 ^ n2922;
  assign n49500 = n49499 ^ n44278;
  assign n49501 = n49500 ^ n38515;
  assign n49498 = n49461 ^ n49448;
  assign n49502 = n49501 ^ n49498;
  assign n49504 = n47587 ^ n3237;
  assign n49505 = n49504 ^ n44095;
  assign n49506 = n49505 ^ n38520;
  assign n49503 = n49447 ^ n49398;
  assign n49507 = n49506 ^ n49503;
  assign n49511 = n49446 ^ n49399;
  assign n49508 = n47413 ^ n39940;
  assign n49509 = n49508 ^ n43490;
  assign n49510 = n49509 ^ n38525;
  assign n49512 = n49511 ^ n49510;
  assign n49516 = n49445 ^ n49400;
  assign n49513 = n47417 ^ n39944;
  assign n49514 = n49513 ^ n43932;
  assign n49515 = n49514 ^ n3083;
  assign n49517 = n49516 ^ n49515;
  assign n49521 = n49444 ^ n49402;
  assign n49518 = n47574 ^ n40060;
  assign n49519 = n49518 ^ n43937;
  assign n49520 = n49519 ^ n2573;
  assign n49522 = n49521 ^ n49520;
  assign n49678 = n49677 ^ n49526;
  assign n49679 = n49527 & ~n49678;
  assign n49680 = n49679 ^ n49525;
  assign n49681 = n49680 ^ n49521;
  assign n49682 = n49522 & ~n49681;
  assign n49683 = n49682 ^ n49520;
  assign n49684 = n49683 ^ n49516;
  assign n49685 = n49517 & ~n49684;
  assign n49686 = n49685 ^ n49515;
  assign n49687 = n49686 ^ n49511;
  assign n49688 = ~n49512 & n49687;
  assign n49689 = n49688 ^ n49510;
  assign n49690 = n49689 ^ n49506;
  assign n49691 = n49507 & ~n49690;
  assign n49692 = n49691 ^ n49503;
  assign n49693 = n49692 ^ n49498;
  assign n49694 = ~n49502 & n49693;
  assign n49695 = n49694 ^ n49501;
  assign n49696 = n49695 ^ n49496;
  assign n49697 = ~n49497 & n49696;
  assign n49698 = n49697 ^ n49495;
  assign n49487 = n49476 ^ n49471;
  assign n49488 = ~n49472 & n49487;
  assign n49489 = n49488 ^ n46411;
  assign n49490 = n49489 ^ n46403;
  assign n49483 = n49470 ^ n49467;
  assign n49484 = ~n49468 & ~n49483;
  assign n49485 = n49484 ^ n49470;
  assign n49479 = n48448 ^ n47101;
  assign n49480 = n49479 ^ n47781;
  assign n49482 = n49481 ^ n49480;
  assign n49486 = n49485 ^ n49482;
  assign n49491 = n49490 ^ n49486;
  assign n49478 = ~n49462 & n49477;
  assign n49492 = n49491 ^ n49478;
  assign n49699 = n49698 ^ n49492;
  assign n49703 = n49702 ^ n49699;
  assign n49841 = n49200 ^ n47816;
  assign n49842 = n49841 ^ n48270;
  assign n49843 = ~n49703 & n49842;
  assign n49846 = n49845 ^ n49843;
  assign n49824 = n47758 ^ n40087;
  assign n49825 = n49824 ^ n44269;
  assign n49826 = n49825 ^ n38504;
  assign n49820 = n49702 ^ n49492;
  assign n49821 = n49699 & ~n49820;
  assign n49822 = n49821 ^ n49702;
  assign n49775 = n49486 ^ n46403;
  assign n49776 = n49489 ^ n49486;
  assign n49777 = ~n49775 & n49776;
  assign n49778 = n49777 ^ n46403;
  assign n49756 = n47779 ^ n47096;
  assign n49757 = n49756 ^ n48451;
  assign n49754 = n49138 ^ n49110;
  assign n49751 = n49485 ^ n49481;
  assign n49752 = n49482 & n49751;
  assign n49753 = n49752 ^ n49480;
  assign n49755 = n49754 ^ n49753;
  assign n49773 = n49757 ^ n49755;
  assign n49774 = n49773 ^ n46401;
  assign n49787 = n49778 ^ n49774;
  assign n49786 = ~n49478 & ~n49491;
  assign n49819 = n49787 ^ n49786;
  assign n49823 = n49822 ^ n49819;
  assign n49847 = n49826 ^ n49823;
  assign n49848 = n49847 ^ n49845;
  assign n49849 = ~n49846 & ~n49848;
  assign n49850 = n49849 ^ n49843;
  assign n49827 = n49826 ^ n49819;
  assign n49828 = n49823 & ~n49827;
  assign n49829 = n49828 ^ n49826;
  assign n49815 = n47747 ^ n39925;
  assign n49816 = n49815 ^ n44263;
  assign n49817 = n49816 ^ n1745;
  assign n49839 = n49829 ^ n49817;
  assign n49779 = n49778 ^ n49773;
  assign n49780 = ~n49774 & ~n49779;
  assign n49781 = n49780 ^ n46401;
  assign n49758 = n49757 ^ n49754;
  assign n49759 = ~n49755 & n49758;
  assign n49760 = n49759 ^ n49757;
  assign n49747 = n48443 ^ n47092;
  assign n49748 = n49747 ^ n47775;
  assign n49770 = n49760 ^ n49748;
  assign n49771 = n49770 ^ n49749;
  assign n49772 = n49771 ^ n46395;
  assign n49789 = n49781 ^ n49772;
  assign n49788 = ~n49786 & n49787;
  assign n49814 = n49789 ^ n49788;
  assign n49840 = n49839 ^ n49814;
  assign n49851 = n49850 ^ n49840;
  assign n49852 = n48909 ^ n48486;
  assign n49853 = n49852 ^ n47645;
  assign n49854 = n49853 ^ n49840;
  assign n49855 = ~n49851 & ~n49854;
  assign n49856 = n49855 ^ n49853;
  assign n49837 = n49218 ^ n48264;
  assign n49838 = n49837 ^ n47641;
  assign n49857 = n49856 ^ n49838;
  assign n49818 = n49817 ^ n49814;
  assign n49830 = n49829 ^ n49814;
  assign n49831 = n49818 & ~n49830;
  assign n49832 = n49831 ^ n49817;
  assign n49810 = n47768 ^ n39920;
  assign n49811 = n49810 ^ n44258;
  assign n49812 = n49811 ^ n38497;
  assign n49790 = n49788 & n49789;
  assign n49782 = n49781 ^ n49771;
  assign n49783 = n49772 & n49782;
  assign n49784 = n49783 ^ n46395;
  assign n49764 = n47657 ^ n46975;
  assign n49765 = n49764 ^ n48439;
  assign n49767 = n49766 ^ n49765;
  assign n49750 = n49749 ^ n49748;
  assign n49761 = n49760 ^ n49749;
  assign n49762 = n49750 & n49761;
  assign n49763 = n49762 ^ n49748;
  assign n49768 = n49767 ^ n49763;
  assign n49769 = n49768 ^ n46158;
  assign n49785 = n49784 ^ n49769;
  assign n49809 = n49790 ^ n49785;
  assign n49813 = n49812 ^ n49809;
  assign n49858 = n49832 ^ n49813;
  assign n49859 = n49858 ^ n49856;
  assign n49860 = ~n49857 & ~n49859;
  assign n49861 = n49860 ^ n49838;
  assign n49833 = n49832 ^ n49812;
  assign n49834 = ~n49813 & ~n49833;
  assign n49835 = n49834 ^ n49809;
  assign n49805 = n49766 ^ n49763;
  assign n49806 = ~n49767 & ~n49805;
  assign n49807 = n49806 ^ n49765;
  assign n49799 = n49784 ^ n49768;
  assign n49800 = ~n49769 & ~n49799;
  assign n49801 = n49800 ^ n46158;
  assign n49796 = n49147 ^ n49098;
  assign n49795 = n49063 ^ n47655;
  assign n49797 = n49796 ^ n49795;
  assign n49792 = n47741 ^ n39915;
  assign n49793 = n49792 ^ n44310;
  assign n49794 = n49793 ^ n38492;
  assign n49798 = n49797 ^ n49794;
  assign n49802 = n49801 ^ n49798;
  assign n49791 = ~n49785 & ~n49790;
  assign n49803 = n49802 ^ n49791;
  assign n49804 = n49803 ^ n48435;
  assign n49808 = n49807 ^ n49804;
  assign n49836 = n49835 ^ n49808;
  assign n49862 = n49861 ^ n49836;
  assign n49863 = n48904 ^ n47833;
  assign n49864 = n49863 ^ n48496;
  assign n49865 = n49864 ^ n49836;
  assign n49866 = ~n49862 & ~n49865;
  assign n49867 = n49866 ^ n49864;
  assign n49868 = n49867 ^ n49745;
  assign n49869 = ~n49746 & ~n49868;
  assign n49870 = n49869 ^ n49744;
  assign n49871 = n49870 ^ n49741;
  assign n49872 = n49742 & ~n49871;
  assign n49873 = n49872 ^ n49739;
  assign n49737 = n49612 ^ n49609;
  assign n49874 = n49873 ^ n49737;
  assign n49875 = n48891 ^ n47626;
  assign n49876 = n49875 ^ n48255;
  assign n49877 = n49876 ^ n49737;
  assign n49878 = ~n49874 & ~n49877;
  assign n49879 = n49878 ^ n49876;
  assign n49880 = n49879 ^ n49735;
  assign n49881 = ~n49736 & n49880;
  assign n49882 = n49881 ^ n49734;
  assign n49732 = n49619 ^ n49594;
  assign n49883 = n49882 ^ n49732;
  assign n49884 = n48886 ^ n47617;
  assign n49885 = n49884 ^ n48601;
  assign n49886 = n49885 ^ n49732;
  assign n49887 = n49883 & n49886;
  assign n49888 = n49887 ^ n49885;
  assign n49889 = n49888 ^ n49728;
  assign n49890 = n49731 & n49889;
  assign n49891 = n49890 ^ n49730;
  assign n49727 = n49629 ^ n49588;
  assign n49892 = n49891 ^ n49727;
  assign n49893 = n48664 ^ n47609;
  assign n49894 = n49893 ^ n48876;
  assign n49895 = n49894 ^ n49727;
  assign n49896 = ~n49892 & n49895;
  assign n49897 = n49896 ^ n49894;
  assign n49898 = n49897 ^ n49725;
  assign n49899 = ~n49726 & n49898;
  assign n49900 = n49899 ^ n49724;
  assign n49902 = n49901 ^ n49900;
  assign n49903 = n48879 ^ n47607;
  assign n49904 = n49903 ^ n48861;
  assign n49905 = n49904 ^ n49901;
  assign n49906 = ~n49902 & n49905;
  assign n49907 = n49906 ^ n49904;
  assign n49908 = n49907 ^ n49721;
  assign n49909 = ~n49722 & n49908;
  assign n49910 = n49909 ^ n49720;
  assign n49912 = n49911 ^ n49910;
  assign n49913 = n48852 ^ n47876;
  assign n49914 = n49913 ^ n48869;
  assign n49915 = n49914 ^ n49911;
  assign n49916 = n49912 & ~n49915;
  assign n49917 = n49916 ^ n49914;
  assign n49919 = n49918 ^ n49917;
  assign n49920 = n48862 ^ n47999;
  assign n49921 = n49920 ^ n48846;
  assign n49922 = n49921 ^ n49918;
  assign n49923 = ~n49919 & n49922;
  assign n49924 = n49923 ^ n49921;
  assign n49717 = n49649 ^ n49559;
  assign n49718 = n49717 ^ n49556;
  assign n49925 = n49924 ^ n49718;
  assign n49926 = n48855 ^ n48239;
  assign n49927 = n49926 ^ n48840;
  assign n49928 = n49927 ^ n49718;
  assign n49929 = n49925 & n49928;
  assign n49930 = n49929 ^ n49927;
  assign n49931 = n49930 ^ n49715;
  assign n49932 = n49716 & n49931;
  assign n49933 = n49932 ^ n49714;
  assign n49934 = n49933 ^ n49709;
  assign n49935 = n49712 & n49934;
  assign n49936 = n49935 ^ n49711;
  assign n49708 = n49662 ^ n49549;
  assign n49937 = n49936 ^ n49708;
  assign n49938 = n49449 ^ n48837;
  assign n49939 = n49938 ^ n48289;
  assign n49940 = n49939 ^ n49708;
  assign n49941 = n49937 & ~n49940;
  assign n49942 = n49941 ^ n49939;
  assign n50058 = n49944 ^ n49942;
  assign n50059 = n49947 & n50058;
  assign n50060 = n50059 ^ n49946;
  assign n50122 = n50061 ^ n50060;
  assign n50123 = ~n50064 & ~n50122;
  assign n50124 = n50123 ^ n50063;
  assign n50121 = n49671 ^ n49537;
  assign n50125 = n50124 ^ n50121;
  assign n50119 = n49754 ^ n48976;
  assign n50120 = n50119 ^ n48284;
  assign n50133 = n50121 ^ n50120;
  assign n50134 = n50125 & n50133;
  assign n50135 = n50134 ^ n50120;
  assign n50340 = n50136 ^ n50135;
  assign n50341 = ~n50139 & ~n50340;
  assign n50342 = n50341 ^ n50138;
  assign n50347 = n50346 ^ n50342;
  assign n50348 = n50347 ^ n47104;
  assign n50140 = n50139 ^ n50135;
  assign n50141 = n50140 ^ n46902;
  assign n50126 = n50125 ^ n50120;
  assign n50127 = n50126 ^ n47713;
  assign n50065 = n50064 ^ n50060;
  assign n50066 = n50065 ^ n47694;
  assign n49948 = n49947 ^ n49942;
  assign n49949 = n49948 ^ n47680;
  assign n49950 = n49939 ^ n49937;
  assign n49951 = n49950 ^ n47664;
  assign n49952 = n49933 ^ n49712;
  assign n49953 = n49952 ^ n47206;
  assign n49954 = n49930 ^ n49714;
  assign n49955 = n49954 ^ n49715;
  assign n49956 = n49955 ^ n46907;
  assign n49957 = n49927 ^ n49925;
  assign n49958 = n49957 ^ n46910;
  assign n49959 = n49921 ^ n49919;
  assign n49960 = n49959 ^ n46915;
  assign n49961 = n49914 ^ n49912;
  assign n49962 = n49961 ^ n47187;
  assign n49966 = n49897 ^ n49724;
  assign n49967 = n49966 ^ n49725;
  assign n49968 = n49967 ^ n46926;
  assign n49969 = n49894 ^ n49892;
  assign n49970 = n49969 ^ n46930;
  assign n49971 = n49888 ^ n49731;
  assign n49972 = n49971 ^ n46935;
  assign n49973 = n49885 ^ n49883;
  assign n49974 = n49973 ^ n46936;
  assign n49975 = n49879 ^ n49736;
  assign n49976 = n49975 ^ n46940;
  assign n49977 = n49876 ^ n49874;
  assign n49978 = n49977 ^ n46941;
  assign n49979 = n49870 ^ n49742;
  assign n49980 = n49979 ^ n46945;
  assign n49981 = n49867 ^ n49746;
  assign n49982 = n49981 ^ n46950;
  assign n49984 = n49853 ^ n49851;
  assign n49985 = n49984 ^ n46957;
  assign n49986 = n49842 ^ n49703;
  assign n49987 = ~n46968 & ~n49986;
  assign n49988 = n49987 ^ n46962;
  assign n49989 = n49847 ^ n49846;
  assign n49990 = n49989 ^ n49987;
  assign n49991 = n49988 & ~n49990;
  assign n49992 = n49991 ^ n46962;
  assign n49993 = n49992 ^ n49984;
  assign n49994 = n49985 & n49993;
  assign n49995 = n49994 ^ n46957;
  assign n49983 = n49858 ^ n49857;
  assign n49996 = n49995 ^ n49983;
  assign n49997 = n49983 ^ n46956;
  assign n49998 = n49996 & ~n49997;
  assign n49999 = n49998 ^ n46956;
  assign n50000 = n49999 ^ n46955;
  assign n50001 = n49864 ^ n49862;
  assign n50002 = n50001 ^ n49999;
  assign n50003 = n50000 & ~n50002;
  assign n50004 = n50003 ^ n46955;
  assign n50005 = n50004 ^ n49981;
  assign n50006 = ~n49982 & n50005;
  assign n50007 = n50006 ^ n46950;
  assign n50008 = n50007 ^ n49979;
  assign n50009 = n49980 & n50008;
  assign n50010 = n50009 ^ n46945;
  assign n50011 = n50010 ^ n49977;
  assign n50012 = n49978 & n50011;
  assign n50013 = n50012 ^ n46941;
  assign n50014 = n50013 ^ n49975;
  assign n50015 = n49976 & n50014;
  assign n50016 = n50015 ^ n46940;
  assign n50017 = n50016 ^ n49973;
  assign n50018 = n49974 & n50017;
  assign n50019 = n50018 ^ n46936;
  assign n50020 = n50019 ^ n49971;
  assign n50021 = ~n49972 & n50020;
  assign n50022 = n50021 ^ n46935;
  assign n50023 = n50022 ^ n49969;
  assign n50024 = ~n49970 & ~n50023;
  assign n50025 = n50024 ^ n46930;
  assign n50026 = n50025 ^ n49967;
  assign n50027 = ~n49968 & ~n50026;
  assign n50028 = n50027 ^ n46926;
  assign n49965 = n49904 ^ n49902;
  assign n50029 = n50028 ^ n49965;
  assign n50030 = n49965 ^ n46922;
  assign n50031 = ~n50029 & ~n50030;
  assign n50032 = n50031 ^ n46922;
  assign n49963 = n49907 ^ n49720;
  assign n49964 = n49963 ^ n49721;
  assign n50033 = n50032 ^ n49964;
  assign n50034 = n49964 ^ n46917;
  assign n50035 = ~n50033 & ~n50034;
  assign n50036 = n50035 ^ n46917;
  assign n50037 = n50036 ^ n49961;
  assign n50038 = n49962 & n50037;
  assign n50039 = n50038 ^ n47187;
  assign n50040 = n50039 ^ n49959;
  assign n50041 = n49960 & n50040;
  assign n50042 = n50041 ^ n46915;
  assign n50043 = n50042 ^ n49957;
  assign n50044 = n49958 & ~n50043;
  assign n50045 = n50044 ^ n46910;
  assign n50046 = n50045 ^ n49955;
  assign n50047 = n49956 & n50046;
  assign n50048 = n50047 ^ n46907;
  assign n50049 = n50048 ^ n49952;
  assign n50050 = ~n49953 & n50049;
  assign n50051 = n50050 ^ n47206;
  assign n50052 = n50051 ^ n49950;
  assign n50053 = ~n49951 & n50052;
  assign n50054 = n50053 ^ n47664;
  assign n50055 = n50054 ^ n49948;
  assign n50056 = ~n49949 & ~n50055;
  assign n50057 = n50056 ^ n47680;
  assign n50116 = n50065 ^ n50057;
  assign n50117 = n50066 & n50116;
  assign n50118 = n50117 ^ n47694;
  assign n50130 = n50126 ^ n50118;
  assign n50131 = ~n50127 & ~n50130;
  assign n50132 = n50131 ^ n47713;
  assign n50337 = n50140 ^ n50132;
  assign n50338 = ~n50141 & n50337;
  assign n50339 = n50338 ^ n46902;
  assign n50349 = n50348 ^ n50339;
  assign n50067 = n50066 ^ n50057;
  assign n50068 = n50051 ^ n49951;
  assign n50069 = n50036 ^ n47187;
  assign n50070 = n50069 ^ n49961;
  assign n50071 = n50025 ^ n49968;
  assign n50072 = n49989 ^ n49988;
  assign n50073 = n49992 ^ n49985;
  assign n50074 = ~n50072 & ~n50073;
  assign n50075 = n49996 ^ n46956;
  assign n50076 = ~n50074 & n50075;
  assign n50077 = n50001 ^ n46955;
  assign n50078 = n50077 ^ n49999;
  assign n50079 = ~n50076 & n50078;
  assign n50080 = n50004 ^ n49982;
  assign n50081 = ~n50079 & n50080;
  assign n50082 = n50007 ^ n49980;
  assign n50083 = ~n50081 & n50082;
  assign n50084 = n50010 ^ n46941;
  assign n50085 = n50084 ^ n49977;
  assign n50086 = n50083 & ~n50085;
  assign n50087 = n50013 ^ n49976;
  assign n50088 = n50086 & n50087;
  assign n50089 = n50016 ^ n46936;
  assign n50090 = n50089 ^ n49973;
  assign n50091 = ~n50088 & n50090;
  assign n50092 = n50019 ^ n49972;
  assign n50093 = n50091 & n50092;
  assign n50094 = n50022 ^ n46930;
  assign n50095 = n50094 ^ n49969;
  assign n50096 = n50093 & n50095;
  assign n50097 = ~n50071 & n50096;
  assign n50098 = n50029 ^ n46922;
  assign n50099 = n50097 & n50098;
  assign n50100 = n50033 ^ n46917;
  assign n50101 = ~n50099 & n50100;
  assign n50102 = n50070 & n50101;
  assign n50103 = n50039 ^ n49960;
  assign n50104 = ~n50102 & n50103;
  assign n50105 = n50042 ^ n46910;
  assign n50106 = n50105 ^ n49957;
  assign n50107 = ~n50104 & n50106;
  assign n50108 = n50045 ^ n49956;
  assign n50109 = ~n50107 & ~n50108;
  assign n50110 = n50048 ^ n49953;
  assign n50111 = n50109 & ~n50110;
  assign n50112 = ~n50068 & n50111;
  assign n50113 = n50054 ^ n49949;
  assign n50114 = ~n50112 & n50113;
  assign n50115 = n50067 & n50114;
  assign n50128 = n50127 ^ n50118;
  assign n50129 = ~n50115 & ~n50128;
  assign n50142 = n50141 ^ n50132;
  assign n50336 = n50129 & n50142;
  assign n50350 = n50349 ^ n50336;
  assign n50333 = n48232 ^ n40737;
  assign n50334 = n50333 ^ n3119;
  assign n50335 = n50334 ^ n2828;
  assign n50351 = n50350 ^ n50335;
  assign n50143 = n50142 ^ n50129;
  assign n49705 = n47602 ^ n40742;
  assign n49706 = n49705 ^ n2738;
  assign n49707 = n49706 ^ n3117;
  assign n50144 = n50143 ^ n49707;
  assign n50148 = n50128 ^ n50115;
  assign n50145 = n48053 ^ n3095;
  assign n50146 = n50145 ^ n44979;
  assign n50147 = n50146 ^ n2730;
  assign n50149 = n50148 ^ n50147;
  assign n50154 = n50113 ^ n50112;
  assign n50151 = n48063 ^ n40784;
  assign n50152 = n50151 ^ n44956;
  assign n50153 = n50152 ^ n39301;
  assign n50155 = n50154 ^ n50153;
  assign n50159 = n50111 ^ n50068;
  assign n50156 = n48067 ^ n40752;
  assign n50157 = n50156 ^ n44966;
  assign n50158 = n50157 ^ n39231;
  assign n50160 = n50159 ^ n50158;
  assign n50165 = n50108 ^ n50107;
  assign n50162 = n48073 ^ n40762;
  assign n50163 = n50162 ^ n1486;
  assign n50164 = n50163 ^ n39238;
  assign n50166 = n50165 ^ n50164;
  assign n50171 = n50103 ^ n50102;
  assign n50168 = n48080 ^ n1264;
  assign n50169 = n50168 ^ n44552;
  assign n50170 = n50169 ^ n1460;
  assign n50172 = n50171 ^ n50170;
  assign n50176 = n50101 ^ n50070;
  assign n50173 = n48085 ^ n1246;
  assign n50174 = n50173 ^ n44557;
  assign n50175 = n50174 ^ n39275;
  assign n50177 = n50176 ^ n50175;
  assign n50179 = n48091 ^ n3341;
  assign n50180 = n50179 ^ n44562;
  assign n50181 = n50180 ^ n39247;
  assign n50178 = n50100 ^ n50099;
  assign n50182 = n50181 ^ n50178;
  assign n50186 = n50098 ^ n50097;
  assign n50183 = n48095 ^ n40394;
  assign n50184 = n50183 ^ n44567;
  assign n50185 = n50184 ^ n39252;
  assign n50187 = n50186 ^ n50185;
  assign n50191 = n50096 ^ n50071;
  assign n50188 = n48100 ^ n40302;
  assign n50189 = n50188 ^ n44572;
  assign n50190 = n50189 ^ n39257;
  assign n50192 = n50191 ^ n50190;
  assign n50197 = n50092 ^ n50091;
  assign n50194 = n48110 ^ n40311;
  assign n50195 = n50194 ^ n44652;
  assign n50196 = n50195 ^ n38755;
  assign n50198 = n50197 ^ n50196;
  assign n50203 = n50087 ^ n50086;
  assign n50200 = n48120 ^ n40318;
  assign n50201 = n50200 ^ n44642;
  assign n50202 = n50201 ^ n38761;
  assign n50204 = n50203 ^ n50202;
  assign n50211 = n50082 ^ n50081;
  assign n50208 = n48130 ^ n40328;
  assign n50209 = n50208 ^ n44632;
  assign n50210 = n50209 ^ n38770;
  assign n50212 = n50211 ^ n50210;
  assign n50222 = n50075 ^ n50074;
  assign n50219 = n48145 ^ n40338;
  assign n50220 = n50219 ^ n44606;
  assign n50221 = n50220 ^ n38781;
  assign n50223 = n50222 ^ n50221;
  assign n50227 = n50073 ^ n50072;
  assign n50224 = n48153 ^ n40342;
  assign n50225 = n50224 ^ n44610;
  assign n50226 = n50225 ^ n38787;
  assign n50228 = n50227 ^ n50226;
  assign n50234 = n48149 ^ n40345;
  assign n50235 = n50234 ^ n44613;
  assign n50236 = n50235 ^ n2066;
  assign n50229 = n48381 ^ n40828;
  assign n50230 = n50229 ^ n1940;
  assign n50231 = n50230 ^ n39196;
  assign n50232 = n49986 ^ n46968;
  assign n50233 = n50231 & n50232;
  assign n50237 = n50236 ^ n50233;
  assign n50238 = n50233 ^ n50072;
  assign n50239 = n50237 & n50238;
  assign n50240 = n50239 ^ n50236;
  assign n50241 = n50240 ^ n50227;
  assign n50242 = ~n50228 & n50241;
  assign n50243 = n50242 ^ n50226;
  assign n50244 = n50243 ^ n50222;
  assign n50245 = ~n50223 & n50244;
  assign n50246 = n50245 ^ n50221;
  assign n50216 = n48140 ^ n40359;
  assign n50217 = n50216 ^ n44600;
  assign n50218 = n50217 ^ n38799;
  assign n50247 = n50246 ^ n50218;
  assign n50248 = n50078 ^ n50076;
  assign n50249 = n50248 ^ n50246;
  assign n50250 = n50247 & ~n50249;
  assign n50251 = n50250 ^ n50218;
  assign n50213 = n48135 ^ n40333;
  assign n50214 = n50213 ^ n44595;
  assign n50215 = n50214 ^ n38775;
  assign n50252 = n50251 ^ n50215;
  assign n50253 = n50080 ^ n50079;
  assign n50254 = n50253 ^ n50251;
  assign n50255 = n50252 & n50254;
  assign n50256 = n50255 ^ n50215;
  assign n50257 = n50256 ^ n50211;
  assign n50258 = n50212 & ~n50257;
  assign n50259 = n50258 ^ n50210;
  assign n50205 = n48125 ^ n40323;
  assign n50206 = n50205 ^ n44590;
  assign n50207 = n50206 ^ n38766;
  assign n50260 = n50259 ^ n50207;
  assign n50261 = n50085 ^ n50083;
  assign n50262 = n50261 ^ n50259;
  assign n50263 = n50260 & ~n50262;
  assign n50264 = n50263 ^ n50207;
  assign n50265 = n50264 ^ n50203;
  assign n50266 = ~n50204 & n50265;
  assign n50267 = n50266 ^ n50202;
  assign n50199 = n50090 ^ n50088;
  assign n50268 = n50267 ^ n50199;
  assign n50269 = n48116 ^ n40378;
  assign n50270 = n50269 ^ n44584;
  assign n50271 = n50270 ^ n38818;
  assign n50272 = n50271 ^ n50199;
  assign n50273 = n50268 & ~n50272;
  assign n50274 = n50273 ^ n50271;
  assign n50275 = n50274 ^ n50197;
  assign n50276 = n50198 & ~n50275;
  assign n50277 = n50276 ^ n50196;
  assign n50193 = n50095 ^ n50093;
  assign n50278 = n50277 ^ n50193;
  assign n50279 = n48105 ^ n40306;
  assign n50280 = n50279 ^ n44577;
  assign n50281 = n50280 ^ n788;
  assign n50282 = n50281 ^ n50193;
  assign n50283 = ~n50278 & n50282;
  assign n50284 = n50283 ^ n50281;
  assign n50285 = n50284 ^ n50191;
  assign n50286 = ~n50192 & n50285;
  assign n50287 = n50286 ^ n50190;
  assign n50288 = n50287 ^ n50186;
  assign n50289 = n50187 & ~n50288;
  assign n50290 = n50289 ^ n50185;
  assign n50291 = n50290 ^ n50178;
  assign n50292 = n50182 & ~n50291;
  assign n50293 = n50292 ^ n50181;
  assign n50294 = n50293 ^ n50176;
  assign n50295 = ~n50177 & n50294;
  assign n50296 = n50295 ^ n50175;
  assign n50297 = n50296 ^ n50171;
  assign n50298 = ~n50172 & n50297;
  assign n50299 = n50298 ^ n50170;
  assign n50167 = n50106 ^ n50104;
  assign n50300 = n50299 ^ n50167;
  assign n1441 = n1428 ^ n1362;
  assign n1469 = n1468 ^ n1441;
  assign n1476 = n1475 ^ n1469;
  assign n50301 = n50167 ^ n1476;
  assign n50302 = ~n50300 & n50301;
  assign n50303 = n50302 ^ n1476;
  assign n50304 = n50303 ^ n50165;
  assign n50305 = n50166 & ~n50304;
  assign n50306 = n50305 ^ n50164;
  assign n50161 = n50110 ^ n50109;
  assign n50307 = n50306 ^ n50161;
  assign n50308 = n48211 ^ n40757;
  assign n50309 = n50308 ^ n44117;
  assign n50310 = n50309 ^ n39291;
  assign n50311 = n50310 ^ n50161;
  assign n50312 = n50307 & ~n50311;
  assign n50313 = n50312 ^ n50310;
  assign n50314 = n50313 ^ n50159;
  assign n50315 = ~n50160 & n50314;
  assign n50316 = n50315 ^ n50158;
  assign n50317 = n50316 ^ n50154;
  assign n50318 = n50155 & ~n50317;
  assign n50319 = n50318 ^ n50153;
  assign n50150 = n50114 ^ n50067;
  assign n50320 = n50319 ^ n50150;
  assign n50321 = n48058 ^ n2624;
  assign n50322 = n50321 ^ n44951;
  assign n50323 = n50322 ^ n3203;
  assign n50324 = n50323 ^ n50150;
  assign n50325 = n50320 & ~n50324;
  assign n50326 = n50325 ^ n50323;
  assign n50327 = n50326 ^ n50148;
  assign n50328 = n50149 & ~n50327;
  assign n50329 = n50328 ^ n50147;
  assign n50330 = n50329 ^ n50143;
  assign n50331 = n50144 & ~n50330;
  assign n50332 = n50331 ^ n49707;
  assign n50486 = n50350 ^ n50332;
  assign n50487 = n50351 & ~n50486;
  assign n50488 = n50487 ^ n50335;
  assign n50419 = n50347 ^ n50339;
  assign n50420 = n50348 & n50419;
  assign n50421 = n50420 ^ n47104;
  assign n50391 = n48451 ^ n47793;
  assign n50392 = n50391 ^ n49796;
  assign n50387 = n50343 ^ n50342;
  assign n50388 = n50346 & ~n50387;
  assign n50389 = n50388 ^ n50345;
  assign n50386 = n49680 ^ n49522;
  assign n50390 = n50389 ^ n50386;
  assign n50417 = n50392 ^ n50390;
  assign n50418 = n50417 ^ n47111;
  assign n50434 = n50421 ^ n50418;
  assign n50433 = ~n50336 & n50349;
  assign n50485 = n50434 ^ n50433;
  assign n50489 = n50488 ^ n50485;
  assign n50490 = n48407 ^ n40803;
  assign n50491 = n50490 ^ n44943;
  assign n50492 = n50491 ^ n39320;
  assign n50493 = n50492 ^ n50485;
  assign n50494 = n50489 & ~n50493;
  assign n50495 = n50494 ^ n50492;
  assign n50435 = ~n50433 & n50434;
  assign n50422 = n50421 ^ n50417;
  assign n50423 = n50418 & ~n50422;
  assign n50424 = n50423 ^ n47111;
  assign n50397 = n48443 ^ n47781;
  assign n50398 = n50397 ^ n49178;
  assign n50393 = n50392 ^ n50386;
  assign n50394 = ~n50390 & n50393;
  assign n50395 = n50394 ^ n50392;
  assign n50384 = n49683 ^ n49515;
  assign n50385 = n50384 ^ n49516;
  assign n50396 = n50395 ^ n50385;
  assign n50415 = n50398 ^ n50396;
  assign n50416 = n50415 ^ n47101;
  assign n50432 = n50424 ^ n50416;
  assign n50480 = n50435 ^ n50432;
  assign n50484 = n50483 ^ n50480;
  assign n50522 = n50495 ^ n50484;
  assign n50643 = n50524 ^ n50522;
  assign n50644 = ~n47816 & n50643;
  assign n50645 = n50644 ^ n47648;
  assign n50525 = ~n50522 & ~n50524;
  assign n50519 = n49741 ^ n49218;
  assign n50520 = n50519 ^ n48269;
  assign n50646 = n50525 ^ n50520;
  assign n50496 = n50495 ^ n50480;
  assign n50497 = ~n50484 & n50496;
  assign n50498 = n50497 ^ n50483;
  assign n50425 = n50424 ^ n50415;
  assign n50426 = n50416 & ~n50425;
  assign n50427 = n50426 ^ n47101;
  assign n50403 = n48439 ^ n47779;
  assign n50404 = n50403 ^ n49185;
  assign n50399 = n50398 ^ n50385;
  assign n50400 = ~n50396 & n50399;
  assign n50401 = n50400 ^ n50398;
  assign n50383 = n49686 ^ n49512;
  assign n50402 = n50401 ^ n50383;
  assign n50413 = n50404 ^ n50402;
  assign n50414 = n50413 ^ n47096;
  assign n50437 = n50427 ^ n50414;
  assign n50436 = ~n50432 & ~n50435;
  assign n50478 = n50437 ^ n50436;
  assign n50475 = n48398 ^ n40726;
  assign n50476 = n50475 ^ n44999;
  assign n50477 = n50476 ^ n39212;
  assign n50479 = n50478 ^ n50477;
  assign n50518 = n50498 ^ n50479;
  assign n50647 = n50646 ^ n50518;
  assign n50648 = n50647 ^ n50644;
  assign n50649 = n50645 & ~n50648;
  assign n50650 = n50649 ^ n47648;
  assign n50530 = n49737 ^ n48904;
  assign n50531 = n50530 ^ n48486;
  assign n50521 = n50520 ^ n50518;
  assign n50526 = n50525 ^ n50518;
  assign n50527 = ~n50521 & n50526;
  assign n50528 = n50527 ^ n50525;
  assign n50499 = n50498 ^ n50478;
  assign n50500 = n50479 & ~n50499;
  assign n50501 = n50500 ^ n50477;
  assign n50438 = ~n50436 & ~n50437;
  assign n50428 = n50427 ^ n50413;
  assign n50429 = ~n50414 & n50428;
  assign n50430 = n50429 ^ n47096;
  assign n50409 = n48435 ^ n47775;
  assign n50410 = n50409 ^ n49190;
  assign n50405 = n50404 ^ n50383;
  assign n50406 = n50402 & ~n50405;
  assign n50407 = n50406 ^ n50404;
  assign n50382 = n49689 ^ n49507;
  assign n50408 = n50407 ^ n50382;
  assign n50411 = n50410 ^ n50408;
  assign n50412 = n50411 ^ n47092;
  assign n50431 = n50430 ^ n50412;
  assign n50473 = n50438 ^ n50431;
  assign n50470 = n48392 ^ n40816;
  assign n50471 = n50470 ^ n44932;
  assign n50472 = n50471 ^ n39207;
  assign n50474 = n50473 ^ n50472;
  assign n50517 = n50501 ^ n50474;
  assign n50529 = n50528 ^ n50517;
  assign n50642 = n50531 ^ n50529;
  assign n50651 = n50650 ^ n50642;
  assign n50652 = n50642 ^ n47645;
  assign n50653 = n50651 & ~n50652;
  assign n50654 = n50653 ^ n47645;
  assign n50532 = n50531 ^ n50517;
  assign n50533 = ~n50529 & ~n50532;
  assign n50534 = n50533 ^ n50531;
  assign n50514 = n49735 ^ n48900;
  assign n50515 = n50514 ^ n48264;
  assign n50506 = n48428 ^ n1802;
  assign n50507 = n50506 ^ n44927;
  assign n50508 = n50507 ^ n39202;
  assign n50502 = n50501 ^ n50473;
  assign n50503 = n50474 & ~n50502;
  assign n50504 = n50503 ^ n50472;
  assign n50449 = n50430 ^ n50411;
  assign n50450 = n50412 & n50449;
  assign n50451 = n50450 ^ n47092;
  assign n50443 = n50410 ^ n50382;
  assign n50444 = ~n50408 & ~n50443;
  assign n50445 = n50444 ^ n50410;
  assign n50442 = n49692 ^ n49502;
  assign n50446 = n50445 ^ n50442;
  assign n50440 = n48467 ^ n47657;
  assign n50441 = n50440 ^ n49171;
  assign n50447 = n50446 ^ n50441;
  assign n50448 = n50447 ^ n46975;
  assign n50452 = n50451 ^ n50448;
  assign n50439 = n50431 & n50438;
  assign n50469 = n50452 ^ n50439;
  assign n50505 = n50504 ^ n50469;
  assign n50513 = n50508 ^ n50505;
  assign n50516 = n50515 ^ n50513;
  assign n50640 = n50534 ^ n50516;
  assign n50641 = n50640 ^ n47641;
  assign n50721 = n50654 ^ n50641;
  assign n50718 = n50647 ^ n50645;
  assign n50719 = n50651 ^ n47645;
  assign n50720 = ~n50718 & n50719;
  assign n50817 = n50721 ^ n50720;
  assign n50814 = n48734 ^ n41040;
  assign n50815 = n50814 ^ n45378;
  assign n50816 = n50815 ^ n2352;
  assign n50818 = n50817 ^ n50816;
  assign n50822 = n50643 ^ n47816;
  assign n50823 = n49061 ^ n2013;
  assign n50824 = n50823 ^ n45639;
  assign n50825 = n50824 ^ n40102;
  assign n50826 = ~n50822 & n50825;
  assign n50819 = n48738 ^ n41044;
  assign n50820 = n50819 ^ n45381;
  assign n50821 = n50820 ^ n2185;
  assign n50827 = n50826 ^ n50821;
  assign n50828 = n50826 ^ n50718;
  assign n50829 = n50827 & n50828;
  assign n50830 = n50829 ^ n50821;
  assign n2160 = n2159 ^ n2111;
  assign n2194 = n2193 ^ n2160;
  assign n2204 = n2203 ^ n2194;
  assign n50831 = n50830 ^ n2204;
  assign n50832 = n50719 ^ n50718;
  assign n50833 = n50832 ^ n50830;
  assign n50834 = n50831 & ~n50833;
  assign n50835 = n50834 ^ n2204;
  assign n50836 = n50835 ^ n50817;
  assign n50837 = n50818 & ~n50836;
  assign n50838 = n50837 ^ n50816;
  assign n50722 = ~n50720 & ~n50721;
  assign n50655 = n50654 ^ n50640;
  assign n50656 = ~n50641 & n50655;
  assign n50657 = n50656 ^ n47641;
  assign n50539 = n49732 ^ n48895;
  assign n50540 = n50539 ^ n48496;
  assign n50535 = n50534 ^ n50513;
  assign n50536 = n50516 & n50535;
  assign n50537 = n50536 ^ n50515;
  assign n50509 = n50508 ^ n50469;
  assign n50510 = ~n50505 & n50509;
  assign n50511 = n50510 ^ n50508;
  assign n50462 = n50451 ^ n50447;
  assign n50463 = n50448 & n50462;
  assign n50464 = n50463 ^ n46975;
  assign n50465 = n50464 ^ n46973;
  assign n50460 = n49695 ^ n49497;
  assign n50456 = n50442 ^ n50441;
  assign n50457 = ~n50446 & ~n50456;
  assign n50458 = n50457 ^ n50441;
  assign n50454 = n48275 ^ n47655;
  assign n50455 = n50454 ^ n49167;
  assign n50459 = n50458 ^ n50455;
  assign n50461 = n50460 ^ n50459;
  assign n50466 = n50465 ^ n50461;
  assign n50453 = ~n50439 & n50452;
  assign n50467 = n50466 ^ n50453;
  assign n50379 = n48387 ^ n45012;
  assign n50380 = n50379 ^ n40717;
  assign n50381 = n50380 ^ n1932;
  assign n50468 = n50467 ^ n50381;
  assign n50512 = n50511 ^ n50468;
  assign n50538 = n50537 ^ n50512;
  assign n50638 = n50540 ^ n50538;
  assign n50639 = n50638 ^ n47833;
  assign n50717 = n50657 ^ n50639;
  assign n50812 = n50722 ^ n50717;
  assign n50809 = n48752 ^ n41036;
  assign n50810 = n50809 ^ n2363;
  assign n50811 = n50810 ^ n39423;
  assign n50813 = n50812 ^ n50811;
  assign n51262 = n50838 ^ n50813;
  assign n50969 = n50835 ^ n50818;
  assign n50967 = n49911 ^ n48882;
  assign n50363 = n50264 ^ n50202;
  assign n50364 = n50363 ^ n50203;
  assign n50968 = n50967 ^ n50364;
  assign n50970 = n50969 ^ n50968;
  assign n50576 = n50256 ^ n50210;
  assign n50577 = n50576 ^ n50211;
  assign n50975 = n50577 ^ n49237;
  assign n50976 = n50975 ^ n49901;
  assign n50973 = n50821 ^ n50718;
  assign n50974 = n50973 ^ n50826;
  assign n50977 = n50976 ^ n50974;
  assign n50568 = n50253 ^ n50215;
  assign n50569 = n50568 ^ n50251;
  assign n50979 = n50569 ^ n48891;
  assign n50980 = n50979 ^ n49725;
  assign n50978 = n50825 ^ n50822;
  assign n50981 = n50980 ^ n50978;
  assign n51209 = n49086 ^ n41429;
  assign n51210 = n51209 ^ n45650;
  assign n51211 = n51210 ^ n39920;
  assign n51029 = n49703 ^ n49190;
  assign n51030 = n51029 ^ n48443;
  assign n50987 = n50442 ^ n48448;
  assign n50988 = n50987 ^ n49178;
  assign n50986 = n50313 ^ n50160;
  assign n50989 = n50988 ^ n50986;
  assign n50991 = n50382 ^ n49796;
  assign n50992 = n50991 ^ n49066;
  assign n50990 = n50310 ^ n50307;
  assign n50993 = n50992 ^ n50990;
  assign n50995 = n50385 ^ n48250;
  assign n50996 = n50995 ^ n49749;
  assign n50944 = n50300 ^ n1476;
  assign n50997 = n50996 ^ n50944;
  assign n50998 = n50386 ^ n48833;
  assign n50999 = n50998 ^ n49754;
  assign n50949 = n50296 ^ n50170;
  assign n50950 = n50949 ^ n50171;
  assign n51000 = n50999 ^ n50950;
  assign n50752 = n49467 ^ n48843;
  assign n50753 = n50752 ^ n50136;
  assign n50750 = n50290 ^ n50181;
  assign n50751 = n50750 ^ n50178;
  assign n50754 = n50753 ^ n50751;
  assign n50609 = n50061 ^ n48830;
  assign n50610 = n50609 ^ n48855;
  assign n50608 = n50284 ^ n50192;
  assign n50611 = n50610 ^ n50608;
  assign n50355 = n49944 ^ n48835;
  assign n50356 = n50355 ^ n48862;
  assign n50354 = n50281 ^ n50278;
  assign n50357 = n50356 ^ n50354;
  assign n50361 = n50271 ^ n50268;
  assign n50359 = n49709 ^ n48873;
  assign n50360 = n50359 ^ n48846;
  assign n50362 = n50361 ^ n50360;
  assign n50372 = n50236 ^ n50072;
  assign n50373 = n50372 ^ n50233;
  assign n50370 = n49727 ^ n49237;
  assign n50371 = n50370 ^ n48258;
  assign n50374 = n50373 ^ n50371;
  assign n50377 = n50232 ^ n50231;
  assign n50375 = n49728 ^ n48262;
  assign n50376 = n50375 ^ n48891;
  assign n50378 = n50377 ^ n50376;
  assign n50541 = n50540 ^ n50512;
  assign n50542 = n50538 & ~n50541;
  assign n50543 = n50542 ^ n50540;
  assign n50544 = n50543 ^ n50377;
  assign n50545 = ~n50378 & ~n50544;
  assign n50546 = n50545 ^ n50376;
  assign n50547 = n50546 ^ n50373;
  assign n50548 = ~n50374 & ~n50547;
  assign n50549 = n50548 ^ n50371;
  assign n50369 = n50240 ^ n50228;
  assign n50550 = n50549 ^ n50369;
  assign n50551 = n48886 ^ n48255;
  assign n50552 = n50551 ^ n49725;
  assign n50553 = n50552 ^ n50369;
  assign n50554 = n50550 & n50553;
  assign n50555 = n50554 ^ n50552;
  assign n50367 = n50243 ^ n50221;
  assign n50368 = n50367 ^ n50222;
  assign n50556 = n50555 ^ n50368;
  assign n50557 = n48882 ^ n48518;
  assign n50558 = n50557 ^ n49901;
  assign n50559 = n50558 ^ n50368;
  assign n50560 = ~n50556 & ~n50559;
  assign n50561 = n50560 ^ n50558;
  assign n50366 = n50248 ^ n50247;
  assign n50562 = n50561 ^ n50366;
  assign n50563 = n48876 ^ n48601;
  assign n50564 = n50563 ^ n49721;
  assign n50565 = n50564 ^ n50366;
  assign n50566 = ~n50562 & n50565;
  assign n50567 = n50566 ^ n50564;
  assign n50570 = n50569 ^ n50567;
  assign n50571 = n49911 ^ n48645;
  assign n50572 = n50571 ^ n48867;
  assign n50573 = n50572 ^ n50569;
  assign n50574 = n50570 & n50573;
  assign n50575 = n50574 ^ n50572;
  assign n50578 = n50577 ^ n50575;
  assign n50579 = n49918 ^ n48664;
  assign n50580 = n50579 ^ n48861;
  assign n50581 = n50580 ^ n50577;
  assign n50582 = n50578 & ~n50581;
  assign n50583 = n50582 ^ n50580;
  assign n50365 = n50261 ^ n50260;
  assign n50584 = n50583 ^ n50365;
  assign n50585 = n48858 ^ n48821;
  assign n50586 = n50585 ^ n49718;
  assign n50587 = n50586 ^ n50365;
  assign n50588 = n50584 & n50587;
  assign n50589 = n50588 ^ n50586;
  assign n50590 = n50589 ^ n50364;
  assign n50591 = n48879 ^ n48852;
  assign n50592 = n50591 ^ n49715;
  assign n50593 = n50592 ^ n50364;
  assign n50594 = n50590 & ~n50593;
  assign n50595 = n50594 ^ n50592;
  assign n50596 = n50595 ^ n50361;
  assign n50597 = ~n50362 & n50596;
  assign n50598 = n50597 ^ n50360;
  assign n50358 = n50274 ^ n50198;
  assign n50599 = n50598 ^ n50358;
  assign n50600 = n49708 ^ n48840;
  assign n50601 = n50600 ^ n48869;
  assign n50602 = n50601 ^ n50358;
  assign n50603 = ~n50599 & ~n50602;
  assign n50604 = n50603 ^ n50601;
  assign n50605 = n50604 ^ n50354;
  assign n50606 = n50357 & n50605;
  assign n50607 = n50606 ^ n50356;
  assign n50703 = n50608 ^ n50607;
  assign n50704 = ~n50611 & n50703;
  assign n50705 = n50704 ^ n50610;
  assign n50702 = n50287 ^ n50187;
  assign n50706 = n50705 ^ n50702;
  assign n50700 = n49449 ^ n48849;
  assign n50701 = n50700 ^ n50121;
  assign n50747 = n50702 ^ n50701;
  assign n50748 = ~n50706 & ~n50747;
  assign n50749 = n50748 ^ n50701;
  assign n50922 = n50751 ^ n50749;
  assign n50923 = n50754 & n50922;
  assign n50924 = n50923 ^ n50753;
  assign n50920 = n50293 ^ n50175;
  assign n50921 = n50920 ^ n50176;
  assign n50925 = n50924 ^ n50921;
  assign n50918 = n50343 ^ n48837;
  assign n50919 = n50918 ^ n49481;
  assign n51001 = n50921 ^ n50919;
  assign n51002 = n50925 & n51001;
  assign n51003 = n51002 ^ n50919;
  assign n51004 = n51003 ^ n50950;
  assign n51005 = ~n51000 & ~n51004;
  assign n51006 = n51005 ^ n50999;
  assign n51007 = n51006 ^ n50944;
  assign n51008 = ~n50997 & ~n51007;
  assign n51009 = n51008 ^ n50996;
  assign n50994 = n50303 ^ n50166;
  assign n51010 = n51009 ^ n50994;
  assign n51011 = n49766 ^ n48976;
  assign n51012 = n51011 ^ n50383;
  assign n51013 = n51012 ^ n50994;
  assign n51014 = n51010 & ~n51013;
  assign n51015 = n51014 ^ n51012;
  assign n51016 = n51015 ^ n50990;
  assign n51017 = n50993 & ~n51016;
  assign n51018 = n51017 ^ n50992;
  assign n51019 = n51018 ^ n50986;
  assign n51020 = ~n50989 & ~n51019;
  assign n51021 = n51020 ^ n50988;
  assign n50938 = n50316 ^ n50155;
  assign n51022 = n51021 ^ n50938;
  assign n51023 = n50460 ^ n48451;
  assign n51024 = n51023 ^ n49185;
  assign n51025 = n51024 ^ n50938;
  assign n51026 = ~n51022 & ~n51025;
  assign n51027 = n51026 ^ n51024;
  assign n50985 = n50323 ^ n50320;
  assign n51028 = n51027 ^ n50985;
  assign n51053 = n51030 ^ n51028;
  assign n51054 = n51053 ^ n47781;
  assign n51055 = n51024 ^ n51022;
  assign n51056 = n51055 ^ n47793;
  assign n51057 = n51018 ^ n50989;
  assign n51058 = n51057 ^ n47785;
  assign n51059 = n51015 ^ n50993;
  assign n51060 = n51059 ^ n47598;
  assign n51061 = n51012 ^ n51010;
  assign n51062 = n51061 ^ n48284;
  assign n51063 = n51006 ^ n50997;
  assign n51064 = n51063 ^ n48318;
  assign n51065 = n51003 ^ n51000;
  assign n51066 = n51065 ^ n48311;
  assign n50926 = n50925 ^ n50919;
  assign n50927 = n50926 ^ n48289;
  assign n50755 = n50754 ^ n50749;
  assign n50756 = n50755 ^ n48293;
  assign n50707 = n50706 ^ n50701;
  assign n50708 = n50707 ^ n48297;
  assign n50612 = n50611 ^ n50607;
  assign n50613 = n50612 ^ n48239;
  assign n50614 = n50604 ^ n50357;
  assign n50615 = n50614 ^ n47999;
  assign n50616 = n50601 ^ n50599;
  assign n50617 = n50616 ^ n47876;
  assign n50618 = n50595 ^ n50362;
  assign n50619 = n50618 ^ n47603;
  assign n50620 = n50592 ^ n50590;
  assign n50621 = n50620 ^ n47607;
  assign n50622 = n50586 ^ n50584;
  assign n50623 = n50622 ^ n47608;
  assign n50624 = n50580 ^ n50578;
  assign n50625 = n50624 ^ n47609;
  assign n50626 = n50572 ^ n50570;
  assign n50627 = n50626 ^ n47613;
  assign n50628 = n50564 ^ n50562;
  assign n50629 = n50628 ^ n47617;
  assign n50630 = n50558 ^ n50556;
  assign n50631 = n50630 ^ n47621;
  assign n50632 = n50552 ^ n50550;
  assign n50633 = n50632 ^ n47626;
  assign n50634 = n50546 ^ n50374;
  assign n50635 = n50634 ^ n47632;
  assign n50636 = n50543 ^ n50378;
  assign n50637 = n50636 ^ n47634;
  assign n50658 = n50657 ^ n50638;
  assign n50659 = ~n50639 & n50658;
  assign n50660 = n50659 ^ n47833;
  assign n50661 = n50660 ^ n50636;
  assign n50662 = n50637 & n50661;
  assign n50663 = n50662 ^ n47634;
  assign n50664 = n50663 ^ n50634;
  assign n50665 = n50635 & n50664;
  assign n50666 = n50665 ^ n47632;
  assign n50667 = n50666 ^ n50632;
  assign n50668 = ~n50633 & ~n50667;
  assign n50669 = n50668 ^ n47626;
  assign n50670 = n50669 ^ n50630;
  assign n50671 = ~n50631 & n50670;
  assign n50672 = n50671 ^ n47621;
  assign n50673 = n50672 ^ n50628;
  assign n50674 = n50629 & n50673;
  assign n50675 = n50674 ^ n47617;
  assign n50676 = n50675 ^ n50626;
  assign n50677 = ~n50627 & ~n50676;
  assign n50678 = n50677 ^ n47613;
  assign n50679 = n50678 ^ n50624;
  assign n50680 = ~n50625 & n50679;
  assign n50681 = n50680 ^ n47609;
  assign n50682 = n50681 ^ n50622;
  assign n50683 = n50623 & ~n50682;
  assign n50684 = n50683 ^ n47608;
  assign n50685 = n50684 ^ n50620;
  assign n50686 = n50621 & ~n50685;
  assign n50687 = n50686 ^ n47607;
  assign n50688 = n50687 ^ n50618;
  assign n50689 = n50619 & ~n50688;
  assign n50690 = n50689 ^ n47603;
  assign n50691 = n50690 ^ n50616;
  assign n50692 = ~n50617 & ~n50691;
  assign n50693 = n50692 ^ n47876;
  assign n50694 = n50693 ^ n50614;
  assign n50695 = n50615 & n50694;
  assign n50696 = n50695 ^ n47999;
  assign n50697 = n50696 ^ n50612;
  assign n50698 = n50613 & ~n50697;
  assign n50699 = n50698 ^ n48239;
  assign n50744 = n50707 ^ n50699;
  assign n50745 = ~n50708 & ~n50744;
  assign n50746 = n50745 ^ n48297;
  assign n50915 = n50755 ^ n50746;
  assign n50916 = ~n50756 & n50915;
  assign n50917 = n50916 ^ n48293;
  assign n51067 = n50926 ^ n50917;
  assign n51068 = ~n50927 & ~n51067;
  assign n51069 = n51068 ^ n48289;
  assign n51070 = n51069 ^ n51065;
  assign n51071 = ~n51066 & n51070;
  assign n51072 = n51071 ^ n48311;
  assign n51073 = n51072 ^ n51063;
  assign n51074 = ~n51064 & ~n51073;
  assign n51075 = n51074 ^ n48318;
  assign n51076 = n51075 ^ n51061;
  assign n51077 = n51062 & ~n51076;
  assign n51078 = n51077 ^ n48284;
  assign n51079 = n51078 ^ n51059;
  assign n51080 = n51060 & n51079;
  assign n51081 = n51080 ^ n47598;
  assign n51082 = n51081 ^ n51057;
  assign n51083 = ~n51058 & n51082;
  assign n51084 = n51083 ^ n47785;
  assign n51085 = n51084 ^ n51055;
  assign n51086 = n51056 & ~n51085;
  assign n51087 = n51086 ^ n47793;
  assign n51088 = n51087 ^ n51053;
  assign n51089 = n51054 & n51088;
  assign n51090 = n51089 ^ n47781;
  assign n51035 = n49847 ^ n49171;
  assign n51036 = n51035 ^ n48439;
  assign n51031 = n51030 ^ n50985;
  assign n51032 = ~n51028 & ~n51031;
  assign n51033 = n51032 ^ n51030;
  assign n50984 = n50326 ^ n50149;
  assign n51034 = n51033 ^ n50984;
  assign n51051 = n51036 ^ n51034;
  assign n51052 = n51051 ^ n47779;
  assign n51099 = n51090 ^ n51052;
  assign n51100 = n51084 ^ n51056;
  assign n51101 = n51072 ^ n51064;
  assign n50709 = n50708 ^ n50699;
  assign n50710 = n50696 ^ n50613;
  assign n50711 = n50684 ^ n50621;
  assign n50712 = n50678 ^ n50625;
  assign n50713 = n50669 ^ n50631;
  assign n50714 = n50666 ^ n50633;
  assign n50715 = n50663 ^ n50635;
  assign n50716 = n50660 ^ n50637;
  assign n50723 = n50717 & ~n50722;
  assign n50724 = n50716 & ~n50723;
  assign n50725 = n50715 & ~n50724;
  assign n50726 = n50714 & n50725;
  assign n50727 = ~n50713 & n50726;
  assign n50728 = n50672 ^ n50629;
  assign n50729 = ~n50727 & ~n50728;
  assign n50730 = n50675 ^ n50627;
  assign n50731 = n50729 & ~n50730;
  assign n50732 = n50712 & n50731;
  assign n50733 = n50681 ^ n50623;
  assign n50734 = n50732 & ~n50733;
  assign n50735 = ~n50711 & n50734;
  assign n50736 = n50687 ^ n50619;
  assign n50737 = ~n50735 & n50736;
  assign n50738 = n50690 ^ n50617;
  assign n50739 = n50737 & ~n50738;
  assign n50740 = n50693 ^ n50615;
  assign n50741 = ~n50739 & n50740;
  assign n50742 = n50710 & ~n50741;
  assign n50743 = n50709 & ~n50742;
  assign n50757 = n50756 ^ n50746;
  assign n50914 = n50743 & ~n50757;
  assign n50928 = n50927 ^ n50917;
  assign n51102 = n50914 & ~n50928;
  assign n51103 = n51069 ^ n51066;
  assign n51104 = ~n51102 & ~n51103;
  assign n51105 = ~n51101 & n51104;
  assign n51106 = n51075 ^ n51062;
  assign n51107 = ~n51105 & n51106;
  assign n51108 = n51078 ^ n51060;
  assign n51109 = n51107 & n51108;
  assign n51110 = n51081 ^ n51058;
  assign n51111 = ~n51109 & ~n51110;
  assign n51112 = ~n51100 & ~n51111;
  assign n51113 = n51087 ^ n51054;
  assign n51114 = ~n51112 & n51113;
  assign n51115 = n51099 & ~n51114;
  assign n51091 = n51090 ^ n51051;
  assign n51092 = n51052 & ~n51091;
  assign n51093 = n51092 ^ n47779;
  assign n51041 = n49167 ^ n48435;
  assign n51042 = n51041 ^ n49840;
  assign n51037 = n51036 ^ n50984;
  assign n51038 = ~n51034 & n51037;
  assign n51039 = n51038 ^ n51036;
  assign n50933 = n50329 ^ n50144;
  assign n51040 = n51039 ^ n50933;
  assign n51049 = n51042 ^ n51040;
  assign n51050 = n51049 ^ n47775;
  assign n51098 = n51093 ^ n51050;
  assign n51139 = n51115 ^ n51098;
  assign n51136 = n49157 ^ n41433;
  assign n51137 = n51136 ^ n45655;
  assign n51138 = n51137 ^ n39925;
  assign n51140 = n51139 ^ n51138;
  assign n51145 = n51113 ^ n51112;
  assign n51142 = n49096 ^ n41444;
  assign n51143 = n51142 ^ n45665;
  assign n51144 = n51143 ^ n39930;
  assign n51146 = n51145 ^ n51144;
  assign n51147 = n51111 ^ n51100;
  assign n2895 = n2894 ^ n2870;
  assign n2932 = n2931 ^ n2895;
  assign n2939 = n2938 ^ n2932;
  assign n51148 = n51147 ^ n2939;
  assign n51152 = n51110 ^ n51109;
  assign n51149 = n49103 ^ n3135;
  assign n51150 = n51149 ^ n3239;
  assign n51151 = n51150 ^ n2922;
  assign n51153 = n51152 ^ n51151;
  assign n51158 = n51106 ^ n51105;
  assign n51155 = n49113 ^ n3215;
  assign n51156 = n51155 ^ n45469;
  assign n51157 = n51156 ^ n39940;
  assign n51159 = n51158 ^ n51157;
  assign n51164 = n51103 ^ n51102;
  assign n51161 = n49124 ^ n41460;
  assign n51162 = n51161 ^ n45459;
  assign n51163 = n51162 ^ n40060;
  assign n51165 = n51164 ^ n51163;
  assign n50929 = n50928 ^ n50914;
  assign n50911 = n48811 ^ n41510;
  assign n50912 = n50911 ^ n45311;
  assign n50913 = n50912 ^ n39950;
  assign n50930 = n50929 ^ n50913;
  assign n50762 = n50742 ^ n50709;
  assign n50759 = n48671 ^ n41471;
  assign n50760 = n50759 ^ n45322;
  assign n50761 = n50760 ^ n39956;
  assign n50763 = n50762 ^ n50761;
  assign n50768 = n50740 ^ n50739;
  assign n50765 = n48681 ^ n41478;
  assign n50766 = n50765 ^ n45331;
  assign n50767 = n50766 ^ n39967;
  assign n50769 = n50768 ^ n50767;
  assign n50773 = n50738 ^ n50737;
  assign n50770 = n48686 ^ n41487;
  assign n50771 = n50770 ^ n45334;
  assign n50772 = n50771 ^ n1124;
  assign n50774 = n50773 ^ n50772;
  assign n50778 = n50736 ^ n50735;
  assign n50775 = n48691 ^ n41096;
  assign n50776 = n50775 ^ n995;
  assign n50777 = n50776 ^ n39973;
  assign n50779 = n50778 ^ n50777;
  assign n50783 = n50734 ^ n50711;
  assign n50780 = n48696 ^ n41090;
  assign n50781 = n50780 ^ n45339;
  assign n50782 = n50781 ^ n984;
  assign n50784 = n50783 ^ n50782;
  assign n50787 = n48781 ^ n41005;
  assign n50788 = n50787 ^ n45421;
  assign n50789 = n50788 ^ n39985;
  assign n50786 = n50731 ^ n50712;
  assign n50790 = n50789 ^ n50786;
  assign n50792 = n48774 ^ n41010;
  assign n50793 = n50792 ^ n45351;
  assign n50794 = n50793 ^ n39990;
  assign n50791 = n50730 ^ n50729;
  assign n50795 = n50794 ^ n50791;
  assign n50800 = n50726 ^ n50713;
  assign n50797 = n48714 ^ n41016;
  assign n50798 = n50797 ^ n45360;
  assign n50799 = n50798 ^ n39999;
  assign n50801 = n50800 ^ n50799;
  assign n50806 = n50724 ^ n50715;
  assign n50803 = n48724 ^ n41025;
  assign n50804 = n50803 ^ n45402;
  assign n50805 = n50804 ^ n39432;
  assign n50807 = n50806 ^ n50805;
  assign n50839 = n50838 ^ n50812;
  assign n50840 = n50813 & ~n50839;
  assign n50841 = n50840 ^ n50811;
  assign n50808 = n50723 ^ n50716;
  assign n50842 = n50841 ^ n50808;
  assign n50843 = n48729 ^ n41031;
  assign n50844 = n50843 ^ n45372;
  assign n50845 = n50844 ^ n39406;
  assign n50846 = n50845 ^ n50808;
  assign n50847 = n50842 & ~n50846;
  assign n50848 = n50847 ^ n50845;
  assign n50849 = n50848 ^ n50806;
  assign n50850 = n50807 & ~n50849;
  assign n50851 = n50850 ^ n50805;
  assign n50802 = n50725 ^ n50714;
  assign n50852 = n50851 ^ n50802;
  assign n50853 = n48718 ^ n41020;
  assign n50854 = n50853 ^ n45365;
  assign n50855 = n50854 ^ n40004;
  assign n50856 = n50855 ^ n50802;
  assign n50857 = n50852 & ~n50856;
  assign n50858 = n50857 ^ n50855;
  assign n50859 = n50858 ^ n50800;
  assign n50860 = n50801 & ~n50859;
  assign n50861 = n50860 ^ n50799;
  assign n50796 = n50728 ^ n50727;
  assign n50862 = n50861 ^ n50796;
  assign n50863 = n48709 ^ n41073;
  assign n50864 = n50863 ^ n45355;
  assign n50865 = n50864 ^ n39995;
  assign n50866 = n50865 ^ n50796;
  assign n50867 = ~n50862 & n50866;
  assign n50868 = n50867 ^ n50865;
  assign n50869 = n50868 ^ n50791;
  assign n50870 = ~n50795 & n50869;
  assign n50871 = n50870 ^ n50794;
  assign n50872 = n50871 ^ n50786;
  assign n50873 = n50790 & ~n50872;
  assign n50874 = n50873 ^ n50789;
  assign n50785 = n50733 ^ n50732;
  assign n50875 = n50874 ^ n50785;
  assign n50876 = n48702 ^ n848;
  assign n50877 = n50876 ^ n45345;
  assign n50878 = n50877 ^ n39980;
  assign n50879 = n50878 ^ n50785;
  assign n50880 = n50875 & ~n50879;
  assign n50881 = n50880 ^ n50878;
  assign n50882 = n50881 ^ n50783;
  assign n50883 = ~n50784 & n50882;
  assign n50884 = n50883 ^ n50782;
  assign n50885 = n50884 ^ n50778;
  assign n50886 = n50779 & ~n50885;
  assign n50887 = n50886 ^ n50777;
  assign n50888 = n50887 ^ n50773;
  assign n50889 = n50774 & ~n50888;
  assign n50890 = n50889 ^ n50772;
  assign n50891 = n50890 ^ n50768;
  assign n50892 = ~n50769 & n50891;
  assign n50893 = n50892 ^ n50767;
  assign n50764 = n50741 ^ n50710;
  assign n50894 = n50893 ^ n50764;
  assign n50895 = n48676 ^ n41497;
  assign n50896 = n50895 ^ n45326;
  assign n50897 = n50896 ^ n39962;
  assign n50898 = n50897 ^ n50764;
  assign n50899 = ~n50894 & n50898;
  assign n50900 = n50899 ^ n50897;
  assign n50901 = n50900 ^ n50762;
  assign n50902 = ~n50763 & n50901;
  assign n50903 = n50902 ^ n50761;
  assign n50758 = n50757 ^ n50743;
  assign n50904 = n50903 ^ n50758;
  assign n50905 = n48254 ^ n41467;
  assign n50906 = n50905 ^ n45316;
  assign n50907 = n50906 ^ n40050;
  assign n50908 = n50907 ^ n50758;
  assign n50909 = n50904 & ~n50908;
  assign n50910 = n50909 ^ n50907;
  assign n51166 = n50929 ^ n50910;
  assign n51167 = ~n50930 & n51166;
  assign n51168 = n51167 ^ n50913;
  assign n51169 = n51168 ^ n51164;
  assign n51170 = ~n51165 & n51169;
  assign n51171 = n51170 ^ n51163;
  assign n51160 = n51104 ^ n51101;
  assign n51172 = n51171 ^ n51160;
  assign n51173 = n49118 ^ n41455;
  assign n51174 = n51173 ^ n45305;
  assign n51175 = n51174 ^ n39944;
  assign n51176 = n51175 ^ n51160;
  assign n51177 = ~n51172 & n51176;
  assign n51178 = n51177 ^ n51175;
  assign n51179 = n51178 ^ n51158;
  assign n51180 = ~n51159 & n51179;
  assign n51181 = n51180 ^ n51157;
  assign n51154 = n51108 ^ n51107;
  assign n51182 = n51181 ^ n51154;
  assign n51183 = n49108 ^ n2796;
  assign n51184 = n51183 ^ n45300;
  assign n51185 = n51184 ^ n3237;
  assign n51186 = n51185 ^ n51154;
  assign n51187 = ~n51182 & n51186;
  assign n51188 = n51187 ^ n51185;
  assign n51189 = n51188 ^ n51152;
  assign n51190 = ~n51153 & n51189;
  assign n51191 = n51190 ^ n51151;
  assign n51192 = n51191 ^ n51147;
  assign n51193 = n51148 & ~n51192;
  assign n51194 = n51193 ^ n2939;
  assign n51195 = n51194 ^ n51145;
  assign n51196 = n51146 & ~n51195;
  assign n51197 = n51196 ^ n51144;
  assign n51141 = n51114 ^ n51099;
  assign n51198 = n51197 ^ n51141;
  assign n51199 = n49092 ^ n41439;
  assign n51200 = n51199 ^ n45660;
  assign n51201 = n51200 ^ n40087;
  assign n51202 = n51201 ^ n51141;
  assign n51203 = n51198 & ~n51202;
  assign n51204 = n51203 ^ n51201;
  assign n51205 = n51204 ^ n51139;
  assign n51206 = ~n51140 & n51205;
  assign n51207 = n51206 ^ n51138;
  assign n51116 = ~n51098 & n51115;
  assign n51094 = n51093 ^ n51049;
  assign n51095 = ~n51050 & ~n51094;
  assign n51096 = n51095 ^ n47775;
  assign n51043 = n51042 ^ n50933;
  assign n51044 = ~n51040 & n51043;
  assign n51045 = n51044 ^ n51042;
  assign n50352 = n50351 ^ n50332;
  assign n51046 = n51045 ^ n50352;
  assign n50982 = n49858 ^ n48467;
  assign n50983 = n50982 ^ n49200;
  assign n51047 = n51046 ^ n50983;
  assign n51048 = n51047 ^ n47657;
  assign n51097 = n51096 ^ n51048;
  assign n51135 = n51116 ^ n51097;
  assign n51208 = n51207 ^ n51135;
  assign n51218 = n51211 ^ n51208;
  assign n51216 = n49728 ^ n48900;
  assign n51217 = n51216 ^ n50368;
  assign n51219 = n51218 ^ n51217;
  assign n51225 = n50373 ^ n49735;
  assign n51226 = n51225 ^ n49218;
  assign n51221 = n51194 ^ n51146;
  assign n51222 = n49737 ^ n48909;
  assign n51223 = n51222 ^ n50377;
  assign n51224 = n51221 & ~n51223;
  assign n51227 = n51226 ^ n51224;
  assign n51228 = n51201 ^ n51198;
  assign n51229 = n51228 ^ n51226;
  assign n51230 = ~n51227 & ~n51229;
  assign n51231 = n51230 ^ n51224;
  assign n51220 = n51204 ^ n51140;
  assign n51232 = n51231 ^ n51220;
  assign n51233 = n49732 ^ n48904;
  assign n51234 = n51233 ^ n50369;
  assign n51235 = n51234 ^ n51220;
  assign n51236 = n51232 & ~n51235;
  assign n51237 = n51236 ^ n51234;
  assign n51238 = n51237 ^ n51218;
  assign n51239 = ~n51219 & n51238;
  assign n51240 = n51239 ^ n51217;
  assign n51212 = n51211 ^ n51135;
  assign n51213 = n51208 & ~n51212;
  assign n51214 = n51213 ^ n51211;
  assign n51130 = n51096 ^ n51047;
  assign n51131 = ~n51048 & ~n51130;
  assign n51132 = n51131 ^ n47657;
  assign n51126 = n50983 ^ n50352;
  assign n51127 = ~n51046 & ~n51126;
  assign n51128 = n51127 ^ n50983;
  assign n51120 = n49080 ^ n41424;
  assign n51121 = n51120 ^ n45645;
  assign n51122 = n51121 ^ n39915;
  assign n51123 = n51122 ^ n50454;
  assign n51119 = n50492 ^ n50489;
  assign n51124 = n51123 ^ n51119;
  assign n51118 = n49836 ^ n49208;
  assign n51125 = n51124 ^ n51118;
  assign n51129 = n51128 ^ n51125;
  assign n51133 = n51132 ^ n51129;
  assign n51117 = ~n51097 & ~n51116;
  assign n51134 = n51133 ^ n51117;
  assign n51215 = n51214 ^ n51134;
  assign n51241 = n51240 ^ n51215;
  assign n51242 = n49727 ^ n48895;
  assign n51243 = n51242 ^ n50366;
  assign n51244 = n51243 ^ n51215;
  assign n51245 = n51241 & n51244;
  assign n51246 = n51245 ^ n51243;
  assign n51247 = n51246 ^ n50978;
  assign n51248 = ~n50981 & ~n51247;
  assign n51249 = n51248 ^ n50980;
  assign n51250 = n51249 ^ n50974;
  assign n51251 = ~n50977 & n51250;
  assign n51252 = n51251 ^ n50976;
  assign n50971 = n50832 ^ n2204;
  assign n50972 = n50971 ^ n50830;
  assign n51253 = n51252 ^ n50972;
  assign n51254 = n49721 ^ n48886;
  assign n51255 = n51254 ^ n50365;
  assign n51256 = n51255 ^ n50972;
  assign n51257 = ~n51253 & n51256;
  assign n51258 = n51257 ^ n51255;
  assign n51259 = n51258 ^ n50969;
  assign n51260 = ~n50970 & ~n51259;
  assign n51261 = n51260 ^ n50968;
  assign n51263 = n51262 ^ n51261;
  assign n51264 = n50361 ^ n48876;
  assign n51265 = n51264 ^ n49918;
  assign n51266 = n51265 ^ n51262;
  assign n51267 = n51263 & n51266;
  assign n51268 = n51267 ^ n51265;
  assign n50965 = n50845 ^ n50842;
  assign n50963 = n49718 ^ n48867;
  assign n50964 = n50963 ^ n50358;
  assign n50966 = n50965 ^ n50964;
  assign n51371 = n51268 ^ n50966;
  assign n51372 = n51371 ^ n48645;
  assign n51373 = n51265 ^ n51263;
  assign n51374 = n51373 ^ n48601;
  assign n51375 = n51258 ^ n50970;
  assign n51376 = n51375 ^ n48518;
  assign n51377 = n51255 ^ n51253;
  assign n51378 = n51377 ^ n48255;
  assign n51379 = n51249 ^ n50977;
  assign n51380 = n51379 ^ n48258;
  assign n51381 = n51246 ^ n50981;
  assign n51382 = n51381 ^ n48262;
  assign n51383 = n51243 ^ n51241;
  assign n51384 = n51383 ^ n48496;
  assign n51385 = n51237 ^ n51219;
  assign n51386 = n51385 ^ n48264;
  assign n51387 = n51234 ^ n51232;
  assign n51388 = n51387 ^ n48486;
  assign n51389 = n51223 ^ n51221;
  assign n51390 = ~n48270 & ~n51389;
  assign n51391 = n51390 ^ n48269;
  assign n51392 = n51228 ^ n51227;
  assign n51393 = n51392 ^ n51390;
  assign n51394 = n51391 & ~n51393;
  assign n51395 = n51394 ^ n48269;
  assign n51396 = n51395 ^ n51387;
  assign n51397 = ~n51388 & n51396;
  assign n51398 = n51397 ^ n48486;
  assign n51399 = n51398 ^ n51385;
  assign n51400 = ~n51386 & n51399;
  assign n51401 = n51400 ^ n48264;
  assign n51402 = n51401 ^ n51383;
  assign n51403 = n51384 & ~n51402;
  assign n51404 = n51403 ^ n48496;
  assign n51405 = n51404 ^ n51381;
  assign n51406 = ~n51382 & ~n51405;
  assign n51407 = n51406 ^ n48262;
  assign n51408 = n51407 ^ n51379;
  assign n51409 = ~n51380 & ~n51408;
  assign n51410 = n51409 ^ n48258;
  assign n51411 = n51410 ^ n51377;
  assign n51412 = ~n51378 & ~n51411;
  assign n51413 = n51412 ^ n48255;
  assign n51414 = n51413 ^ n51375;
  assign n51415 = n51376 & ~n51414;
  assign n51416 = n51415 ^ n48518;
  assign n51417 = n51416 ^ n51373;
  assign n51418 = ~n51374 & ~n51417;
  assign n51419 = n51418 ^ n48601;
  assign n51420 = n51419 ^ n51371;
  assign n51421 = n51372 & ~n51420;
  assign n51422 = n51421 ^ n48645;
  assign n51273 = n49715 ^ n48861;
  assign n51274 = n51273 ^ n50354;
  assign n51269 = n51268 ^ n50965;
  assign n51270 = n50966 & n51269;
  assign n51271 = n51270 ^ n50964;
  assign n50962 = n50848 ^ n50807;
  assign n51272 = n51271 ^ n50962;
  assign n51369 = n51274 ^ n51272;
  assign n51370 = n51369 ^ n48664;
  assign n51494 = n51422 ^ n51370;
  assign n51475 = n51419 ^ n51372;
  assign n51476 = n51416 ^ n51374;
  assign n51477 = n51413 ^ n51376;
  assign n51478 = n51410 ^ n51378;
  assign n51479 = n51398 ^ n51386;
  assign n51480 = n51392 ^ n51391;
  assign n51481 = n51395 ^ n51388;
  assign n51482 = ~n51480 & n51481;
  assign n51483 = ~n51479 & ~n51482;
  assign n51484 = n51401 ^ n51384;
  assign n51485 = ~n51483 & ~n51484;
  assign n51486 = n51404 ^ n51382;
  assign n51487 = ~n51485 & ~n51486;
  assign n51488 = n51407 ^ n51380;
  assign n51489 = ~n51487 & ~n51488;
  assign n51490 = n51478 & n51489;
  assign n51491 = n51477 & n51490;
  assign n51492 = n51476 & ~n51491;
  assign n51493 = n51475 & n51492;
  assign n51579 = n51494 ^ n51493;
  assign n51576 = n49568 ^ n45959;
  assign n51577 = n51576 ^ n42209;
  assign n51578 = n51577 ^ n40306;
  assign n51580 = n51579 ^ n51578;
  assign n51584 = n51492 ^ n51475;
  assign n51581 = n49571 ^ n42214;
  assign n51582 = n51581 ^ n45965;
  assign n51583 = n51582 ^ n40311;
  assign n51585 = n51584 ^ n51583;
  assign n51590 = n51490 ^ n51477;
  assign n51587 = n49581 ^ n41676;
  assign n51588 = n51587 ^ n45975;
  assign n51589 = n51588 ^ n40318;
  assign n51591 = n51590 ^ n51589;
  assign n51596 = n51488 ^ n51487;
  assign n51593 = n49626 ^ n41687;
  assign n51594 = n51593 ^ n45985;
  assign n51595 = n51594 ^ n40328;
  assign n51597 = n51596 ^ n51595;
  assign n51602 = n51484 ^ n51483;
  assign n51599 = n41712 ^ n2397;
  assign n51600 = n51599 ^ n46012;
  assign n51601 = n51600 ^ n40359;
  assign n51603 = n51602 ^ n51601;
  assign n51607 = n51482 ^ n51479;
  assign n51604 = n49612 ^ n2299;
  assign n51605 = n51604 ^ n45991;
  assign n51606 = n51605 ^ n40338;
  assign n51608 = n51607 ^ n51606;
  assign n51612 = n51481 ^ n51480;
  assign n51609 = n49604 ^ n2281;
  assign n51610 = n51609 ^ n45996;
  assign n51611 = n51610 ^ n40342;
  assign n51613 = n51612 ^ n51611;
  assign n51617 = n49794 ^ n42312;
  assign n51618 = n51617 ^ n46296;
  assign n51619 = n51618 ^ n40828;
  assign n51620 = n51389 ^ n48270;
  assign n51621 = n51619 & n51620;
  assign n51614 = n49600 ^ n41698;
  assign n51615 = n51614 ^ n46000;
  assign n51616 = n51615 ^ n40345;
  assign n51622 = n51621 ^ n51616;
  assign n51623 = n51621 ^ n51480;
  assign n51624 = n51622 & n51623;
  assign n51625 = n51624 ^ n51616;
  assign n51626 = n51625 ^ n51612;
  assign n51627 = n51613 & ~n51626;
  assign n51628 = n51627 ^ n51611;
  assign n51629 = n51628 ^ n51607;
  assign n51630 = n51608 & ~n51629;
  assign n51631 = n51630 ^ n51606;
  assign n51632 = n51631 ^ n51602;
  assign n51633 = ~n51603 & n51632;
  assign n51634 = n51633 ^ n51601;
  assign n51598 = n51486 ^ n51485;
  assign n51635 = n51634 ^ n51598;
  assign n51636 = n49592 ^ n41692;
  assign n51637 = n51636 ^ n46019;
  assign n51638 = n51637 ^ n40333;
  assign n51639 = n51638 ^ n51598;
  assign n51640 = ~n51635 & n51639;
  assign n51641 = n51640 ^ n51638;
  assign n51642 = n51641 ^ n51596;
  assign n51643 = ~n51597 & n51642;
  assign n51644 = n51643 ^ n51595;
  assign n51592 = n51489 ^ n51478;
  assign n51645 = n51644 ^ n51592;
  assign n51646 = n49586 ^ n41681;
  assign n51647 = n51646 ^ n45979;
  assign n51648 = n51647 ^ n40323;
  assign n51649 = n51648 ^ n51592;
  assign n51650 = n51645 & ~n51649;
  assign n51651 = n51650 ^ n51648;
  assign n51652 = n51651 ^ n51590;
  assign n51653 = ~n51591 & n51652;
  assign n51654 = n51653 ^ n51589;
  assign n51586 = n51491 ^ n51476;
  assign n51655 = n51654 ^ n51586;
  assign n51656 = n49576 ^ n41119;
  assign n51657 = n51656 ^ n45970;
  assign n51658 = n51657 ^ n40378;
  assign n51659 = n51658 ^ n51586;
  assign n51660 = n51655 & ~n51659;
  assign n51661 = n51660 ^ n51658;
  assign n51662 = n51661 ^ n51584;
  assign n51663 = n51585 & ~n51662;
  assign n51664 = n51663 ^ n51583;
  assign n51665 = n51664 ^ n51579;
  assign n51666 = n51580 & ~n51665;
  assign n51667 = n51666 ^ n51578;
  assign n51495 = n51493 & n51494;
  assign n51423 = n51422 ^ n51369;
  assign n51424 = n51370 & ~n51423;
  assign n51425 = n51424 ^ n48664;
  assign n51275 = n51274 ^ n50962;
  assign n51276 = n51272 & ~n51275;
  assign n51277 = n51276 ^ n51274;
  assign n50960 = n50855 ^ n50852;
  assign n50958 = n50608 ^ n48858;
  assign n50959 = n50958 ^ n49709;
  assign n50961 = n50960 ^ n50959;
  assign n51367 = n51277 ^ n50961;
  assign n51368 = n51367 ^ n48821;
  assign n51474 = n51425 ^ n51368;
  assign n51574 = n51495 ^ n51474;
  assign n51571 = n49563 ^ n42204;
  assign n51572 = n51571 ^ n45954;
  assign n51573 = n51572 ^ n40302;
  assign n51575 = n51574 ^ n51573;
  assign n51755 = n51667 ^ n51575;
  assign n50946 = n50878 ^ n50875;
  assign n53363 = n51755 ^ n50946;
  assign n51729 = n51168 ^ n51165;
  assign n51727 = n49847 ^ n49185;
  assign n51728 = n51727 ^ n51119;
  assign n51730 = n51729 ^ n51728;
  assign n50935 = n50907 ^ n50904;
  assign n50932 = n50460 ^ n49796;
  assign n50934 = n50933 ^ n50932;
  assign n50936 = n50935 ^ n50934;
  assign n51335 = n50900 ^ n50763;
  assign n51328 = n50897 ^ n50894;
  assign n50940 = n50890 ^ n50767;
  assign n50941 = n50940 ^ n50768;
  assign n50937 = n50383 ^ n49754;
  assign n50939 = n50938 ^ n50937;
  assign n50942 = n50941 ^ n50939;
  assign n51318 = n50887 ^ n50774;
  assign n51311 = n50884 ^ n50779;
  assign n51304 = n50881 ^ n50784;
  assign n50943 = n50136 ^ n48830;
  assign n50945 = n50944 ^ n50943;
  assign n50947 = n50946 ^ n50945;
  assign n50952 = n50871 ^ n50790;
  assign n50948 = n50121 ^ n48835;
  assign n50951 = n50950 ^ n50948;
  assign n50953 = n50952 ^ n50951;
  assign n51291 = n50868 ^ n50795;
  assign n50956 = n50865 ^ n50862;
  assign n50954 = n49944 ^ n48846;
  assign n50955 = n50954 ^ n50751;
  assign n50957 = n50956 ^ n50955;
  assign n51281 = n50858 ^ n50801;
  assign n51278 = n51277 ^ n50960;
  assign n51279 = ~n50961 & ~n51278;
  assign n51280 = n51279 ^ n50959;
  assign n51282 = n51281 ^ n51280;
  assign n51283 = n49708 ^ n48852;
  assign n51284 = n51283 ^ n50702;
  assign n51285 = n51284 ^ n51281;
  assign n51286 = ~n51282 & n51285;
  assign n51287 = n51286 ^ n51284;
  assign n51288 = n51287 ^ n50956;
  assign n51289 = n50957 & ~n51288;
  assign n51290 = n51289 ^ n50955;
  assign n51292 = n51291 ^ n51290;
  assign n51293 = n50061 ^ n48840;
  assign n51294 = n51293 ^ n50921;
  assign n51295 = n51294 ^ n51291;
  assign n51296 = n51292 & ~n51295;
  assign n51297 = n51296 ^ n51294;
  assign n51298 = n51297 ^ n50952;
  assign n51299 = n50953 & ~n51298;
  assign n51300 = n51299 ^ n50951;
  assign n51301 = n51300 ^ n50946;
  assign n51302 = n50947 & n51301;
  assign n51303 = n51302 ^ n50945;
  assign n51305 = n51304 ^ n51303;
  assign n51306 = n50343 ^ n49449;
  assign n51307 = n51306 ^ n50994;
  assign n51308 = n51307 ^ n51304;
  assign n51309 = ~n51305 & n51308;
  assign n51310 = n51309 ^ n51307;
  assign n51312 = n51311 ^ n51310;
  assign n51313 = n50386 ^ n49467;
  assign n51314 = n51313 ^ n50990;
  assign n51315 = n51314 ^ n51311;
  assign n51316 = n51312 & n51315;
  assign n51317 = n51316 ^ n51314;
  assign n51319 = n51318 ^ n51317;
  assign n51320 = n50385 ^ n49481;
  assign n51321 = n51320 ^ n50986;
  assign n51322 = n51321 ^ n51318;
  assign n51323 = ~n51319 & n51322;
  assign n51324 = n51323 ^ n51321;
  assign n51325 = n51324 ^ n50939;
  assign n51326 = ~n50942 & ~n51325;
  assign n51327 = n51326 ^ n50941;
  assign n51329 = n51328 ^ n51327;
  assign n51330 = n50382 ^ n49749;
  assign n51331 = n51330 ^ n50985;
  assign n51332 = n51331 ^ n51328;
  assign n51333 = n51329 & ~n51332;
  assign n51334 = n51333 ^ n51331;
  assign n51336 = n51335 ^ n51334;
  assign n51337 = n50442 ^ n49766;
  assign n51338 = n51337 ^ n50984;
  assign n51339 = n51338 ^ n51335;
  assign n51340 = ~n51336 & n51339;
  assign n51341 = n51340 ^ n51338;
  assign n51342 = n51341 ^ n50934;
  assign n51343 = n50936 & ~n51342;
  assign n51344 = n51343 ^ n50935;
  assign n50931 = n50930 ^ n50910;
  assign n51345 = n51344 ^ n50931;
  assign n49704 = n49703 ^ n49178;
  assign n50353 = n50352 ^ n49704;
  assign n51724 = n50931 ^ n50353;
  assign n51725 = ~n51345 & n51724;
  assign n51726 = n51725 ^ n50353;
  assign n51731 = n51730 ^ n51726;
  assign n51840 = n51731 ^ n48451;
  assign n51347 = n51338 ^ n51336;
  assign n51348 = n51347 ^ n48976;
  assign n51349 = n51331 ^ n51329;
  assign n51350 = n51349 ^ n48250;
  assign n51353 = n51314 ^ n51312;
  assign n51354 = n51353 ^ n48843;
  assign n51355 = n51307 ^ n51305;
  assign n51356 = n51355 ^ n48849;
  assign n51357 = n51300 ^ n50947;
  assign n51358 = n51357 ^ n48855;
  assign n51359 = n51297 ^ n50953;
  assign n51360 = n51359 ^ n48862;
  assign n51361 = n51294 ^ n51292;
  assign n51362 = n51361 ^ n48869;
  assign n51363 = n51287 ^ n50957;
  assign n51364 = n51363 ^ n48873;
  assign n51365 = n51284 ^ n51282;
  assign n51366 = n51365 ^ n48879;
  assign n51426 = n51425 ^ n51367;
  assign n51427 = ~n51368 & ~n51426;
  assign n51428 = n51427 ^ n48821;
  assign n51429 = n51428 ^ n51365;
  assign n51430 = n51366 & n51429;
  assign n51431 = n51430 ^ n48879;
  assign n51432 = n51431 ^ n51363;
  assign n51433 = ~n51364 & ~n51432;
  assign n51434 = n51433 ^ n48873;
  assign n51435 = n51434 ^ n51361;
  assign n51436 = ~n51362 & ~n51435;
  assign n51437 = n51436 ^ n48869;
  assign n51438 = n51437 ^ n51359;
  assign n51439 = ~n51360 & ~n51438;
  assign n51440 = n51439 ^ n48862;
  assign n51441 = n51440 ^ n51357;
  assign n51442 = ~n51358 & n51441;
  assign n51443 = n51442 ^ n48855;
  assign n51444 = n51443 ^ n51355;
  assign n51445 = n51356 & ~n51444;
  assign n51446 = n51445 ^ n48849;
  assign n51447 = n51446 ^ n51353;
  assign n51448 = ~n51354 & ~n51447;
  assign n51449 = n51448 ^ n48843;
  assign n51352 = n51321 ^ n51319;
  assign n51450 = n51449 ^ n51352;
  assign n51451 = n51352 ^ n48837;
  assign n51452 = ~n51450 & n51451;
  assign n51453 = n51452 ^ n48837;
  assign n51351 = n51324 ^ n50942;
  assign n51454 = n51453 ^ n51351;
  assign n51455 = n51351 ^ n48833;
  assign n51456 = n51454 & n51455;
  assign n51457 = n51456 ^ n48833;
  assign n51458 = n51457 ^ n51349;
  assign n51459 = ~n51350 & n51458;
  assign n51460 = n51459 ^ n48250;
  assign n51461 = n51460 ^ n51347;
  assign n51462 = ~n51348 & ~n51461;
  assign n51463 = n51462 ^ n48976;
  assign n51464 = n51463 ^ n49066;
  assign n51465 = n51341 ^ n50936;
  assign n51466 = n51465 ^ n51463;
  assign n51467 = ~n51464 & n51466;
  assign n51468 = n51467 ^ n49066;
  assign n51346 = n51345 ^ n50353;
  assign n51469 = n51468 ^ n51346;
  assign n51720 = n51346 ^ n48448;
  assign n51721 = ~n51469 & n51720;
  assign n51722 = n51721 ^ n48448;
  assign n51841 = n51731 ^ n51722;
  assign n51842 = n51840 & ~n51841;
  assign n51843 = n51842 ^ n48451;
  assign n51813 = n51728 ^ n51726;
  assign n51814 = n51730 & ~n51813;
  assign n51815 = n51814 ^ n51729;
  assign n51811 = n51175 ^ n51172;
  assign n51809 = n49840 ^ n49190;
  assign n51810 = n51809 ^ n50522;
  assign n51812 = n51811 ^ n51810;
  assign n51839 = n51815 ^ n51812;
  assign n51844 = n51843 ^ n51839;
  assign n51845 = n51843 ^ n48443;
  assign n51846 = ~n51844 & ~n51845;
  assign n51847 = n51846 ^ n48443;
  assign n51816 = n51815 ^ n51810;
  assign n51817 = n51812 & n51816;
  assign n51818 = n51817 ^ n51811;
  assign n51807 = n51178 ^ n51159;
  assign n51805 = n49858 ^ n49171;
  assign n51806 = n51805 ^ n50518;
  assign n51808 = n51807 ^ n51806;
  assign n51837 = n51818 ^ n51808;
  assign n51838 = n51837 ^ n48439;
  assign n51856 = n51847 ^ n51838;
  assign n51857 = n51844 ^ n48443;
  assign n51723 = n51722 ^ n48451;
  assign n51732 = n51731 ^ n51723;
  assign n51470 = n51469 ^ n48448;
  assign n51471 = n51460 ^ n51348;
  assign n51472 = n51434 ^ n51362;
  assign n51473 = n51431 ^ n51364;
  assign n51496 = ~n51474 & n51495;
  assign n51497 = n51428 ^ n51366;
  assign n51498 = n51496 & ~n51497;
  assign n51499 = n51473 & ~n51498;
  assign n51500 = ~n51472 & n51499;
  assign n51501 = n51437 ^ n51360;
  assign n51502 = ~n51500 & ~n51501;
  assign n51503 = n51440 ^ n51358;
  assign n51504 = ~n51502 & ~n51503;
  assign n51505 = n51443 ^ n51356;
  assign n51506 = ~n51504 & ~n51505;
  assign n51507 = n51446 ^ n51354;
  assign n51508 = n51506 & n51507;
  assign n51509 = n51450 ^ n48837;
  assign n51510 = n51508 & n51509;
  assign n51511 = n51454 ^ n48833;
  assign n51512 = ~n51510 & ~n51511;
  assign n51513 = n51457 ^ n48250;
  assign n51514 = n51513 ^ n51349;
  assign n51515 = n51512 & ~n51514;
  assign n51516 = n51471 & ~n51515;
  assign n51517 = n51465 ^ n51464;
  assign n51518 = n51516 & n51517;
  assign n51733 = n51470 & ~n51518;
  assign n51858 = ~n51732 & ~n51733;
  assign n51859 = ~n51857 & ~n51858;
  assign n51860 = ~n51856 & ~n51859;
  assign n51848 = n51847 ^ n51837;
  assign n51849 = ~n51838 & ~n51848;
  assign n51850 = n51849 ^ n48439;
  assign n51824 = n49836 ^ n49167;
  assign n51825 = n51824 ^ n50517;
  assign n51822 = n51185 ^ n51182;
  assign n51819 = n51818 ^ n51807;
  assign n51820 = n51808 & n51819;
  assign n51821 = n51820 ^ n51806;
  assign n51823 = n51822 ^ n51821;
  assign n51835 = n51825 ^ n51823;
  assign n51836 = n51835 ^ n48435;
  assign n51855 = n51850 ^ n51836;
  assign n51886 = n51860 ^ n51855;
  assign n51883 = n49826 ^ n42300;
  assign n51884 = n51883 ^ n46321;
  assign n51885 = n51884 ^ n40816;
  assign n51887 = n51886 ^ n51885;
  assign n51889 = n49702 ^ n42293;
  assign n51890 = n51889 ^ n46325;
  assign n51891 = n51890 ^ n40726;
  assign n51888 = n51859 ^ n51856;
  assign n51892 = n51891 ^ n51888;
  assign n51894 = n49495 ^ n3010;
  assign n51895 = n51894 ^ n46330;
  assign n51896 = n51895 ^ n40731;
  assign n51893 = n51858 ^ n51857;
  assign n51897 = n51896 ^ n51893;
  assign n51735 = n49501 ^ n2995;
  assign n51736 = n51735 ^ n46336;
  assign n51737 = n51736 ^ n40803;
  assign n51734 = n51733 ^ n51732;
  assign n51738 = n51737 ^ n51734;
  assign n51523 = n51517 ^ n51516;
  assign n51520 = n49510 ^ n42166;
  assign n51521 = n51520 ^ n46345;
  assign n51522 = n51521 ^ n40742;
  assign n51524 = n51523 ^ n51522;
  assign n51526 = n49515 ^ n42170;
  assign n51527 = n51526 ^ n46351;
  assign n51528 = n51527 ^ n3095;
  assign n51525 = n51515 ^ n51471;
  assign n51529 = n51528 ^ n51525;
  assign n51533 = n51514 ^ n51512;
  assign n51530 = n49520 ^ n42175;
  assign n51531 = n51530 ^ n46355;
  assign n51532 = n51531 ^ n2624;
  assign n51534 = n51533 ^ n51532;
  assign n51538 = n51511 ^ n51510;
  assign n51535 = n49525 ^ n42180;
  assign n51536 = n51535 ^ n45500;
  assign n51537 = n51536 ^ n40784;
  assign n51539 = n51538 ^ n51537;
  assign n51541 = n49531 ^ n42185;
  assign n51542 = n51541 ^ n45929;
  assign n51543 = n51542 ^ n40752;
  assign n51540 = n51509 ^ n51508;
  assign n51544 = n51543 ^ n51540;
  assign n51549 = n51505 ^ n51504;
  assign n51546 = n49540 ^ n42192;
  assign n51547 = n51546 ^ n1439;
  assign n51548 = n51547 ^ n40762;
  assign n51550 = n51549 ^ n51548;
  assign n51554 = n51503 ^ n51502;
  assign n51551 = n49545 ^ n42251;
  assign n51552 = n51551 ^ n46059;
  assign n51553 = n51552 ^ n1428;
  assign n51555 = n51554 ^ n51553;
  assign n51559 = n51499 ^ n51472;
  assign n51556 = n49659 ^ n42241;
  assign n51557 = n51556 ^ n45940;
  assign n51558 = n51557 ^ n1246;
  assign n51560 = n51559 ^ n51558;
  assign n51564 = n51498 ^ n51473;
  assign n51561 = n49553 ^ n1068;
  assign n51562 = n51561 ^ n45944;
  assign n51563 = n51562 ^ n3341;
  assign n51565 = n51564 ^ n51563;
  assign n51566 = n51497 ^ n51496;
  assign n51570 = n51569 ^ n51566;
  assign n51668 = n51667 ^ n51574;
  assign n51669 = ~n51575 & n51668;
  assign n51670 = n51669 ^ n51573;
  assign n51671 = n51670 ^ n51569;
  assign n51672 = ~n51570 & ~n51671;
  assign n51673 = n51672 ^ n51566;
  assign n51674 = n51673 ^ n51564;
  assign n51675 = n51565 & n51674;
  assign n51676 = n51675 ^ n51563;
  assign n51677 = n51676 ^ n51559;
  assign n51678 = n51560 & ~n51677;
  assign n51679 = n51678 ^ n51558;
  assign n1218 = n1217 ^ n1169;
  assign n1255 = n1254 ^ n1218;
  assign n1265 = n1264 ^ n1255;
  assign n51680 = n51679 ^ n1265;
  assign n51681 = n51501 ^ n51500;
  assign n51682 = n51681 ^ n51679;
  assign n51683 = n51680 & ~n51682;
  assign n51684 = n51683 ^ n1265;
  assign n51685 = n51684 ^ n51554;
  assign n51686 = ~n51555 & n51685;
  assign n51687 = n51686 ^ n51553;
  assign n51688 = n51687 ^ n51549;
  assign n51689 = n51550 & ~n51688;
  assign n51690 = n51689 ^ n51548;
  assign n51545 = n51507 ^ n51506;
  assign n51691 = n51690 ^ n51545;
  assign n51692 = n49535 ^ n42261;
  assign n51693 = n51692 ^ n46069;
  assign n51694 = n51693 ^ n40757;
  assign n51695 = n51694 ^ n51545;
  assign n51696 = ~n51691 & n51695;
  assign n51697 = n51696 ^ n51694;
  assign n51698 = n51697 ^ n51543;
  assign n51699 = n51544 & ~n51698;
  assign n51700 = n51699 ^ n51540;
  assign n51701 = n51700 ^ n51538;
  assign n51702 = ~n51539 & n51701;
  assign n51703 = n51702 ^ n51537;
  assign n51704 = n51703 ^ n51533;
  assign n51705 = n51534 & ~n51704;
  assign n51706 = n51705 ^ n51532;
  assign n51707 = n51706 ^ n51528;
  assign n51708 = ~n51529 & ~n51707;
  assign n51709 = n51708 ^ n51525;
  assign n51710 = n51709 ^ n51523;
  assign n51711 = n51524 & n51710;
  assign n51712 = n51711 ^ n51522;
  assign n51519 = n51518 ^ n51470;
  assign n51713 = n51712 ^ n51519;
  assign n51714 = n49506 ^ n42160;
  assign n51715 = n51714 ^ n46340;
  assign n51716 = n51715 ^ n40737;
  assign n51717 = n51716 ^ n51519;
  assign n51718 = ~n51713 & n51717;
  assign n51719 = n51718 ^ n51716;
  assign n51898 = n51737 ^ n51719;
  assign n51899 = n51738 & ~n51898;
  assign n51900 = n51899 ^ n51734;
  assign n51901 = n51900 ^ n51896;
  assign n51902 = ~n51897 & ~n51901;
  assign n51903 = n51902 ^ n51893;
  assign n51904 = n51903 ^ n51891;
  assign n51905 = n51892 & n51904;
  assign n51906 = n51905 ^ n51888;
  assign n51907 = n51906 ^ n51886;
  assign n51908 = n51887 & ~n51907;
  assign n51909 = n51908 ^ n51885;
  assign n51879 = n49817 ^ n42150;
  assign n51880 = n51879 ^ n46315;
  assign n51881 = n51880 ^ n1802;
  assign n51861 = n51855 & n51860;
  assign n51851 = n51850 ^ n51835;
  assign n51852 = ~n51836 & n51851;
  assign n51853 = n51852 ^ n48435;
  assign n51831 = n51188 ^ n51153;
  assign n51829 = n49745 ^ n49200;
  assign n51830 = n51829 ^ n50513;
  assign n51832 = n51831 ^ n51830;
  assign n51826 = n51825 ^ n51822;
  assign n51827 = n51823 & ~n51826;
  assign n51828 = n51827 ^ n51825;
  assign n51833 = n51832 ^ n51828;
  assign n51834 = n51833 ^ n48467;
  assign n51854 = n51853 ^ n51834;
  assign n51878 = n51861 ^ n51854;
  assign n51882 = n51881 ^ n51878;
  assign n51937 = n51909 ^ n51882;
  assign n51919 = n51906 ^ n51885;
  assign n51920 = n51919 ^ n51886;
  assign n51917 = n50366 ^ n49732;
  assign n51918 = n51917 ^ n50972;
  assign n51921 = n51920 ^ n51918;
  assign n51926 = n50368 ^ n49735;
  assign n51927 = n51926 ^ n50974;
  assign n51922 = n51900 ^ n51897;
  assign n51923 = n50369 ^ n49737;
  assign n51924 = n51923 ^ n50978;
  assign n51925 = ~n51922 & n51924;
  assign n51928 = n51927 ^ n51925;
  assign n51929 = n51903 ^ n51892;
  assign n51930 = n51929 ^ n51927;
  assign n51931 = n51928 & n51930;
  assign n51932 = n51931 ^ n51925;
  assign n51933 = n51932 ^ n51920;
  assign n51934 = n51921 & ~n51933;
  assign n51935 = n51934 ^ n51918;
  assign n51915 = n50569 ^ n49728;
  assign n51916 = n51915 ^ n50969;
  assign n51936 = n51935 ^ n51916;
  assign n52024 = n51937 ^ n51936;
  assign n52025 = n52024 ^ n48900;
  assign n52026 = n51932 ^ n51921;
  assign n52027 = n52026 ^ n48904;
  assign n52028 = n51924 ^ n51922;
  assign n52029 = ~n48909 & ~n52028;
  assign n52030 = n52029 ^ n49218;
  assign n52031 = n51929 ^ n51928;
  assign n52032 = n52031 ^ n52029;
  assign n52033 = n52030 & n52032;
  assign n52034 = n52033 ^ n49218;
  assign n52035 = n52034 ^ n52026;
  assign n52036 = ~n52027 & ~n52035;
  assign n52037 = n52036 ^ n48904;
  assign n52038 = n52037 ^ n52024;
  assign n52039 = ~n52025 & ~n52038;
  assign n52040 = n52039 ^ n48900;
  assign n52110 = n52040 ^ n48895;
  assign n51938 = n51937 ^ n51935;
  assign n51939 = n51936 & n51938;
  assign n51940 = n51939 ^ n51916;
  assign n51910 = n51909 ^ n51881;
  assign n51911 = ~n51882 & ~n51910;
  assign n51912 = n51911 ^ n51878;
  assign n51872 = n51853 ^ n51833;
  assign n51873 = ~n51834 & ~n51872;
  assign n51874 = n51873 ^ n48467;
  assign n51870 = n51191 ^ n51148;
  assign n51866 = n51830 ^ n51828;
  assign n51867 = ~n51832 & n51866;
  assign n51868 = n51867 ^ n51828;
  assign n51864 = n49741 ^ n49208;
  assign n51865 = n51864 ^ n50512;
  assign n51869 = n51868 ^ n51865;
  assign n51871 = n51870 ^ n51869;
  assign n51875 = n51874 ^ n51871;
  assign n51876 = n51875 ^ n48275;
  assign n51862 = ~n51854 & ~n51861;
  assign n51802 = n49812 ^ n42146;
  assign n51803 = n51802 ^ n46391;
  assign n51804 = n51803 ^ n40717;
  assign n51863 = n51862 ^ n51804;
  assign n51877 = n51876 ^ n51863;
  assign n51913 = n51912 ^ n51877;
  assign n51800 = n50577 ^ n49727;
  assign n51801 = n51800 ^ n51262;
  assign n51914 = n51913 ^ n51801;
  assign n52022 = n51940 ^ n51914;
  assign n52111 = n52110 ^ n52022;
  assign n52112 = n52037 ^ n52025;
  assign n52113 = n52031 ^ n52030;
  assign n52114 = n52034 ^ n48904;
  assign n52115 = n52114 ^ n52026;
  assign n52116 = n52113 & n52115;
  assign n52117 = n52112 & ~n52116;
  assign n52118 = ~n52111 & ~n52117;
  assign n52023 = n52022 ^ n48895;
  assign n52041 = n52040 ^ n52022;
  assign n52042 = n52023 & ~n52041;
  assign n52043 = n52042 ^ n48895;
  assign n51945 = n50365 ^ n49725;
  assign n51946 = n51945 ^ n50965;
  assign n51941 = n51940 ^ n51913;
  assign n51942 = n51914 & n51941;
  assign n51943 = n51942 ^ n51801;
  assign n51799 = n51620 ^ n51619;
  assign n51944 = n51943 ^ n51799;
  assign n52021 = n51946 ^ n51944;
  assign n52044 = n52043 ^ n52021;
  assign n52119 = n52044 ^ n48891;
  assign n52120 = ~n52118 & ~n52119;
  assign n52045 = n52021 ^ n48891;
  assign n52046 = ~n52044 & ~n52045;
  assign n52047 = n52046 ^ n48891;
  assign n52121 = n52047 ^ n49237;
  assign n51951 = n50364 ^ n49901;
  assign n51952 = n51951 ^ n50962;
  assign n51947 = n51946 ^ n51799;
  assign n51948 = n51944 & ~n51947;
  assign n51949 = n51948 ^ n51946;
  assign n51797 = n51616 ^ n51480;
  assign n51798 = n51797 ^ n51621;
  assign n51950 = n51949 ^ n51798;
  assign n52019 = n51952 ^ n51950;
  assign n52122 = n52121 ^ n52019;
  assign n52123 = ~n52120 & ~n52122;
  assign n52020 = n52019 ^ n49237;
  assign n52048 = n52047 ^ n52019;
  assign n52049 = ~n52020 & n52048;
  assign n52050 = n52049 ^ n49237;
  assign n51953 = n51952 ^ n51798;
  assign n51954 = ~n51950 & ~n51953;
  assign n51955 = n51954 ^ n51952;
  assign n51795 = n51625 ^ n51613;
  assign n51793 = n50361 ^ n49721;
  assign n51794 = n51793 ^ n50960;
  assign n51796 = n51795 ^ n51794;
  assign n52018 = n51955 ^ n51796;
  assign n52051 = n52050 ^ n52018;
  assign n52124 = n52051 ^ n48886;
  assign n52125 = n52123 & n52124;
  assign n52052 = n52018 ^ n48886;
  assign n52053 = n52051 & n52052;
  assign n52054 = n52053 ^ n48886;
  assign n51956 = n51955 ^ n51795;
  assign n51957 = n51796 & ~n51956;
  assign n51958 = n51957 ^ n51794;
  assign n51791 = n51628 ^ n51608;
  assign n51789 = n50358 ^ n49911;
  assign n51790 = n51789 ^ n51281;
  assign n51792 = n51791 ^ n51790;
  assign n52017 = n51958 ^ n51792;
  assign n52055 = n52054 ^ n52017;
  assign n52126 = n52055 ^ n48882;
  assign n52127 = n52125 & ~n52126;
  assign n52056 = n52017 ^ n48882;
  assign n52057 = ~n52055 & n52056;
  assign n52058 = n52057 ^ n48882;
  assign n51959 = n51958 ^ n51791;
  assign n51960 = n51792 & ~n51959;
  assign n51961 = n51960 ^ n51790;
  assign n51785 = n50354 ^ n49918;
  assign n51786 = n51785 ^ n50956;
  assign n52014 = n51961 ^ n51786;
  assign n51787 = n51631 ^ n51603;
  assign n52015 = n52014 ^ n51787;
  assign n52016 = n52015 ^ n48876;
  assign n52109 = n52058 ^ n52016;
  assign n52197 = n52127 ^ n52109;
  assign n52194 = n50202 ^ n42502;
  assign n52195 = n52194 ^ n46756;
  assign n52196 = n52195 ^ n41073;
  assign n52198 = n52197 ^ n52196;
  assign n52202 = n52126 ^ n52125;
  assign n52199 = n50207 ^ n42560;
  assign n52200 = n52199 ^ n46761;
  assign n52201 = n52200 ^ n41016;
  assign n52203 = n52202 ^ n52201;
  assign n52207 = n52124 ^ n52123;
  assign n52204 = n50210 ^ n42508;
  assign n52205 = n52204 ^ n46765;
  assign n52206 = n52205 ^ n41020;
  assign n52208 = n52207 ^ n52206;
  assign n52212 = n52122 ^ n52120;
  assign n52209 = n50215 ^ n42550;
  assign n52210 = n52209 ^ n46770;
  assign n52211 = n52210 ^ n41025;
  assign n52213 = n52212 ^ n52211;
  assign n52218 = n52117 ^ n52111;
  assign n52215 = n50221 ^ n42518;
  assign n52216 = n52215 ^ n46795;
  assign n52217 = n52216 ^ n41036;
  assign n52219 = n52218 ^ n52217;
  assign n52223 = n52116 ^ n52112;
  assign n52220 = n50226 ^ n42523;
  assign n52221 = n52220 ^ n46787;
  assign n52222 = n52221 ^ n41040;
  assign n52224 = n52223 ^ n52222;
  assign n52233 = n50231 ^ n42529;
  assign n52234 = n52233 ^ n2024;
  assign n52235 = n52234 ^ n41044;
  assign n52228 = n52028 ^ n48909;
  assign n52229 = n50381 ^ n42849;
  assign n52230 = n52229 ^ n47041;
  assign n52231 = n52230 ^ n2013;
  assign n52232 = n52228 & n52231;
  assign n52236 = n52235 ^ n52232;
  assign n52237 = n52232 ^ n52113;
  assign n52238 = n52236 & ~n52237;
  assign n52239 = n52238 ^ n52235;
  assign n52225 = n50236 ^ n42533;
  assign n52226 = n52225 ^ n46777;
  assign n52227 = n52226 ^ n2159;
  assign n52240 = n52239 ^ n52227;
  assign n52241 = n52115 ^ n52113;
  assign n52242 = n52241 ^ n52239;
  assign n52243 = n52240 & n52242;
  assign n52244 = n52243 ^ n52227;
  assign n52245 = n52244 ^ n52223;
  assign n52246 = ~n52224 & n52245;
  assign n52247 = n52246 ^ n52222;
  assign n52248 = n52247 ^ n52218;
  assign n52249 = ~n52219 & n52248;
  assign n52250 = n52249 ^ n52217;
  assign n52214 = n52119 ^ n52118;
  assign n52251 = n52250 ^ n52214;
  assign n52252 = n50218 ^ n42513;
  assign n52253 = n52252 ^ n46802;
  assign n52254 = n52253 ^ n41031;
  assign n52255 = n52254 ^ n52214;
  assign n52256 = ~n52251 & n52255;
  assign n52257 = n52256 ^ n52254;
  assign n52258 = n52257 ^ n52212;
  assign n52259 = ~n52213 & n52258;
  assign n52260 = n52259 ^ n52211;
  assign n52261 = n52260 ^ n52207;
  assign n52262 = ~n52208 & n52261;
  assign n52263 = n52262 ^ n52206;
  assign n52264 = n52263 ^ n52202;
  assign n52265 = n52203 & ~n52264;
  assign n52266 = n52265 ^ n52201;
  assign n52267 = n52266 ^ n52197;
  assign n52268 = ~n52198 & n52267;
  assign n52269 = n52268 ^ n52196;
  assign n52190 = n50271 ^ n42570;
  assign n52191 = n52190 ^ n46751;
  assign n52192 = n52191 ^ n41010;
  assign n52375 = n52269 ^ n52192;
  assign n52128 = n52109 & ~n52127;
  assign n51788 = n51787 ^ n51786;
  assign n51962 = n51961 ^ n51787;
  assign n51963 = n51788 & n51962;
  assign n51964 = n51963 ^ n51786;
  assign n51783 = n51638 ^ n51635;
  assign n51781 = n50608 ^ n49718;
  assign n51782 = n51781 ^ n51291;
  assign n51784 = n51783 ^ n51782;
  assign n52063 = n51964 ^ n51784;
  assign n52107 = n52063 ^ n48867;
  assign n52059 = n52058 ^ n52015;
  assign n52060 = n52016 & ~n52059;
  assign n52061 = n52060 ^ n48876;
  assign n52108 = n52107 ^ n52061;
  assign n52189 = n52128 ^ n52108;
  assign n52376 = n52375 ^ n52189;
  assign n53364 = n53363 ^ n52376;
  assign n52636 = n50969 ^ n50368;
  assign n52637 = n52636 ^ n51798;
  assign n52631 = n50972 ^ n50369;
  assign n52632 = n52631 ^ n51799;
  assign n52320 = n50984 ^ n50383;
  assign n52321 = n52320 ^ n51729;
  assign n52318 = n51681 ^ n1265;
  assign n52319 = n52318 ^ n51679;
  assign n52322 = n52321 ^ n52319;
  assign n51746 = n50938 ^ n50386;
  assign n51747 = n51746 ^ n50935;
  assign n51745 = n51673 ^ n51565;
  assign n51748 = n51747 ^ n51745;
  assign n51750 = n50986 ^ n50343;
  assign n51751 = n51750 ^ n51335;
  assign n51749 = n51670 ^ n51570;
  assign n51752 = n51751 ^ n51749;
  assign n51753 = n50990 ^ n50136;
  assign n51754 = n51753 ^ n51328;
  assign n51756 = n51755 ^ n51754;
  assign n51758 = n50994 ^ n50121;
  assign n51759 = n51758 ^ n50941;
  assign n51757 = n51664 ^ n51580;
  assign n51760 = n51759 ^ n51757;
  assign n51763 = n51661 ^ n51585;
  assign n51761 = n50944 ^ n50061;
  assign n51762 = n51761 ^ n51318;
  assign n51764 = n51763 ^ n51762;
  assign n51766 = n50950 ^ n49944;
  assign n51767 = n51766 ^ n51311;
  assign n51765 = n51658 ^ n51655;
  assign n51768 = n51767 ^ n51765;
  assign n51771 = n51651 ^ n51591;
  assign n51769 = n50921 ^ n49708;
  assign n51770 = n51769 ^ n51304;
  assign n51772 = n51771 ^ n51770;
  assign n51774 = n50751 ^ n49709;
  assign n51775 = n51774 ^ n50946;
  assign n51773 = n51648 ^ n51645;
  assign n51776 = n51775 ^ n51773;
  assign n51779 = n51641 ^ n51597;
  assign n51777 = n50702 ^ n49715;
  assign n51778 = n51777 ^ n50952;
  assign n51780 = n51779 ^ n51778;
  assign n51965 = n51964 ^ n51782;
  assign n51966 = n51784 & n51965;
  assign n51967 = n51966 ^ n51783;
  assign n51968 = n51967 ^ n51779;
  assign n51969 = n51780 & n51968;
  assign n51970 = n51969 ^ n51778;
  assign n51971 = n51970 ^ n51775;
  assign n51972 = n51776 & ~n51971;
  assign n51973 = n51972 ^ n51773;
  assign n51974 = n51973 ^ n51771;
  assign n51975 = n51772 & ~n51974;
  assign n51976 = n51975 ^ n51770;
  assign n51977 = n51976 ^ n51765;
  assign n51978 = ~n51768 & ~n51977;
  assign n51979 = n51978 ^ n51767;
  assign n51980 = n51979 ^ n51763;
  assign n51981 = ~n51764 & ~n51980;
  assign n51982 = n51981 ^ n51762;
  assign n51983 = n51982 ^ n51757;
  assign n51984 = n51760 & n51983;
  assign n51985 = n51984 ^ n51759;
  assign n51986 = n51985 ^ n51755;
  assign n51987 = ~n51756 & n51986;
  assign n51988 = n51987 ^ n51754;
  assign n51989 = n51988 ^ n51749;
  assign n51990 = ~n51752 & n51989;
  assign n51991 = n51990 ^ n51751;
  assign n51992 = n51991 ^ n51747;
  assign n51993 = n51748 & n51992;
  assign n51994 = n51993 ^ n51745;
  assign n51744 = n51676 ^ n51560;
  assign n51995 = n51994 ^ n51744;
  assign n51742 = n50985 ^ n50385;
  assign n51743 = n51742 ^ n50931;
  assign n52315 = n51744 ^ n51743;
  assign n52316 = n51995 & n52315;
  assign n52317 = n52316 ^ n51743;
  assign n52323 = n52322 ^ n52317;
  assign n52324 = n52323 ^ n49754;
  assign n51997 = n51991 ^ n51748;
  assign n51998 = n51997 ^ n49467;
  assign n52000 = n51985 ^ n51754;
  assign n52001 = n52000 ^ n51755;
  assign n52002 = n52001 ^ n48830;
  assign n52003 = n51982 ^ n51760;
  assign n52004 = n52003 ^ n48835;
  assign n52005 = n51979 ^ n51762;
  assign n52006 = n52005 ^ n51763;
  assign n52007 = n52006 ^ n48840;
  assign n52008 = n51976 ^ n51768;
  assign n52009 = n52008 ^ n48846;
  assign n52010 = n51973 ^ n51772;
  assign n52011 = n52010 ^ n48852;
  assign n52012 = n51967 ^ n51780;
  assign n52013 = n52012 ^ n48861;
  assign n52062 = n52061 ^ n48867;
  assign n52064 = n52063 ^ n52061;
  assign n52065 = ~n52062 & n52064;
  assign n52066 = n52065 ^ n48867;
  assign n52067 = n52066 ^ n52012;
  assign n52068 = n52013 & n52067;
  assign n52069 = n52068 ^ n48861;
  assign n52070 = n52069 ^ n48858;
  assign n52071 = n51970 ^ n51776;
  assign n52072 = n52071 ^ n52069;
  assign n52073 = ~n52070 & n52072;
  assign n52074 = n52073 ^ n48858;
  assign n52075 = n52074 ^ n52010;
  assign n52076 = n52011 & ~n52075;
  assign n52077 = n52076 ^ n48852;
  assign n52078 = n52077 ^ n52008;
  assign n52079 = ~n52009 & n52078;
  assign n52080 = n52079 ^ n48846;
  assign n52081 = n52080 ^ n52006;
  assign n52082 = ~n52007 & ~n52081;
  assign n52083 = n52082 ^ n48840;
  assign n52084 = n52083 ^ n52003;
  assign n52085 = ~n52004 & n52084;
  assign n52086 = n52085 ^ n48835;
  assign n52087 = n52086 ^ n52001;
  assign n52088 = ~n52002 & n52087;
  assign n52089 = n52088 ^ n48830;
  assign n51999 = n51988 ^ n51752;
  assign n52090 = n52089 ^ n51999;
  assign n52091 = n51999 ^ n49449;
  assign n52092 = n52090 & n52091;
  assign n52093 = n52092 ^ n49449;
  assign n52094 = n52093 ^ n51997;
  assign n52095 = ~n51998 & n52094;
  assign n52096 = n52095 ^ n49467;
  assign n51996 = n51995 ^ n51743;
  assign n52097 = n52096 ^ n51996;
  assign n52312 = n51996 ^ n49481;
  assign n52313 = ~n52097 & n52312;
  assign n52314 = n52313 ^ n49481;
  assign n52325 = n52324 ^ n52314;
  assign n52098 = n52097 ^ n49481;
  assign n52099 = n52090 ^ n49449;
  assign n52100 = n52086 ^ n52002;
  assign n52101 = n52077 ^ n48846;
  assign n52102 = n52101 ^ n52008;
  assign n52103 = n52071 ^ n48858;
  assign n52104 = n52103 ^ n52069;
  assign n52105 = n52066 ^ n48861;
  assign n52106 = n52105 ^ n52012;
  assign n52129 = n52108 & n52128;
  assign n52130 = ~n52106 & n52129;
  assign n52131 = n52104 & n52130;
  assign n52132 = n52074 ^ n48852;
  assign n52133 = n52132 ^ n52010;
  assign n52134 = n52131 & ~n52133;
  assign n52135 = ~n52102 & ~n52134;
  assign n52136 = n52080 ^ n52007;
  assign n52137 = n52135 & ~n52136;
  assign n52138 = n52083 ^ n52004;
  assign n52139 = ~n52137 & ~n52138;
  assign n52140 = n52100 & ~n52139;
  assign n52141 = n52099 & ~n52140;
  assign n52142 = n52093 ^ n49467;
  assign n52143 = n52142 ^ n51997;
  assign n52144 = n52141 & n52143;
  assign n52326 = ~n52098 & n52144;
  assign n52493 = ~n52325 & ~n52326;
  assign n52468 = n52323 ^ n52314;
  assign n52469 = ~n52324 & n52468;
  assign n52470 = n52469 ^ n49754;
  assign n52430 = n52319 ^ n52317;
  assign n52431 = n52322 & ~n52430;
  assign n52432 = n52431 ^ n52321;
  assign n52428 = n51684 ^ n51555;
  assign n52426 = n50933 ^ n50382;
  assign n52427 = n52426 ^ n51811;
  assign n52429 = n52428 ^ n52427;
  assign n52467 = n52432 ^ n52429;
  assign n52471 = n52470 ^ n52467;
  assign n52494 = n52471 ^ n49749;
  assign n52495 = n52493 & ~n52494;
  assign n52472 = n52467 ^ n49749;
  assign n52473 = ~n52471 & ~n52472;
  assign n52474 = n52473 ^ n49749;
  assign n52496 = n52474 ^ n49766;
  assign n52433 = n52432 ^ n52427;
  assign n52434 = ~n52429 & ~n52433;
  assign n52435 = n52434 ^ n52428;
  assign n52423 = n50442 ^ n50352;
  assign n52424 = n52423 ^ n51807;
  assign n52365 = n51687 ^ n51550;
  assign n52425 = n52424 ^ n52365;
  assign n52465 = n52435 ^ n52425;
  assign n52497 = n52496 ^ n52465;
  assign n52498 = ~n52495 & ~n52497;
  assign n52466 = n52465 ^ n49766;
  assign n52475 = n52474 ^ n52465;
  assign n52476 = ~n52466 & n52475;
  assign n52477 = n52476 ^ n49766;
  assign n52436 = n52435 ^ n52365;
  assign n52437 = n52425 & n52436;
  assign n52438 = n52437 ^ n52424;
  assign n52420 = n51119 ^ n50460;
  assign n52421 = n52420 ^ n51822;
  assign n52358 = n51694 ^ n51691;
  assign n52422 = n52421 ^ n52358;
  assign n52463 = n52438 ^ n52422;
  assign n52464 = n52463 ^ n49796;
  assign n52499 = n52477 ^ n52464;
  assign n52500 = n52498 & n52499;
  assign n52478 = n52477 ^ n52463;
  assign n52479 = n52464 & ~n52478;
  assign n52480 = n52479 ^ n49796;
  assign n52439 = n52438 ^ n52358;
  assign n52440 = n52422 & ~n52439;
  assign n52441 = n52440 ^ n52421;
  assign n52417 = n50522 ^ n49703;
  assign n52418 = n52417 ^ n51831;
  assign n52354 = n51697 ^ n51544;
  assign n52419 = n52418 ^ n52354;
  assign n52461 = n52441 ^ n52419;
  assign n52462 = n52461 ^ n49178;
  assign n52492 = n52480 ^ n52462;
  assign n52576 = n52500 ^ n52492;
  assign n52573 = n49707 ^ n42949;
  assign n52574 = n52573 ^ n2804;
  assign n52575 = n52574 ^ n3135;
  assign n52577 = n52576 ^ n52575;
  assign n52581 = n52499 ^ n52498;
  assign n52578 = n50147 ^ n3107;
  assign n52579 = n52578 ^ n46692;
  assign n52580 = n52579 ^ n2796;
  assign n52582 = n52581 ^ n52580;
  assign n52587 = n52494 ^ n52493;
  assign n52584 = n50153 ^ n42894;
  assign n52585 = n52584 ^ n46702;
  assign n52586 = n52585 ^ n41455;
  assign n52588 = n52587 ^ n52586;
  assign n52327 = n52326 ^ n52325;
  assign n52309 = n50158 ^ n42899;
  assign n52310 = n52309 ^ n46707;
  assign n52311 = n52310 ^ n41460;
  assign n52328 = n52327 ^ n52311;
  assign n52149 = n52143 ^ n52141;
  assign n52146 = n50164 ^ n42908;
  assign n52147 = n52146 ^ n46718;
  assign n52148 = n52147 ^ n41467;
  assign n52150 = n52149 ^ n52148;
  assign n52154 = n52140 ^ n52099;
  assign n52151 = n42913 ^ n1476;
  assign n52152 = n52151 ^ n46722;
  assign n52153 = n52152 ^ n41471;
  assign n52155 = n52154 ^ n52153;
  assign n52159 = n52139 ^ n52100;
  assign n52156 = n50170 ^ n1372;
  assign n52157 = n52156 ^ n46850;
  assign n52158 = n52157 ^ n41497;
  assign n52160 = n52159 ^ n52158;
  assign n52164 = n52138 ^ n52137;
  assign n52161 = n50175 ^ n1354;
  assign n52162 = n52161 ^ n46729;
  assign n52163 = n52162 ^ n41478;
  assign n52165 = n52164 ^ n52163;
  assign n52169 = n52136 ^ n52135;
  assign n52166 = n50181 ^ n3350;
  assign n52167 = n52166 ^ n46733;
  assign n52168 = n52167 ^ n41487;
  assign n52170 = n52169 ^ n52168;
  assign n52174 = n52134 ^ n52102;
  assign n52171 = n50185 ^ n42481;
  assign n52172 = n52171 ^ n46738;
  assign n52173 = n52172 ^ n41096;
  assign n52175 = n52174 ^ n52173;
  assign n52179 = n52133 ^ n52131;
  assign n52176 = n50190 ^ n42486;
  assign n52177 = n52176 ^ n46743;
  assign n52178 = n52177 ^ n41090;
  assign n52180 = n52179 ^ n52178;
  assign n52187 = n52129 ^ n52106;
  assign n52184 = n50196 ^ n42495;
  assign n52185 = n52184 ^ n46824;
  assign n52186 = n52185 ^ n41005;
  assign n52188 = n52187 ^ n52186;
  assign n52193 = n52192 ^ n52189;
  assign n52270 = n52269 ^ n52189;
  assign n52271 = n52193 & ~n52270;
  assign n52272 = n52271 ^ n52192;
  assign n52273 = n52272 ^ n52187;
  assign n52274 = ~n52188 & n52273;
  assign n52275 = n52274 ^ n52186;
  assign n52181 = n50281 ^ n42490;
  assign n52182 = n52181 ^ n46831;
  assign n52183 = n52182 ^ n848;
  assign n52276 = n52275 ^ n52183;
  assign n52277 = n52130 ^ n52104;
  assign n52278 = n52277 ^ n52275;
  assign n52279 = n52276 & ~n52278;
  assign n52280 = n52279 ^ n52183;
  assign n52281 = n52280 ^ n52179;
  assign n52282 = ~n52180 & n52281;
  assign n52283 = n52282 ^ n52178;
  assign n52284 = n52283 ^ n52174;
  assign n52285 = ~n52175 & n52284;
  assign n52286 = n52285 ^ n52173;
  assign n52287 = n52286 ^ n52169;
  assign n52288 = n52170 & ~n52287;
  assign n52289 = n52288 ^ n52168;
  assign n52290 = n52289 ^ n52164;
  assign n52291 = n52165 & ~n52290;
  assign n52292 = n52291 ^ n52163;
  assign n52293 = n52292 ^ n52159;
  assign n52294 = n52160 & ~n52293;
  assign n52295 = n52294 ^ n52158;
  assign n52296 = n52295 ^ n52154;
  assign n52297 = ~n52155 & n52296;
  assign n52298 = n52297 ^ n52153;
  assign n52299 = n52298 ^ n52149;
  assign n52300 = n52150 & ~n52299;
  assign n52301 = n52300 ^ n52148;
  assign n52145 = n52144 ^ n52098;
  assign n52302 = n52301 ^ n52145;
  assign n52303 = n50310 ^ n42904;
  assign n52304 = n52303 ^ n46712;
  assign n52305 = n52304 ^ n41510;
  assign n52306 = n52305 ^ n52145;
  assign n52307 = n52302 & ~n52306;
  assign n52308 = n52307 ^ n52305;
  assign n52589 = n52327 ^ n52308;
  assign n52590 = ~n52328 & n52589;
  assign n52591 = n52590 ^ n52311;
  assign n52592 = n52591 ^ n52587;
  assign n52593 = n52588 & ~n52592;
  assign n52594 = n52593 ^ n52586;
  assign n52583 = n52497 ^ n52495;
  assign n52595 = n52594 ^ n52583;
  assign n52596 = n50323 ^ n2681;
  assign n52597 = n52596 ^ n46697;
  assign n52598 = n52597 ^ n3215;
  assign n52599 = n52598 ^ n52583;
  assign n52600 = ~n52595 & n52599;
  assign n52601 = n52600 ^ n52598;
  assign n52602 = n52601 ^ n52581;
  assign n52603 = n52582 & ~n52602;
  assign n52604 = n52603 ^ n52580;
  assign n52605 = n52604 ^ n52576;
  assign n52606 = n52577 & ~n52605;
  assign n52607 = n52606 ^ n52575;
  assign n52570 = n50335 ^ n42885;
  assign n52571 = n52570 ^ n3137;
  assign n52572 = n52571 ^ n2894;
  assign n52608 = n52607 ^ n52572;
  assign n52501 = n52492 & ~n52500;
  assign n52481 = n52480 ^ n52461;
  assign n52482 = ~n52462 & n52481;
  assign n52483 = n52482 ^ n49178;
  assign n52446 = n50518 ^ n49847;
  assign n52447 = n52446 ^ n51870;
  assign n52442 = n52441 ^ n52354;
  assign n52443 = ~n52419 & ~n52442;
  assign n52444 = n52443 ^ n52418;
  assign n52347 = n51700 ^ n51539;
  assign n52445 = n52444 ^ n52347;
  assign n52459 = n52447 ^ n52445;
  assign n52460 = n52459 ^ n49185;
  assign n52491 = n52483 ^ n52460;
  assign n52609 = n52501 ^ n52491;
  assign n52610 = n52609 ^ n52607;
  assign n52611 = n52608 & n52610;
  assign n52612 = n52611 ^ n52572;
  assign n52566 = n50492 ^ n42880;
  assign n52567 = n52566 ^ n46883;
  assign n52568 = n52567 ^ n41444;
  assign n52633 = n52612 ^ n52568;
  assign n52484 = n52483 ^ n52459;
  assign n52485 = n52460 & n52484;
  assign n52486 = n52485 ^ n49185;
  assign n52448 = n52447 ^ n52347;
  assign n52449 = ~n52445 & n52448;
  assign n52450 = n52449 ^ n52447;
  assign n52414 = n50517 ^ n49840;
  assign n52415 = n52414 ^ n51221;
  assign n52456 = n52450 ^ n52415;
  assign n52342 = n51703 ^ n51534;
  assign n52457 = n52456 ^ n52342;
  assign n52458 = n52457 ^ n49190;
  assign n52503 = n52486 ^ n52458;
  assign n52502 = n52491 & ~n52501;
  assign n52565 = n52503 ^ n52502;
  assign n52634 = n52633 ^ n52565;
  assign n52635 = ~n52632 & n52634;
  assign n52638 = n52637 ^ n52635;
  assign n52569 = n52568 ^ n52565;
  assign n52613 = n52612 ^ n52565;
  assign n52614 = n52569 & ~n52613;
  assign n52615 = n52614 ^ n52568;
  assign n52504 = ~n52502 & n52503;
  assign n52487 = n52486 ^ n52457;
  assign n52488 = n52458 & ~n52487;
  assign n52489 = n52488 ^ n49190;
  assign n52416 = n52415 ^ n52342;
  assign n52451 = n52450 ^ n52342;
  assign n52452 = n52416 & n52451;
  assign n52453 = n52452 ^ n52415;
  assign n52411 = n50513 ^ n49858;
  assign n52412 = n52411 ^ n51228;
  assign n52337 = n51706 ^ n51529;
  assign n52413 = n52412 ^ n52337;
  assign n52454 = n52453 ^ n52413;
  assign n52455 = n52454 ^ n49171;
  assign n52490 = n52489 ^ n52455;
  assign n52560 = n52504 ^ n52490;
  assign n52564 = n52563 ^ n52560;
  assign n52639 = n52615 ^ n52564;
  assign n52640 = n52639 ^ n52637;
  assign n52641 = n52638 & n52640;
  assign n52642 = n52641 ^ n52635;
  assign n52628 = n51262 ^ n50366;
  assign n52629 = n52628 ^ n51795;
  assign n52795 = n52642 ^ n52629;
  assign n52616 = n52615 ^ n52560;
  assign n52617 = ~n52564 & n52616;
  assign n52618 = n52617 ^ n52563;
  assign n52556 = n50477 ^ n42874;
  assign n52557 = n52556 ^ n47069;
  assign n52558 = n52557 ^ n41433;
  assign n52626 = n52618 ^ n52558;
  assign n52513 = n52489 ^ n52454;
  assign n52514 = ~n52455 & ~n52513;
  assign n52515 = n52514 ^ n49171;
  assign n52509 = n52453 ^ n52412;
  assign n52510 = ~n52413 & ~n52509;
  assign n52511 = n52510 ^ n52337;
  assign n52506 = n50512 ^ n49836;
  assign n52507 = n52506 ^ n51220;
  assign n52334 = n51709 ^ n51524;
  assign n52508 = n52507 ^ n52334;
  assign n52512 = n52511 ^ n52508;
  assign n52516 = n52515 ^ n52512;
  assign n52517 = n52516 ^ n49167;
  assign n52505 = n52490 & ~n52504;
  assign n52555 = n52517 ^ n52505;
  assign n52627 = n52626 ^ n52555;
  assign n52796 = n52795 ^ n52627;
  assign n52797 = n52796 ^ n49732;
  assign n52798 = n52634 ^ n52632;
  assign n52799 = n49737 & ~n52798;
  assign n52800 = n52799 ^ n49735;
  assign n52801 = n52639 ^ n52638;
  assign n52802 = n52801 ^ n52799;
  assign n52803 = n52800 & n52802;
  assign n52804 = n52803 ^ n49735;
  assign n52805 = n52804 ^ n52796;
  assign n52806 = ~n52797 & n52805;
  assign n52807 = n52806 ^ n49732;
  assign n52559 = n52558 ^ n52555;
  assign n52619 = n52618 ^ n52555;
  assign n52620 = ~n52559 & n52619;
  assign n52621 = n52620 ^ n52558;
  assign n52527 = n52512 ^ n49167;
  assign n52528 = ~n52516 & ~n52527;
  assign n52529 = n52528 ^ n49167;
  assign n52523 = n50377 ^ n49745;
  assign n52524 = n52523 ^ n51218;
  assign n52522 = n51716 ^ n51713;
  assign n52525 = n52524 ^ n52522;
  assign n52519 = n52511 ^ n52334;
  assign n52520 = ~n52508 & ~n52519;
  assign n52521 = n52520 ^ n52507;
  assign n52526 = n52525 ^ n52521;
  assign n52530 = n52529 ^ n52526;
  assign n52531 = n52530 ^ n49200;
  assign n52518 = n52505 & ~n52517;
  assign n52553 = n52531 ^ n52518;
  assign n52550 = n50472 ^ n42868;
  assign n52551 = n52550 ^ n47063;
  assign n52552 = n52551 ^ n41429;
  assign n52554 = n52553 ^ n52552;
  assign n52649 = n52621 ^ n52554;
  assign n52646 = n50965 ^ n50569;
  assign n52647 = n52646 ^ n51791;
  assign n52793 = n52649 ^ n52647;
  assign n52630 = n52629 ^ n52627;
  assign n52643 = n52642 ^ n52627;
  assign n52644 = ~n52630 & n52643;
  assign n52645 = n52644 ^ n52629;
  assign n52794 = n52793 ^ n52645;
  assign n52808 = n52807 ^ n52794;
  assign n52897 = n52808 ^ n49728;
  assign n52894 = n52801 ^ n52800;
  assign n52895 = n52804 ^ n52797;
  assign n52896 = n52894 & n52895;
  assign n53055 = n52897 ^ n52896;
  assign n2256 = n2255 ^ n2204;
  assign n2290 = n2289 ^ n2256;
  assign n2300 = n2299 ^ n2290;
  assign n53056 = n53055 ^ n2300;
  assign n53060 = n52895 ^ n52894;
  assign n53057 = n50821 ^ n43362;
  assign n53058 = n53057 ^ n47481;
  assign n53059 = n53058 ^ n2281;
  assign n53061 = n53060 ^ n53059;
  assign n53065 = n51122 ^ n43622;
  assign n53066 = n53065 ^ n47737;
  assign n53067 = n53066 ^ n42312;
  assign n53068 = n52798 ^ n49737;
  assign n53069 = n53067 & ~n53068;
  assign n53062 = n50825 ^ n2100;
  assign n53063 = n53062 ^ n47476;
  assign n53064 = n53063 ^ n41698;
  assign n53070 = n53069 ^ n53064;
  assign n53071 = n53069 ^ n52894;
  assign n53072 = n53070 & ~n53071;
  assign n53073 = n53072 ^ n53064;
  assign n53074 = n53073 ^ n53060;
  assign n53075 = ~n53061 & n53074;
  assign n53076 = n53075 ^ n53059;
  assign n53077 = n53076 ^ n53055;
  assign n53078 = n53056 & ~n53077;
  assign n53079 = n53078 ^ n2300;
  assign n53051 = n50816 ^ n43356;
  assign n53052 = n53051 ^ n47471;
  assign n53053 = n53052 ^ n41712;
  assign n53226 = n53079 ^ n53053;
  assign n52654 = n50962 ^ n50577;
  assign n52655 = n52654 ^ n51787;
  assign n52648 = n52647 ^ n52645;
  assign n52650 = n52649 ^ n52645;
  assign n52651 = n52648 & ~n52650;
  assign n52652 = n52651 ^ n52647;
  assign n52622 = n52621 ^ n52553;
  assign n52623 = n52554 & ~n52622;
  assign n52624 = n52623 ^ n52552;
  assign n52543 = n52526 ^ n49200;
  assign n52544 = n52530 & n52543;
  assign n52545 = n52544 ^ n49200;
  assign n52546 = n52545 ^ n49208;
  assign n52539 = n52524 ^ n52521;
  assign n52540 = ~n52525 & n52539;
  assign n52541 = n52540 ^ n52521;
  assign n52536 = n50373 ^ n49741;
  assign n52537 = n52536 ^ n51215;
  assign n51739 = n51738 ^ n51719;
  assign n52538 = n52537 ^ n51739;
  assign n52542 = n52541 ^ n52538;
  assign n52547 = n52546 ^ n52542;
  assign n52533 = n50508 ^ n1868;
  assign n52534 = n52533 ^ n47059;
  assign n52535 = n52534 ^ n41424;
  assign n52548 = n52547 ^ n52535;
  assign n52532 = ~n52518 & n52531;
  assign n52549 = n52548 ^ n52532;
  assign n52625 = n52624 ^ n52549;
  assign n52653 = n52652 ^ n52625;
  assign n52813 = n52655 ^ n52653;
  assign n52809 = n52794 ^ n49728;
  assign n52810 = ~n52808 & ~n52809;
  assign n52811 = n52810 ^ n49728;
  assign n52812 = n52811 ^ n49727;
  assign n52899 = n52813 ^ n52812;
  assign n52898 = ~n52896 & ~n52897;
  assign n53050 = n52899 ^ n52898;
  assign n53227 = n53226 ^ n53050;
  assign n53224 = n51757 ^ n50952;
  assign n52693 = n52266 ^ n52198;
  assign n53225 = n53224 ^ n52693;
  assign n53228 = n53227 ^ n53225;
  assign n53231 = n53076 ^ n2300;
  assign n53232 = n53231 ^ n53055;
  assign n52380 = n52263 ^ n52203;
  assign n53229 = n52380 ^ n51291;
  assign n53230 = n53229 ^ n51763;
  assign n53233 = n53232 ^ n53230;
  assign n53236 = n53073 ^ n53059;
  assign n53237 = n53236 ^ n53060;
  assign n53234 = n51765 ^ n50956;
  assign n52683 = n52260 ^ n52208;
  assign n53235 = n53234 ^ n52683;
  assign n53238 = n53237 ^ n53235;
  assign n53241 = n53064 ^ n52894;
  assign n53242 = n53241 ^ n53069;
  assign n52384 = n52257 ^ n52211;
  assign n52385 = n52384 ^ n52212;
  assign n53239 = n52385 ^ n51281;
  assign n53240 = n53239 ^ n51771;
  assign n53243 = n53242 ^ n53240;
  assign n53246 = n53068 ^ n53067;
  assign n52389 = n52254 ^ n52251;
  assign n53244 = n52389 ^ n50960;
  assign n53245 = n53244 ^ n51773;
  assign n53247 = n53246 ^ n53245;
  assign n53169 = n52598 ^ n52595;
  assign n53167 = n51218 ^ n50513;
  assign n53168 = n53167 ^ n51929;
  assign n53170 = n53169 ^ n53168;
  assign n52747 = n52591 ^ n52588;
  assign n52744 = n51922 ^ n50517;
  assign n52745 = n52744 ^ n51220;
  assign n53171 = n52747 ^ n52745;
  assign n52329 = n52328 ^ n52308;
  assign n51740 = n51739 ^ n50518;
  assign n51741 = n51740 ^ n51228;
  assign n52330 = n52329 ^ n51741;
  assign n52333 = n51870 ^ n51119;
  assign n52335 = n52334 ^ n52333;
  assign n52332 = n52298 ^ n52150;
  assign n52336 = n52335 ^ n52332;
  assign n52340 = n52295 ^ n52155;
  assign n52338 = n52337 ^ n50352;
  assign n52339 = n52338 ^ n51831;
  assign n52341 = n52340 ^ n52339;
  assign n52345 = n52292 ^ n52160;
  assign n52343 = n52342 ^ n50933;
  assign n52344 = n52343 ^ n51822;
  assign n52346 = n52345 ^ n52344;
  assign n52350 = n52289 ^ n52163;
  assign n52351 = n52350 ^ n52164;
  assign n52348 = n52347 ^ n51807;
  assign n52349 = n52348 ^ n50984;
  assign n52352 = n52351 ^ n52349;
  assign n52356 = n52286 ^ n52170;
  assign n52353 = n51811 ^ n50985;
  assign n52355 = n52354 ^ n52353;
  assign n52357 = n52356 ^ n52355;
  assign n52361 = n52283 ^ n52173;
  assign n52362 = n52361 ^ n52174;
  assign n52359 = n52358 ^ n50938;
  assign n52360 = n52359 ^ n51729;
  assign n52363 = n52362 ^ n52360;
  assign n52367 = n52280 ^ n52180;
  assign n52364 = n50986 ^ n50931;
  assign n52366 = n52365 ^ n52364;
  assign n52368 = n52367 ^ n52366;
  assign n52706 = n52277 ^ n52183;
  assign n52707 = n52706 ^ n52275;
  assign n52371 = n52272 ^ n52188;
  assign n52369 = n52319 ^ n51335;
  assign n52370 = n52369 ^ n50994;
  assign n52372 = n52371 ^ n52370;
  assign n52373 = n51328 ^ n50944;
  assign n52374 = n52373 ^ n51744;
  assign n52377 = n52376 ^ n52374;
  assign n52378 = n51749 ^ n51318;
  assign n52379 = n52378 ^ n50921;
  assign n52381 = n52380 ^ n52379;
  assign n52382 = n51304 ^ n50702;
  assign n52383 = n52382 ^ n51757;
  assign n52386 = n52385 ^ n52383;
  assign n52387 = n50946 ^ n50608;
  assign n52388 = n52387 ^ n51763;
  assign n52390 = n52389 ^ n52388;
  assign n52393 = n52247 ^ n52217;
  assign n52394 = n52393 ^ n52218;
  assign n52391 = n50952 ^ n50354;
  assign n52392 = n52391 ^ n51765;
  assign n52395 = n52394 ^ n52392;
  assign n52399 = n50956 ^ n50361;
  assign n52400 = n52399 ^ n51773;
  assign n52398 = n52241 ^ n52240;
  assign n52401 = n52400 ^ n52398;
  assign n52404 = n51281 ^ n50364;
  assign n52405 = n52404 ^ n51779;
  assign n52402 = n52235 ^ n52113;
  assign n52403 = n52402 ^ n52232;
  assign n52406 = n52405 ^ n52403;
  assign n52409 = n52231 ^ n52228;
  assign n52407 = n50960 ^ n50365;
  assign n52408 = n52407 ^ n51783;
  assign n52410 = n52409 ^ n52408;
  assign n52656 = n52655 ^ n52625;
  assign n52657 = n52653 & n52656;
  assign n52658 = n52657 ^ n52655;
  assign n52659 = n52658 ^ n52409;
  assign n52660 = ~n52410 & n52659;
  assign n52661 = n52660 ^ n52408;
  assign n52662 = n52661 ^ n52403;
  assign n52663 = n52406 & n52662;
  assign n52664 = n52663 ^ n52405;
  assign n52665 = n52664 ^ n52400;
  assign n52666 = ~n52401 & ~n52665;
  assign n52667 = n52666 ^ n52398;
  assign n52396 = n52244 ^ n52222;
  assign n52397 = n52396 ^ n52223;
  assign n52668 = n52667 ^ n52397;
  assign n52669 = n51291 ^ n50358;
  assign n52670 = n52669 ^ n51771;
  assign n52671 = n52670 ^ n52397;
  assign n52672 = ~n52668 & ~n52671;
  assign n52673 = n52672 ^ n52670;
  assign n52674 = n52673 ^ n52394;
  assign n52675 = n52395 & n52674;
  assign n52676 = n52675 ^ n52392;
  assign n52677 = n52676 ^ n52389;
  assign n52678 = n52390 & n52677;
  assign n52679 = n52678 ^ n52388;
  assign n52680 = n52679 ^ n52383;
  assign n52681 = n52386 & n52680;
  assign n52682 = n52681 ^ n52385;
  assign n52684 = n52683 ^ n52682;
  assign n52685 = n51311 ^ n50751;
  assign n52686 = n52685 ^ n51755;
  assign n52687 = n52686 ^ n52683;
  assign n52688 = ~n52684 & n52687;
  assign n52689 = n52688 ^ n52686;
  assign n52690 = n52689 ^ n52380;
  assign n52691 = n52381 & n52690;
  assign n52692 = n52691 ^ n52379;
  assign n52694 = n52693 ^ n52692;
  assign n52695 = n51745 ^ n50941;
  assign n52696 = n52695 ^ n50950;
  assign n52697 = n52696 ^ n52693;
  assign n52698 = n52694 & n52697;
  assign n52699 = n52698 ^ n52696;
  assign n52700 = n52699 ^ n52376;
  assign n52701 = n52377 & n52700;
  assign n52702 = n52701 ^ n52374;
  assign n52703 = n52702 ^ n52370;
  assign n52704 = n52372 & n52703;
  assign n52705 = n52704 ^ n52371;
  assign n52708 = n52707 ^ n52705;
  assign n52709 = n52428 ^ n50990;
  assign n52710 = n52709 ^ n50935;
  assign n52711 = n52710 ^ n52707;
  assign n52712 = n52708 & ~n52711;
  assign n52713 = n52712 ^ n52710;
  assign n52714 = n52713 ^ n52367;
  assign n52715 = ~n52368 & ~n52714;
  assign n52716 = n52715 ^ n52366;
  assign n52717 = n52716 ^ n52362;
  assign n52718 = n52363 & n52717;
  assign n52719 = n52718 ^ n52360;
  assign n52720 = n52719 ^ n52355;
  assign n52721 = ~n52357 & ~n52720;
  assign n52722 = n52721 ^ n52356;
  assign n52723 = n52722 ^ n52351;
  assign n52724 = n52352 & ~n52723;
  assign n52725 = n52724 ^ n52349;
  assign n52726 = n52725 ^ n52345;
  assign n52727 = n52346 & ~n52726;
  assign n52728 = n52727 ^ n52344;
  assign n52729 = n52728 ^ n52340;
  assign n52730 = ~n52341 & n52729;
  assign n52731 = n52730 ^ n52339;
  assign n52732 = n52731 ^ n52335;
  assign n52733 = n52336 & ~n52732;
  assign n52734 = n52733 ^ n52332;
  assign n52331 = n52305 ^ n52302;
  assign n52735 = n52734 ^ n52331;
  assign n52736 = n51221 ^ n50522;
  assign n52737 = n52736 ^ n52522;
  assign n52738 = n52737 ^ n52331;
  assign n52739 = n52735 & n52738;
  assign n52740 = n52739 ^ n52737;
  assign n52741 = n52740 ^ n52329;
  assign n52742 = n52330 & ~n52741;
  assign n52743 = n52742 ^ n51741;
  assign n53172 = n52747 ^ n52743;
  assign n53173 = n53171 & n53172;
  assign n53174 = n53173 ^ n52745;
  assign n53264 = n53174 ^ n53169;
  assign n53265 = n53170 & ~n53264;
  assign n53266 = n53265 ^ n53168;
  assign n53261 = n51920 ^ n51215;
  assign n53262 = n53261 ^ n50512;
  assign n53276 = n53266 ^ n53262;
  assign n53260 = n52601 ^ n52582;
  assign n53277 = n53276 ^ n53260;
  assign n53278 = n53277 ^ n49836;
  assign n53175 = n53174 ^ n53170;
  assign n53176 = n53175 ^ n49858;
  assign n52750 = n52740 ^ n52330;
  assign n52751 = n52750 ^ n49847;
  assign n52752 = n52737 ^ n52735;
  assign n52753 = n52752 ^ n49703;
  assign n52754 = n52731 ^ n52336;
  assign n52755 = n52754 ^ n50460;
  assign n52756 = n52728 ^ n52339;
  assign n52757 = n52756 ^ n52340;
  assign n52758 = n52757 ^ n50442;
  assign n52759 = n52725 ^ n52346;
  assign n52760 = n52759 ^ n50382;
  assign n52761 = n52722 ^ n52349;
  assign n52762 = n52761 ^ n52351;
  assign n52763 = n52762 ^ n50383;
  assign n52764 = n52719 ^ n52357;
  assign n52765 = n52764 ^ n50385;
  assign n52766 = n52716 ^ n52363;
  assign n52767 = n52766 ^ n50386;
  assign n52768 = n52713 ^ n52366;
  assign n52769 = n52768 ^ n52367;
  assign n52770 = n52769 ^ n50343;
  assign n52772 = n52702 ^ n52372;
  assign n52773 = n52772 ^ n50121;
  assign n52774 = n52699 ^ n52377;
  assign n52775 = n52774 ^ n50061;
  assign n52776 = n52696 ^ n52694;
  assign n52777 = n52776 ^ n49944;
  assign n52778 = n52689 ^ n52379;
  assign n52779 = n52778 ^ n52380;
  assign n52780 = n52779 ^ n49708;
  assign n52781 = n52686 ^ n52684;
  assign n52782 = n52781 ^ n49709;
  assign n52783 = n52679 ^ n52386;
  assign n52784 = n52783 ^ n49715;
  assign n52787 = n52673 ^ n52395;
  assign n52788 = n52787 ^ n49918;
  assign n52789 = n52670 ^ n52668;
  assign n52790 = n52789 ^ n49911;
  assign n52791 = n52661 ^ n52406;
  assign n52792 = n52791 ^ n49901;
  assign n52814 = n52813 ^ n52811;
  assign n52815 = n52812 & n52814;
  assign n52816 = n52815 ^ n49727;
  assign n52817 = n52816 ^ n49725;
  assign n52818 = n52658 ^ n52410;
  assign n52819 = n52818 ^ n52816;
  assign n52820 = ~n52817 & n52819;
  assign n52821 = n52820 ^ n49725;
  assign n52822 = n52821 ^ n52791;
  assign n52823 = n52792 & n52822;
  assign n52824 = n52823 ^ n49901;
  assign n52825 = n52824 ^ n49721;
  assign n52826 = n52664 ^ n52401;
  assign n52827 = n52826 ^ n52824;
  assign n52828 = ~n52825 & ~n52827;
  assign n52829 = n52828 ^ n49721;
  assign n52830 = n52829 ^ n52789;
  assign n52831 = n52790 & ~n52830;
  assign n52832 = n52831 ^ n49911;
  assign n52833 = n52832 ^ n52787;
  assign n52834 = ~n52788 & ~n52833;
  assign n52835 = n52834 ^ n49918;
  assign n52785 = n52676 ^ n52388;
  assign n52786 = n52785 ^ n52389;
  assign n52836 = n52835 ^ n52786;
  assign n52837 = n52786 ^ n49718;
  assign n52838 = ~n52836 & ~n52837;
  assign n52839 = n52838 ^ n49718;
  assign n52840 = n52839 ^ n52783;
  assign n52841 = ~n52784 & ~n52840;
  assign n52842 = n52841 ^ n49715;
  assign n52843 = n52842 ^ n52781;
  assign n52844 = ~n52782 & ~n52843;
  assign n52845 = n52844 ^ n49709;
  assign n52846 = n52845 ^ n52779;
  assign n52847 = n52780 & n52846;
  assign n52848 = n52847 ^ n49708;
  assign n52849 = n52848 ^ n52776;
  assign n52850 = ~n52777 & n52849;
  assign n52851 = n52850 ^ n49944;
  assign n52852 = n52851 ^ n52774;
  assign n52853 = n52775 & ~n52852;
  assign n52854 = n52853 ^ n50061;
  assign n52855 = n52854 ^ n52772;
  assign n52856 = ~n52773 & n52855;
  assign n52857 = n52856 ^ n50121;
  assign n52771 = n52710 ^ n52708;
  assign n52858 = n52857 ^ n52771;
  assign n52859 = n52771 ^ n50136;
  assign n52860 = n52858 & ~n52859;
  assign n52861 = n52860 ^ n50136;
  assign n52862 = n52861 ^ n52769;
  assign n52863 = n52770 & n52862;
  assign n52864 = n52863 ^ n50343;
  assign n52865 = n52864 ^ n52766;
  assign n52866 = n52767 & ~n52865;
  assign n52867 = n52866 ^ n50386;
  assign n52868 = n52867 ^ n52764;
  assign n52869 = n52765 & ~n52868;
  assign n52870 = n52869 ^ n50385;
  assign n52871 = n52870 ^ n52762;
  assign n52872 = ~n52763 & ~n52871;
  assign n52873 = n52872 ^ n50383;
  assign n52874 = n52873 ^ n52759;
  assign n52875 = n52760 & n52874;
  assign n52876 = n52875 ^ n50382;
  assign n52877 = n52876 ^ n52757;
  assign n52878 = n52758 & n52877;
  assign n52879 = n52878 ^ n50442;
  assign n52880 = n52879 ^ n52754;
  assign n52881 = ~n52755 & n52880;
  assign n52882 = n52881 ^ n50460;
  assign n52883 = n52882 ^ n52752;
  assign n52884 = ~n52753 & n52883;
  assign n52885 = n52884 ^ n49703;
  assign n52886 = n52885 ^ n52750;
  assign n52887 = n52751 & ~n52886;
  assign n52888 = n52887 ^ n49847;
  assign n53163 = n52888 ^ n49840;
  assign n52746 = n52745 ^ n52743;
  assign n52748 = n52747 ^ n52746;
  assign n53164 = n52888 ^ n52748;
  assign n53165 = ~n53163 & ~n53164;
  assign n53166 = n53165 ^ n49840;
  assign n53279 = n53175 ^ n53166;
  assign n53280 = ~n53176 & ~n53279;
  assign n53281 = n53280 ^ n49858;
  assign n53282 = n53281 ^ n53277;
  assign n53283 = n53278 & n53282;
  assign n53284 = n53283 ^ n49836;
  assign n53263 = n53262 ^ n53260;
  assign n53267 = n53266 ^ n53260;
  assign n53268 = n53263 & ~n53267;
  assign n53269 = n53268 ^ n53262;
  assign n53258 = n52604 ^ n52577;
  assign n53256 = n51937 ^ n50978;
  assign n53257 = n53256 ^ n50377;
  assign n53259 = n53258 ^ n53257;
  assign n53274 = n53269 ^ n53259;
  assign n53275 = n53274 ^ n49745;
  assign n53293 = n53284 ^ n53275;
  assign n53177 = n53176 ^ n53166;
  assign n52749 = n52748 ^ n49840;
  assign n52889 = n52888 ^ n52749;
  assign n52890 = n52876 ^ n52758;
  assign n52891 = n52867 ^ n52765;
  assign n52892 = n52826 ^ n52825;
  assign n52893 = n52818 ^ n52817;
  assign n52900 = ~n52898 & ~n52899;
  assign n52901 = ~n52893 & ~n52900;
  assign n52902 = n52821 ^ n52792;
  assign n52903 = ~n52901 & ~n52902;
  assign n52904 = ~n52892 & n52903;
  assign n52905 = n52829 ^ n49911;
  assign n52906 = n52905 ^ n52789;
  assign n52907 = n52904 & ~n52906;
  assign n52908 = n52832 ^ n52788;
  assign n52909 = ~n52907 & ~n52908;
  assign n52910 = n52836 ^ n49718;
  assign n52911 = n52909 & n52910;
  assign n52912 = n52839 ^ n52784;
  assign n52913 = n52911 & ~n52912;
  assign n52914 = n52842 ^ n52782;
  assign n52915 = n52913 & n52914;
  assign n52916 = n52845 ^ n52780;
  assign n52917 = n52915 & n52916;
  assign n52918 = n52848 ^ n49944;
  assign n52919 = n52918 ^ n52776;
  assign n52920 = ~n52917 & ~n52919;
  assign n52921 = n52851 ^ n50061;
  assign n52922 = n52921 ^ n52774;
  assign n52923 = n52920 & n52922;
  assign n52924 = n52854 ^ n50121;
  assign n52925 = n52924 ^ n52772;
  assign n52926 = ~n52923 & n52925;
  assign n52927 = n52858 ^ n50136;
  assign n52928 = ~n52926 & ~n52927;
  assign n52929 = n52861 ^ n52770;
  assign n52930 = ~n52928 & ~n52929;
  assign n52931 = n52864 ^ n52767;
  assign n52932 = n52930 & n52931;
  assign n52933 = n52891 & n52932;
  assign n52934 = n52870 ^ n52763;
  assign n52935 = ~n52933 & n52934;
  assign n52936 = n52873 ^ n52760;
  assign n52937 = n52935 & n52936;
  assign n52938 = n52890 & ~n52937;
  assign n52939 = n52879 ^ n50460;
  assign n52940 = n52939 ^ n52754;
  assign n52941 = n52938 & n52940;
  assign n52942 = n52882 ^ n52753;
  assign n52943 = ~n52941 & ~n52942;
  assign n52944 = n52885 ^ n52751;
  assign n52945 = ~n52943 & ~n52944;
  assign n53178 = ~n52889 & ~n52945;
  assign n53290 = ~n53177 & ~n53178;
  assign n53291 = n53281 ^ n53278;
  assign n53292 = n53290 & ~n53291;
  assign n53300 = n53293 ^ n53292;
  assign n53297 = n51138 ^ n43632;
  assign n53298 = n53297 ^ n47768;
  assign n53299 = n53298 ^ n42150;
  assign n53301 = n53300 ^ n53299;
  assign n53305 = n53291 ^ n53290;
  assign n53302 = n51201 ^ n42300;
  assign n53303 = n53302 ^ n47747;
  assign n53304 = n53303 ^ n43637;
  assign n53306 = n53305 ^ n53304;
  assign n53179 = n53178 ^ n53177;
  assign n53160 = n51144 ^ n43651;
  assign n53161 = n53160 ^ n47758;
  assign n53162 = n53161 ^ n42293;
  assign n53180 = n53179 ^ n53162;
  assign n52946 = n52945 ^ n52889;
  assign n2967 = n2966 ^ n2939;
  assign n3004 = n3003 ^ n2967;
  assign n3011 = n3010 ^ n3004;
  assign n52947 = n52946 ^ n3011;
  assign n52954 = n52942 ^ n52941;
  assign n52951 = n51185 ^ n2862;
  assign n52952 = n52951 ^ n47407;
  assign n52953 = n52952 ^ n42160;
  assign n52955 = n52954 ^ n52953;
  assign n52957 = n51157 ^ n3227;
  assign n52958 = n52957 ^ n47587;
  assign n52959 = n52958 ^ n42166;
  assign n52956 = n52940 ^ n52938;
  assign n52960 = n52959 ^ n52956;
  assign n52964 = n52937 ^ n52890;
  assign n52961 = n51175 ^ n43456;
  assign n52962 = n52961 ^ n47413;
  assign n52963 = n52962 ^ n42170;
  assign n52965 = n52964 ^ n52963;
  assign n52969 = n52936 ^ n52935;
  assign n52966 = n47417 ^ n43292;
  assign n52967 = n52966 ^ n51163;
  assign n52968 = n52967 ^ n42175;
  assign n52970 = n52969 ^ n52968;
  assign n52974 = n52934 ^ n52933;
  assign n52971 = n50913 ^ n43297;
  assign n52972 = n52971 ^ n47574;
  assign n52973 = n52972 ^ n42180;
  assign n52975 = n52974 ^ n52973;
  assign n52979 = n52932 ^ n52891;
  assign n52976 = n50907 ^ n43303;
  assign n52977 = n52976 ^ n47567;
  assign n52978 = n52977 ^ n42185;
  assign n52980 = n52979 ^ n52978;
  assign n52982 = n50761 ^ n43307;
  assign n52983 = n52982 ^ n47560;
  assign n52984 = n52983 ^ n42261;
  assign n52981 = n52931 ^ n52930;
  assign n52985 = n52984 ^ n52981;
  assign n52989 = n52929 ^ n52928;
  assign n52986 = n50897 ^ n43437;
  assign n52987 = n52986 ^ n47553;
  assign n52988 = n52987 ^ n42192;
  assign n52990 = n52989 ^ n52988;
  assign n52994 = n52927 ^ n52926;
  assign n52991 = n50767 ^ n43430;
  assign n52992 = n52991 ^ n47546;
  assign n52993 = n52992 ^ n42251;
  assign n52995 = n52994 ^ n52993;
  assign n52999 = n52925 ^ n52923;
  assign n52996 = n50772 ^ n43314;
  assign n52997 = n52996 ^ n47427;
  assign n52998 = n52997 ^ n1217;
  assign n53000 = n52999 ^ n52998;
  assign n53004 = n52922 ^ n52920;
  assign n53001 = n50777 ^ n43319;
  assign n53002 = n53001 ^ n1079;
  assign n53003 = n53002 ^ n42241;
  assign n53005 = n53004 ^ n53003;
  assign n53010 = n52916 ^ n52915;
  assign n53007 = n50878 ^ n914;
  assign n53008 = n53007 ^ n47530;
  assign n53009 = n53008 ^ n42231;
  assign n53011 = n53010 ^ n53009;
  assign n53013 = n50789 ^ n43332;
  assign n53014 = n53013 ^ n47521;
  assign n53015 = n53014 ^ n42204;
  assign n53012 = n52914 ^ n52913;
  assign n53016 = n53015 ^ n53012;
  assign n53020 = n52912 ^ n52911;
  assign n53017 = n50794 ^ n43408;
  assign n53018 = n53017 ^ n47441;
  assign n53019 = n53018 ^ n42209;
  assign n53021 = n53020 ^ n53019;
  assign n53023 = n50865 ^ n43401;
  assign n53024 = n53023 ^ n47445;
  assign n53025 = n53024 ^ n42214;
  assign n53022 = n52910 ^ n52909;
  assign n53026 = n53025 ^ n53022;
  assign n53030 = n52908 ^ n52907;
  assign n53027 = n50799 ^ n43339;
  assign n53028 = n53027 ^ n47450;
  assign n53029 = n53028 ^ n41119;
  assign n53031 = n53030 ^ n53029;
  assign n53035 = n52906 ^ n52904;
  assign n53032 = n50855 ^ n43391;
  assign n53033 = n53032 ^ n47455;
  assign n53034 = n53033 ^ n41676;
  assign n53036 = n53035 ^ n53034;
  assign n53040 = n52903 ^ n52892;
  assign n53037 = n50805 ^ n43344;
  assign n53038 = n53037 ^ n47461;
  assign n53039 = n53038 ^ n41681;
  assign n53041 = n53040 ^ n53039;
  assign n53043 = n50845 ^ n43381;
  assign n53044 = n53043 ^ n47466;
  assign n53045 = n53044 ^ n41687;
  assign n53042 = n52902 ^ n52901;
  assign n53046 = n53045 ^ n53042;
  assign n53054 = n53053 ^ n53050;
  assign n53080 = n53079 ^ n53050;
  assign n53081 = ~n53054 & n53080;
  assign n53082 = n53081 ^ n53053;
  assign n53047 = n50811 ^ n43351;
  assign n53048 = n53047 ^ n47497;
  assign n53049 = n53048 ^ n41692;
  assign n53083 = n53082 ^ n53049;
  assign n53084 = n52900 ^ n52893;
  assign n53085 = n53084 ^ n53082;
  assign n53086 = n53083 & ~n53085;
  assign n53087 = n53086 ^ n53049;
  assign n53088 = n53087 ^ n53042;
  assign n53089 = ~n53046 & n53088;
  assign n53090 = n53089 ^ n53045;
  assign n53091 = n53090 ^ n53040;
  assign n53092 = n53041 & ~n53091;
  assign n53093 = n53092 ^ n53039;
  assign n53094 = n53093 ^ n53035;
  assign n53095 = n53036 & ~n53094;
  assign n53096 = n53095 ^ n53034;
  assign n53097 = n53096 ^ n53030;
  assign n53098 = n53031 & ~n53097;
  assign n53099 = n53098 ^ n53029;
  assign n53100 = n53099 ^ n53022;
  assign n53101 = n53026 & ~n53100;
  assign n53102 = n53101 ^ n53025;
  assign n53103 = n53102 ^ n53020;
  assign n53104 = ~n53021 & n53103;
  assign n53105 = n53104 ^ n53019;
  assign n53106 = n53105 ^ n53012;
  assign n53107 = n53016 & ~n53106;
  assign n53108 = n53107 ^ n53015;
  assign n53109 = n53108 ^ n53010;
  assign n53110 = n53011 & ~n53109;
  assign n53111 = n53110 ^ n53009;
  assign n53006 = n52919 ^ n52917;
  assign n53112 = n53111 ^ n53006;
  assign n53113 = n50782 ^ n43324;
  assign n53114 = n53113 ^ n47434;
  assign n53115 = n53114 ^ n1068;
  assign n53116 = n53115 ^ n53006;
  assign n53117 = n53112 & ~n53116;
  assign n53118 = n53117 ^ n53115;
  assign n53119 = n53118 ^ n53004;
  assign n53120 = ~n53005 & n53119;
  assign n53121 = n53120 ^ n53003;
  assign n53122 = n53121 ^ n52999;
  assign n53123 = ~n53000 & n53122;
  assign n53124 = n53123 ^ n52998;
  assign n53125 = n53124 ^ n52994;
  assign n53126 = ~n52995 & n53125;
  assign n53127 = n53126 ^ n52993;
  assign n53128 = n53127 ^ n52989;
  assign n53129 = n52990 & ~n53128;
  assign n53130 = n53129 ^ n52988;
  assign n53131 = n53130 ^ n52984;
  assign n53132 = n52985 & ~n53131;
  assign n53133 = n53132 ^ n52981;
  assign n53134 = n53133 ^ n52979;
  assign n53135 = n52980 & ~n53134;
  assign n53136 = n53135 ^ n52978;
  assign n53137 = n53136 ^ n52974;
  assign n53138 = n52975 & ~n53137;
  assign n53139 = n53138 ^ n52973;
  assign n53140 = n53139 ^ n52969;
  assign n53141 = ~n52970 & n53140;
  assign n53142 = n53141 ^ n52968;
  assign n53143 = n53142 ^ n52964;
  assign n53144 = ~n52965 & n53143;
  assign n53145 = n53144 ^ n52963;
  assign n53146 = n53145 ^ n52959;
  assign n53147 = n52960 & ~n53146;
  assign n53148 = n53147 ^ n52956;
  assign n53149 = n53148 ^ n52954;
  assign n53150 = ~n52955 & n53149;
  assign n53151 = n53150 ^ n52953;
  assign n52948 = n51151 ^ n43483;
  assign n52949 = n52948 ^ n47401;
  assign n52950 = n52949 ^ n2995;
  assign n53152 = n53151 ^ n52950;
  assign n53153 = n52944 ^ n52943;
  assign n53154 = n53153 ^ n53151;
  assign n53155 = n53152 & ~n53154;
  assign n53156 = n53155 ^ n52950;
  assign n53157 = n53156 ^ n52946;
  assign n53158 = ~n52947 & n53157;
  assign n53159 = n53158 ^ n3011;
  assign n53307 = n53179 ^ n53159;
  assign n53308 = n53180 & ~n53307;
  assign n53309 = n53308 ^ n53162;
  assign n53310 = n53309 ^ n53305;
  assign n53311 = ~n53306 & n53310;
  assign n53312 = n53311 ^ n53304;
  assign n53313 = n53312 ^ n53300;
  assign n53314 = n53301 & ~n53313;
  assign n53315 = n53314 ^ n53299;
  assign n53294 = ~n53292 & n53293;
  assign n53285 = n53284 ^ n53274;
  assign n53286 = ~n53275 & ~n53285;
  assign n53287 = n53286 ^ n49745;
  assign n53270 = n53269 ^ n53258;
  assign n53271 = n53259 & ~n53270;
  assign n53272 = n53271 ^ n53257;
  assign n53254 = n52609 ^ n52608;
  assign n53253 = n52536 ^ n50974;
  assign n53255 = n53254 ^ n53253;
  assign n53273 = n53272 ^ n53255;
  assign n53288 = n53287 ^ n53273;
  assign n53289 = n53288 ^ n51913;
  assign n53295 = n53294 ^ n53289;
  assign n53250 = n51211 ^ n43627;
  assign n53251 = n53250 ^ n47741;
  assign n53252 = n53251 ^ n42146;
  assign n53296 = n53295 ^ n53252;
  assign n53316 = n53315 ^ n53296;
  assign n53248 = n51779 ^ n50962;
  assign n53249 = n53248 ^ n52394;
  assign n53317 = n53316 ^ n53249;
  assign n53320 = n52397 ^ n50965;
  assign n53321 = n53320 ^ n51783;
  assign n53318 = n53312 ^ n53299;
  assign n53319 = n53318 ^ n53300;
  assign n53322 = n53321 ^ n53319;
  assign n53325 = n53309 ^ n53304;
  assign n53326 = n53325 ^ n53305;
  assign n53323 = n52398 ^ n51787;
  assign n53324 = n53323 ^ n51262;
  assign n53327 = n53326 ^ n53324;
  assign n53332 = n52403 ^ n50969;
  assign n53333 = n53332 ^ n51791;
  assign n53328 = n53156 ^ n52947;
  assign n53329 = n51795 ^ n50972;
  assign n53330 = n53329 ^ n52409;
  assign n53331 = ~n53328 & n53330;
  assign n53334 = n53333 ^ n53331;
  assign n53181 = n53180 ^ n53159;
  assign n53335 = n53333 ^ n53181;
  assign n53336 = n53334 & ~n53335;
  assign n53337 = n53336 ^ n53331;
  assign n53338 = n53337 ^ n53326;
  assign n53339 = ~n53327 & n53338;
  assign n53340 = n53339 ^ n53324;
  assign n53341 = n53340 ^ n53321;
  assign n53342 = n53322 & ~n53341;
  assign n53343 = n53342 ^ n53319;
  assign n53344 = n53343 ^ n53316;
  assign n53345 = ~n53317 & n53344;
  assign n53346 = n53345 ^ n53249;
  assign n53347 = n53346 ^ n53246;
  assign n53348 = ~n53247 & n53347;
  assign n53349 = n53348 ^ n53245;
  assign n53350 = n53349 ^ n53242;
  assign n53351 = n53243 & ~n53350;
  assign n53352 = n53351 ^ n53240;
  assign n53353 = n53352 ^ n53237;
  assign n53354 = ~n53238 & n53353;
  assign n53355 = n53354 ^ n53235;
  assign n53356 = n53355 ^ n53232;
  assign n53357 = ~n53233 & ~n53356;
  assign n53358 = n53357 ^ n53230;
  assign n53359 = n53358 ^ n53227;
  assign n53360 = n53228 & ~n53359;
  assign n53361 = n53360 ^ n53225;
  assign n53223 = n53084 ^ n53083;
  assign n53362 = n53361 ^ n53223;
  assign n53432 = n53364 ^ n53362;
  assign n53433 = n53432 ^ n50608;
  assign n53437 = n53349 ^ n53243;
  assign n53438 = n53437 ^ n50364;
  assign n53439 = n53346 ^ n53245;
  assign n53440 = n53439 ^ n53246;
  assign n53441 = n53440 ^ n50365;
  assign n53442 = n53343 ^ n53317;
  assign n53443 = n53442 ^ n50577;
  assign n53444 = n53340 ^ n53322;
  assign n53445 = n53444 ^ n50569;
  assign n53446 = n53337 ^ n53324;
  assign n53447 = n53446 ^ n53326;
  assign n53448 = n53447 ^ n50366;
  assign n53449 = n53330 ^ n53328;
  assign n53450 = ~n50369 & ~n53449;
  assign n53451 = n53450 ^ n50368;
  assign n53452 = n53334 ^ n53181;
  assign n53453 = n53452 ^ n53450;
  assign n53454 = ~n53451 & ~n53453;
  assign n53455 = n53454 ^ n50368;
  assign n53456 = n53455 ^ n53447;
  assign n53457 = ~n53448 & ~n53456;
  assign n53458 = n53457 ^ n50366;
  assign n53459 = n53458 ^ n53444;
  assign n53460 = ~n53445 & ~n53459;
  assign n53461 = n53460 ^ n50569;
  assign n53462 = n53461 ^ n53442;
  assign n53463 = ~n53443 & ~n53462;
  assign n53464 = n53463 ^ n50577;
  assign n53465 = n53464 ^ n53440;
  assign n53466 = ~n53441 & n53465;
  assign n53467 = n53466 ^ n50365;
  assign n53468 = n53467 ^ n53437;
  assign n53469 = ~n53438 & ~n53468;
  assign n53470 = n53469 ^ n50364;
  assign n53436 = n53352 ^ n53238;
  assign n53471 = n53470 ^ n53436;
  assign n53472 = n53436 ^ n50361;
  assign n53473 = ~n53471 & n53472;
  assign n53474 = n53473 ^ n50361;
  assign n53475 = n53474 ^ n50358;
  assign n53476 = n53355 ^ n53233;
  assign n53477 = n53476 ^ n53474;
  assign n53478 = ~n53475 & ~n53477;
  assign n53479 = n53478 ^ n50358;
  assign n53434 = n53358 ^ n53225;
  assign n53435 = n53434 ^ n53227;
  assign n53480 = n53479 ^ n53435;
  assign n53481 = n53435 ^ n50354;
  assign n53482 = n53480 & ~n53481;
  assign n53483 = n53482 ^ n50354;
  assign n53484 = n53483 ^ n53432;
  assign n53485 = n53433 & n53484;
  assign n53486 = n53485 ^ n50608;
  assign n53365 = n53364 ^ n53223;
  assign n53366 = n53362 & n53365;
  assign n53367 = n53366 ^ n53364;
  assign n53220 = n51749 ^ n51304;
  assign n53221 = n53220 ^ n52371;
  assign n53219 = n53087 ^ n53046;
  assign n53222 = n53221 ^ n53219;
  assign n53431 = n53367 ^ n53222;
  assign n53487 = n53486 ^ n53431;
  assign n53488 = n53431 ^ n50702;
  assign n53489 = n53487 & n53488;
  assign n53490 = n53489 ^ n50702;
  assign n53368 = n53367 ^ n53221;
  assign n53369 = n53222 & n53368;
  assign n53370 = n53369 ^ n53219;
  assign n53217 = n53090 ^ n53041;
  assign n53215 = n51745 ^ n51311;
  assign n53216 = n53215 ^ n52707;
  assign n53218 = n53217 ^ n53216;
  assign n53430 = n53370 ^ n53218;
  assign n53491 = n53490 ^ n53430;
  assign n53492 = n53430 ^ n50751;
  assign n53493 = ~n53491 & n53492;
  assign n53494 = n53493 ^ n50751;
  assign n53371 = n53370 ^ n53217;
  assign n53372 = ~n53218 & n53371;
  assign n53373 = n53372 ^ n53216;
  assign n53213 = n53093 ^ n53036;
  assign n53211 = n52367 ^ n51318;
  assign n53212 = n53211 ^ n51744;
  assign n53214 = n53213 ^ n53212;
  assign n53428 = n53373 ^ n53214;
  assign n53429 = n53428 ^ n50921;
  assign n53550 = n53494 ^ n53429;
  assign n53525 = n53487 ^ n50702;
  assign n53526 = n53464 ^ n53441;
  assign n53527 = n53452 ^ n53451;
  assign n53528 = n53455 ^ n53448;
  assign n53529 = n53527 & ~n53528;
  assign n53530 = n53458 ^ n53445;
  assign n53531 = ~n53529 & ~n53530;
  assign n53532 = n53461 ^ n53443;
  assign n53533 = ~n53531 & ~n53532;
  assign n53534 = ~n53526 & ~n53533;
  assign n53535 = n53467 ^ n50364;
  assign n53536 = n53535 ^ n53437;
  assign n53537 = ~n53534 & n53536;
  assign n53538 = n53471 ^ n50361;
  assign n53539 = n53537 & n53538;
  assign n53540 = n53476 ^ n50358;
  assign n53541 = n53540 ^ n53474;
  assign n53542 = n53539 & ~n53541;
  assign n53543 = n53480 ^ n50354;
  assign n53544 = ~n53542 & ~n53543;
  assign n53545 = n53483 ^ n53433;
  assign n53546 = n53544 & n53545;
  assign n53547 = ~n53525 & n53546;
  assign n53548 = n53491 ^ n50751;
  assign n53549 = n53547 & n53548;
  assign n53593 = n53550 ^ n53549;
  assign n53590 = n51573 ^ n43967;
  assign n53591 = n53590 ^ n48095;
  assign n53592 = n53591 ^ n42486;
  assign n53594 = n53593 ^ n53592;
  assign n53599 = n53546 ^ n53525;
  assign n53596 = n51583 ^ n43977;
  assign n53597 = n53596 ^ n48105;
  assign n53598 = n53597 ^ n42495;
  assign n53600 = n53599 ^ n53598;
  assign n53602 = n51658 ^ n44046;
  assign n53603 = n53602 ^ n48110;
  assign n53604 = n53603 ^ n42570;
  assign n53601 = n53545 ^ n53544;
  assign n53605 = n53604 ^ n53601;
  assign n53609 = n53543 ^ n53542;
  assign n53606 = n51589 ^ n44039;
  assign n53607 = n53606 ^ n48116;
  assign n53608 = n53607 ^ n42502;
  assign n53610 = n53609 ^ n53608;
  assign n53614 = n53541 ^ n53539;
  assign n53611 = n51648 ^ n44032;
  assign n53612 = n53611 ^ n48120;
  assign n53613 = n53612 ^ n42560;
  assign n53615 = n53614 ^ n53613;
  assign n53617 = n51595 ^ n43986;
  assign n53618 = n53617 ^ n48125;
  assign n53619 = n53618 ^ n42508;
  assign n53616 = n53538 ^ n53537;
  assign n53620 = n53619 ^ n53616;
  assign n53622 = n51638 ^ n44022;
  assign n53623 = n53622 ^ n48130;
  assign n53624 = n53623 ^ n42550;
  assign n53621 = n53536 ^ n53534;
  assign n53625 = n53624 ^ n53621;
  assign n53639 = n51804 ^ n44243;
  assign n53640 = n53639 ^ n48381;
  assign n53641 = n53640 ^ n42849;
  assign n53642 = n53449 ^ n50369;
  assign n53643 = n53641 & n53642;
  assign n53636 = n51619 ^ n44003;
  assign n53637 = n53636 ^ n48149;
  assign n53638 = n53637 ^ n42529;
  assign n53644 = n53643 ^ n53638;
  assign n53645 = n53643 ^ n53527;
  assign n53646 = n53644 & ~n53645;
  assign n53647 = n53646 ^ n53638;
  assign n53633 = n51616 ^ n44000;
  assign n53634 = n53633 ^ n48153;
  assign n53635 = n53634 ^ n42533;
  assign n53648 = n53647 ^ n53635;
  assign n53649 = n53528 ^ n53527;
  assign n53650 = n53649 ^ n53647;
  assign n53651 = n53648 & ~n53650;
  assign n53652 = n53651 ^ n53635;
  assign n53630 = n51611 ^ n2389;
  assign n53631 = n53630 ^ n48145;
  assign n53632 = n53631 ^ n42523;
  assign n53653 = n53652 ^ n53632;
  assign n53654 = n53530 ^ n53529;
  assign n53655 = n53654 ^ n53652;
  assign n53656 = n53653 & ~n53655;
  assign n53657 = n53656 ^ n53632;
  assign n53627 = n51606 ^ n2407;
  assign n53628 = n53627 ^ n48140;
  assign n53629 = n53628 ^ n42518;
  assign n53658 = n53657 ^ n53629;
  assign n53659 = n53532 ^ n53531;
  assign n53660 = n53659 ^ n53657;
  assign n53661 = n53658 & n53660;
  assign n53662 = n53661 ^ n53629;
  assign n53626 = n53533 ^ n53526;
  assign n53663 = n53662 ^ n53626;
  assign n53664 = n51601 ^ n43991;
  assign n53665 = n53664 ^ n48135;
  assign n53666 = n53665 ^ n42513;
  assign n53667 = n53666 ^ n53626;
  assign n53668 = ~n53663 & n53667;
  assign n53669 = n53668 ^ n53666;
  assign n53670 = n53669 ^ n53624;
  assign n53671 = n53625 & ~n53670;
  assign n53672 = n53671 ^ n53621;
  assign n53673 = n53672 ^ n53619;
  assign n53674 = ~n53620 & ~n53673;
  assign n53675 = n53674 ^ n53616;
  assign n53676 = n53675 ^ n53614;
  assign n53677 = n53615 & n53676;
  assign n53678 = n53677 ^ n53613;
  assign n53679 = n53678 ^ n53609;
  assign n53680 = n53610 & ~n53679;
  assign n53681 = n53680 ^ n53608;
  assign n53682 = n53681 ^ n53604;
  assign n53683 = n53605 & ~n53682;
  assign n53684 = n53683 ^ n53601;
  assign n53685 = n53684 ^ n53599;
  assign n53686 = ~n53600 & n53685;
  assign n53687 = n53686 ^ n53598;
  assign n53595 = n53548 ^ n53547;
  assign n53688 = n53687 ^ n53595;
  assign n53689 = n51578 ^ n43973;
  assign n53690 = n53689 ^ n48100;
  assign n53691 = n53690 ^ n42490;
  assign n53692 = n53691 ^ n53595;
  assign n53693 = ~n53688 & n53692;
  assign n53694 = n53693 ^ n53691;
  assign n53695 = n53694 ^ n53593;
  assign n53696 = ~n53594 & n53695;
  assign n53697 = n53696 ^ n53592;
  assign n53551 = n53549 & ~n53550;
  assign n53495 = n53494 ^ n53428;
  assign n53496 = ~n53429 & ~n53495;
  assign n53497 = n53496 ^ n50921;
  assign n53378 = n52362 ^ n52319;
  assign n53379 = n53378 ^ n50941;
  assign n53374 = n53373 ^ n53213;
  assign n53375 = ~n53214 & n53374;
  assign n53376 = n53375 ^ n53212;
  assign n53210 = n53096 ^ n53031;
  assign n53377 = n53376 ^ n53210;
  assign n53426 = n53379 ^ n53377;
  assign n53427 = n53426 ^ n50950;
  assign n53524 = n53497 ^ n53427;
  assign n53589 = n53551 ^ n53524;
  assign n53698 = n53697 ^ n53589;
  assign n54128 = n53701 ^ n53698;
  assign n54120 = n53694 ^ n53592;
  assign n54121 = n54120 ^ n53593;
  assign n53821 = n52365 ^ n52340;
  assign n53408 = n53121 ^ n52998;
  assign n53409 = n53408 ^ n52999;
  assign n53822 = n53821 ^ n53409;
  assign n53820 = n53684 ^ n53600;
  assign n53823 = n53822 ^ n53820;
  assign n53826 = n53681 ^ n53605;
  assign n53189 = n53118 ^ n53003;
  assign n53190 = n53189 ^ n53004;
  assign n53824 = n53190 ^ n52428;
  assign n53825 = n53824 ^ n52345;
  assign n53827 = n53826 ^ n53825;
  assign n53830 = n53678 ^ n53610;
  assign n53828 = n52351 ^ n52319;
  assign n53194 = n53115 ^ n53112;
  assign n53829 = n53828 ^ n53194;
  assign n53831 = n53830 ^ n53829;
  assign n53383 = n53099 ^ n53025;
  assign n53384 = n53383 ^ n53022;
  assign n53837 = n53384 ^ n52707;
  assign n53838 = n53837 ^ n51755;
  assign n53836 = n53666 ^ n53663;
  assign n53839 = n53838 ^ n53836;
  assign n53841 = n53210 ^ n52371;
  assign n53842 = n53841 ^ n51757;
  assign n53840 = n53659 ^ n53658;
  assign n53843 = n53842 ^ n53840;
  assign n53846 = n53654 ^ n53632;
  assign n53847 = n53846 ^ n53652;
  assign n53844 = n52376 ^ n51763;
  assign n53845 = n53844 ^ n53213;
  assign n53848 = n53847 ^ n53845;
  assign n53851 = n53649 ^ n53635;
  assign n53852 = n53851 ^ n53647;
  assign n53849 = n52693 ^ n51765;
  assign n53850 = n53849 ^ n53217;
  assign n53853 = n53852 ^ n53850;
  assign n53856 = n53638 ^ n53527;
  assign n53857 = n53856 ^ n53643;
  assign n53854 = n53219 ^ n52380;
  assign n53855 = n53854 ^ n51771;
  assign n53858 = n53857 ^ n53855;
  assign n53861 = n53642 ^ n53641;
  assign n53859 = n52683 ^ n51773;
  assign n53860 = n53859 ^ n53223;
  assign n53862 = n53861 ^ n53860;
  assign n53865 = n51920 ^ n51220;
  assign n53866 = n53865 ^ n52634;
  assign n53802 = n53139 ^ n52970;
  assign n53867 = n53866 ^ n53802;
  assign n53868 = n53254 ^ n51228;
  assign n53869 = n53868 ^ n51929;
  assign n53808 = n53136 ^ n52973;
  assign n53809 = n53808 ^ n52974;
  assign n53870 = n53869 ^ n53809;
  assign n53742 = n52334 ^ n51822;
  assign n53743 = n53742 ^ n52747;
  assign n53741 = n53124 ^ n52995;
  assign n53744 = n53743 ^ n53741;
  assign n53406 = n52337 ^ n51807;
  assign n53407 = n53406 ^ n52329;
  assign n53410 = n53409 ^ n53407;
  assign n53187 = n52342 ^ n51811;
  assign n53188 = n53187 ^ n52331;
  assign n53191 = n53190 ^ n53188;
  assign n53192 = n52347 ^ n52332;
  assign n53193 = n53192 ^ n51729;
  assign n53195 = n53194 ^ n53193;
  assign n53197 = n52340 ^ n50931;
  assign n53198 = n53197 ^ n52354;
  assign n53196 = n53108 ^ n53011;
  assign n53199 = n53198 ^ n53196;
  assign n53202 = n53105 ^ n53015;
  assign n53203 = n53202 ^ n53012;
  assign n53200 = n52358 ^ n52345;
  assign n53201 = n53200 ^ n50935;
  assign n53204 = n53203 ^ n53201;
  assign n53207 = n52351 ^ n51335;
  assign n53208 = n53207 ^ n52365;
  assign n53205 = n53102 ^ n53019;
  assign n53206 = n53205 ^ n53020;
  assign n53209 = n53208 ^ n53206;
  assign n53380 = n53379 ^ n53210;
  assign n53381 = n53377 & n53380;
  assign n53382 = n53381 ^ n53379;
  assign n53385 = n53384 ^ n53382;
  assign n53386 = n52428 ^ n52356;
  assign n53387 = n53386 ^ n51328;
  assign n53388 = n53387 ^ n53384;
  assign n53389 = ~n53385 & ~n53388;
  assign n53390 = n53389 ^ n53387;
  assign n53391 = n53390 ^ n53206;
  assign n53392 = n53209 & ~n53391;
  assign n53393 = n53392 ^ n53208;
  assign n53394 = n53393 ^ n53203;
  assign n53395 = ~n53204 & n53394;
  assign n53396 = n53395 ^ n53201;
  assign n53397 = n53396 ^ n53196;
  assign n53398 = n53199 & n53397;
  assign n53399 = n53398 ^ n53198;
  assign n53400 = n53399 ^ n53194;
  assign n53401 = ~n53195 & n53400;
  assign n53402 = n53401 ^ n53193;
  assign n53403 = n53402 ^ n53190;
  assign n53404 = n53191 & n53403;
  assign n53405 = n53404 ^ n53188;
  assign n53738 = n53407 ^ n53405;
  assign n53739 = n53410 & ~n53738;
  assign n53740 = n53739 ^ n53409;
  assign n53766 = n53741 ^ n53740;
  assign n53767 = n53744 & ~n53766;
  assign n53768 = n53767 ^ n53743;
  assign n53763 = n52522 ^ n51831;
  assign n53764 = n53763 ^ n53169;
  assign n53872 = n53768 ^ n53764;
  assign n53762 = n53127 ^ n52990;
  assign n53873 = n53768 ^ n53762;
  assign n53874 = n53872 & n53873;
  assign n53875 = n53874 ^ n53764;
  assign n53871 = n53130 ^ n52985;
  assign n53876 = n53875 ^ n53871;
  assign n53877 = n51870 ^ n51739;
  assign n53878 = n53877 ^ n53260;
  assign n53879 = n53878 ^ n53871;
  assign n53880 = n53876 & n53879;
  assign n53881 = n53880 ^ n53878;
  assign n53814 = n53133 ^ n52978;
  assign n53815 = n53814 ^ n52979;
  assign n53882 = n53881 ^ n53815;
  assign n53883 = n53258 ^ n51221;
  assign n53884 = n53883 ^ n51922;
  assign n53885 = n53884 ^ n53815;
  assign n53886 = ~n53882 & ~n53885;
  assign n53887 = n53886 ^ n53884;
  assign n53888 = n53887 ^ n53809;
  assign n53889 = ~n53870 & n53888;
  assign n53890 = n53889 ^ n53869;
  assign n53922 = n53890 ^ n53866;
  assign n53923 = n53867 & ~n53922;
  assign n53924 = n53923 ^ n53802;
  assign n53797 = n53142 ^ n52965;
  assign n53925 = n53924 ^ n53797;
  assign n53926 = n51937 ^ n51218;
  assign n53927 = n53926 ^ n52639;
  assign n53938 = n53927 ^ n53797;
  assign n53939 = ~n53925 & n53938;
  assign n53940 = n53939 ^ n53927;
  assign n53935 = n52627 ^ n51913;
  assign n53936 = n53935 ^ n51215;
  assign n53791 = n53145 ^ n52960;
  assign n53937 = n53936 ^ n53791;
  assign n53941 = n53940 ^ n53937;
  assign n53942 = n53941 ^ n50512;
  assign n53891 = n53890 ^ n53867;
  assign n53892 = n53891 ^ n50517;
  assign n53893 = n53887 ^ n53869;
  assign n53894 = n53893 ^ n53809;
  assign n53895 = n53894 ^ n50518;
  assign n53765 = n53764 ^ n53762;
  assign n53769 = n53768 ^ n53765;
  assign n53898 = n53769 ^ n50352;
  assign n53745 = n53744 ^ n53740;
  assign n53746 = n53745 ^ n50933;
  assign n53412 = n53402 ^ n53191;
  assign n53413 = n53412 ^ n50985;
  assign n53414 = n53399 ^ n53195;
  assign n53415 = n53414 ^ n50938;
  assign n53416 = n53396 ^ n53198;
  assign n53417 = n53416 ^ n53196;
  assign n53418 = n53417 ^ n50986;
  assign n53419 = n53393 ^ n53204;
  assign n53420 = n53419 ^ n50990;
  assign n53421 = n53390 ^ n53208;
  assign n53422 = n53421 ^ n53206;
  assign n53423 = n53422 ^ n50994;
  assign n53424 = n53387 ^ n53385;
  assign n53425 = n53424 ^ n50944;
  assign n53498 = n53497 ^ n53426;
  assign n53499 = n53427 & ~n53498;
  assign n53500 = n53499 ^ n50950;
  assign n53501 = n53500 ^ n53424;
  assign n53502 = ~n53425 & ~n53501;
  assign n53503 = n53502 ^ n50944;
  assign n53504 = n53503 ^ n53422;
  assign n53505 = ~n53423 & n53504;
  assign n53506 = n53505 ^ n50994;
  assign n53507 = n53506 ^ n53419;
  assign n53508 = ~n53420 & ~n53507;
  assign n53509 = n53508 ^ n50990;
  assign n53510 = n53509 ^ n53417;
  assign n53511 = n53418 & ~n53510;
  assign n53512 = n53511 ^ n50986;
  assign n53513 = n53512 ^ n53414;
  assign n53514 = ~n53415 & ~n53513;
  assign n53515 = n53514 ^ n50938;
  assign n53516 = n53515 ^ n53412;
  assign n53517 = ~n53413 & ~n53516;
  assign n53518 = n53517 ^ n50985;
  assign n53519 = n53518 ^ n50984;
  assign n53411 = n53410 ^ n53405;
  assign n53735 = n53518 ^ n53411;
  assign n53736 = ~n53519 & ~n53735;
  assign n53737 = n53736 ^ n50984;
  assign n53758 = n53745 ^ n53737;
  assign n53759 = ~n53746 & n53758;
  assign n53760 = n53759 ^ n50933;
  assign n53899 = n53769 ^ n53760;
  assign n53900 = n53898 & ~n53899;
  assign n53901 = n53900 ^ n50352;
  assign n53897 = n53878 ^ n53876;
  assign n53902 = n53901 ^ n53897;
  assign n53903 = n53897 ^ n51119;
  assign n53904 = n53902 & n53903;
  assign n53905 = n53904 ^ n51119;
  assign n53896 = n53884 ^ n53882;
  assign n53906 = n53905 ^ n53896;
  assign n53907 = n53896 ^ n50522;
  assign n53908 = ~n53906 & n53907;
  assign n53909 = n53908 ^ n50522;
  assign n53910 = n53909 ^ n53894;
  assign n53911 = n53895 & n53910;
  assign n53912 = n53911 ^ n50518;
  assign n53929 = n53912 ^ n53891;
  assign n53930 = ~n53892 & n53929;
  assign n53931 = n53930 ^ n50517;
  assign n53928 = n53927 ^ n53925;
  assign n53932 = n53931 ^ n53928;
  assign n53943 = n53928 ^ n50513;
  assign n53944 = n53932 & ~n53943;
  assign n53945 = n53944 ^ n50513;
  assign n53956 = n53945 ^ n53941;
  assign n53957 = ~n53942 & ~n53956;
  assign n53958 = n53957 ^ n50512;
  assign n53951 = n53940 ^ n53791;
  assign n53952 = ~n53937 & n53951;
  assign n53953 = n53952 ^ n53936;
  assign n53948 = n52649 ^ n50978;
  assign n53949 = n53948 ^ n51799;
  assign n53786 = n53148 ^ n52953;
  assign n53787 = n53786 ^ n52954;
  assign n53950 = n53949 ^ n53787;
  assign n53954 = n53953 ^ n53950;
  assign n53955 = n53954 ^ n50377;
  assign n53959 = n53958 ^ n53955;
  assign n53913 = n53912 ^ n53892;
  assign n53747 = n53746 ^ n53737;
  assign n53520 = n53519 ^ n53411;
  assign n53521 = n53515 ^ n50985;
  assign n53522 = n53521 ^ n53412;
  assign n53523 = n53509 ^ n53418;
  assign n53552 = n53524 & ~n53551;
  assign n53553 = n53500 ^ n53425;
  assign n53554 = n53552 & ~n53553;
  assign n53555 = n53503 ^ n50994;
  assign n53556 = n53555 ^ n53422;
  assign n53557 = ~n53554 & ~n53556;
  assign n53558 = n53506 ^ n50990;
  assign n53559 = n53558 ^ n53419;
  assign n53560 = ~n53557 & n53559;
  assign n53561 = ~n53523 & ~n53560;
  assign n53562 = n53512 ^ n53415;
  assign n53563 = n53561 & n53562;
  assign n53564 = ~n53522 & n53563;
  assign n53748 = ~n53520 & ~n53564;
  assign n53757 = n53747 & n53748;
  assign n53761 = n53760 ^ n50352;
  assign n53770 = n53769 ^ n53761;
  assign n53914 = ~n53757 & n53770;
  assign n53915 = n53902 ^ n51119;
  assign n53916 = n53914 & n53915;
  assign n53917 = n53906 ^ n50522;
  assign n53918 = ~n53916 & n53917;
  assign n53919 = n53909 ^ n53895;
  assign n53920 = ~n53918 & ~n53919;
  assign n53921 = n53913 & ~n53920;
  assign n53933 = n53932 ^ n50513;
  assign n53934 = ~n53921 & ~n53933;
  assign n53946 = n53945 ^ n53942;
  assign n53947 = n53934 & ~n53946;
  assign n53981 = n53959 ^ n53947;
  assign n53978 = n51885 ^ n44258;
  assign n53979 = n53978 ^ n48428;
  assign n53980 = n53979 ^ n42868;
  assign n53982 = n53981 ^ n53980;
  assign n53984 = n51891 ^ n44263;
  assign n53985 = n53984 ^ n48392;
  assign n53986 = n53985 ^ n42874;
  assign n53983 = n53946 ^ n53934;
  assign n53987 = n53986 ^ n53983;
  assign n53991 = n53933 ^ n53921;
  assign n53988 = n51896 ^ n44269;
  assign n53989 = n53988 ^ n48398;
  assign n53990 = n53989 ^ n42962;
  assign n53992 = n53991 ^ n53990;
  assign n53996 = n53920 ^ n53913;
  assign n53993 = n51737 ^ n44273;
  assign n53994 = n53993 ^ n48403;
  assign n53995 = n53994 ^ n42880;
  assign n53997 = n53996 ^ n53995;
  assign n54001 = n53919 ^ n53918;
  assign n53998 = n51716 ^ n44289;
  assign n53999 = n53998 ^ n48407;
  assign n54000 = n53999 ^ n42885;
  assign n54002 = n54001 ^ n54000;
  assign n53771 = n53770 ^ n53757;
  assign n53753 = n51532 ^ n43490;
  assign n53754 = n53753 ^ n48053;
  assign n53755 = n53754 ^ n2681;
  assign n54005 = n53771 ^ n53755;
  assign n53569 = n53563 ^ n53522;
  assign n53566 = n51694 ^ n44080;
  assign n53567 = n53566 ^ n48067;
  assign n53568 = n53567 ^ n42904;
  assign n53570 = n53569 ^ n53568;
  assign n53574 = n53562 ^ n53561;
  assign n53571 = n51548 ^ n43944;
  assign n53572 = n53571 ^ n48211;
  assign n53573 = n53572 ^ n42908;
  assign n53575 = n53574 ^ n53573;
  assign n53577 = n51553 ^ n43949;
  assign n53578 = n53577 ^ n48073;
  assign n53579 = n53578 ^ n42913;
  assign n53576 = n53560 ^ n53523;
  assign n53580 = n53579 ^ n53576;
  assign n53581 = n53559 ^ n53557;
  assign n1326 = n1325 ^ n1265;
  assign n1363 = n1362 ^ n1326;
  assign n1373 = n1372 ^ n1363;
  assign n53582 = n53581 ^ n1373;
  assign n53585 = n51563 ^ n1158;
  assign n53586 = n53585 ^ n48085;
  assign n53587 = n53586 ^ n3350;
  assign n53584 = n53553 ^ n53552;
  assign n53588 = n53587 ^ n53584;
  assign n53702 = n53701 ^ n53589;
  assign n53703 = ~n53698 & n53702;
  assign n53704 = n53703 ^ n53701;
  assign n53705 = n53704 ^ n53587;
  assign n53706 = n53588 & ~n53705;
  assign n53707 = n53706 ^ n53584;
  assign n53583 = n53556 ^ n53554;
  assign n53708 = n53707 ^ n53583;
  assign n53709 = n51558 ^ n43955;
  assign n53710 = n53709 ^ n48080;
  assign n53711 = n53710 ^ n1354;
  assign n53712 = n53711 ^ n53583;
  assign n53713 = ~n53708 & n53712;
  assign n53714 = n53713 ^ n53711;
  assign n53715 = n53714 ^ n53581;
  assign n53716 = n53582 & ~n53715;
  assign n53717 = n53716 ^ n1373;
  assign n53718 = n53717 ^ n53576;
  assign n53719 = n53580 & ~n53718;
  assign n53720 = n53719 ^ n53579;
  assign n53721 = n53720 ^ n53574;
  assign n53722 = n53575 & ~n53721;
  assign n53723 = n53722 ^ n53573;
  assign n53724 = n53723 ^ n53569;
  assign n53725 = ~n53570 & n53724;
  assign n53726 = n53725 ^ n53568;
  assign n53565 = n53564 ^ n53520;
  assign n53727 = n53726 ^ n53565;
  assign n53728 = n51543 ^ n43937;
  assign n53729 = n53728 ^ n48063;
  assign n53730 = n53729 ^ n42899;
  assign n53731 = n53730 ^ n53565;
  assign n53732 = n53727 & ~n53731;
  assign n53733 = n53732 ^ n53730;
  assign n53184 = n51537 ^ n43932;
  assign n53185 = n53184 ^ n48058;
  assign n53186 = n53185 ^ n42894;
  assign n53734 = n53733 ^ n53186;
  assign n53749 = n53748 ^ n53747;
  assign n53750 = n53749 ^ n53733;
  assign n53751 = n53734 & n53750;
  assign n53752 = n53751 ^ n53186;
  assign n54006 = n53771 ^ n53752;
  assign n54007 = ~n54005 & n54006;
  assign n54008 = n54007 ^ n53755;
  assign n54004 = n53915 ^ n53914;
  assign n54009 = n54008 ^ n54004;
  assign n54010 = n51528 ^ n44095;
  assign n54011 = n54010 ^ n47602;
  assign n54012 = n54011 ^ n3107;
  assign n54013 = n54012 ^ n54004;
  assign n54014 = ~n54009 & n54013;
  assign n54015 = n54014 ^ n54012;
  assign n54003 = n53917 ^ n53916;
  assign n54016 = n54015 ^ n54003;
  assign n54017 = n51522 ^ n44278;
  assign n54018 = n54017 ^ n48232;
  assign n54019 = n54018 ^ n42949;
  assign n54020 = n54019 ^ n54003;
  assign n54021 = ~n54016 & n54020;
  assign n54022 = n54021 ^ n54019;
  assign n54023 = n54022 ^ n54001;
  assign n54024 = n54002 & ~n54023;
  assign n54025 = n54024 ^ n54000;
  assign n54026 = n54025 ^ n53996;
  assign n54027 = n53997 & ~n54026;
  assign n54028 = n54027 ^ n53995;
  assign n54029 = n54028 ^ n53991;
  assign n54030 = n53992 & ~n54029;
  assign n54031 = n54030 ^ n53990;
  assign n54032 = n54031 ^ n53986;
  assign n54033 = ~n53987 & ~n54032;
  assign n54034 = n54033 ^ n53983;
  assign n54035 = n54034 ^ n53981;
  assign n54036 = ~n53982 & ~n54035;
  assign n54037 = n54036 ^ n53980;
  assign n53972 = n53958 ^ n53954;
  assign n53973 = ~n53955 & ~n53972;
  assign n53974 = n53973 ^ n50377;
  assign n53966 = n53953 ^ n53787;
  assign n53967 = n53950 & ~n53966;
  assign n53968 = n53967 ^ n53949;
  assign n53778 = n53153 ^ n52950;
  assign n53779 = n53778 ^ n53151;
  assign n53969 = n53968 ^ n53779;
  assign n53964 = n51798 ^ n50974;
  assign n53965 = n53964 ^ n52625;
  assign n53970 = n53969 ^ n53965;
  assign n53971 = n53970 ^ n50373;
  assign n53975 = n53974 ^ n53971;
  assign n53961 = n51881 ^ n44310;
  assign n53962 = n53961 ^ n48387;
  assign n53963 = n53962 ^ n1868;
  assign n53976 = n53975 ^ n53963;
  assign n53960 = ~n53947 & ~n53959;
  assign n53977 = n53976 ^ n53960;
  assign n54038 = n54037 ^ n53977;
  assign n53863 = n53227 ^ n52385;
  assign n53864 = n53863 ^ n51779;
  assign n54039 = n54038 ^ n53864;
  assign n54042 = n54034 ^ n53982;
  assign n54040 = n53232 ^ n52389;
  assign n54041 = n54040 ^ n51783;
  assign n54043 = n54042 ^ n54041;
  assign n54048 = n54028 ^ n53992;
  assign n54046 = n53242 ^ n51791;
  assign n54047 = n54046 ^ n52397;
  assign n54049 = n54048 ^ n54047;
  assign n54050 = n53246 ^ n52398;
  assign n54051 = n54050 ^ n51795;
  assign n54052 = n54025 ^ n53995;
  assign n54053 = n54052 ^ n53996;
  assign n54054 = n54051 & n54053;
  assign n54055 = n54054 ^ n54048;
  assign n54056 = n54049 & n54055;
  assign n54057 = n54056 ^ n54054;
  assign n54044 = n53237 ^ n52394;
  assign n54045 = n54044 ^ n51787;
  assign n54058 = n54057 ^ n54045;
  assign n54059 = n54031 ^ n53987;
  assign n54060 = n54059 ^ n54057;
  assign n54061 = ~n54058 & n54060;
  assign n54062 = n54061 ^ n54045;
  assign n54063 = n54062 ^ n54042;
  assign n54064 = n54043 & n54063;
  assign n54065 = n54064 ^ n54041;
  assign n54066 = n54065 ^ n54038;
  assign n54067 = n54039 & n54066;
  assign n54068 = n54067 ^ n53864;
  assign n54069 = n54068 ^ n53861;
  assign n54070 = n53862 & n54069;
  assign n54071 = n54070 ^ n53860;
  assign n54072 = n54071 ^ n53857;
  assign n54073 = n53858 & ~n54072;
  assign n54074 = n54073 ^ n53855;
  assign n54075 = n54074 ^ n53852;
  assign n54076 = n53853 & ~n54075;
  assign n54077 = n54076 ^ n53850;
  assign n54078 = n54077 ^ n53847;
  assign n54079 = n53848 & ~n54078;
  assign n54080 = n54079 ^ n53845;
  assign n54081 = n54080 ^ n53840;
  assign n54082 = n53843 & n54081;
  assign n54083 = n54082 ^ n53842;
  assign n54084 = n54083 ^ n53836;
  assign n54085 = ~n53839 & n54084;
  assign n54086 = n54085 ^ n53838;
  assign n53835 = n53669 ^ n53625;
  assign n54087 = n54086 ^ n53835;
  assign n54088 = n53206 ^ n52367;
  assign n54089 = n54088 ^ n51749;
  assign n54090 = n54089 ^ n53835;
  assign n54091 = n54087 & ~n54090;
  assign n54092 = n54091 ^ n54089;
  assign n53834 = n53672 ^ n53620;
  assign n54093 = n54092 ^ n53834;
  assign n54094 = n52362 ^ n51745;
  assign n54095 = n54094 ^ n53203;
  assign n54096 = n54095 ^ n53834;
  assign n54097 = ~n54093 & ~n54096;
  assign n54098 = n54097 ^ n54095;
  assign n53832 = n53675 ^ n53613;
  assign n53833 = n53832 ^ n53614;
  assign n54099 = n54098 ^ n53833;
  assign n54100 = n52356 ^ n51744;
  assign n54101 = n54100 ^ n53196;
  assign n54102 = n54101 ^ n53833;
  assign n54103 = n54099 & ~n54102;
  assign n54104 = n54103 ^ n54101;
  assign n54105 = n54104 ^ n53830;
  assign n54106 = ~n53831 & ~n54105;
  assign n54107 = n54106 ^ n53829;
  assign n54108 = n54107 ^ n53826;
  assign n54109 = n53827 & n54108;
  assign n54110 = n54109 ^ n53825;
  assign n54111 = n54110 ^ n53820;
  assign n54112 = ~n53823 & n54111;
  assign n54113 = n54112 ^ n53822;
  assign n53819 = n53691 ^ n53688;
  assign n54114 = n54113 ^ n53819;
  assign n54115 = n53741 ^ n52358;
  assign n54116 = n54115 ^ n52332;
  assign n54117 = n54116 ^ n53819;
  assign n54118 = ~n54114 & ~n54117;
  assign n54119 = n54118 ^ n54116;
  assign n54122 = n54121 ^ n54119;
  assign n54123 = n52354 ^ n52331;
  assign n54124 = n54123 ^ n53762;
  assign n54125 = n54124 ^ n54121;
  assign n54126 = ~n54122 & n54125;
  assign n54127 = n54126 ^ n54124;
  assign n54129 = n54128 ^ n54127;
  assign n54130 = n53871 ^ n52329;
  assign n54131 = n54130 ^ n52347;
  assign n54132 = n54131 ^ n54128;
  assign n54133 = n54129 & n54132;
  assign n54134 = n54133 ^ n54131;
  assign n53816 = n53815 ^ n52342;
  assign n53817 = n53816 ^ n52747;
  assign n54166 = n54134 ^ n53817;
  assign n53813 = n53704 ^ n53588;
  assign n54167 = n54166 ^ n53813;
  assign n54168 = n54167 ^ n51811;
  assign n54169 = n54131 ^ n54129;
  assign n54170 = n54169 ^ n51729;
  assign n54171 = n54124 ^ n54122;
  assign n54172 = n54171 ^ n50931;
  assign n54173 = n54116 ^ n54114;
  assign n54174 = n54173 ^ n50935;
  assign n54175 = n54110 ^ n53823;
  assign n54176 = n54175 ^ n51335;
  assign n54177 = n54107 ^ n53825;
  assign n54178 = n54177 ^ n53826;
  assign n54179 = n54178 ^ n51328;
  assign n54180 = n54104 ^ n53831;
  assign n54181 = n54180 ^ n50941;
  assign n54182 = n54101 ^ n54099;
  assign n54183 = n54182 ^ n51318;
  assign n54184 = n54095 ^ n54093;
  assign n54185 = n54184 ^ n51311;
  assign n54186 = n54089 ^ n54087;
  assign n54187 = n54186 ^ n51304;
  assign n54189 = n54080 ^ n53842;
  assign n54190 = n54189 ^ n53840;
  assign n54191 = n54190 ^ n50952;
  assign n54194 = n54074 ^ n53853;
  assign n54195 = n54194 ^ n50956;
  assign n54196 = n54071 ^ n53858;
  assign n54197 = n54196 ^ n51281;
  assign n54198 = n54068 ^ n53862;
  assign n54199 = n54198 ^ n50960;
  assign n54202 = n54062 ^ n54043;
  assign n54203 = n54202 ^ n50965;
  assign n54206 = n54053 ^ n54051;
  assign n54207 = n50972 & n54206;
  assign n54208 = n54207 ^ n50969;
  assign n54209 = n54054 ^ n54047;
  assign n54210 = n54209 ^ n54048;
  assign n54211 = n54210 ^ n54207;
  assign n54212 = n54208 & n54211;
  assign n54213 = n54212 ^ n50969;
  assign n54204 = n54059 ^ n54045;
  assign n54205 = n54204 ^ n54057;
  assign n54214 = n54213 ^ n54205;
  assign n54215 = n54205 ^ n51262;
  assign n54216 = ~n54214 & n54215;
  assign n54217 = n54216 ^ n51262;
  assign n54218 = n54217 ^ n54202;
  assign n54219 = n54203 & n54218;
  assign n54220 = n54219 ^ n50965;
  assign n54200 = n54065 ^ n53864;
  assign n54201 = n54200 ^ n54038;
  assign n54221 = n54220 ^ n54201;
  assign n54222 = n54201 ^ n50962;
  assign n54223 = n54221 & n54222;
  assign n54224 = n54223 ^ n50962;
  assign n54225 = n54224 ^ n54198;
  assign n54226 = n54199 & n54225;
  assign n54227 = n54226 ^ n50960;
  assign n54228 = n54227 ^ n54196;
  assign n54229 = n54197 & n54228;
  assign n54230 = n54229 ^ n51281;
  assign n54231 = n54230 ^ n54194;
  assign n54232 = n54195 & ~n54231;
  assign n54233 = n54232 ^ n50956;
  assign n54192 = n54077 ^ n53845;
  assign n54193 = n54192 ^ n53847;
  assign n54234 = n54233 ^ n54193;
  assign n54235 = n54193 ^ n51291;
  assign n54236 = ~n54234 & ~n54235;
  assign n54237 = n54236 ^ n51291;
  assign n54238 = n54237 ^ n54190;
  assign n54239 = n54191 & n54238;
  assign n54240 = n54239 ^ n50952;
  assign n54188 = n54083 ^ n53839;
  assign n54241 = n54240 ^ n54188;
  assign n54242 = n54240 ^ n50946;
  assign n54243 = ~n54241 & ~n54242;
  assign n54244 = n54243 ^ n50946;
  assign n54245 = n54244 ^ n54186;
  assign n54246 = ~n54187 & n54245;
  assign n54247 = n54246 ^ n51304;
  assign n54248 = n54247 ^ n54184;
  assign n54249 = n54185 & n54248;
  assign n54250 = n54249 ^ n51311;
  assign n54251 = n54250 ^ n54182;
  assign n54252 = ~n54183 & n54251;
  assign n54253 = n54252 ^ n51318;
  assign n54254 = n54253 ^ n54180;
  assign n54255 = n54181 & n54254;
  assign n54256 = n54255 ^ n50941;
  assign n54257 = n54256 ^ n54178;
  assign n54258 = ~n54179 & ~n54257;
  assign n54259 = n54258 ^ n51328;
  assign n54260 = n54259 ^ n54175;
  assign n54261 = n54176 & n54260;
  assign n54262 = n54261 ^ n51335;
  assign n54263 = n54262 ^ n54173;
  assign n54264 = n54174 & ~n54263;
  assign n54265 = n54264 ^ n50935;
  assign n54266 = n54265 ^ n54171;
  assign n54267 = n54172 & ~n54266;
  assign n54268 = n54267 ^ n50931;
  assign n54269 = n54268 ^ n54169;
  assign n54270 = n54170 & ~n54269;
  assign n54271 = n54270 ^ n51729;
  assign n54272 = n54271 ^ n54167;
  assign n54273 = n54168 & n54272;
  assign n54274 = n54273 ^ n51811;
  assign n53818 = n53817 ^ n53813;
  assign n54135 = n54134 ^ n53813;
  assign n54136 = n53818 & ~n54135;
  assign n54137 = n54136 ^ n53817;
  assign n53810 = n53809 ^ n53169;
  assign n53811 = n53810 ^ n52337;
  assign n53807 = n53711 ^ n53708;
  assign n53812 = n53811 ^ n53807;
  assign n54165 = n54137 ^ n53812;
  assign n54275 = n54274 ^ n54165;
  assign n54276 = n54165 ^ n51807;
  assign n54277 = n54275 & n54276;
  assign n54278 = n54277 ^ n51807;
  assign n54279 = n54278 ^ n51822;
  assign n54138 = n54137 ^ n53811;
  assign n54139 = ~n53812 & n54138;
  assign n54140 = n54139 ^ n53807;
  assign n53805 = n53714 ^ n53582;
  assign n53803 = n53802 ^ n53260;
  assign n53804 = n53803 ^ n52334;
  assign n53806 = n53805 ^ n53804;
  assign n54280 = n54140 ^ n53806;
  assign n54281 = n54280 ^ n54278;
  assign n54282 = ~n54279 & n54281;
  assign n54283 = n54282 ^ n51822;
  assign n54141 = n54140 ^ n53805;
  assign n54142 = n53806 & ~n54141;
  assign n54143 = n54142 ^ n53804;
  assign n53799 = n53717 ^ n53579;
  assign n53800 = n53799 ^ n53576;
  assign n53796 = n53258 ^ n52522;
  assign n53798 = n53797 ^ n53796;
  assign n53801 = n53800 ^ n53798;
  assign n54164 = n54143 ^ n53801;
  assign n54284 = n54283 ^ n54164;
  assign n54306 = n54284 ^ n51831;
  assign n54307 = n54275 ^ n51807;
  assign n54308 = n54265 ^ n50931;
  assign n54309 = n54308 ^ n54171;
  assign n54310 = n54262 ^ n50935;
  assign n54311 = n54310 ^ n54173;
  assign n54312 = n54230 ^ n54195;
  assign n54313 = n54214 ^ n51262;
  assign n54314 = n54210 ^ n54208;
  assign n54315 = ~n54313 & n54314;
  assign n54316 = n54217 ^ n54203;
  assign n54317 = ~n54315 & n54316;
  assign n54318 = n54221 ^ n50962;
  assign n54319 = ~n54317 & n54318;
  assign n54320 = n54224 ^ n54199;
  assign n54321 = ~n54319 & n54320;
  assign n54322 = n54227 ^ n54197;
  assign n54323 = ~n54321 & n54322;
  assign n54324 = ~n54312 & n54323;
  assign n54325 = n54234 ^ n51291;
  assign n54326 = n54324 & n54325;
  assign n54327 = n54237 ^ n54191;
  assign n54328 = ~n54326 & ~n54327;
  assign n54329 = n54241 ^ n50946;
  assign n54330 = n54328 & ~n54329;
  assign n54331 = n54244 ^ n51304;
  assign n54332 = n54331 ^ n54186;
  assign n54333 = n54330 & n54332;
  assign n54334 = n54247 ^ n51311;
  assign n54335 = n54334 ^ n54184;
  assign n54336 = n54333 & ~n54335;
  assign n54337 = n54250 ^ n51318;
  assign n54338 = n54337 ^ n54182;
  assign n54339 = n54336 & ~n54338;
  assign n54340 = n54253 ^ n50941;
  assign n54341 = n54340 ^ n54180;
  assign n54342 = ~n54339 & ~n54341;
  assign n54343 = n54256 ^ n51328;
  assign n54344 = n54343 ^ n54178;
  assign n54345 = n54342 & ~n54344;
  assign n54346 = n54259 ^ n54176;
  assign n54347 = ~n54345 & n54346;
  assign n54348 = n54311 & ~n54347;
  assign n54349 = ~n54309 & ~n54348;
  assign n54350 = n54268 ^ n51729;
  assign n54351 = n54350 ^ n54169;
  assign n54352 = n54349 & ~n54351;
  assign n54353 = n54271 ^ n54168;
  assign n54354 = n54352 & ~n54353;
  assign n54355 = ~n54307 & ~n54354;
  assign n54356 = n54280 ^ n51822;
  assign n54357 = n54356 ^ n54278;
  assign n54358 = n54355 & n54357;
  assign n54359 = n54306 & ~n54358;
  assign n54285 = n54164 ^ n51831;
  assign n54286 = n54284 & n54285;
  assign n54287 = n54286 ^ n51831;
  assign n54360 = n54287 ^ n51870;
  assign n54144 = n54143 ^ n53800;
  assign n54145 = ~n53801 & ~n54144;
  assign n54146 = n54145 ^ n53798;
  assign n53794 = n53720 ^ n53575;
  assign n53792 = n53791 ^ n53254;
  assign n53793 = n53792 ^ n51739;
  assign n53795 = n53794 ^ n53793;
  assign n54162 = n54146 ^ n53795;
  assign n54361 = n54360 ^ n54162;
  assign n54362 = n54359 & ~n54361;
  assign n54147 = n54146 ^ n53794;
  assign n54148 = ~n53795 & n54147;
  assign n54149 = n54148 ^ n53793;
  assign n53788 = n53787 ^ n51922;
  assign n53789 = n53788 ^ n52634;
  assign n53784 = n53723 ^ n53568;
  assign n53785 = n53784 ^ n53569;
  assign n53790 = n53789 ^ n53785;
  assign n54292 = n54149 ^ n53790;
  assign n54163 = n54162 ^ n51870;
  assign n54288 = n54287 ^ n54162;
  assign n54289 = n54163 & n54288;
  assign n54290 = n54289 ^ n51870;
  assign n54291 = n54290 ^ n51221;
  assign n54363 = n54292 ^ n54291;
  assign n54364 = ~n54362 & ~n54363;
  assign n54293 = n54292 ^ n54290;
  assign n54294 = n54291 & ~n54293;
  assign n54295 = n54294 ^ n51221;
  assign n54150 = n54149 ^ n53789;
  assign n54151 = ~n53790 & n54150;
  assign n54152 = n54151 ^ n53785;
  assign n53782 = n53730 ^ n53727;
  assign n53780 = n53779 ^ n51929;
  assign n53781 = n53780 ^ n52639;
  assign n53783 = n53782 ^ n53781;
  assign n54161 = n54152 ^ n53783;
  assign n54296 = n54295 ^ n54161;
  assign n54365 = n54296 ^ n51228;
  assign n54366 = ~n54364 & ~n54365;
  assign n54153 = n54152 ^ n53782;
  assign n54154 = ~n53783 & ~n54153;
  assign n54155 = n54154 ^ n53781;
  assign n53776 = n53749 ^ n53734;
  assign n53774 = n52627 ^ n51920;
  assign n53775 = n53774 ^ n53328;
  assign n53777 = n53776 ^ n53775;
  assign n54301 = n54155 ^ n53777;
  assign n54367 = n54301 ^ n51220;
  assign n54297 = n54161 ^ n51228;
  assign n54298 = ~n54296 & ~n54297;
  assign n54299 = n54298 ^ n51228;
  assign n54368 = n54367 ^ n54299;
  assign n54369 = ~n54366 & n54368;
  assign n54300 = n54299 ^ n51220;
  assign n54302 = n54301 ^ n54299;
  assign n54303 = n54300 & ~n54302;
  assign n54304 = n54303 ^ n51220;
  assign n54156 = n54155 ^ n53776;
  assign n54157 = ~n53777 & n54156;
  assign n54158 = n54157 ^ n53775;
  assign n53756 = n53755 ^ n53752;
  assign n53772 = n53771 ^ n53756;
  assign n53182 = n53181 ^ n51937;
  assign n53183 = n53182 ^ n52649;
  assign n53773 = n53772 ^ n53183;
  assign n54159 = n54158 ^ n53773;
  assign n54160 = n54159 ^ n51218;
  assign n54305 = n54304 ^ n54160;
  assign n54388 = n54369 ^ n54305;
  assign n54385 = n52568 ^ n44999;
  assign n54386 = n54385 ^ n49092;
  assign n54387 = n54386 ^ n43651;
  assign n54389 = n54388 ^ n54387;
  assign n54393 = n54368 ^ n54366;
  assign n54390 = n52572 ^ n44938;
  assign n54391 = n54390 ^ n49096;
  assign n54392 = n54391 ^ n2966;
  assign n54394 = n54393 ^ n54392;
  assign n54396 = n52575 ^ n44943;
  assign n54397 = n54396 ^ n2870;
  assign n54398 = n54397 ^ n43483;
  assign n54395 = n54365 ^ n54364;
  assign n54399 = n54398 ^ n54395;
  assign n54403 = n54363 ^ n54362;
  assign n54400 = n52580 ^ n3119;
  assign n54401 = n54400 ^ n49103;
  assign n54402 = n54401 ^ n2862;
  assign n54404 = n54403 ^ n54402;
  assign n54407 = n52586 ^ n44979;
  assign n54408 = n54407 ^ n49113;
  assign n54409 = n54408 ^ n43456;
  assign n54406 = n54358 ^ n54306;
  assign n54410 = n54409 ^ n54406;
  assign n54415 = n54354 ^ n54307;
  assign n54412 = n52305 ^ n44956;
  assign n54413 = n54412 ^ n49124;
  assign n54414 = n54413 ^ n43297;
  assign n54416 = n54415 ^ n54414;
  assign n54421 = n54351 ^ n54349;
  assign n54418 = n52153 ^ n44117;
  assign n54419 = n54418 ^ n48254;
  assign n54420 = n54419 ^ n43307;
  assign n54422 = n54421 ^ n54420;
  assign n54424 = n52158 ^ n1486;
  assign n54425 = n54424 ^ n48671;
  assign n54426 = n54425 ^ n43437;
  assign n54423 = n54348 ^ n54309;
  assign n54427 = n54426 ^ n54423;
  assign n54429 = n52163 ^ n1468;
  assign n54430 = n54429 ^ n48676;
  assign n54431 = n54430 ^ n43430;
  assign n54428 = n54347 ^ n54311;
  assign n54432 = n54431 ^ n54428;
  assign n54436 = n54346 ^ n54345;
  assign n54433 = n52168 ^ n44552;
  assign n54434 = n54433 ^ n48681;
  assign n54435 = n54434 ^ n43314;
  assign n54437 = n54436 ^ n54435;
  assign n54441 = n54344 ^ n54342;
  assign n54438 = n52173 ^ n44557;
  assign n54439 = n54438 ^ n48686;
  assign n54440 = n54439 ^ n43319;
  assign n54442 = n54441 ^ n54440;
  assign n54446 = n54341 ^ n54339;
  assign n54443 = n52178 ^ n44562;
  assign n54444 = n54443 ^ n48691;
  assign n54445 = n54444 ^ n43324;
  assign n54447 = n54446 ^ n54445;
  assign n54451 = n54338 ^ n54336;
  assign n54448 = n52183 ^ n44567;
  assign n54449 = n54448 ^ n48696;
  assign n54450 = n54449 ^ n914;
  assign n54452 = n54451 ^ n54450;
  assign n54460 = n54329 ^ n54328;
  assign n54457 = n52196 ^ n44652;
  assign n54458 = n54457 ^ n48774;
  assign n54459 = n54458 ^ n43401;
  assign n54461 = n54460 ^ n54459;
  assign n54467 = n54323 ^ n54312;
  assign n54464 = n52211 ^ n44590;
  assign n54465 = n54464 ^ n48718;
  assign n54466 = n54465 ^ n43344;
  assign n54468 = n54467 ^ n54466;
  assign n54470 = n52254 ^ n44632;
  assign n54471 = n54470 ^ n48724;
  assign n54472 = n54471 ^ n43381;
  assign n54469 = n54322 ^ n54321;
  assign n54473 = n54472 ^ n54469;
  assign n54479 = n54316 ^ n54315;
  assign n54476 = n52227 ^ n44606;
  assign n54477 = n54476 ^ n48734;
  assign n54478 = n54477 ^ n2255;
  assign n54480 = n54479 ^ n54478;
  assign n54487 = n52535 ^ n1940;
  assign n54488 = n54487 ^ n49061;
  assign n54489 = n54488 ^ n43622;
  assign n54490 = n54206 ^ n50972;
  assign n54491 = n54489 & n54490;
  assign n54484 = n52231 ^ n44613;
  assign n54485 = n54484 ^ n48738;
  assign n54486 = n54485 ^ n2100;
  assign n54492 = n54491 ^ n54486;
  assign n54493 = n54491 ^ n54314;
  assign n54494 = n54492 & ~n54493;
  assign n54495 = n54494 ^ n54486;
  assign n54481 = n52235 ^ n44610;
  assign n54482 = n54481 ^ n2111;
  assign n54483 = n54482 ^ n43362;
  assign n54496 = n54495 ^ n54483;
  assign n54497 = n54314 ^ n54313;
  assign n54498 = n54497 ^ n54495;
  assign n54499 = n54496 & ~n54498;
  assign n54500 = n54499 ^ n54483;
  assign n54501 = n54500 ^ n54479;
  assign n54502 = ~n54480 & n54501;
  assign n54503 = n54502 ^ n54478;
  assign n54475 = n54318 ^ n54317;
  assign n54504 = n54503 ^ n54475;
  assign n54505 = n52222 ^ n44600;
  assign n54506 = n54505 ^ n48752;
  assign n54507 = n54506 ^ n43356;
  assign n54508 = n54507 ^ n54475;
  assign n54509 = ~n54504 & n54508;
  assign n54510 = n54509 ^ n54507;
  assign n54474 = n54320 ^ n54319;
  assign n54511 = n54510 ^ n54474;
  assign n54512 = n52217 ^ n44595;
  assign n54513 = n54512 ^ n48729;
  assign n54514 = n54513 ^ n43351;
  assign n54515 = n54514 ^ n54474;
  assign n54516 = n54511 & ~n54515;
  assign n54517 = n54516 ^ n54514;
  assign n54518 = n54517 ^ n54472;
  assign n54519 = n54473 & ~n54518;
  assign n54520 = n54519 ^ n54469;
  assign n54521 = n54520 ^ n54467;
  assign n54522 = n54468 & ~n54521;
  assign n54523 = n54522 ^ n54466;
  assign n54463 = n54325 ^ n54324;
  assign n54524 = n54523 ^ n54463;
  assign n54525 = n52206 ^ n44642;
  assign n54526 = n54525 ^ n48714;
  assign n54527 = n54526 ^ n43391;
  assign n54528 = n54527 ^ n54463;
  assign n54529 = n54524 & ~n54528;
  assign n54530 = n54529 ^ n54527;
  assign n54462 = n54327 ^ n54326;
  assign n54531 = n54530 ^ n54462;
  assign n54532 = n52201 ^ n44584;
  assign n54533 = n54532 ^ n48709;
  assign n54534 = n54533 ^ n43339;
  assign n54535 = n54534 ^ n54530;
  assign n54536 = ~n54531 & n54535;
  assign n54537 = n54536 ^ n54534;
  assign n54538 = n54537 ^ n54460;
  assign n54539 = ~n54461 & n54538;
  assign n54540 = n54539 ^ n54459;
  assign n54454 = n52192 ^ n44577;
  assign n54455 = n54454 ^ n48781;
  assign n54456 = n54455 ^ n43408;
  assign n54541 = n54540 ^ n54456;
  assign n54542 = n54332 ^ n54330;
  assign n54543 = n54542 ^ n54456;
  assign n54544 = ~n54541 & n54543;
  assign n54545 = n54544 ^ n54542;
  assign n54453 = n54335 ^ n54333;
  assign n54546 = n54545 ^ n54453;
  assign n54547 = n52186 ^ n44572;
  assign n54548 = n54547 ^ n48702;
  assign n54549 = n54548 ^ n43332;
  assign n54550 = n54549 ^ n54453;
  assign n54551 = n54546 & ~n54550;
  assign n54552 = n54551 ^ n54549;
  assign n54553 = n54552 ^ n54451;
  assign n54554 = ~n54452 & n54553;
  assign n54555 = n54554 ^ n54450;
  assign n54556 = n54555 ^ n54446;
  assign n54557 = ~n54447 & n54556;
  assign n54558 = n54557 ^ n54445;
  assign n54559 = n54558 ^ n54441;
  assign n54560 = n54442 & ~n54559;
  assign n54561 = n54560 ^ n54440;
  assign n54562 = n54561 ^ n54436;
  assign n54563 = ~n54437 & n54562;
  assign n54564 = n54563 ^ n54435;
  assign n54565 = n54564 ^ n54428;
  assign n54566 = n54432 & ~n54565;
  assign n54567 = n54566 ^ n54431;
  assign n54568 = n54567 ^ n54426;
  assign n54569 = n54427 & ~n54568;
  assign n54570 = n54569 ^ n54423;
  assign n54571 = n54570 ^ n54421;
  assign n54572 = ~n54422 & n54571;
  assign n54573 = n54572 ^ n54420;
  assign n54417 = n54353 ^ n54352;
  assign n54574 = n54573 ^ n54417;
  assign n54575 = n52148 ^ n44966;
  assign n54576 = n54575 ^ n48811;
  assign n54577 = n54576 ^ n43303;
  assign n54578 = n54577 ^ n54417;
  assign n54579 = n54574 & ~n54578;
  assign n54580 = n54579 ^ n54577;
  assign n54581 = n54580 ^ n54415;
  assign n54582 = ~n54416 & n54581;
  assign n54583 = n54582 ^ n54414;
  assign n54411 = n54357 ^ n54355;
  assign n54584 = n54583 ^ n54411;
  assign n54585 = n52311 ^ n44951;
  assign n54586 = n54585 ^ n49118;
  assign n54587 = n54586 ^ n43292;
  assign n54588 = n54587 ^ n54411;
  assign n54589 = n54584 & ~n54588;
  assign n54590 = n54589 ^ n54587;
  assign n54591 = n54590 ^ n54409;
  assign n54592 = ~n54410 & ~n54591;
  assign n54593 = n54592 ^ n54406;
  assign n54405 = n54361 ^ n54359;
  assign n54594 = n54593 ^ n54405;
  assign n54595 = n52598 ^ n2738;
  assign n54596 = n54595 ^ n49108;
  assign n54597 = n54596 ^ n3227;
  assign n54598 = n54597 ^ n54405;
  assign n54599 = ~n54594 & ~n54598;
  assign n54600 = n54599 ^ n54597;
  assign n54601 = n54600 ^ n54403;
  assign n54602 = ~n54404 & n54601;
  assign n54603 = n54602 ^ n54402;
  assign n54604 = n54603 ^ n54398;
  assign n54605 = n54399 & ~n54604;
  assign n54606 = n54605 ^ n54395;
  assign n54607 = n54606 ^ n54393;
  assign n54608 = n54394 & ~n54607;
  assign n54609 = n54608 ^ n54392;
  assign n54610 = n54609 ^ n54388;
  assign n54611 = ~n54389 & n54610;
  assign n54612 = n54611 ^ n54387;
  assign n54379 = n54304 ^ n54159;
  assign n54380 = ~n54160 & n54379;
  assign n54381 = n54380 ^ n51218;
  assign n54382 = n54381 ^ n51215;
  assign n54375 = n54158 ^ n53772;
  assign n54376 = n53773 & n54375;
  assign n54377 = n54376 ^ n53183;
  assign n54372 = n52625 ^ n51913;
  assign n54373 = n54372 ^ n53326;
  assign n54371 = n54012 ^ n54009;
  assign n54374 = n54373 ^ n54371;
  assign n54378 = n54377 ^ n54374;
  assign n54383 = n54382 ^ n54378;
  assign n54370 = n54305 & ~n54369;
  assign n54384 = n54383 ^ n54370;
  assign n54613 = n54612 ^ n54384;
  assign n54656 = n54616 ^ n54613;
  assign n56060 = n54656 ^ n54038;
  assign n56061 = n56060 ^ n53316;
  assign n55181 = n52968 ^ n45469;
  assign n55182 = n55181 ^ n49515;
  assign n55183 = n55182 ^ n43490;
  assign n54822 = n54549 ^ n54546;
  assign n54820 = n53871 ^ n52332;
  assign n54821 = n54820 ^ n53805;
  assign n54823 = n54822 ^ n54821;
  assign n54826 = n54542 ^ n54541;
  assign n54824 = n53762 ^ n52340;
  assign n54825 = n54824 ^ n53807;
  assign n54827 = n54826 ^ n54825;
  assign n54828 = n53813 ^ n52345;
  assign n54829 = n54828 ^ n53741;
  assign n54773 = n54537 ^ n54459;
  assign n54774 = n54773 ^ n54460;
  assign n54830 = n54829 ^ n54774;
  assign n54831 = n54128 ^ n53409;
  assign n54832 = n54831 ^ n52351;
  assign n54777 = n54534 ^ n54531;
  assign n54833 = n54832 ^ n54777;
  assign n54836 = n54527 ^ n54524;
  assign n54834 = n53190 ^ n52356;
  assign n54835 = n54834 ^ n54121;
  assign n54837 = n54836 ^ n54835;
  assign n54840 = n53819 ^ n53194;
  assign n54841 = n54840 ^ n52362;
  assign n54838 = n54520 ^ n54466;
  assign n54839 = n54838 ^ n54467;
  assign n54842 = n54841 ^ n54839;
  assign n54845 = n54517 ^ n54473;
  assign n54843 = n53820 ^ n52367;
  assign n54844 = n54843 ^ n53196;
  assign n54846 = n54845 ^ n54844;
  assign n54849 = n54514 ^ n54511;
  assign n54847 = n53203 ^ n52707;
  assign n54848 = n54847 ^ n53826;
  assign n54850 = n54849 ^ n54848;
  assign n54853 = n54507 ^ n54504;
  assign n54851 = n53830 ^ n52371;
  assign n54852 = n54851 ^ n53206;
  assign n54854 = n54853 ^ n54852;
  assign n54857 = n54500 ^ n54478;
  assign n54858 = n54857 ^ n54479;
  assign n54855 = n53833 ^ n53384;
  assign n54856 = n54855 ^ n52376;
  assign n54859 = n54858 ^ n54856;
  assign n54862 = n54497 ^ n54483;
  assign n54863 = n54862 ^ n54495;
  assign n54860 = n53210 ^ n52693;
  assign n54861 = n54860 ^ n53834;
  assign n54864 = n54863 ^ n54861;
  assign n54867 = n54486 ^ n54314;
  assign n54868 = n54867 ^ n54491;
  assign n54865 = n53835 ^ n52380;
  assign n54866 = n54865 ^ n53213;
  assign n54869 = n54868 ^ n54866;
  assign n54761 = n54490 ^ n54489;
  assign n54759 = n53836 ^ n53217;
  assign n54760 = n54759 ^ n52683;
  assign n54762 = n54761 ^ n54760;
  assign n54637 = n54370 & n54383;
  assign n54631 = n54378 ^ n51215;
  assign n54632 = n54381 ^ n54378;
  assign n54633 = ~n54631 & n54632;
  assign n54634 = n54633 ^ n51215;
  assign n54626 = n54377 ^ n54373;
  assign n54627 = ~n54374 & ~n54626;
  assign n54628 = n54627 ^ n54371;
  assign n54624 = n52409 ^ n51799;
  assign n54625 = n54624 ^ n53319;
  assign n54629 = n54628 ^ n54625;
  assign n54623 = n54019 ^ n54016;
  assign n54630 = n54629 ^ n54623;
  assign n54635 = n54634 ^ n54630;
  assign n54636 = n54635 ^ n50978;
  assign n54638 = n54637 ^ n54636;
  assign n54620 = n52558 ^ n44927;
  assign n54621 = n54620 ^ n49086;
  assign n54622 = n54621 ^ n43632;
  assign n54639 = n54638 ^ n54622;
  assign n54617 = n54616 ^ n54384;
  assign n54618 = ~n54613 & n54617;
  assign n54619 = n54618 ^ n54616;
  assign n54706 = n54638 ^ n54619;
  assign n54707 = ~n54639 & n54706;
  assign n54708 = n54707 ^ n54622;
  assign n54701 = n54630 ^ n50978;
  assign n54702 = n54635 & ~n54701;
  assign n54703 = n54702 ^ n50978;
  assign n54696 = n54625 ^ n54623;
  assign n54697 = n54628 ^ n54623;
  assign n54698 = n54696 & ~n54697;
  assign n54699 = n54698 ^ n54625;
  assign n54690 = ~n54636 & ~n54637;
  assign n54691 = n54690 ^ n43627;
  assign n54692 = n54691 ^ n52552;
  assign n54687 = n54022 ^ n54002;
  assign n54688 = n54687 ^ n52403;
  assign n54689 = n54688 ^ n45012;
  assign n54693 = n54692 ^ n54689;
  assign n54694 = n54693 ^ n49080;
  assign n54695 = n54694 ^ n53964;
  assign n54700 = n54699 ^ n54695;
  assign n54704 = n54703 ^ n54700;
  assign n54705 = n54704 ^ n53316;
  assign n54709 = n54708 ^ n54705;
  assign n54684 = n53840 ^ n52385;
  assign n54685 = n54684 ^ n53219;
  assign n54755 = n54709 ^ n54685;
  assign n54649 = n53232 ^ n52397;
  assign n54650 = n54649 ^ n53857;
  assign n54644 = n54606 ^ n54392;
  assign n54645 = n54644 ^ n54393;
  assign n54646 = n53861 ^ n52398;
  assign n54647 = n54646 ^ n53237;
  assign n54648 = n54645 & n54647;
  assign n54651 = n54650 ^ n54648;
  assign n54652 = n54609 ^ n54389;
  assign n54653 = n54652 ^ n54650;
  assign n54654 = ~n54651 & ~n54653;
  assign n54655 = n54654 ^ n54648;
  assign n54657 = n54656 ^ n54655;
  assign n54658 = n53852 ^ n52394;
  assign n54659 = n54658 ^ n53227;
  assign n54660 = n54659 ^ n54656;
  assign n54661 = ~n54657 & n54660;
  assign n54662 = n54661 ^ n54659;
  assign n54641 = n53223 ^ n52389;
  assign n54642 = n54641 ^ n53847;
  assign n54680 = n54662 ^ n54642;
  assign n54640 = n54639 ^ n54619;
  assign n54681 = n54662 ^ n54640;
  assign n54682 = n54680 & n54681;
  assign n54683 = n54682 ^ n54642;
  assign n54756 = n54709 ^ n54683;
  assign n54757 = ~n54755 & ~n54756;
  assign n54758 = n54757 ^ n54685;
  assign n54870 = n54761 ^ n54758;
  assign n54871 = ~n54762 & n54870;
  assign n54872 = n54871 ^ n54760;
  assign n54873 = n54872 ^ n54868;
  assign n54874 = n54869 & n54873;
  assign n54875 = n54874 ^ n54866;
  assign n54876 = n54875 ^ n54863;
  assign n54877 = n54864 & ~n54876;
  assign n54878 = n54877 ^ n54861;
  assign n54879 = n54878 ^ n54858;
  assign n54880 = n54859 & n54879;
  assign n54881 = n54880 ^ n54856;
  assign n54882 = n54881 ^ n54853;
  assign n54883 = n54854 & n54882;
  assign n54884 = n54883 ^ n54852;
  assign n54885 = n54884 ^ n54849;
  assign n54886 = ~n54850 & n54885;
  assign n54887 = n54886 ^ n54848;
  assign n54888 = n54887 ^ n54845;
  assign n54889 = n54846 & ~n54888;
  assign n54890 = n54889 ^ n54844;
  assign n54891 = n54890 ^ n54841;
  assign n54892 = n54842 & ~n54891;
  assign n54893 = n54892 ^ n54839;
  assign n54894 = n54893 ^ n54836;
  assign n54895 = ~n54837 & n54894;
  assign n54896 = n54895 ^ n54835;
  assign n54897 = n54896 ^ n54777;
  assign n54898 = ~n54833 & ~n54897;
  assign n54899 = n54898 ^ n54832;
  assign n54900 = n54899 ^ n54829;
  assign n54901 = n54830 & ~n54900;
  assign n54902 = n54901 ^ n54774;
  assign n54903 = n54902 ^ n54826;
  assign n54904 = ~n54827 & n54903;
  assign n54905 = n54904 ^ n54825;
  assign n54906 = n54905 ^ n54822;
  assign n54907 = ~n54823 & ~n54906;
  assign n54908 = n54907 ^ n54821;
  assign n54819 = n54552 ^ n54452;
  assign n54909 = n54908 ^ n54819;
  assign n54910 = n53800 ^ n52331;
  assign n54911 = n54910 ^ n53815;
  assign n54912 = n54911 ^ n54819;
  assign n54913 = n54909 & n54912;
  assign n54914 = n54913 ^ n54911;
  assign n54816 = n53809 ^ n53794;
  assign n54817 = n54816 ^ n52329;
  assign n54815 = n54555 ^ n54447;
  assign n54818 = n54817 ^ n54815;
  assign n54971 = n54914 ^ n54818;
  assign n54972 = n54971 ^ n52347;
  assign n54973 = n54911 ^ n54909;
  assign n54974 = n54973 ^ n52354;
  assign n54975 = n54905 ^ n54821;
  assign n54976 = n54975 ^ n54822;
  assign n54977 = n54976 ^ n52358;
  assign n54978 = n54902 ^ n54827;
  assign n54979 = n54978 ^ n52365;
  assign n54980 = n54899 ^ n54830;
  assign n54981 = n54980 ^ n52428;
  assign n54982 = n54896 ^ n54833;
  assign n54983 = n54982 ^ n52319;
  assign n54984 = n54893 ^ n54837;
  assign n54985 = n54984 ^ n51744;
  assign n54986 = n54887 ^ n54846;
  assign n54987 = n54986 ^ n51749;
  assign n54989 = n54881 ^ n54852;
  assign n54990 = n54989 ^ n54853;
  assign n54991 = n54990 ^ n51757;
  assign n54992 = n54878 ^ n54859;
  assign n54993 = n54992 ^ n51763;
  assign n54996 = n54872 ^ n54866;
  assign n54997 = n54996 ^ n54868;
  assign n54998 = n54997 ^ n51771;
  assign n54686 = n54685 ^ n54683;
  assign n54710 = n54709 ^ n54686;
  assign n54711 = n54710 ^ n51779;
  assign n54643 = n54642 ^ n54640;
  assign n54663 = n54662 ^ n54643;
  assign n54664 = n54663 ^ n51783;
  assign n54665 = n54659 ^ n54657;
  assign n54666 = n54665 ^ n51787;
  assign n54667 = n54647 ^ n54645;
  assign n54668 = n51795 & n54667;
  assign n54669 = n54668 ^ n51791;
  assign n54670 = n54652 ^ n54651;
  assign n54671 = n54670 ^ n54668;
  assign n54672 = n54669 & ~n54671;
  assign n54673 = n54672 ^ n51791;
  assign n54674 = n54673 ^ n54665;
  assign n54675 = ~n54666 & ~n54674;
  assign n54676 = n54675 ^ n51787;
  assign n54677 = n54676 ^ n54663;
  assign n54678 = ~n54664 & ~n54677;
  assign n54679 = n54678 ^ n51783;
  assign n54764 = n54710 ^ n54679;
  assign n54765 = n54711 & n54764;
  assign n54766 = n54765 ^ n51779;
  assign n54763 = n54762 ^ n54758;
  assign n54767 = n54766 ^ n54763;
  assign n54999 = n54763 ^ n51773;
  assign n55000 = n54767 & ~n54999;
  assign n55001 = n55000 ^ n51773;
  assign n55002 = n55001 ^ n54997;
  assign n55003 = n54998 & ~n55002;
  assign n55004 = n55003 ^ n51771;
  assign n54994 = n54875 ^ n54861;
  assign n54995 = n54994 ^ n54863;
  assign n55005 = n55004 ^ n54995;
  assign n55006 = n54995 ^ n51765;
  assign n55007 = n55005 & ~n55006;
  assign n55008 = n55007 ^ n51765;
  assign n55009 = n55008 ^ n54992;
  assign n55010 = n54993 & n55009;
  assign n55011 = n55010 ^ n51763;
  assign n55012 = n55011 ^ n54990;
  assign n55013 = ~n54991 & n55012;
  assign n55014 = n55013 ^ n51757;
  assign n54988 = n54884 ^ n54850;
  assign n55015 = n55014 ^ n54988;
  assign n55016 = n54988 ^ n51755;
  assign n55017 = n55015 & n55016;
  assign n55018 = n55017 ^ n51755;
  assign n55019 = n55018 ^ n54986;
  assign n55020 = ~n54987 & n55019;
  assign n55021 = n55020 ^ n51749;
  assign n55022 = n55021 ^ n51745;
  assign n55023 = n54890 ^ n54842;
  assign n55024 = n55023 ^ n55021;
  assign n55025 = n55022 & n55024;
  assign n55026 = n55025 ^ n51745;
  assign n55027 = n55026 ^ n54984;
  assign n55028 = ~n54985 & ~n55027;
  assign n55029 = n55028 ^ n51744;
  assign n55030 = n55029 ^ n54982;
  assign n55031 = ~n54983 & n55030;
  assign n55032 = n55031 ^ n52319;
  assign n55033 = n55032 ^ n54980;
  assign n55034 = n54981 & n55033;
  assign n55035 = n55034 ^ n52428;
  assign n55036 = n55035 ^ n54978;
  assign n55037 = n54979 & n55036;
  assign n55038 = n55037 ^ n52365;
  assign n55039 = n55038 ^ n54976;
  assign n55040 = n54977 & ~n55039;
  assign n55041 = n55040 ^ n52358;
  assign n55042 = n55041 ^ n54973;
  assign n55043 = n54974 & ~n55042;
  assign n55044 = n55043 ^ n52354;
  assign n55045 = n55044 ^ n54971;
  assign n55046 = n54972 & n55045;
  assign n55047 = n55046 ^ n52347;
  assign n55077 = n55047 ^ n52342;
  assign n54919 = n53785 ^ n52747;
  assign n54920 = n54919 ^ n53802;
  assign n54915 = n54914 ^ n54815;
  assign n54916 = n54818 & ~n54915;
  assign n54917 = n54916 ^ n54817;
  assign n54814 = n54558 ^ n54442;
  assign n54918 = n54917 ^ n54814;
  assign n54969 = n54920 ^ n54918;
  assign n55078 = n55077 ^ n54969;
  assign n55079 = n55032 ^ n54981;
  assign n55080 = n55026 ^ n54985;
  assign n55081 = n55023 ^ n51745;
  assign n55082 = n55081 ^ n55021;
  assign n55083 = n55015 ^ n51755;
  assign n54712 = n54711 ^ n54679;
  assign n54713 = n54670 ^ n54669;
  assign n54714 = n54673 ^ n54666;
  assign n54715 = ~n54713 & n54714;
  assign n54716 = n54676 ^ n54664;
  assign n54717 = ~n54715 & n54716;
  assign n54754 = ~n54712 & ~n54717;
  assign n54768 = n54767 ^ n51773;
  assign n55084 = ~n54754 & n54768;
  assign n55085 = n55001 ^ n54998;
  assign n55086 = ~n55084 & n55085;
  assign n55087 = n55005 ^ n51765;
  assign n55088 = n55086 & ~n55087;
  assign n55089 = n55008 ^ n54993;
  assign n55090 = n55088 & n55089;
  assign n55091 = n55011 ^ n54991;
  assign n55092 = ~n55090 & ~n55091;
  assign n55093 = n55083 & n55092;
  assign n55094 = n55018 ^ n54987;
  assign n55095 = n55093 & n55094;
  assign n55096 = n55082 & n55095;
  assign n55097 = n55080 & n55096;
  assign n55098 = n55029 ^ n54983;
  assign n55099 = ~n55097 & n55098;
  assign n55100 = ~n55079 & n55099;
  assign n55101 = n55035 ^ n54979;
  assign n55102 = ~n55100 & ~n55101;
  assign n55103 = n55038 ^ n54977;
  assign n55104 = ~n55102 & ~n55103;
  assign n55105 = n55041 ^ n54974;
  assign n55106 = ~n55104 & n55105;
  assign n55107 = n55044 ^ n54972;
  assign n55108 = n55106 & n55107;
  assign n55109 = n55078 & n55108;
  assign n54970 = n54969 ^ n52342;
  assign n55048 = n55047 ^ n54969;
  assign n55049 = ~n54970 & ~n55048;
  assign n55050 = n55049 ^ n52342;
  assign n54921 = n54920 ^ n54814;
  assign n54922 = n54918 & n54921;
  assign n54923 = n54922 ^ n54920;
  assign n54811 = n53782 ^ n53169;
  assign n54812 = n54811 ^ n53797;
  assign n54967 = n54923 ^ n54812;
  assign n54810 = n54561 ^ n54437;
  assign n54968 = n54967 ^ n54810;
  assign n55051 = n55050 ^ n54968;
  assign n55110 = n55051 ^ n52337;
  assign n55111 = ~n55109 & ~n55110;
  assign n55052 = n54968 ^ n52337;
  assign n55053 = n55051 & n55052;
  assign n55054 = n55053 ^ n52337;
  assign n54813 = n54812 ^ n54810;
  assign n54924 = n54923 ^ n54810;
  assign n54925 = ~n54813 & n54924;
  assign n54926 = n54925 ^ n54812;
  assign n54808 = n54564 ^ n54432;
  assign n54806 = n53791 ^ n53260;
  assign n54807 = n54806 ^ n53776;
  assign n54809 = n54808 ^ n54807;
  assign n54965 = n54926 ^ n54809;
  assign n54966 = n54965 ^ n52334;
  assign n55112 = n55054 ^ n54966;
  assign n55113 = n55111 & n55112;
  assign n55055 = n55054 ^ n54965;
  assign n55056 = n54966 & ~n55055;
  assign n55057 = n55056 ^ n52334;
  assign n54931 = n53787 ^ n53258;
  assign n54932 = n54931 ^ n53772;
  assign n54927 = n54926 ^ n54808;
  assign n54928 = ~n54809 & ~n54927;
  assign n54929 = n54928 ^ n54807;
  assign n54805 = n54567 ^ n54427;
  assign n54930 = n54929 ^ n54805;
  assign n54964 = n54932 ^ n54930;
  assign n55058 = n55057 ^ n54964;
  assign n55076 = n55058 ^ n52522;
  assign n55180 = n55113 ^ n55076;
  assign n55184 = n55183 ^ n55180;
  assign n55188 = n55112 ^ n55111;
  assign n55185 = n52973 ^ n45305;
  assign n55186 = n55185 ^ n49520;
  assign n55187 = n55186 ^ n43932;
  assign n55189 = n55188 ^ n55187;
  assign n55193 = n55110 ^ n55109;
  assign n55190 = n52978 ^ n45459;
  assign n55191 = n55190 ^ n49525;
  assign n55192 = n55191 ^ n43937;
  assign n55194 = n55193 ^ n55192;
  assign n55198 = n55108 ^ n55078;
  assign n55195 = n52984 ^ n45311;
  assign n55196 = n55195 ^ n49531;
  assign n55197 = n55196 ^ n44080;
  assign n55199 = n55198 ^ n55197;
  assign n55203 = n55107 ^ n55106;
  assign n55200 = n52988 ^ n45316;
  assign n55201 = n55200 ^ n49535;
  assign n55202 = n55201 ^ n43944;
  assign n55204 = n55203 ^ n55202;
  assign n55208 = n55105 ^ n55104;
  assign n55205 = n52993 ^ n45322;
  assign n55206 = n55205 ^ n49540;
  assign n55207 = n55206 ^ n43949;
  assign n55209 = n55208 ^ n55207;
  assign n55213 = n55103 ^ n55102;
  assign n55210 = n52998 ^ n45326;
  assign n55211 = n55210 ^ n49545;
  assign n55212 = n55211 ^ n1325;
  assign n55214 = n55213 ^ n55212;
  assign n55218 = n55101 ^ n55100;
  assign n55215 = n53003 ^ n45331;
  assign n55216 = n55215 ^ n1169;
  assign n55217 = n55216 ^ n43955;
  assign n55219 = n55218 ^ n55217;
  assign n55223 = n55099 ^ n55079;
  assign n55220 = n53115 ^ n45334;
  assign n55221 = n55220 ^ n49659;
  assign n55222 = n55221 ^ n1158;
  assign n55224 = n55223 ^ n55222;
  assign n55228 = n55098 ^ n55097;
  assign n55225 = n53009 ^ n995;
  assign n55226 = n55225 ^ n49553;
  assign n55227 = n55226 ^ n43963;
  assign n55229 = n55228 ^ n55227;
  assign n55233 = n55096 ^ n55080;
  assign n55230 = n53015 ^ n45339;
  assign n55231 = n55230 ^ n49559;
  assign n55232 = n55231 ^ n43967;
  assign n55234 = n55233 ^ n55232;
  assign n55238 = n55095 ^ n55082;
  assign n55235 = n53019 ^ n49563;
  assign n55236 = n55235 ^ n45345;
  assign n55237 = n55236 ^ n43973;
  assign n55239 = n55238 ^ n55237;
  assign n55241 = n53025 ^ n45421;
  assign n55242 = n55241 ^ n49568;
  assign n55243 = n55242 ^ n43977;
  assign n55240 = n55094 ^ n55093;
  assign n55244 = n55243 ^ n55240;
  assign n55248 = n55092 ^ n55083;
  assign n55245 = n53029 ^ n45351;
  assign n55246 = n55245 ^ n49571;
  assign n55247 = n55246 ^ n44046;
  assign n55249 = n55248 ^ n55247;
  assign n55253 = n55091 ^ n55090;
  assign n55250 = n53034 ^ n45355;
  assign n55251 = n55250 ^ n49576;
  assign n55252 = n55251 ^ n44039;
  assign n55254 = n55253 ^ n55252;
  assign n55256 = n53039 ^ n45360;
  assign n55257 = n55256 ^ n49581;
  assign n55258 = n55257 ^ n44032;
  assign n55255 = n55089 ^ n55088;
  assign n55259 = n55258 ^ n55255;
  assign n55264 = n55085 ^ n55084;
  assign n55261 = n53049 ^ n45402;
  assign n55262 = n55261 ^ n49626;
  assign n55263 = n55262 ^ n44022;
  assign n55265 = n55264 ^ n55263;
  assign n54769 = n54768 ^ n54754;
  assign n54751 = n53053 ^ n45372;
  assign n54752 = n54751 ^ n49592;
  assign n54753 = n54752 ^ n43991;
  assign n54770 = n54769 ^ n54753;
  assign n54718 = n54717 ^ n54712;
  assign n2364 = n2363 ^ n2300;
  assign n2398 = n2397 ^ n2364;
  assign n2408 = n2407 ^ n2398;
  assign n54719 = n54718 ^ n2408;
  assign n54727 = n53252 ^ n45639;
  assign n54728 = n54727 ^ n49794;
  assign n54729 = n54728 ^ n44243;
  assign n54730 = n54667 ^ n51795;
  assign n54731 = n54729 & n54730;
  assign n54724 = n53067 ^ n45381;
  assign n54725 = n54724 ^ n49600;
  assign n54726 = n54725 ^ n44003;
  assign n54732 = n54731 ^ n54726;
  assign n54733 = n54731 ^ n54713;
  assign n54734 = n54732 & n54733;
  assign n54735 = n54734 ^ n54726;
  assign n54723 = n54714 ^ n54713;
  assign n54736 = n54735 ^ n54723;
  assign n54737 = n53064 ^ n2193;
  assign n54738 = n54737 ^ n49604;
  assign n54739 = n54738 ^ n44000;
  assign n54740 = n54739 ^ n54735;
  assign n54741 = ~n54736 & n54740;
  assign n54742 = n54741 ^ n54739;
  assign n54720 = n53059 ^ n45378;
  assign n54721 = n54720 ^ n49612;
  assign n54722 = n54721 ^ n2389;
  assign n54743 = n54742 ^ n54722;
  assign n54744 = n54716 ^ n54715;
  assign n54745 = n54744 ^ n54742;
  assign n54746 = n54743 & n54745;
  assign n54747 = n54746 ^ n54722;
  assign n54748 = n54747 ^ n54718;
  assign n54749 = ~n54719 & n54748;
  assign n54750 = n54749 ^ n2408;
  assign n55266 = n54769 ^ n54750;
  assign n55267 = ~n54770 & n55266;
  assign n55268 = n55267 ^ n54753;
  assign n55269 = n55268 ^ n55264;
  assign n55270 = n55265 & ~n55269;
  assign n55271 = n55270 ^ n55263;
  assign n55260 = n55087 ^ n55086;
  assign n55272 = n55271 ^ n55260;
  assign n55273 = n53045 ^ n45365;
  assign n55274 = n55273 ^ n49586;
  assign n55275 = n55274 ^ n43986;
  assign n55276 = n55275 ^ n55260;
  assign n55277 = ~n55272 & n55276;
  assign n55278 = n55277 ^ n55275;
  assign n55279 = n55278 ^ n55258;
  assign n55280 = ~n55259 & ~n55279;
  assign n55281 = n55280 ^ n55255;
  assign n55282 = n55281 ^ n55253;
  assign n55283 = n55254 & n55282;
  assign n55284 = n55283 ^ n55252;
  assign n55285 = n55284 ^ n55248;
  assign n55286 = n55249 & ~n55285;
  assign n55287 = n55286 ^ n55247;
  assign n55288 = n55287 ^ n55243;
  assign n55289 = n55244 & ~n55288;
  assign n55290 = n55289 ^ n55240;
  assign n55291 = n55290 ^ n55238;
  assign n55292 = n55239 & ~n55291;
  assign n55293 = n55292 ^ n55237;
  assign n55294 = n55293 ^ n55233;
  assign n55295 = n55234 & ~n55294;
  assign n55296 = n55295 ^ n55232;
  assign n55297 = n55296 ^ n55228;
  assign n55298 = n55229 & ~n55297;
  assign n55299 = n55298 ^ n55227;
  assign n55300 = n55299 ^ n55223;
  assign n55301 = n55224 & ~n55300;
  assign n55302 = n55301 ^ n55222;
  assign n55303 = n55302 ^ n55218;
  assign n55304 = n55219 & ~n55303;
  assign n55305 = n55304 ^ n55217;
  assign n55306 = n55305 ^ n55213;
  assign n55307 = ~n55214 & n55306;
  assign n55308 = n55307 ^ n55212;
  assign n55309 = n55308 ^ n55208;
  assign n55310 = ~n55209 & n55309;
  assign n55311 = n55310 ^ n55207;
  assign n55312 = n55311 ^ n55203;
  assign n55313 = n55204 & ~n55312;
  assign n55314 = n55313 ^ n55202;
  assign n55315 = n55314 ^ n55198;
  assign n55316 = n55199 & ~n55315;
  assign n55317 = n55316 ^ n55197;
  assign n55318 = n55317 ^ n55193;
  assign n55319 = ~n55194 & n55318;
  assign n55320 = n55319 ^ n55192;
  assign n55321 = n55320 ^ n55188;
  assign n55322 = ~n55189 & n55321;
  assign n55323 = n55322 ^ n55187;
  assign n55324 = n55323 ^ n55183;
  assign n55325 = ~n55184 & ~n55324;
  assign n55326 = n55325 ^ n55180;
  assign n55059 = n54964 ^ n52522;
  assign n55060 = ~n55058 & ~n55059;
  assign n55061 = n55060 ^ n52522;
  assign n54933 = n54932 ^ n54805;
  assign n54934 = n54930 & n54933;
  assign n54935 = n54934 ^ n54932;
  assign n54802 = n54570 ^ n54420;
  assign n54803 = n54802 ^ n54421;
  assign n54800 = n54371 ^ n53779;
  assign n54801 = n54800 ^ n53254;
  assign n54804 = n54803 ^ n54801;
  assign n54962 = n54935 ^ n54804;
  assign n54963 = n54962 ^ n51739;
  assign n55115 = n55061 ^ n54963;
  assign n55114 = n55076 & ~n55113;
  assign n55178 = n55115 ^ n55114;
  assign n55175 = n52963 ^ n45300;
  assign n55176 = n55175 ^ n49510;
  assign n55177 = n55176 ^ n44095;
  assign n55179 = n55178 ^ n55177;
  assign n56059 = n55326 ^ n55179;
  assign n56062 = n56061 ^ n56059;
  assign n56041 = n55323 ^ n55184;
  assign n56039 = n54042 ^ n53319;
  assign n56040 = n56039 ^ n54652;
  assign n56042 = n56041 ^ n56040;
  assign n56014 = n55320 ^ n55189;
  assign n56012 = n54059 ^ n53326;
  assign n56013 = n56012 ^ n54645;
  assign n56015 = n56014 ^ n56013;
  assign n55963 = n54053 ^ n53328;
  assign n55143 = n54600 ^ n54404;
  assign n55964 = n55963 ^ n55143;
  assign n55961 = n55314 ^ n55197;
  assign n55962 = n55961 ^ n55198;
  assign n55965 = n55964 ^ n55962;
  assign n55909 = n55308 ^ n55207;
  assign n55910 = n55909 ^ n55208;
  assign n54792 = n54590 ^ n54410;
  assign n55907 = n54792 ^ n53787;
  assign n55908 = n55907 ^ n54623;
  assign n55911 = n55910 ^ n55908;
  assign n55887 = n55305 ^ n55212;
  assign n55888 = n55887 ^ n55213;
  assign n54796 = n54587 ^ n54584;
  assign n55885 = n54796 ^ n53791;
  assign n55886 = n55885 ^ n54371;
  assign n55889 = n55888 ^ n55886;
  assign n54945 = n54580 ^ n54416;
  assign n55865 = n54945 ^ n53797;
  assign n55866 = n55865 ^ n53772;
  assign n55864 = n55302 ^ n55219;
  assign n55867 = n55866 ^ n55864;
  assign n55814 = n55296 ^ n55227;
  assign n55815 = n55814 ^ n55228;
  assign n55812 = n54803 ^ n53782;
  assign n55813 = n55812 ^ n53809;
  assign n55816 = n55815 ^ n55813;
  assign n55614 = n55293 ^ n55234;
  assign n55612 = n53815 ^ n53785;
  assign n55613 = n55612 ^ n54805;
  assign n55615 = n55614 ^ n55613;
  assign n55595 = n54808 ^ n53871;
  assign n55596 = n55595 ^ n53794;
  assign n55594 = n55290 ^ n55239;
  assign n55597 = n55596 ^ n55594;
  assign n55585 = n55287 ^ n55244;
  assign n55583 = n54810 ^ n53800;
  assign n55584 = n55583 ^ n53762;
  assign n55586 = n55585 ^ n55584;
  assign n55556 = n55281 ^ n55252;
  assign n55557 = n55556 ^ n55253;
  assign n55554 = n54815 ^ n53807;
  assign n55555 = n55554 ^ n53409;
  assign n55558 = n55557 ^ n55555;
  assign n55542 = n55278 ^ n55259;
  assign n55539 = n54819 ^ n53190;
  assign n55540 = n55539 ^ n53813;
  assign n55550 = n55542 ^ n55540;
  assign n54780 = n54747 ^ n54719;
  assign n54778 = n54777 ^ n53820;
  assign n54779 = n54778 ^ n53206;
  assign n54781 = n54780 ^ n54779;
  assign n55371 = n54853 ^ n53835;
  assign n55372 = n55371 ^ n53219;
  assign n55327 = n55326 ^ n55178;
  assign n55328 = n55179 & n55327;
  assign n55329 = n55328 ^ n55177;
  assign n55062 = n55061 ^ n54962;
  assign n55063 = n54963 & ~n55062;
  assign n55064 = n55063 ^ n51739;
  assign n54940 = n54577 ^ n54573;
  assign n54941 = n54940 ^ n54417;
  assign n54936 = n54935 ^ n54803;
  assign n54937 = n54804 & n54936;
  assign n54938 = n54937 ^ n54801;
  assign n54798 = n54623 ^ n52634;
  assign n54799 = n54798 ^ n53328;
  assign n54939 = n54938 ^ n54799;
  assign n54960 = n54941 ^ n54939;
  assign n54961 = n54960 ^ n51922;
  assign n55117 = n55064 ^ n54961;
  assign n55116 = n55114 & n55115;
  assign n55174 = n55117 ^ n55116;
  assign n55330 = n55329 ^ n55174;
  assign n55331 = n52959 ^ n3239;
  assign n55332 = n55331 ^ n49506;
  assign n55333 = n55332 ^ n44278;
  assign n55334 = n55333 ^ n55174;
  assign n55335 = n55330 & ~n55334;
  assign n55336 = n55335 ^ n55333;
  assign n55065 = n55064 ^ n54960;
  assign n55066 = n54961 & n55065;
  assign n55067 = n55066 ^ n51922;
  assign n54947 = n54687 ^ n52639;
  assign n54948 = n54947 ^ n53181;
  assign n54942 = n54941 ^ n54799;
  assign n54943 = n54939 & ~n54942;
  assign n54944 = n54943 ^ n54938;
  assign n54946 = n54945 ^ n54944;
  assign n54958 = n54948 ^ n54946;
  assign n54959 = n54958 ^ n51929;
  assign n55119 = n55067 ^ n54959;
  assign n55118 = ~n55116 & ~n55117;
  assign n55173 = n55119 ^ n55118;
  assign n55337 = n55336 ^ n55173;
  assign n55338 = n52953 ^ n2931;
  assign n55339 = n55338 ^ n49501;
  assign n55340 = n55339 ^ n44289;
  assign n55341 = n55340 ^ n55173;
  assign n55342 = ~n55337 & n55341;
  assign n55343 = n55342 ^ n55340;
  assign n55170 = n52950 ^ n45665;
  assign n55171 = n55170 ^ n49495;
  assign n55172 = n55171 ^ n44273;
  assign n55344 = n55343 ^ n55172;
  assign n55068 = n55067 ^ n54958;
  assign n55069 = n54959 & ~n55068;
  assign n55070 = n55069 ^ n51929;
  assign n54949 = n54948 ^ n54945;
  assign n54950 = ~n54946 & n54949;
  assign n54951 = n54950 ^ n54948;
  assign n54794 = n53326 ^ n52627;
  assign n54795 = n54794 ^ n54053;
  assign n54797 = n54796 ^ n54795;
  assign n54956 = n54951 ^ n54797;
  assign n54957 = n54956 ^ n51920;
  assign n55121 = n55070 ^ n54957;
  assign n55120 = ~n55118 & ~n55119;
  assign n55345 = n55121 ^ n55120;
  assign n55346 = n55345 ^ n55343;
  assign n55347 = n55344 & ~n55346;
  assign n55348 = n55347 ^ n55172;
  assign n55122 = ~n55120 & n55121;
  assign n55071 = n55070 ^ n54956;
  assign n55072 = n54957 & n55071;
  assign n55073 = n55072 ^ n51920;
  assign n54952 = n54951 ^ n54796;
  assign n54953 = ~n54797 & ~n54952;
  assign n54954 = n54953 ^ n54795;
  assign n54790 = n54048 ^ n53319;
  assign n54791 = n54790 ^ n52649;
  assign n54793 = n54792 ^ n54791;
  assign n54955 = n54954 ^ n54793;
  assign n55074 = n55073 ^ n54955;
  assign n55075 = n55074 ^ n51937;
  assign n55169 = n55122 ^ n55075;
  assign n55349 = n55348 ^ n55169;
  assign n55350 = n45660 ^ n3011;
  assign n55351 = n55350 ^ n49702;
  assign n55352 = n55351 ^ n44269;
  assign n55353 = n55352 ^ n55169;
  assign n55354 = n55349 & ~n55353;
  assign n55355 = n55354 ^ n55352;
  assign n55132 = n54955 ^ n51937;
  assign n55133 = n55074 & n55132;
  assign n55134 = n55133 ^ n51937;
  assign n55128 = n54954 ^ n54792;
  assign n55129 = ~n54793 & n55128;
  assign n55130 = n55129 ^ n54791;
  assign n55126 = n54597 ^ n54594;
  assign n55124 = n54059 ^ n53316;
  assign n55125 = n55124 ^ n52625;
  assign n55127 = n55126 ^ n55125;
  assign n55131 = n55130 ^ n55127;
  assign n55135 = n55134 ^ n55131;
  assign n55136 = n55135 ^ n51913;
  assign n55123 = n55075 & ~n55122;
  assign n55168 = n55136 ^ n55123;
  assign n55356 = n55355 ^ n55168;
  assign n55357 = n53162 ^ n45655;
  assign n55358 = n55357 ^ n49826;
  assign n55359 = n55358 ^ n44263;
  assign n55360 = n55359 ^ n55168;
  assign n55361 = n55356 & ~n55360;
  assign n55362 = n55361 ^ n55359;
  assign n55147 = n55131 ^ n51913;
  assign n55148 = ~n55135 & n55147;
  assign n55149 = n55148 ^ n51913;
  assign n55140 = n55130 ^ n55126;
  assign n55141 = ~n55127 & ~n55140;
  assign n55142 = n55141 ^ n55125;
  assign n55144 = n55143 ^ n55142;
  assign n55138 = n53246 ^ n52409;
  assign n55139 = n55138 ^ n54042;
  assign n55145 = n55144 ^ n55139;
  assign n55146 = n55145 ^ n51799;
  assign n55150 = n55149 ^ n55146;
  assign n55137 = n55123 & ~n55136;
  assign n55167 = n55150 ^ n55137;
  assign n55363 = n55362 ^ n55167;
  assign n55364 = n53304 ^ n45650;
  assign n55365 = n55364 ^ n49817;
  assign n55366 = n55365 ^ n44258;
  assign n55367 = n55366 ^ n55167;
  assign n55368 = n55363 & ~n55367;
  assign n55369 = n55368 ^ n55366;
  assign n55162 = n55149 ^ n55145;
  assign n55163 = ~n55146 & ~n55162;
  assign n55164 = n55163 ^ n51799;
  assign n55157 = n55143 ^ n55139;
  assign n55158 = ~n55144 & n55157;
  assign n55159 = n55158 ^ n55139;
  assign n55155 = n54603 ^ n54399;
  assign n55153 = n54038 ^ n53242;
  assign n55154 = n55153 ^ n52403;
  assign n55156 = n55155 ^ n55154;
  assign n55160 = n55159 ^ n55156;
  assign n55161 = n55160 ^ n51798;
  assign n55165 = n55164 ^ n55161;
  assign n55151 = ~n55137 & ~n55150;
  assign n54787 = n53299 ^ n45645;
  assign n54788 = n54787 ^ n49812;
  assign n54789 = n54788 ^ n44310;
  assign n55152 = n55151 ^ n54789;
  assign n55166 = n55165 ^ n55152;
  assign n55370 = n55369 ^ n55166;
  assign n55373 = n55372 ^ n55370;
  assign n55381 = n53847 ^ n53232;
  assign n55382 = n55381 ^ n54868;
  assign n55376 = n55345 ^ n55172;
  assign n55377 = n55376 ^ n55343;
  assign n55378 = n54761 ^ n53852;
  assign n55379 = n55378 ^ n53237;
  assign n55380 = n55377 & ~n55379;
  assign n55383 = n55382 ^ n55380;
  assign n55384 = n55352 ^ n55349;
  assign n55385 = n55384 ^ n55382;
  assign n55386 = n55383 & n55385;
  assign n55387 = n55386 ^ n55380;
  assign n55375 = n55359 ^ n55356;
  assign n55388 = n55387 ^ n55375;
  assign n55389 = n54863 ^ n53227;
  assign n55390 = n55389 ^ n53840;
  assign n55391 = n55390 ^ n55375;
  assign n55392 = n55388 & ~n55391;
  assign n55393 = n55392 ^ n55390;
  assign n55374 = n55366 ^ n55363;
  assign n55394 = n55393 ^ n55374;
  assign n55395 = n53836 ^ n53223;
  assign n55396 = n55395 ^ n54858;
  assign n55397 = n55396 ^ n55374;
  assign n55398 = n55394 & n55397;
  assign n55399 = n55398 ^ n55396;
  assign n55400 = n55399 ^ n55370;
  assign n55401 = n55373 & ~n55400;
  assign n55402 = n55401 ^ n55372;
  assign n54786 = n54730 ^ n54729;
  assign n55403 = n55402 ^ n54786;
  assign n55404 = n54849 ^ n53834;
  assign n55405 = n55404 ^ n53217;
  assign n55406 = n55405 ^ n54786;
  assign n55407 = n55403 & n55406;
  assign n55408 = n55407 ^ n55405;
  assign n54784 = n54726 ^ n54713;
  assign n54785 = n54784 ^ n54731;
  assign n55409 = n55408 ^ n54785;
  assign n55410 = n54845 ^ n53213;
  assign n55411 = n55410 ^ n53833;
  assign n55412 = n55411 ^ n54785;
  assign n55413 = n55409 & n55412;
  assign n55414 = n55413 ^ n55411;
  assign n54783 = n54739 ^ n54736;
  assign n55415 = n55414 ^ n54783;
  assign n55416 = n53830 ^ n53210;
  assign n55417 = n55416 ^ n54839;
  assign n55418 = n55417 ^ n54783;
  assign n55419 = n55415 & n55418;
  assign n55420 = n55419 ^ n55417;
  assign n54782 = n54744 ^ n54743;
  assign n55421 = n55420 ^ n54782;
  assign n55422 = n54836 ^ n53384;
  assign n55423 = n55422 ^ n53826;
  assign n55424 = n55423 ^ n54782;
  assign n55425 = n55421 & n55424;
  assign n55426 = n55425 ^ n55423;
  assign n55427 = n55426 ^ n54780;
  assign n55428 = ~n54781 & ~n55427;
  assign n55429 = n55428 ^ n54779;
  assign n54772 = n53819 ^ n53203;
  assign n54775 = n54774 ^ n54772;
  assign n55509 = n55429 ^ n54775;
  assign n54771 = n54770 ^ n54750;
  assign n55510 = n55429 ^ n54771;
  assign n55511 = ~n55509 & n55510;
  assign n55512 = n55511 ^ n54775;
  assign n55508 = n55268 ^ n55265;
  assign n55513 = n55512 ^ n55508;
  assign n55506 = n54826 ^ n54121;
  assign n55507 = n55506 ^ n53196;
  assign n55525 = n55508 ^ n55507;
  assign n55526 = n55513 & ~n55525;
  assign n55527 = n55526 ^ n55507;
  assign n55524 = n55275 ^ n55272;
  assign n55528 = n55527 ^ n55524;
  assign n55522 = n54822 ^ n54128;
  assign n55523 = n55522 ^ n53194;
  assign n55536 = n55524 ^ n55523;
  assign n55537 = n55528 & n55536;
  assign n55538 = n55537 ^ n55523;
  assign n55551 = n55542 ^ n55538;
  assign n55552 = ~n55550 & n55551;
  assign n55553 = n55552 ^ n55540;
  assign n55569 = n55557 ^ n55553;
  assign n55570 = ~n55558 & n55569;
  assign n55571 = n55570 ^ n55555;
  assign n55568 = n55284 ^ n55249;
  assign n55572 = n55571 ^ n55568;
  assign n55566 = n54814 ^ n53805;
  assign n55567 = n55566 ^ n53741;
  assign n55580 = n55568 ^ n55567;
  assign n55581 = ~n55572 & ~n55580;
  assign n55582 = n55581 ^ n55567;
  assign n55591 = n55585 ^ n55582;
  assign n55592 = ~n55586 & n55591;
  assign n55593 = n55592 ^ n55584;
  assign n55609 = n55596 ^ n55593;
  assign n55610 = n55597 & n55609;
  assign n55611 = n55610 ^ n55594;
  assign n55809 = n55614 ^ n55611;
  assign n55810 = ~n55615 & ~n55809;
  assign n55811 = n55810 ^ n55613;
  assign n55837 = n55815 ^ n55811;
  assign n55838 = n55816 & n55837;
  assign n55839 = n55838 ^ n55813;
  assign n55836 = n55299 ^ n55224;
  assign n55840 = n55839 ^ n55836;
  assign n55834 = n54941 ^ n53802;
  assign n55835 = n55834 ^ n53776;
  assign n55861 = n55836 ^ n55835;
  assign n55862 = ~n55840 & ~n55861;
  assign n55863 = n55862 ^ n55835;
  assign n55882 = n55866 ^ n55863;
  assign n55883 = ~n55867 & ~n55882;
  assign n55884 = n55883 ^ n55864;
  assign n55904 = n55888 ^ n55884;
  assign n55905 = n55889 & n55904;
  assign n55906 = n55905 ^ n55886;
  assign n55939 = n55910 ^ n55906;
  assign n55940 = ~n55911 & ~n55939;
  assign n55941 = n55940 ^ n55908;
  assign n55938 = n55311 ^ n55204;
  assign n55942 = n55941 ^ n55938;
  assign n55936 = n55126 ^ n53779;
  assign n55937 = n55936 ^ n54687;
  assign n55958 = n55938 ^ n55937;
  assign n55959 = ~n55942 & n55958;
  assign n55960 = n55959 ^ n55937;
  assign n55991 = n55964 ^ n55960;
  assign n55992 = n55965 & ~n55991;
  assign n55993 = n55992 ^ n55962;
  assign n55989 = n55317 ^ n55192;
  assign n55990 = n55989 ^ n55193;
  assign n55994 = n55993 ^ n55990;
  assign n55987 = n55155 ^ n53181;
  assign n55988 = n55987 ^ n54048;
  assign n56009 = n55990 ^ n55988;
  assign n56010 = n55994 & ~n56009;
  assign n56011 = n56010 ^ n55988;
  assign n56036 = n56014 ^ n56011;
  assign n56037 = ~n56015 & n56036;
  assign n56038 = n56037 ^ n56013;
  assign n56056 = n56041 ^ n56038;
  assign n56057 = n56042 & n56056;
  assign n56058 = n56057 ^ n56040;
  assign n56089 = n56061 ^ n56058;
  assign n56090 = ~n56062 & n56089;
  assign n56091 = n56090 ^ n56059;
  assign n56087 = n55333 ^ n55330;
  assign n56085 = n54640 ^ n53246;
  assign n56086 = n56085 ^ n53861;
  assign n56088 = n56087 ^ n56086;
  assign n56092 = n56091 ^ n56088;
  assign n56093 = n56092 ^ n52409;
  assign n56063 = n56062 ^ n56058;
  assign n56064 = n56063 ^ n52625;
  assign n56043 = n56042 ^ n56038;
  assign n56044 = n56043 ^ n52649;
  assign n56016 = n56015 ^ n56011;
  assign n56017 = n56016 ^ n52627;
  assign n55995 = n55994 ^ n55988;
  assign n55996 = n55995 ^ n52639;
  assign n55943 = n55942 ^ n55937;
  assign n55944 = n55943 ^ n53254;
  assign n55890 = n55889 ^ n55884;
  assign n55891 = n55890 ^ n53260;
  assign n55868 = n55867 ^ n55863;
  assign n55869 = n55868 ^ n53169;
  assign n55841 = n55840 ^ n55835;
  assign n55842 = n55841 ^ n52747;
  assign n55817 = n55816 ^ n55811;
  assign n55818 = n55817 ^ n52329;
  assign n55616 = n55615 ^ n55611;
  assign n55617 = n55616 ^ n52331;
  assign n55587 = n55586 ^ n55582;
  assign n55588 = n55587 ^ n52340;
  assign n55573 = n55572 ^ n55567;
  assign n55574 = n55573 ^ n52345;
  assign n55559 = n55558 ^ n55553;
  assign n55560 = n55559 ^ n52351;
  assign n55541 = n55540 ^ n55538;
  assign n55543 = n55542 ^ n55541;
  assign n55544 = n55543 ^ n52356;
  assign n55529 = n55528 ^ n55523;
  assign n55532 = n55529 ^ n52362;
  assign n55514 = n55513 ^ n55507;
  assign n55515 = n55514 ^ n52367;
  assign n55431 = n55426 ^ n54781;
  assign n55432 = n55431 ^ n52371;
  assign n55433 = n55423 ^ n55421;
  assign n55434 = n55433 ^ n52376;
  assign n55435 = n55417 ^ n55415;
  assign n55436 = n55435 ^ n52693;
  assign n55437 = n55411 ^ n55409;
  assign n55438 = n55437 ^ n52380;
  assign n55440 = n55399 ^ n55372;
  assign n55441 = n55440 ^ n55370;
  assign n55442 = n55441 ^ n52385;
  assign n55443 = n55396 ^ n55394;
  assign n55444 = n55443 ^ n52389;
  assign n55445 = n55390 ^ n55388;
  assign n55446 = n55445 ^ n52394;
  assign n55447 = n55379 ^ n55377;
  assign n55448 = ~n52398 & ~n55447;
  assign n55449 = n55448 ^ n52397;
  assign n55450 = n55384 ^ n55383;
  assign n55451 = n55450 ^ n55448;
  assign n55452 = ~n55449 & n55451;
  assign n55453 = n55452 ^ n52397;
  assign n55454 = n55453 ^ n55445;
  assign n55455 = n55446 & ~n55454;
  assign n55456 = n55455 ^ n52394;
  assign n55457 = n55456 ^ n55443;
  assign n55458 = n55444 & n55457;
  assign n55459 = n55458 ^ n52389;
  assign n55460 = n55459 ^ n55441;
  assign n55461 = n55442 & n55460;
  assign n55462 = n55461 ^ n52385;
  assign n55439 = n55405 ^ n55403;
  assign n55463 = n55462 ^ n55439;
  assign n55464 = n55439 ^ n52683;
  assign n55465 = ~n55463 & n55464;
  assign n55466 = n55465 ^ n52683;
  assign n55467 = n55466 ^ n55437;
  assign n55468 = n55438 & n55467;
  assign n55469 = n55468 ^ n52380;
  assign n55470 = n55469 ^ n55435;
  assign n55471 = n55436 & n55470;
  assign n55472 = n55471 ^ n52693;
  assign n55473 = n55472 ^ n55433;
  assign n55474 = n55434 & n55473;
  assign n55475 = n55474 ^ n52376;
  assign n55476 = n55475 ^ n55431;
  assign n55477 = ~n55432 & ~n55476;
  assign n55478 = n55477 ^ n52371;
  assign n54776 = n54775 ^ n54771;
  assign n55430 = n55429 ^ n54776;
  assign n55479 = n55478 ^ n55430;
  assign n55503 = n55430 ^ n52707;
  assign n55504 = n55479 & n55503;
  assign n55505 = n55504 ^ n52707;
  assign n55518 = n55514 ^ n55505;
  assign n55519 = ~n55515 & ~n55518;
  assign n55520 = n55519 ^ n52367;
  assign n55533 = n55529 ^ n55520;
  assign n55534 = n55532 & ~n55533;
  assign n55535 = n55534 ^ n52362;
  assign n55547 = n55543 ^ n55535;
  assign n55548 = ~n55544 & ~n55547;
  assign n55549 = n55548 ^ n52356;
  assign n55563 = n55559 ^ n55549;
  assign n55564 = ~n55560 & n55563;
  assign n55565 = n55564 ^ n52351;
  assign n55577 = n55573 ^ n55565;
  assign n55578 = ~n55574 & n55577;
  assign n55579 = n55578 ^ n52345;
  assign n55600 = n55587 ^ n55579;
  assign n55601 = ~n55588 & ~n55600;
  assign n55602 = n55601 ^ n52340;
  assign n55605 = n55602 ^ n52332;
  assign n55598 = n55597 ^ n55593;
  assign n55606 = n55602 ^ n55598;
  assign n55607 = ~n55605 & ~n55606;
  assign n55608 = n55607 ^ n52332;
  assign n55806 = n55616 ^ n55608;
  assign n55807 = n55617 & n55806;
  assign n55808 = n55807 ^ n52331;
  assign n55831 = n55817 ^ n55808;
  assign n55832 = n55818 & ~n55831;
  assign n55833 = n55832 ^ n52329;
  assign n55858 = n55841 ^ n55833;
  assign n55859 = ~n55842 & ~n55858;
  assign n55860 = n55859 ^ n52747;
  assign n55879 = n55868 ^ n55860;
  assign n55880 = n55869 & ~n55879;
  assign n55881 = n55880 ^ n53169;
  assign n55913 = n55890 ^ n55881;
  assign n55914 = n55891 & ~n55913;
  assign n55915 = n55914 ^ n53260;
  assign n55912 = n55911 ^ n55906;
  assign n55916 = n55915 ^ n55912;
  assign n55933 = n55912 ^ n53258;
  assign n55934 = ~n55916 & n55933;
  assign n55935 = n55934 ^ n53258;
  assign n55967 = n55943 ^ n55935;
  assign n55968 = ~n55944 & ~n55967;
  assign n55969 = n55968 ^ n53254;
  assign n55966 = n55965 ^ n55960;
  assign n55970 = n55969 ^ n55966;
  assign n55984 = n55966 ^ n52634;
  assign n55985 = n55970 & n55984;
  assign n55986 = n55985 ^ n52634;
  assign n56006 = n55995 ^ n55986;
  assign n56007 = n55996 & n56006;
  assign n56008 = n56007 ^ n52639;
  assign n56033 = n56016 ^ n56008;
  assign n56034 = n56017 & ~n56033;
  assign n56035 = n56034 ^ n52627;
  assign n56053 = n56043 ^ n56035;
  assign n56054 = n56044 & n56053;
  assign n56055 = n56054 ^ n52649;
  assign n56082 = n56063 ^ n56055;
  assign n56083 = ~n56064 & ~n56082;
  assign n56084 = n56083 ^ n52625;
  assign n56094 = n56093 ^ n56084;
  assign n56065 = n56064 ^ n56055;
  assign n55917 = n55916 ^ n53258;
  assign n55870 = n55869 ^ n55860;
  assign n55480 = n55479 ^ n52707;
  assign n55481 = n55456 ^ n52389;
  assign n55482 = n55481 ^ n55443;
  assign n55483 = n55450 ^ n55449;
  assign n55484 = n55453 ^ n55446;
  assign n55485 = ~n55483 & n55484;
  assign n55486 = ~n55482 & ~n55485;
  assign n55487 = n55459 ^ n52385;
  assign n55488 = n55487 ^ n55441;
  assign n55489 = ~n55486 & ~n55488;
  assign n55490 = n55463 ^ n52683;
  assign n55491 = ~n55489 & ~n55490;
  assign n55492 = n55466 ^ n52380;
  assign n55493 = n55492 ^ n55437;
  assign n55494 = ~n55491 & n55493;
  assign n55495 = n55469 ^ n55436;
  assign n55496 = n55494 & ~n55495;
  assign n55497 = n55472 ^ n52376;
  assign n55498 = n55497 ^ n55433;
  assign n55499 = n55496 & n55498;
  assign n55500 = n55475 ^ n55432;
  assign n55501 = ~n55499 & ~n55500;
  assign n55502 = ~n55480 & n55501;
  assign n55516 = n55515 ^ n55505;
  assign n55517 = n55502 & ~n55516;
  assign n55521 = n55520 ^ n52362;
  assign n55530 = n55529 ^ n55521;
  assign n55531 = n55517 & ~n55530;
  assign n55545 = n55544 ^ n55535;
  assign n55546 = n55531 & n55545;
  assign n55561 = n55560 ^ n55549;
  assign n55562 = ~n55546 & n55561;
  assign n55575 = n55574 ^ n55565;
  assign n55576 = n55562 & n55575;
  assign n55589 = n55588 ^ n55579;
  assign n55590 = ~n55576 & ~n55589;
  assign n55599 = n55598 ^ n52332;
  assign n55603 = n55602 ^ n55599;
  assign n55604 = ~n55590 & ~n55603;
  assign n55618 = n55617 ^ n55608;
  assign n55805 = ~n55604 & n55618;
  assign n55819 = n55818 ^ n55808;
  assign n55830 = n55805 & ~n55819;
  assign n55843 = n55842 ^ n55833;
  assign n55871 = n55830 & n55843;
  assign n55878 = ~n55870 & ~n55871;
  assign n55892 = n55891 ^ n55881;
  assign n55918 = n55878 & ~n55892;
  assign n55932 = n55917 & ~n55918;
  assign n55945 = n55944 ^ n55935;
  assign n55957 = n55932 & ~n55945;
  assign n55971 = n55970 ^ n52634;
  assign n55983 = ~n55957 & n55971;
  assign n55997 = n55996 ^ n55986;
  assign n56005 = ~n55983 & n55997;
  assign n56018 = n56017 ^ n56008;
  assign n56032 = ~n56005 & n56018;
  assign n56045 = n56044 ^ n56035;
  assign n56066 = ~n56032 & ~n56045;
  assign n56081 = ~n56065 & n56066;
  assign n56095 = n56094 ^ n56081;
  assign n56077 = n53986 ^ n46315;
  assign n56078 = n56077 ^ n50472;
  assign n56079 = n56078 ^ n44927;
  assign n56118 = n56095 ^ n56079;
  assign n56046 = n56045 ^ n56032;
  assign n56029 = n53995 ^ n46325;
  assign n56030 = n56029 ^ n50483;
  assign n56031 = n56030 ^ n44999;
  assign n56047 = n56046 ^ n56031;
  assign n56020 = n54000 ^ n46330;
  assign n56021 = n56020 ^ n50492;
  assign n56022 = n56021 ^ n44938;
  assign n56019 = n56018 ^ n56005;
  assign n56023 = n56022 ^ n56019;
  assign n55998 = n55997 ^ n55983;
  assign n55979 = n54019 ^ n46336;
  assign n55980 = n55979 ^ n50335;
  assign n55981 = n55980 ^ n44943;
  assign n56001 = n55998 ^ n55981;
  assign n55972 = n55971 ^ n55957;
  assign n55953 = n54012 ^ n46340;
  assign n55954 = n55953 ^ n49707;
  assign n55955 = n55954 ^ n3119;
  assign n55975 = n55972 ^ n55955;
  assign n55946 = n55945 ^ n55932;
  assign n55929 = n53755 ^ n46345;
  assign n55930 = n55929 ^ n50147;
  assign n55931 = n55930 ^ n2738;
  assign n55947 = n55946 ^ n55931;
  assign n55872 = n55871 ^ n55870;
  assign n55854 = n53568 ^ n45500;
  assign n55855 = n55854 ^ n50158;
  assign n55856 = n55855 ^ n44956;
  assign n55894 = n55872 ^ n55856;
  assign n55845 = n53573 ^ n45929;
  assign n55846 = n55845 ^ n50310;
  assign n55847 = n55846 ^ n44966;
  assign n55844 = n55843 ^ n55830;
  assign n55848 = n55847 ^ n55844;
  assign n55821 = n53579 ^ n46069;
  assign n55822 = n55821 ^ n50164;
  assign n55823 = n55822 ^ n44117;
  assign n55820 = n55819 ^ n55805;
  assign n55824 = n55823 ^ n55820;
  assign n55621 = n53711 ^ n1468;
  assign n55622 = n55621 ^ n50170;
  assign n55623 = n55622 ^ n46059;
  assign n55620 = n55603 ^ n55590;
  assign n55624 = n55623 ^ n55620;
  assign n55628 = n55589 ^ n55576;
  assign n55625 = n53587 ^ n1254;
  assign n55626 = n55625 ^ n50175;
  assign n55627 = n55626 ^ n44552;
  assign n55629 = n55628 ^ n55627;
  assign n55631 = n53701 ^ n45940;
  assign n55632 = n55631 ^ n50181;
  assign n55633 = n55632 ^ n44557;
  assign n55630 = n55575 ^ n55562;
  assign n55634 = n55633 ^ n55630;
  assign n55638 = n55561 ^ n55546;
  assign n55635 = n53592 ^ n45944;
  assign n55636 = n55635 ^ n50185;
  assign n55637 = n55636 ^ n44562;
  assign n55639 = n55638 ^ n55637;
  assign n55644 = n55530 ^ n55517;
  assign n55641 = n53598 ^ n45954;
  assign n55642 = n55641 ^ n50281;
  assign n55643 = n55642 ^ n44572;
  assign n55645 = n55644 ^ n55643;
  assign n55649 = n55516 ^ n55502;
  assign n55646 = n53604 ^ n45959;
  assign n55647 = n55646 ^ n50196;
  assign n55648 = n55647 ^ n44577;
  assign n55650 = n55649 ^ n55648;
  assign n55652 = n53608 ^ n45965;
  assign n55653 = n55652 ^ n50271;
  assign n55654 = n55653 ^ n44652;
  assign n55651 = n55501 ^ n55480;
  assign n55655 = n55654 ^ n55651;
  assign n55659 = n55500 ^ n55499;
  assign n55656 = n53613 ^ n45970;
  assign n55657 = n55656 ^ n50202;
  assign n55658 = n55657 ^ n44584;
  assign n55660 = n55659 ^ n55658;
  assign n55664 = n55498 ^ n55496;
  assign n55661 = n53619 ^ n45975;
  assign n55662 = n55661 ^ n50207;
  assign n55663 = n55662 ^ n44642;
  assign n55665 = n55664 ^ n55663;
  assign n55669 = n55495 ^ n55494;
  assign n55666 = n53624 ^ n45979;
  assign n55667 = n55666 ^ n50210;
  assign n55668 = n55667 ^ n44590;
  assign n55670 = n55669 ^ n55668;
  assign n55674 = n55493 ^ n55491;
  assign n55671 = n53666 ^ n50215;
  assign n55672 = n55671 ^ n45985;
  assign n55673 = n55672 ^ n44632;
  assign n55675 = n55674 ^ n55673;
  assign n55679 = n55490 ^ n55489;
  assign n55676 = n53629 ^ n46019;
  assign n55677 = n55676 ^ n50218;
  assign n55678 = n55677 ^ n44595;
  assign n55680 = n55679 ^ n55678;
  assign n55684 = n55488 ^ n55486;
  assign n55681 = n53632 ^ n46012;
  assign n55682 = n55681 ^ n50221;
  assign n55683 = n55682 ^ n44600;
  assign n55685 = n55684 ^ n55683;
  assign n55693 = n53963 ^ n46296;
  assign n55694 = n55693 ^ n50381;
  assign n55695 = n55694 ^ n1940;
  assign n55696 = n55447 ^ n52398;
  assign n55697 = n55695 & n55696;
  assign n55690 = n53641 ^ n46000;
  assign n55691 = n55690 ^ n50231;
  assign n55692 = n55691 ^ n44613;
  assign n55698 = n55697 ^ n55692;
  assign n55699 = n55697 ^ n55483;
  assign n55700 = n55698 & n55699;
  assign n55701 = n55700 ^ n55692;
  assign n55687 = n53638 ^ n45996;
  assign n55688 = n55687 ^ n50236;
  assign n55689 = n55688 ^ n44610;
  assign n55702 = n55701 ^ n55689;
  assign n55703 = n55484 ^ n55483;
  assign n55704 = n55703 ^ n55701;
  assign n55705 = n55702 & ~n55704;
  assign n55706 = n55705 ^ n55689;
  assign n55686 = n55485 ^ n55482;
  assign n55707 = n55706 ^ n55686;
  assign n55708 = n53635 ^ n45991;
  assign n55709 = n55708 ^ n50226;
  assign n55710 = n55709 ^ n44606;
  assign n55711 = n55710 ^ n55686;
  assign n55712 = ~n55707 & n55711;
  assign n55713 = n55712 ^ n55710;
  assign n55714 = n55713 ^ n55684;
  assign n55715 = ~n55685 & n55714;
  assign n55716 = n55715 ^ n55683;
  assign n55717 = n55716 ^ n55679;
  assign n55718 = n55680 & ~n55717;
  assign n55719 = n55718 ^ n55678;
  assign n55720 = n55719 ^ n55674;
  assign n55721 = n55675 & ~n55720;
  assign n55722 = n55721 ^ n55673;
  assign n55723 = n55722 ^ n55669;
  assign n55724 = n55670 & ~n55723;
  assign n55725 = n55724 ^ n55668;
  assign n55726 = n55725 ^ n55664;
  assign n55727 = ~n55665 & n55726;
  assign n55728 = n55727 ^ n55663;
  assign n55729 = n55728 ^ n55659;
  assign n55730 = n55660 & ~n55729;
  assign n55731 = n55730 ^ n55658;
  assign n55732 = n55731 ^ n55654;
  assign n55733 = ~n55655 & ~n55732;
  assign n55734 = n55733 ^ n55651;
  assign n55735 = n55734 ^ n55649;
  assign n55736 = ~n55650 & ~n55735;
  assign n55737 = n55736 ^ n55648;
  assign n55738 = n55737 ^ n55644;
  assign n55739 = ~n55645 & n55738;
  assign n55740 = n55739 ^ n55643;
  assign n55640 = n55545 ^ n55531;
  assign n55741 = n55740 ^ n55640;
  assign n55742 = n53691 ^ n45950;
  assign n55743 = n55742 ^ n50190;
  assign n55744 = n55743 ^ n44567;
  assign n55745 = n55744 ^ n55640;
  assign n55746 = ~n55741 & n55745;
  assign n55747 = n55746 ^ n55744;
  assign n55748 = n55747 ^ n55638;
  assign n55749 = n55639 & ~n55748;
  assign n55750 = n55749 ^ n55637;
  assign n55751 = n55750 ^ n55633;
  assign n55752 = ~n55634 & ~n55751;
  assign n55753 = n55752 ^ n55630;
  assign n55754 = n55753 ^ n55628;
  assign n55755 = n55629 & n55754;
  assign n55756 = n55755 ^ n55627;
  assign n55757 = n55756 ^ n55623;
  assign n55758 = ~n55624 & ~n55757;
  assign n55759 = n55758 ^ n55620;
  assign n55619 = n55618 ^ n55604;
  assign n55760 = n55759 ^ n55619;
  assign n1440 = n1439 ^ n1373;
  assign n1477 = n1476 ^ n1440;
  assign n1487 = n1486 ^ n1477;
  assign n55802 = n55619 ^ n1487;
  assign n55803 = ~n55760 & ~n55802;
  assign n55804 = n55803 ^ n1487;
  assign n55827 = n55823 ^ n55804;
  assign n55828 = ~n55824 & ~n55827;
  assign n55829 = n55828 ^ n55820;
  assign n55851 = n55847 ^ n55829;
  assign n55852 = n55848 & n55851;
  assign n55853 = n55852 ^ n55844;
  assign n55895 = n55872 ^ n55853;
  assign n55896 = ~n55894 & n55895;
  assign n55897 = n55896 ^ n55856;
  assign n55893 = n55892 ^ n55878;
  assign n55898 = n55897 ^ n55893;
  assign n55875 = n53730 ^ n46355;
  assign n55876 = n55875 ^ n50153;
  assign n55877 = n55876 ^ n44951;
  assign n55920 = n55893 ^ n55877;
  assign n55921 = ~n55898 & n55920;
  assign n55922 = n55921 ^ n55877;
  assign n55919 = n55918 ^ n55917;
  assign n55923 = n55922 ^ n55919;
  assign n55901 = n53186 ^ n46351;
  assign n55902 = n55901 ^ n50323;
  assign n55903 = n55902 ^ n44979;
  assign n55926 = n55919 ^ n55903;
  assign n55927 = n55923 & ~n55926;
  assign n55928 = n55927 ^ n55903;
  assign n55950 = n55946 ^ n55928;
  assign n55951 = ~n55947 & n55950;
  assign n55952 = n55951 ^ n55931;
  assign n55976 = n55972 ^ n55952;
  assign n55977 = n55975 & ~n55976;
  assign n55978 = n55977 ^ n55955;
  assign n56002 = n55998 ^ n55978;
  assign n56003 = ~n56001 & n56002;
  assign n56004 = n56003 ^ n55981;
  assign n56026 = n56022 ^ n56004;
  assign n56027 = n56023 & ~n56026;
  assign n56028 = n56027 ^ n56019;
  assign n56068 = n56046 ^ n56028;
  assign n56069 = n56047 & ~n56068;
  assign n56070 = n56069 ^ n56031;
  assign n56067 = n56066 ^ n56065;
  assign n56071 = n56070 ^ n56067;
  assign n56050 = n53990 ^ n46321;
  assign n56051 = n56050 ^ n50477;
  assign n56052 = n56051 ^ n44932;
  assign n56074 = n56067 ^ n56052;
  assign n56075 = n56071 & ~n56074;
  assign n56076 = n56075 ^ n56052;
  assign n56119 = n56095 ^ n56076;
  assign n56120 = n56118 & ~n56119;
  assign n56121 = n56120 ^ n56079;
  assign n56115 = ~n56081 & n56094;
  assign n56109 = n56084 ^ n52409;
  assign n56110 = n56092 ^ n56084;
  assign n56111 = ~n56109 & n56110;
  assign n56112 = n56111 ^ n52409;
  assign n56105 = n56091 ^ n56086;
  assign n56106 = n56088 & ~n56105;
  assign n56107 = n56106 ^ n56091;
  assign n56103 = n55340 ^ n55337;
  assign n56101 = n54709 ^ n53857;
  assign n56102 = n56101 ^ n53242;
  assign n56104 = n56103 ^ n56102;
  assign n56108 = n56107 ^ n56104;
  assign n56113 = n56112 ^ n56108;
  assign n56114 = n56113 ^ n52403;
  assign n56116 = n56115 ^ n56114;
  assign n56098 = n53980 ^ n46391;
  assign n56099 = n56098 ^ n50508;
  assign n56100 = n56099 ^ n45012;
  assign n56117 = n56116 ^ n56100;
  assign n56122 = n56121 ^ n56117;
  assign n55761 = n55760 ^ n1487;
  assign n55762 = n55696 ^ n55695;
  assign n55763 = n55692 ^ n55483;
  assign n55764 = n55763 ^ n55697;
  assign n55765 = n55762 & ~n55764;
  assign n55766 = n55703 ^ n55689;
  assign n55767 = n55766 ^ n55701;
  assign n55768 = n55765 & n55767;
  assign n55769 = n55710 ^ n55707;
  assign n55770 = n55768 & n55769;
  assign n55771 = n55713 ^ n55683;
  assign n55772 = n55771 ^ n55684;
  assign n55773 = n55770 & ~n55772;
  assign n55774 = n55716 ^ n55680;
  assign n55775 = n55773 & n55774;
  assign n55776 = n55719 ^ n55675;
  assign n55777 = n55775 & n55776;
  assign n55778 = n55722 ^ n55668;
  assign n55779 = n55778 ^ n55669;
  assign n55780 = n55777 & n55779;
  assign n55781 = n55725 ^ n55665;
  assign n55782 = ~n55780 & n55781;
  assign n55783 = n55728 ^ n55660;
  assign n55784 = n55782 & ~n55783;
  assign n55785 = n55731 ^ n55655;
  assign n55786 = ~n55784 & ~n55785;
  assign n55787 = n55734 ^ n55650;
  assign n55788 = n55786 & n55787;
  assign n55789 = n55737 ^ n55645;
  assign n55790 = n55788 & ~n55789;
  assign n55791 = n55744 ^ n55741;
  assign n55792 = ~n55790 & ~n55791;
  assign n55793 = n55747 ^ n55639;
  assign n55794 = ~n55792 & n55793;
  assign n55795 = n55750 ^ n55634;
  assign n55796 = n55794 & ~n55795;
  assign n55797 = n55753 ^ n55629;
  assign n55798 = ~n55796 & n55797;
  assign n55799 = n55756 ^ n55624;
  assign n55800 = ~n55798 & ~n55799;
  assign n55801 = ~n55761 & ~n55800;
  assign n55825 = n55824 ^ n55804;
  assign n55826 = ~n55801 & ~n55825;
  assign n55849 = n55848 ^ n55829;
  assign n55850 = n55826 & ~n55849;
  assign n55857 = n55856 ^ n55853;
  assign n55873 = n55872 ^ n55857;
  assign n55874 = n55850 & ~n55873;
  assign n55899 = n55898 ^ n55877;
  assign n55900 = ~n55874 & ~n55899;
  assign n55924 = n55923 ^ n55903;
  assign n55925 = ~n55900 & ~n55924;
  assign n55948 = n55947 ^ n55928;
  assign n55949 = ~n55925 & n55948;
  assign n55956 = n55955 ^ n55952;
  assign n55973 = n55972 ^ n55956;
  assign n55974 = n55949 & ~n55973;
  assign n55982 = n55981 ^ n55978;
  assign n55999 = n55998 ^ n55982;
  assign n56000 = n55974 & n55999;
  assign n56024 = n56023 ^ n56004;
  assign n56025 = ~n56000 & n56024;
  assign n56048 = n56047 ^ n56028;
  assign n56049 = n56025 & n56048;
  assign n56072 = n56071 ^ n56052;
  assign n56073 = ~n56049 & n56072;
  assign n56080 = n56079 ^ n56076;
  assign n56096 = n56095 ^ n56080;
  assign n56097 = n56073 & ~n56096;
  assign n56123 = n56122 ^ n56097;
  assign n56124 = n56096 ^ n56073;
  assign n56125 = n56072 ^ n56049;
  assign n56126 = n56048 ^ n56025;
  assign n56127 = n56024 ^ n56000;
  assign n56128 = n55999 ^ n55974;
  assign n56129 = n55973 ^ n55949;
  assign n56130 = n55948 ^ n55925;
  assign n56131 = n55924 ^ n55900;
  assign n56132 = n55899 ^ n55874;
  assign n56133 = n55873 ^ n55850;
  assign n56134 = n55849 ^ n55826;
  assign n56135 = n55825 ^ n55801;
  assign n56136 = n55800 ^ n55761;
  assign n56137 = n55799 ^ n55798;
  assign n56138 = n55797 ^ n55796;
  assign n56139 = n55795 ^ n55794;
  assign n56140 = n55793 ^ n55792;
  assign n56141 = n55791 ^ n55790;
  assign n56142 = n55789 ^ n55788;
  assign n56143 = n55787 ^ n55786;
  assign n56144 = n55785 ^ n55784;
  assign n56145 = n55783 ^ n55782;
  assign n56146 = n55781 ^ n55780;
  assign n56147 = n55779 ^ n55777;
  assign n56148 = n55776 ^ n55775;
  assign n56149 = n55774 ^ n55773;
  assign n56150 = n55772 ^ n55770;
  assign n56151 = n55769 ^ n55768;
  assign n56152 = n55767 ^ n55765;
  assign n56153 = n55764 ^ n55762;
  assign n56154 = ~n54785 & n54786;
  assign n56155 = n54783 & n56154;
  assign n56156 = n54782 & ~n56155;
  assign n56157 = ~n54780 & ~n56156;
  assign n56158 = ~n54771 & n56157;
  assign n56159 = n55508 & n56158;
  assign n56160 = ~n55524 & ~n56159;
  assign n56161 = n55542 & n56160;
  assign n56162 = n55557 & n56161;
  assign n56163 = n55568 & ~n56162;
  assign n56164 = ~n55585 & ~n56163;
  assign n56165 = n55594 & ~n56164;
  assign n56166 = ~n55614 & ~n56165;
  assign n56167 = n55815 & ~n56166;
  assign n56168 = ~n55836 & ~n56167;
  assign n56169 = ~n55864 & n56168;
  assign n56170 = ~n55888 & ~n56169;
  assign n56171 = n55910 & ~n56170;
  assign n56172 = ~n55938 & n56171;
  assign n56173 = n55962 & ~n56172;
  assign n56174 = ~n55990 & n56173;
  assign n56175 = n56014 & ~n56174;
  assign n56176 = n56041 & n56175;
  assign n56177 = n56059 & n56176;
  assign n56178 = n56087 & n56177;
  assign n56179 = ~n56103 & n56178;
  assign n56180 = ~n55377 & n56179;
  assign n56181 = ~n55384 & ~n56180;
  assign n56182 = n55375 & ~n56181;
  assign n56183 = n55374 & n56182;
  assign n56184 = n56183 ^ n55370;
  assign n56185 = n56182 ^ n55374;
  assign n56186 = n56181 ^ n55375;
  assign n56187 = n56180 ^ n55384;
  assign n56188 = n56179 ^ n55377;
  assign n56189 = n56178 ^ n56103;
  assign n56190 = n56177 ^ n56087;
  assign n56191 = n56176 ^ n56059;
  assign n56192 = n56175 ^ n56041;
  assign n56193 = n56174 ^ n56014;
  assign n56194 = n56173 ^ n55990;
  assign n56195 = n56172 ^ n55962;
  assign n56196 = n56171 ^ n55938;
  assign n56197 = n56170 ^ n55910;
  assign n56198 = n56169 ^ n55888;
  assign n56199 = n56168 ^ n55864;
  assign n56200 = n56167 ^ n55836;
  assign n56201 = n56166 ^ n55815;
  assign n56202 = n56165 ^ n55614;
  assign n56203 = n56164 ^ n55594;
  assign n56204 = n56163 ^ n55585;
  assign n56205 = n56162 ^ n55568;
  assign n56206 = n56161 ^ n55557;
  assign n56207 = n56160 ^ n55542;
  assign n56208 = n56159 ^ n55524;
  assign n56209 = n56158 ^ n55508;
  assign n56210 = n56157 ^ n54771;
  assign n56211 = n56156 ^ n54780;
  assign n56212 = n56155 ^ n54782;
  assign n56213 = n56154 ^ n54783;
  assign n56214 = n54786 ^ n54785;
  assign n56215 = ~n54853 & n54858;
  assign n56216 = n54849 & n56215;
  assign n56217 = ~n54845 & n56216;
  assign n56218 = ~n54839 & n56217;
  assign n56219 = n54836 & n56218;
  assign n56220 = ~n54777 & n56219;
  assign n56221 = ~n54774 & ~n56220;
  assign n56222 = n54826 & n56221;
  assign n56223 = n54822 & ~n56222;
  assign n56224 = n54819 & n56223;
  assign n56225 = n54815 & n56224;
  assign n56226 = n54814 & ~n56225;
  assign n56227 = n54810 & ~n56226;
  assign n56228 = ~n54808 & n56227;
  assign n56229 = n54805 & ~n56228;
  assign n56230 = n54803 & ~n56229;
  assign n56231 = ~n54941 & ~n56230;
  assign n56232 = n54945 & ~n56231;
  assign n56233 = n54796 & n56232;
  assign n56234 = n54792 & n56233;
  assign n56235 = n55126 & ~n56234;
  assign n56236 = n55143 & ~n56235;
  assign n56237 = n55155 & ~n56236;
  assign n56238 = n54645 & n56237;
  assign n56239 = ~n54652 & n56238;
  assign n56240 = ~n54656 & ~n56239;
  assign n56241 = n54640 & n56240;
  assign n56242 = n54709 & ~n56241;
  assign n56243 = n54761 & n56242;
  assign n56244 = n56243 ^ n54868;
  assign n56245 = n56242 ^ n54761;
  assign n56246 = n56241 ^ n54709;
  assign n56247 = n56240 ^ n54640;
  assign n56248 = n56239 ^ n54656;
  assign n56249 = n56238 ^ n54652;
  assign n56250 = n56237 ^ n54645;
  assign n56251 = n56236 ^ n55155;
  assign n56252 = n56235 ^ n55143;
  assign n56253 = n56234 ^ n55126;
  assign n56254 = n56233 ^ n54792;
  assign n56255 = n56232 ^ n54796;
  assign n56256 = n56231 ^ n54945;
  assign n56257 = n56230 ^ n54941;
  assign n56258 = n56229 ^ n54803;
  assign n56259 = n56228 ^ n54805;
  assign n56260 = n56227 ^ n54808;
  assign n56261 = n56226 ^ n54810;
  assign n56262 = n56225 ^ n54814;
  assign n56263 = n56224 ^ n54815;
  assign n56264 = n56223 ^ n54819;
  assign n56265 = n56222 ^ n54822;
  assign n56266 = n56221 ^ n54826;
  assign n56267 = n56220 ^ n54774;
  assign n56268 = n56219 ^ n54777;
  assign n56269 = n56218 ^ n54836;
  assign n56270 = n56217 ^ n54839;
  assign n56271 = n56216 ^ n54845;
  assign n56272 = n56215 ^ n54849;
  assign n56273 = n54858 ^ n54853;
  assign n56274 = n53840 & ~n53847;
  assign n56275 = n53836 & ~n56274;
  assign n56276 = ~n53835 & ~n56275;
  assign n56277 = n53834 & n56276;
  assign n56278 = n53833 & n56277;
  assign n56279 = n53830 & ~n56278;
  assign n56280 = n53826 & n56279;
  assign n56281 = ~n53820 & n56280;
  assign n56282 = ~n53819 & ~n56281;
  assign n56283 = ~n54121 & ~n56282;
  assign n56284 = ~n54128 & ~n56283;
  assign n56285 = n53813 & ~n56284;
  assign n56286 = ~n53807 & ~n56285;
  assign n56287 = n53805 & ~n56286;
  assign n56288 = n53800 & n56287;
  assign n56289 = ~n53794 & ~n56288;
  assign n56290 = ~n53785 & ~n56289;
  assign n56291 = ~n53782 & n56290;
  assign n56292 = n53776 & ~n56291;
  assign n56293 = n53772 & n56292;
  assign n56294 = n54371 & ~n56293;
  assign n56295 = n54623 & n56294;
  assign n56296 = n54687 & n56295;
  assign n56297 = n54053 & n56296;
  assign n56298 = n54048 & n56297;
  assign n56299 = ~n54059 & n56298;
  assign n56300 = ~n54042 & ~n56299;
  assign n56301 = ~n54038 & ~n56300;
  assign n56302 = n53861 & n56301;
  assign n56303 = n56302 ^ n53857;
  assign n56304 = n56301 ^ n53861;
  assign n56305 = n56300 ^ n54038;
  assign n56306 = n56299 ^ n54042;
  assign n56307 = n56298 ^ n54059;
  assign n56308 = n56297 ^ n54048;
  assign n56309 = n56296 ^ n54053;
  assign n56310 = n56295 ^ n54687;
  assign n56311 = n56294 ^ n54623;
  assign n56312 = n56293 ^ n54371;
  assign n56313 = n56292 ^ n53772;
  assign n56314 = n56291 ^ n53776;
  assign n56315 = n56290 ^ n53782;
  assign n56316 = n56289 ^ n53785;
  assign n56317 = n56288 ^ n53794;
  assign n56318 = n56287 ^ n53800;
  assign n56319 = n56286 ^ n53805;
  assign n56320 = n56285 ^ n53807;
  assign n56321 = n56284 ^ n53813;
  assign n56322 = n56283 ^ n54128;
  assign n56323 = n56282 ^ n54121;
  assign n56324 = n56281 ^ n53819;
  assign n56325 = n56280 ^ n53820;
  assign n56326 = n56279 ^ n53826;
  assign n56327 = n56278 ^ n53830;
  assign n56328 = n56277 ^ n53833;
  assign n56329 = n56276 ^ n53834;
  assign n56330 = n56275 ^ n53835;
  assign n56331 = n56274 ^ n53836;
  assign n56332 = n53847 ^ n53840;
  assign n56333 = ~n53217 & n53219;
  assign n56334 = ~n53213 & n56333;
  assign n56335 = ~n53210 & n56334;
  assign n56336 = ~n53384 & n56335;
  assign n56337 = ~n53206 & ~n56336;
  assign n56338 = n53203 & n56337;
  assign n56339 = n53196 & n56338;
  assign n56340 = ~n53194 & n56339;
  assign n56341 = n53190 & ~n56340;
  assign n56342 = n53409 & n56341;
  assign n56343 = n53741 & n56342;
  assign n56344 = n53762 & ~n56343;
  assign n56345 = ~n53871 & ~n56344;
  assign n56346 = n53815 & ~n56345;
  assign n56347 = n53809 & n56346;
  assign n56348 = n53802 & ~n56347;
  assign n56349 = ~n53797 & ~n56348;
  assign n56350 = ~n53791 & ~n56349;
  assign n56351 = n53787 & n56350;
  assign n56352 = ~n53779 & n56351;
  assign n56353 = n53328 & n56352;
  assign n56354 = n53181 & ~n56353;
  assign n56355 = ~n53326 & n56354;
  assign n56356 = n53319 & n56355;
  assign n56357 = ~n53316 & n56356;
  assign n56358 = n53246 & ~n56357;
  assign n56359 = n56358 ^ n53242;
  assign n56360 = n56357 ^ n53246;
  assign n56361 = n56356 ^ n53316;
  assign n56362 = n56355 ^ n53319;
  assign n56363 = n56354 ^ n53326;
  assign n56364 = n56353 ^ n53181;
  assign n56365 = n56352 ^ n53328;
  assign n56366 = n56351 ^ n53779;
  assign n56367 = n56350 ^ n53787;
  assign n56368 = n56349 ^ n53791;
  assign n56369 = n56348 ^ n53797;
  assign n56370 = n56347 ^ n53802;
  assign n56371 = n56346 ^ n53809;
  assign n56372 = n56345 ^ n53815;
  assign n56373 = n56344 ^ n53871;
  assign n56374 = n56343 ^ n53762;
  assign n56375 = n56342 ^ n53741;
  assign n56376 = n56341 ^ n53409;
  assign n56377 = n56340 ^ n53190;
  assign n56378 = n56339 ^ n53194;
  assign n56379 = n56338 ^ n53196;
  assign n56380 = n56337 ^ n53203;
  assign n56381 = n56336 ^ n53206;
  assign n56382 = n56335 ^ n53384;
  assign n56383 = n56334 ^ n53210;
  assign n56384 = n56333 ^ n53213;
  assign n56385 = n53219 ^ n53217;
  assign y0 = n56123;
  assign y1 = n56124;
  assign y2 = n56125;
  assign y3 = n56126;
  assign y4 = ~n56127;
  assign y5 = ~n56128;
  assign y6 = n56129;
  assign y7 = n56130;
  assign y8 = n56131;
  assign y9 = ~n56132;
  assign y10 = ~n56133;
  assign y11 = ~n56134;
  assign y12 = n56135;
  assign y13 = ~n56136;
  assign y14 = n56137;
  assign y15 = n56138;
  assign y16 = ~n56139;
  assign y17 = ~n56140;
  assign y18 = ~n56141;
  assign y19 = ~n56142;
  assign y20 = n56143;
  assign y21 = n56144;
  assign y22 = n56145;
  assign y23 = n56146;
  assign y24 = n56147;
  assign y25 = n56148;
  assign y26 = n56149;
  assign y27 = ~n56150;
  assign y28 = n56151;
  assign y29 = n56152;
  assign y30 = ~n56153;
  assign y31 = ~n55762;
  assign y32 = ~n56184;
  assign y33 = ~n56185;
  assign y34 = n56186;
  assign y35 = n56187;
  assign y36 = n56188;
  assign y37 = n56189;
  assign y38 = ~n56190;
  assign y39 = ~n56191;
  assign y40 = ~n56192;
  assign y41 = n56193;
  assign y42 = ~n56194;
  assign y43 = ~n56195;
  assign y44 = n56196;
  assign y45 = n56197;
  assign y46 = n56198;
  assign y47 = n56199;
  assign y48 = ~n56200;
  assign y49 = ~n56201;
  assign y50 = ~n56202;
  assign y51 = ~n56203;
  assign y52 = ~n56204;
  assign y53 = ~n56205;
  assign y54 = ~n56206;
  assign y55 = ~n56207;
  assign y56 = ~n56208;
  assign y57 = n56209;
  assign y58 = ~n56210;
  assign y59 = n56211;
  assign y60 = n56212;
  assign y61 = n56213;
  assign y62 = ~n56214;
  assign y63 = ~n54786;
  assign y64 = ~n56244;
  assign y65 = n56245;
  assign y66 = ~n56246;
  assign y67 = ~n56247;
  assign y68 = ~n56248;
  assign y69 = ~n56249;
  assign y70 = n56250;
  assign y71 = ~n56251;
  assign y72 = n56252;
  assign y73 = ~n56253;
  assign y74 = ~n56254;
  assign y75 = ~n56255;
  assign y76 = n56256;
  assign y77 = n56257;
  assign y78 = n56258;
  assign y79 = ~n56259;
  assign y80 = n56260;
  assign y81 = n56261;
  assign y82 = ~n56262;
  assign y83 = ~n56263;
  assign y84 = ~n56264;
  assign y85 = n56265;
  assign y86 = n56266;
  assign y87 = n56267;
  assign y88 = n56268;
  assign y89 = ~n56269;
  assign y90 = n56270;
  assign y91 = n56271;
  assign y92 = ~n56272;
  assign y93 = n56273;
  assign y94 = n54858;
  assign y95 = n54863;
  assign y96 = n56303;
  assign y97 = n56304;
  assign y98 = n56305;
  assign y99 = ~n56306;
  assign y100 = ~n56307;
  assign y101 = n56308;
  assign y102 = n56309;
  assign y103 = n56310;
  assign y104 = n56311;
  assign y105 = ~n56312;
  assign y106 = ~n56313;
  assign y107 = n56314;
  assign y108 = ~n56315;
  assign y109 = n56316;
  assign y110 = ~n56317;
  assign y111 = n56318;
  assign y112 = ~n56319;
  assign y113 = ~n56320;
  assign y114 = ~n56321;
  assign y115 = ~n56322;
  assign y116 = n56323;
  assign y117 = ~n56324;
  assign y118 = ~n56325;
  assign y119 = n56326;
  assign y120 = ~n56327;
  assign y121 = ~n56328;
  assign y122 = ~n56329;
  assign y123 = ~n56330;
  assign y124 = ~n56331;
  assign y125 = n56332;
  assign y126 = ~n53847;
  assign y127 = n53852;
  assign y128 = n56359;
  assign y129 = n56360;
  assign y130 = ~n56361;
  assign y131 = n56362;
  assign y132 = ~n56363;
  assign y133 = ~n56364;
  assign y134 = ~n56365;
  assign y135 = n56366;
  assign y136 = ~n56367;
  assign y137 = ~n56368;
  assign y138 = n56369;
  assign y139 = n56370;
  assign y140 = n56371;
  assign y141 = ~n56372;
  assign y142 = ~n56373;
  assign y143 = ~n56374;
  assign y144 = ~n56375;
  assign y145 = ~n56376;
  assign y146 = n56377;
  assign y147 = ~n56378;
  assign y148 = n56379;
  assign y149 = n56380;
  assign y150 = n56381;
  assign y151 = n56382;
  assign y152 = n56383;
  assign y153 = n56384;
  assign y154 = n56385;
  assign y155 = n53219;
  assign y156 = n53223;
  assign y157 = ~n53227;
  assign y158 = n53232;
  assign y159 = ~n53237;
endmodule
