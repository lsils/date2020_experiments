module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 ;
  assign n130 = ~x31 & ~x63 ;
  assign n129 = ~x95 & ~x127 ;
  assign n131 = n130 ^ n129 ;
  assign n274 = x62 ^ x30 ;
  assign n275 = x63 ^ x31 ;
  assign n277 = x60 ^ x28 ;
  assign n279 = x58 ^ x26 ;
  assign n281 = x56 ^ x24 ;
  assign n283 = x54 ^ x22 ;
  assign n285 = x52 ^ x20 ;
  assign n287 = x50 ^ x18 ;
  assign n289 = x48 ^ x16 ;
  assign n291 = x46 ^ x14 ;
  assign n293 = x44 ^ x12 ;
  assign n295 = x42 ^ x10 ;
  assign n297 = x40 ^ x8 ;
  assign n299 = x38 ^ x6 ;
  assign n301 = x36 ^ x4 ;
  assign n303 = x34 ^ x2 ;
  assign n305 = x0 & ~x32 ;
  assign n306 = n305 ^ x34 ;
  assign n304 = x34 ^ x1 ;
  assign n307 = n306 ^ n304 ;
  assign n308 = x33 ^ x1 ;
  assign n309 = n307 & ~n308 ;
  assign n310 = n309 ^ n304 ;
  assign n311 = ~n303 & n310 ;
  assign n312 = n311 ^ x2 ;
  assign n313 = n312 ^ x36 ;
  assign n302 = x36 ^ x3 ;
  assign n314 = n313 ^ n302 ;
  assign n315 = x35 ^ x3 ;
  assign n316 = n314 & ~n315 ;
  assign n317 = n316 ^ n302 ;
  assign n318 = ~n301 & n317 ;
  assign n319 = n318 ^ x4 ;
  assign n320 = n319 ^ x38 ;
  assign n300 = x38 ^ x5 ;
  assign n321 = n320 ^ n300 ;
  assign n322 = x37 ^ x5 ;
  assign n323 = n321 & ~n322 ;
  assign n324 = n323 ^ n300 ;
  assign n325 = ~n299 & n324 ;
  assign n326 = n325 ^ x6 ;
  assign n327 = n326 ^ x40 ;
  assign n298 = x40 ^ x7 ;
  assign n328 = n327 ^ n298 ;
  assign n329 = x39 ^ x7 ;
  assign n330 = n328 & ~n329 ;
  assign n331 = n330 ^ n298 ;
  assign n332 = ~n297 & n331 ;
  assign n333 = n332 ^ x8 ;
  assign n334 = n333 ^ x42 ;
  assign n296 = x42 ^ x9 ;
  assign n335 = n334 ^ n296 ;
  assign n336 = x41 ^ x9 ;
  assign n337 = n335 & ~n336 ;
  assign n338 = n337 ^ n296 ;
  assign n339 = ~n295 & n338 ;
  assign n340 = n339 ^ x10 ;
  assign n341 = n340 ^ x44 ;
  assign n294 = x44 ^ x11 ;
  assign n342 = n341 ^ n294 ;
  assign n343 = x43 ^ x11 ;
  assign n344 = n342 & ~n343 ;
  assign n345 = n344 ^ n294 ;
  assign n346 = ~n293 & n345 ;
  assign n347 = n346 ^ x12 ;
  assign n348 = n347 ^ x46 ;
  assign n292 = x46 ^ x13 ;
  assign n349 = n348 ^ n292 ;
  assign n350 = x45 ^ x13 ;
  assign n351 = n349 & ~n350 ;
  assign n352 = n351 ^ n292 ;
  assign n353 = ~n291 & n352 ;
  assign n354 = n353 ^ x14 ;
  assign n355 = n354 ^ x48 ;
  assign n290 = x48 ^ x15 ;
  assign n356 = n355 ^ n290 ;
  assign n357 = x47 ^ x15 ;
  assign n358 = n356 & ~n357 ;
  assign n359 = n358 ^ n290 ;
  assign n360 = ~n289 & n359 ;
  assign n361 = n360 ^ x16 ;
  assign n362 = n361 ^ x50 ;
  assign n288 = x50 ^ x17 ;
  assign n363 = n362 ^ n288 ;
  assign n364 = x49 ^ x17 ;
  assign n365 = n363 & ~n364 ;
  assign n366 = n365 ^ n288 ;
  assign n367 = ~n287 & n366 ;
  assign n368 = n367 ^ x18 ;
  assign n369 = n368 ^ x52 ;
  assign n286 = x52 ^ x19 ;
  assign n370 = n369 ^ n286 ;
  assign n371 = x51 ^ x19 ;
  assign n372 = n370 & ~n371 ;
  assign n373 = n372 ^ n286 ;
  assign n374 = ~n285 & n373 ;
  assign n375 = n374 ^ x20 ;
  assign n376 = n375 ^ x54 ;
  assign n284 = x54 ^ x21 ;
  assign n377 = n376 ^ n284 ;
  assign n378 = x53 ^ x21 ;
  assign n379 = n377 & ~n378 ;
  assign n380 = n379 ^ n284 ;
  assign n381 = ~n283 & n380 ;
  assign n382 = n381 ^ x22 ;
  assign n383 = n382 ^ x56 ;
  assign n282 = x56 ^ x23 ;
  assign n384 = n383 ^ n282 ;
  assign n385 = x55 ^ x23 ;
  assign n386 = n384 & ~n385 ;
  assign n387 = n386 ^ n282 ;
  assign n388 = ~n281 & n387 ;
  assign n389 = n388 ^ x24 ;
  assign n390 = n389 ^ x58 ;
  assign n280 = x58 ^ x25 ;
  assign n391 = n390 ^ n280 ;
  assign n392 = x57 ^ x25 ;
  assign n393 = n391 & ~n392 ;
  assign n394 = n393 ^ n280 ;
  assign n395 = ~n279 & n394 ;
  assign n396 = n395 ^ x26 ;
  assign n397 = n396 ^ x60 ;
  assign n278 = x60 ^ x27 ;
  assign n398 = n397 ^ n278 ;
  assign n399 = x59 ^ x27 ;
  assign n400 = n398 & ~n399 ;
  assign n401 = n400 ^ n278 ;
  assign n402 = ~n277 & n401 ;
  assign n403 = n402 ^ x28 ;
  assign n404 = n403 ^ x62 ;
  assign n276 = x62 ^ x29 ;
  assign n405 = n404 ^ n276 ;
  assign n406 = x61 ^ x29 ;
  assign n407 = n405 & ~n406 ;
  assign n408 = n407 ^ n276 ;
  assign n409 = ~n274 & n408 ;
  assign n410 = n409 ^ x30 ;
  assign n411 = n410 ^ x63 ;
  assign n412 = ~n275 & n411 ;
  assign n413 = n412 ^ x31 ;
  assign n414 = n274 & ~n413 ;
  assign n415 = n414 ^ x30 ;
  assign n132 = x126 ^ x94 ;
  assign n133 = x127 ^ x95 ;
  assign n135 = x124 ^ x92 ;
  assign n137 = x122 ^ x90 ;
  assign n139 = x120 ^ x88 ;
  assign n141 = x118 ^ x86 ;
  assign n143 = x116 ^ x84 ;
  assign n145 = x114 ^ x82 ;
  assign n147 = x112 ^ x80 ;
  assign n149 = x110 ^ x78 ;
  assign n151 = x108 ^ x76 ;
  assign n153 = x106 ^ x74 ;
  assign n155 = x104 ^ x72 ;
  assign n157 = x102 ^ x70 ;
  assign n159 = x100 ^ x68 ;
  assign n161 = x98 ^ x66 ;
  assign n163 = x64 & ~x96 ;
  assign n164 = n163 ^ x98 ;
  assign n162 = x98 ^ x65 ;
  assign n165 = n164 ^ n162 ;
  assign n166 = x97 ^ x65 ;
  assign n167 = n165 & ~n166 ;
  assign n168 = n167 ^ n162 ;
  assign n169 = ~n161 & n168 ;
  assign n170 = n169 ^ x66 ;
  assign n171 = n170 ^ x100 ;
  assign n160 = x100 ^ x67 ;
  assign n172 = n171 ^ n160 ;
  assign n173 = x99 ^ x67 ;
  assign n174 = n172 & ~n173 ;
  assign n175 = n174 ^ n160 ;
  assign n176 = ~n159 & n175 ;
  assign n177 = n176 ^ x68 ;
  assign n178 = n177 ^ x102 ;
  assign n158 = x102 ^ x69 ;
  assign n179 = n178 ^ n158 ;
  assign n180 = x101 ^ x69 ;
  assign n181 = n179 & ~n180 ;
  assign n182 = n181 ^ n158 ;
  assign n183 = ~n157 & n182 ;
  assign n184 = n183 ^ x70 ;
  assign n185 = n184 ^ x104 ;
  assign n156 = x104 ^ x71 ;
  assign n186 = n185 ^ n156 ;
  assign n187 = x103 ^ x71 ;
  assign n188 = n186 & ~n187 ;
  assign n189 = n188 ^ n156 ;
  assign n190 = ~n155 & n189 ;
  assign n191 = n190 ^ x72 ;
  assign n192 = n191 ^ x106 ;
  assign n154 = x106 ^ x73 ;
  assign n193 = n192 ^ n154 ;
  assign n194 = x105 ^ x73 ;
  assign n195 = n193 & ~n194 ;
  assign n196 = n195 ^ n154 ;
  assign n197 = ~n153 & n196 ;
  assign n198 = n197 ^ x74 ;
  assign n199 = n198 ^ x108 ;
  assign n152 = x108 ^ x75 ;
  assign n200 = n199 ^ n152 ;
  assign n201 = x107 ^ x75 ;
  assign n202 = n200 & ~n201 ;
  assign n203 = n202 ^ n152 ;
  assign n204 = ~n151 & n203 ;
  assign n205 = n204 ^ x76 ;
  assign n206 = n205 ^ x110 ;
  assign n150 = x110 ^ x77 ;
  assign n207 = n206 ^ n150 ;
  assign n208 = x109 ^ x77 ;
  assign n209 = n207 & ~n208 ;
  assign n210 = n209 ^ n150 ;
  assign n211 = ~n149 & n210 ;
  assign n212 = n211 ^ x78 ;
  assign n213 = n212 ^ x112 ;
  assign n148 = x112 ^ x79 ;
  assign n214 = n213 ^ n148 ;
  assign n215 = x111 ^ x79 ;
  assign n216 = n214 & ~n215 ;
  assign n217 = n216 ^ n148 ;
  assign n218 = ~n147 & n217 ;
  assign n219 = n218 ^ x80 ;
  assign n220 = n219 ^ x114 ;
  assign n146 = x114 ^ x81 ;
  assign n221 = n220 ^ n146 ;
  assign n222 = x113 ^ x81 ;
  assign n223 = n221 & ~n222 ;
  assign n224 = n223 ^ n146 ;
  assign n225 = ~n145 & n224 ;
  assign n226 = n225 ^ x82 ;
  assign n227 = n226 ^ x116 ;
  assign n144 = x116 ^ x83 ;
  assign n228 = n227 ^ n144 ;
  assign n229 = x115 ^ x83 ;
  assign n230 = n228 & ~n229 ;
  assign n231 = n230 ^ n144 ;
  assign n232 = ~n143 & n231 ;
  assign n233 = n232 ^ x84 ;
  assign n234 = n233 ^ x118 ;
  assign n142 = x118 ^ x85 ;
  assign n235 = n234 ^ n142 ;
  assign n236 = x117 ^ x85 ;
  assign n237 = n235 & ~n236 ;
  assign n238 = n237 ^ n142 ;
  assign n239 = ~n141 & n238 ;
  assign n240 = n239 ^ x86 ;
  assign n241 = n240 ^ x120 ;
  assign n140 = x120 ^ x87 ;
  assign n242 = n241 ^ n140 ;
  assign n243 = x119 ^ x87 ;
  assign n244 = n242 & ~n243 ;
  assign n245 = n244 ^ n140 ;
  assign n246 = ~n139 & n245 ;
  assign n247 = n246 ^ x88 ;
  assign n248 = n247 ^ x122 ;
  assign n138 = x122 ^ x89 ;
  assign n249 = n248 ^ n138 ;
  assign n250 = x121 ^ x89 ;
  assign n251 = n249 & ~n250 ;
  assign n252 = n251 ^ n138 ;
  assign n253 = ~n137 & n252 ;
  assign n254 = n253 ^ x90 ;
  assign n255 = n254 ^ x124 ;
  assign n136 = x124 ^ x91 ;
  assign n256 = n255 ^ n136 ;
  assign n257 = x123 ^ x91 ;
  assign n258 = n256 & ~n257 ;
  assign n259 = n258 ^ n136 ;
  assign n260 = ~n135 & n259 ;
  assign n261 = n260 ^ x92 ;
  assign n262 = n261 ^ x126 ;
  assign n134 = x126 ^ x93 ;
  assign n263 = n262 ^ n134 ;
  assign n264 = x125 ^ x93 ;
  assign n265 = n263 & ~n264 ;
  assign n266 = n265 ^ n134 ;
  assign n267 = ~n132 & n266 ;
  assign n268 = n267 ^ x94 ;
  assign n269 = n268 ^ x127 ;
  assign n270 = ~n133 & n269 ;
  assign n271 = n270 ^ x95 ;
  assign n272 = n132 & ~n271 ;
  assign n273 = n272 ^ x94 ;
  assign n416 = n415 ^ n273 ;
  assign n419 = n264 & ~n271 ;
  assign n420 = n419 ^ x93 ;
  assign n417 = n406 & ~n413 ;
  assign n418 = n417 ^ x29 ;
  assign n421 = n420 ^ n418 ;
  assign n424 = n135 & ~n271 ;
  assign n425 = n424 ^ x92 ;
  assign n422 = n277 & ~n413 ;
  assign n423 = n422 ^ x28 ;
  assign n426 = n425 ^ n423 ;
  assign n429 = n399 & ~n413 ;
  assign n430 = n429 ^ x27 ;
  assign n427 = n257 & ~n271 ;
  assign n428 = n427 ^ x91 ;
  assign n431 = n430 ^ n428 ;
  assign n434 = n137 & ~n271 ;
  assign n435 = n434 ^ x90 ;
  assign n432 = n279 & ~n413 ;
  assign n433 = n432 ^ x26 ;
  assign n436 = n435 ^ n433 ;
  assign n439 = n392 & ~n413 ;
  assign n440 = n439 ^ x25 ;
  assign n437 = n250 & ~n271 ;
  assign n438 = n437 ^ x89 ;
  assign n441 = n440 ^ n438 ;
  assign n444 = n139 & ~n271 ;
  assign n445 = n444 ^ x88 ;
  assign n442 = n281 & ~n413 ;
  assign n443 = n442 ^ x24 ;
  assign n446 = n445 ^ n443 ;
  assign n449 = n385 & ~n413 ;
  assign n450 = n449 ^ x23 ;
  assign n447 = n243 & ~n271 ;
  assign n448 = n447 ^ x87 ;
  assign n451 = n450 ^ n448 ;
  assign n454 = n141 & ~n271 ;
  assign n455 = n454 ^ x86 ;
  assign n452 = n283 & ~n413 ;
  assign n453 = n452 ^ x22 ;
  assign n456 = n455 ^ n453 ;
  assign n459 = n378 & ~n413 ;
  assign n460 = n459 ^ x21 ;
  assign n457 = n236 & ~n271 ;
  assign n458 = n457 ^ x85 ;
  assign n461 = n460 ^ n458 ;
  assign n464 = n143 & ~n271 ;
  assign n465 = n464 ^ x84 ;
  assign n462 = n285 & ~n413 ;
  assign n463 = n462 ^ x20 ;
  assign n466 = n465 ^ n463 ;
  assign n469 = n371 & ~n413 ;
  assign n470 = n469 ^ x19 ;
  assign n467 = n229 & ~n271 ;
  assign n468 = n467 ^ x83 ;
  assign n471 = n470 ^ n468 ;
  assign n474 = n145 & ~n271 ;
  assign n475 = n474 ^ x82 ;
  assign n472 = n287 & ~n413 ;
  assign n473 = n472 ^ x18 ;
  assign n476 = n475 ^ n473 ;
  assign n479 = n364 & ~n413 ;
  assign n480 = n479 ^ x17 ;
  assign n477 = n222 & ~n271 ;
  assign n478 = n477 ^ x81 ;
  assign n481 = n480 ^ n478 ;
  assign n484 = n147 & ~n271 ;
  assign n485 = n484 ^ x80 ;
  assign n482 = n289 & ~n413 ;
  assign n483 = n482 ^ x16 ;
  assign n486 = n485 ^ n483 ;
  assign n489 = n357 & ~n413 ;
  assign n490 = n489 ^ x15 ;
  assign n487 = n215 & ~n271 ;
  assign n488 = n487 ^ x79 ;
  assign n491 = n490 ^ n488 ;
  assign n494 = n149 & ~n271 ;
  assign n495 = n494 ^ x78 ;
  assign n492 = n291 & ~n413 ;
  assign n493 = n492 ^ x14 ;
  assign n496 = n495 ^ n493 ;
  assign n499 = n350 & ~n413 ;
  assign n500 = n499 ^ x13 ;
  assign n497 = n208 & ~n271 ;
  assign n498 = n497 ^ x77 ;
  assign n501 = n500 ^ n498 ;
  assign n504 = n151 & ~n271 ;
  assign n505 = n504 ^ x76 ;
  assign n502 = n293 & ~n413 ;
  assign n503 = n502 ^ x12 ;
  assign n506 = n505 ^ n503 ;
  assign n509 = n343 & ~n413 ;
  assign n510 = n509 ^ x11 ;
  assign n507 = n201 & ~n271 ;
  assign n508 = n507 ^ x75 ;
  assign n511 = n510 ^ n508 ;
  assign n514 = n153 & ~n271 ;
  assign n515 = n514 ^ x74 ;
  assign n512 = n295 & ~n413 ;
  assign n513 = n512 ^ x10 ;
  assign n516 = n515 ^ n513 ;
  assign n519 = n336 & ~n413 ;
  assign n520 = n519 ^ x9 ;
  assign n517 = n194 & ~n271 ;
  assign n518 = n517 ^ x73 ;
  assign n521 = n520 ^ n518 ;
  assign n524 = n155 & ~n271 ;
  assign n525 = n524 ^ x72 ;
  assign n522 = n297 & ~n413 ;
  assign n523 = n522 ^ x8 ;
  assign n526 = n525 ^ n523 ;
  assign n529 = n329 & ~n413 ;
  assign n530 = n529 ^ x7 ;
  assign n527 = n187 & ~n271 ;
  assign n528 = n527 ^ x71 ;
  assign n531 = n530 ^ n528 ;
  assign n534 = n299 & ~n413 ;
  assign n535 = n534 ^ x6 ;
  assign n532 = n157 & ~n271 ;
  assign n533 = n532 ^ x70 ;
  assign n536 = n535 ^ n533 ;
  assign n539 = n322 & ~n413 ;
  assign n540 = n539 ^ x5 ;
  assign n537 = n180 & ~n271 ;
  assign n538 = n537 ^ x69 ;
  assign n541 = n540 ^ n538 ;
  assign n544 = n159 & ~n271 ;
  assign n545 = n544 ^ x68 ;
  assign n542 = n301 & ~n413 ;
  assign n543 = n542 ^ x4 ;
  assign n546 = n545 ^ n543 ;
  assign n549 = n173 & ~n271 ;
  assign n550 = n549 ^ x67 ;
  assign n547 = n315 & ~n413 ;
  assign n548 = n547 ^ x3 ;
  assign n551 = n550 ^ n548 ;
  assign n554 = n303 & ~n413 ;
  assign n555 = n554 ^ x2 ;
  assign n552 = n161 & ~n271 ;
  assign n553 = n552 ^ x66 ;
  assign n556 = n555 ^ n553 ;
  assign n559 = n308 & ~n413 ;
  assign n560 = n559 ^ x1 ;
  assign n557 = n166 & ~n271 ;
  assign n558 = n557 ^ x65 ;
  assign n561 = n560 ^ n558 ;
  assign n562 = x96 ^ x64 ;
  assign n563 = ~n271 & n562 ;
  assign n564 = n563 ^ x64 ;
  assign n565 = x32 ^ x0 ;
  assign n566 = ~n413 & n565 ;
  assign n567 = n566 ^ x0 ;
  assign n568 = ~n564 & n567 ;
  assign n569 = n568 ^ n560 ;
  assign n570 = ~n561 & n569 ;
  assign n571 = n570 ^ n560 ;
  assign n572 = n571 ^ n555 ;
  assign n573 = ~n556 & n572 ;
  assign n574 = n573 ^ n555 ;
  assign n575 = n574 ^ n550 ;
  assign n576 = ~n551 & ~n575 ;
  assign n577 = n576 ^ n550 ;
  assign n578 = n577 ^ n543 ;
  assign n579 = ~n546 & ~n578 ;
  assign n580 = n579 ^ n543 ;
  assign n581 = n580 ^ n540 ;
  assign n582 = ~n541 & n581 ;
  assign n583 = n582 ^ n540 ;
  assign n584 = n583 ^ n533 ;
  assign n585 = ~n536 & ~n584 ;
  assign n586 = n585 ^ n533 ;
  assign n587 = n586 ^ n530 ;
  assign n588 = ~n531 & ~n587 ;
  assign n589 = n588 ^ n530 ;
  assign n590 = n589 ^ n523 ;
  assign n591 = ~n526 & n590 ;
  assign n592 = n591 ^ n523 ;
  assign n593 = n592 ^ n520 ;
  assign n594 = ~n521 & n593 ;
  assign n595 = n594 ^ n520 ;
  assign n596 = n595 ^ n513 ;
  assign n597 = ~n516 & n596 ;
  assign n598 = n597 ^ n513 ;
  assign n599 = n598 ^ n510 ;
  assign n600 = ~n511 & n599 ;
  assign n601 = n600 ^ n510 ;
  assign n602 = n601 ^ n503 ;
  assign n603 = ~n506 & n602 ;
  assign n604 = n603 ^ n503 ;
  assign n605 = n604 ^ n500 ;
  assign n606 = ~n501 & n605 ;
  assign n607 = n606 ^ n500 ;
  assign n608 = n607 ^ n493 ;
  assign n609 = ~n496 & n608 ;
  assign n610 = n609 ^ n493 ;
  assign n611 = n610 ^ n490 ;
  assign n612 = ~n491 & n611 ;
  assign n613 = n612 ^ n490 ;
  assign n614 = n613 ^ n483 ;
  assign n615 = ~n486 & n614 ;
  assign n616 = n615 ^ n483 ;
  assign n617 = n616 ^ n480 ;
  assign n618 = ~n481 & n617 ;
  assign n619 = n618 ^ n480 ;
  assign n620 = n619 ^ n473 ;
  assign n621 = ~n476 & n620 ;
  assign n622 = n621 ^ n473 ;
  assign n623 = n622 ^ n470 ;
  assign n624 = ~n471 & n623 ;
  assign n625 = n624 ^ n470 ;
  assign n626 = n625 ^ n463 ;
  assign n627 = ~n466 & n626 ;
  assign n628 = n627 ^ n463 ;
  assign n629 = n628 ^ n460 ;
  assign n630 = ~n461 & n629 ;
  assign n631 = n630 ^ n460 ;
  assign n632 = n631 ^ n453 ;
  assign n633 = ~n456 & n632 ;
  assign n634 = n633 ^ n453 ;
  assign n635 = n634 ^ n450 ;
  assign n636 = ~n451 & n635 ;
  assign n637 = n636 ^ n450 ;
  assign n638 = n637 ^ n443 ;
  assign n639 = ~n446 & n638 ;
  assign n640 = n639 ^ n443 ;
  assign n641 = n640 ^ n440 ;
  assign n642 = ~n441 & n641 ;
  assign n643 = n642 ^ n440 ;
  assign n644 = n643 ^ n433 ;
  assign n645 = ~n436 & n644 ;
  assign n646 = n645 ^ n433 ;
  assign n647 = n646 ^ n430 ;
  assign n648 = ~n431 & n647 ;
  assign n649 = n648 ^ n430 ;
  assign n650 = n649 ^ n425 ;
  assign n651 = ~n426 & ~n650 ;
  assign n652 = n651 ^ n425 ;
  assign n653 = n652 ^ n420 ;
  assign n654 = ~n421 & ~n653 ;
  assign n655 = n654 ^ n418 ;
  assign n656 = n655 ^ n415 ;
  assign n657 = ~n416 & ~n656 ;
  assign n658 = n657 ^ n273 ;
  assign n659 = n658 ^ n130 ;
  assign n660 = ~n131 & ~n659 ;
  assign n661 = n660 ^ n129 ;
  assign n662 = n413 ^ n271 ;
  assign n663 = n661 & n662 ;
  assign n664 = n663 ^ n271 ;
  assign n665 = n567 ^ n564 ;
  assign n666 = n661 & n665 ;
  assign n667 = n666 ^ n564 ;
  assign n668 = n561 & n661 ;
  assign n669 = n668 ^ n558 ;
  assign n670 = n556 & n661 ;
  assign n671 = n670 ^ n553 ;
  assign n672 = n551 & n661 ;
  assign n673 = n672 ^ n550 ;
  assign n674 = n546 & n661 ;
  assign n675 = n674 ^ n545 ;
  assign n676 = n541 & n661 ;
  assign n677 = n676 ^ n538 ;
  assign n678 = n536 & n661 ;
  assign n679 = n678 ^ n533 ;
  assign n680 = n531 & ~n661 ;
  assign n681 = n680 ^ n530 ;
  assign n682 = n526 & n661 ;
  assign n683 = n682 ^ n525 ;
  assign n684 = n521 & n661 ;
  assign n685 = n684 ^ n518 ;
  assign n686 = n516 & ~n661 ;
  assign n687 = n686 ^ n513 ;
  assign n688 = n511 & ~n661 ;
  assign n689 = n688 ^ n510 ;
  assign n690 = n506 & n661 ;
  assign n691 = n690 ^ n505 ;
  assign n692 = n501 & n661 ;
  assign n693 = n692 ^ n498 ;
  assign n694 = n496 & ~n661 ;
  assign n695 = n694 ^ n493 ;
  assign n696 = n491 & ~n661 ;
  assign n697 = n696 ^ n490 ;
  assign n698 = n486 & n661 ;
  assign n699 = n698 ^ n485 ;
  assign n700 = n481 & n661 ;
  assign n701 = n700 ^ n478 ;
  assign n702 = n476 & ~n661 ;
  assign n703 = n702 ^ n473 ;
  assign n704 = n471 & ~n661 ;
  assign n705 = n704 ^ n470 ;
  assign n706 = n466 & n661 ;
  assign n707 = n706 ^ n465 ;
  assign n708 = n461 & n661 ;
  assign n709 = n708 ^ n458 ;
  assign n710 = n456 & ~n661 ;
  assign n711 = n710 ^ n453 ;
  assign n712 = n451 & ~n661 ;
  assign n713 = n712 ^ n450 ;
  assign n714 = n446 & n661 ;
  assign n715 = n714 ^ n445 ;
  assign n716 = n441 & n661 ;
  assign n717 = n716 ^ n438 ;
  assign n718 = n436 & ~n661 ;
  assign n719 = n718 ^ n433 ;
  assign n720 = n431 & ~n661 ;
  assign n721 = n720 ^ n430 ;
  assign n722 = n426 & n661 ;
  assign n723 = n722 ^ n425 ;
  assign n724 = n421 & n661 ;
  assign n725 = n724 ^ n420 ;
  assign n726 = n416 & n661 ;
  assign n727 = n726 ^ n273 ;
  assign n728 = n129 & n130 ;
  assign y0 = ~n664 ;
  assign y1 = ~n661 ;
  assign y2 = n667 ;
  assign y3 = n669 ;
  assign y4 = n671 ;
  assign y5 = n673 ;
  assign y6 = n675 ;
  assign y7 = n677 ;
  assign y8 = n679 ;
  assign y9 = n681 ;
  assign y10 = n683 ;
  assign y11 = n685 ;
  assign y12 = n687 ;
  assign y13 = n689 ;
  assign y14 = n691 ;
  assign y15 = n693 ;
  assign y16 = n695 ;
  assign y17 = n697 ;
  assign y18 = n699 ;
  assign y19 = n701 ;
  assign y20 = n703 ;
  assign y21 = n705 ;
  assign y22 = n707 ;
  assign y23 = n709 ;
  assign y24 = n711 ;
  assign y25 = n713 ;
  assign y26 = n715 ;
  assign y27 = n717 ;
  assign y28 = n719 ;
  assign y29 = n721 ;
  assign y30 = n723 ;
  assign y31 = n725 ;
  assign y32 = n727 ;
  assign y33 = ~n728 ;
endmodule
