module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613;
  assign n129 = ~x126 & ~x127;
  assign n130 = x127 ^ x125;
  assign n131 = ~x122 & ~x123;
  assign n132 = x123 ^ x121;
  assign n133 = ~x118 & ~x119;
  assign n134 = x119 ^ x117;
  assign n135 = ~x114 & ~x115;
  assign n136 = x115 ^ x113;
  assign n137 = ~x110 & ~x111;
  assign n138 = x111 ^ x109;
  assign n139 = ~x106 & ~x107;
  assign n140 = x107 ^ x105;
  assign n141 = ~x102 & ~x103;
  assign n142 = x103 ^ x101;
  assign n143 = ~x98 & ~x99;
  assign n144 = x99 ^ x97;
  assign n145 = ~x94 & ~x95;
  assign n146 = x95 ^ x93;
  assign n147 = ~x90 & ~x91;
  assign n148 = x91 ^ x89;
  assign n149 = ~x86 & ~x87;
  assign n150 = x87 ^ x85;
  assign n151 = ~x82 & ~x83;
  assign n152 = x83 ^ x81;
  assign n153 = ~x78 & ~x79;
  assign n154 = x79 ^ x77;
  assign n155 = ~x74 & ~x75;
  assign n156 = x75 ^ x73;
  assign n157 = ~x70 & ~x71;
  assign n158 = x71 ^ x69;
  assign n159 = ~x66 & ~x67;
  assign n160 = x67 ^ x65;
  assign n161 = ~x62 & ~x63;
  assign n162 = x63 ^ x61;
  assign n163 = ~x58 & ~x59;
  assign n164 = x59 ^ x57;
  assign n165 = ~x54 & ~x55;
  assign n166 = x55 ^ x53;
  assign n167 = ~x50 & ~x51;
  assign n168 = x51 ^ x49;
  assign n169 = ~x46 & ~x47;
  assign n170 = x47 ^ x45;
  assign n171 = ~x42 & ~x43;
  assign n172 = x43 ^ x41;
  assign n173 = ~x38 & ~x39;
  assign n174 = x39 ^ x37;
  assign n175 = ~x34 & ~x35;
  assign n176 = x35 ^ x33;
  assign n177 = ~x30 & ~x31;
  assign n178 = x31 ^ x29;
  assign n179 = ~x26 & ~x27;
  assign n180 = x27 ^ x25;
  assign n181 = ~x22 & ~x23;
  assign n182 = x23 ^ x21;
  assign n183 = ~x18 & ~x19;
  assign n184 = x19 ^ x17;
  assign n185 = ~x14 & ~x15;
  assign n186 = x15 ^ x13;
  assign n187 = ~x10 & ~x11;
  assign n188 = x11 ^ x9;
  assign n189 = ~x6 & ~x7;
  assign n190 = x7 ^ x5;
  assign n191 = ~x2 & ~x3;
  assign n192 = x1 & n191;
  assign n193 = n192 ^ x3;
  assign n194 = ~x4 & n193;
  assign n195 = n194 ^ n189;
  assign n196 = n190 & n195;
  assign n197 = n196 ^ n194;
  assign n198 = n189 & n197;
  assign n199 = n198 ^ x7;
  assign n200 = ~x8 & n199;
  assign n201 = n200 ^ n187;
  assign n202 = n188 & n201;
  assign n203 = n202 ^ n200;
  assign n204 = n187 & n203;
  assign n205 = n204 ^ x11;
  assign n206 = ~x12 & n205;
  assign n207 = n206 ^ n185;
  assign n208 = n186 & n207;
  assign n209 = n208 ^ n206;
  assign n210 = n185 & n209;
  assign n211 = n210 ^ x15;
  assign n212 = ~x16 & n211;
  assign n213 = n212 ^ n183;
  assign n214 = n184 & n213;
  assign n215 = n214 ^ n212;
  assign n216 = n183 & n215;
  assign n217 = n216 ^ x19;
  assign n218 = ~x20 & n217;
  assign n219 = n218 ^ n181;
  assign n220 = n182 & n219;
  assign n221 = n220 ^ n218;
  assign n222 = n181 & n221;
  assign n223 = n222 ^ x23;
  assign n224 = ~x24 & n223;
  assign n225 = n224 ^ n179;
  assign n226 = n180 & n225;
  assign n227 = n226 ^ n224;
  assign n228 = n179 & n227;
  assign n229 = n228 ^ x27;
  assign n230 = ~x28 & n229;
  assign n231 = n230 ^ n177;
  assign n232 = n178 & n231;
  assign n233 = n232 ^ n230;
  assign n234 = n177 & n233;
  assign n235 = n234 ^ x31;
  assign n236 = ~x32 & n235;
  assign n237 = n236 ^ n175;
  assign n238 = n176 & n237;
  assign n239 = n238 ^ n236;
  assign n240 = n175 & n239;
  assign n241 = n240 ^ x35;
  assign n242 = ~x36 & n241;
  assign n243 = n242 ^ n173;
  assign n244 = n174 & n243;
  assign n245 = n244 ^ n242;
  assign n246 = n173 & n245;
  assign n247 = n246 ^ x39;
  assign n248 = ~x40 & n247;
  assign n249 = n248 ^ n171;
  assign n250 = n172 & n249;
  assign n251 = n250 ^ n248;
  assign n252 = n171 & n251;
  assign n253 = n252 ^ x43;
  assign n254 = ~x44 & n253;
  assign n255 = n254 ^ n169;
  assign n256 = n170 & n255;
  assign n257 = n256 ^ n254;
  assign n258 = n169 & n257;
  assign n259 = n258 ^ x47;
  assign n260 = ~x48 & n259;
  assign n261 = n260 ^ n167;
  assign n262 = n168 & n261;
  assign n263 = n262 ^ n260;
  assign n264 = n167 & n263;
  assign n265 = n264 ^ x51;
  assign n266 = ~x52 & n265;
  assign n267 = n266 ^ n165;
  assign n268 = n166 & n267;
  assign n269 = n268 ^ n266;
  assign n270 = n165 & n269;
  assign n271 = n270 ^ x55;
  assign n272 = ~x56 & n271;
  assign n273 = n272 ^ n163;
  assign n274 = n164 & n273;
  assign n275 = n274 ^ n272;
  assign n276 = n163 & n275;
  assign n277 = n276 ^ x59;
  assign n278 = ~x60 & n277;
  assign n279 = n278 ^ n161;
  assign n280 = n162 & n279;
  assign n281 = n280 ^ n278;
  assign n282 = n161 & n281;
  assign n283 = n282 ^ x63;
  assign n284 = ~x64 & n283;
  assign n285 = n284 ^ n159;
  assign n286 = n160 & n285;
  assign n287 = n286 ^ n284;
  assign n288 = n159 & n287;
  assign n289 = n288 ^ x67;
  assign n290 = ~x68 & n289;
  assign n291 = n290 ^ n157;
  assign n292 = n158 & n291;
  assign n293 = n292 ^ n290;
  assign n294 = n157 & n293;
  assign n295 = n294 ^ x71;
  assign n296 = ~x72 & n295;
  assign n297 = n296 ^ n155;
  assign n298 = n156 & n297;
  assign n299 = n298 ^ n296;
  assign n300 = n155 & n299;
  assign n301 = n300 ^ x75;
  assign n302 = ~x76 & n301;
  assign n303 = n302 ^ n153;
  assign n304 = n154 & n303;
  assign n305 = n304 ^ n302;
  assign n306 = n153 & n305;
  assign n307 = n306 ^ x79;
  assign n308 = ~x80 & n307;
  assign n309 = n308 ^ n151;
  assign n310 = n152 & n309;
  assign n311 = n310 ^ n308;
  assign n312 = n151 & n311;
  assign n313 = n312 ^ x83;
  assign n314 = ~x84 & n313;
  assign n315 = n314 ^ n149;
  assign n316 = n150 & n315;
  assign n317 = n316 ^ n314;
  assign n318 = n149 & n317;
  assign n319 = n318 ^ x87;
  assign n320 = ~x88 & n319;
  assign n321 = n320 ^ n147;
  assign n322 = n148 & n321;
  assign n323 = n322 ^ n320;
  assign n324 = n147 & n323;
  assign n325 = n324 ^ x91;
  assign n326 = ~x92 & n325;
  assign n327 = n326 ^ n145;
  assign n328 = n146 & n327;
  assign n329 = n328 ^ n326;
  assign n330 = n145 & n329;
  assign n331 = n330 ^ x95;
  assign n332 = ~x96 & n331;
  assign n333 = n332 ^ n143;
  assign n334 = n144 & n333;
  assign n335 = n334 ^ n332;
  assign n336 = n143 & n335;
  assign n337 = n336 ^ x99;
  assign n338 = ~x100 & n337;
  assign n339 = n338 ^ n141;
  assign n340 = n142 & n339;
  assign n341 = n340 ^ n338;
  assign n342 = n141 & n341;
  assign n343 = n342 ^ x103;
  assign n344 = ~x104 & n343;
  assign n345 = n344 ^ n139;
  assign n346 = n140 & n345;
  assign n347 = n346 ^ n344;
  assign n348 = n139 & n347;
  assign n349 = n348 ^ x107;
  assign n350 = ~x108 & n349;
  assign n351 = n350 ^ n137;
  assign n352 = n138 & n351;
  assign n353 = n352 ^ n350;
  assign n354 = n137 & n353;
  assign n355 = n354 ^ x111;
  assign n356 = ~x112 & n355;
  assign n357 = n356 ^ n135;
  assign n358 = n136 & n357;
  assign n359 = n358 ^ n356;
  assign n360 = n135 & n359;
  assign n361 = n360 ^ x115;
  assign n362 = ~x116 & n361;
  assign n363 = n362 ^ n133;
  assign n364 = n134 & n363;
  assign n365 = n364 ^ n362;
  assign n366 = n133 & n365;
  assign n367 = n366 ^ x119;
  assign n368 = ~x120 & n367;
  assign n369 = n368 ^ n131;
  assign n370 = n132 & n369;
  assign n371 = n370 ^ n368;
  assign n372 = n131 & n371;
  assign n373 = n372 ^ x123;
  assign n374 = ~x124 & n373;
  assign n375 = n374 ^ n129;
  assign n376 = n130 & n375;
  assign n377 = n376 ^ n374;
  assign n378 = n129 & n377;
  assign n379 = n378 ^ x127;
  assign n380 = ~x124 & ~x125;
  assign n381 = n129 & n380;
  assign n382 = ~x120 & ~x121;
  assign n383 = ~n133 & n382;
  assign n384 = n131 & ~n383;
  assign n385 = n384 ^ n380;
  assign n386 = n131 & n382;
  assign n387 = ~x116 & ~x117;
  assign n388 = n133 & n387;
  assign n389 = n386 & n388;
  assign n390 = ~x112 & ~x113;
  assign n391 = n135 & n390;
  assign n392 = n389 & n391;
  assign n393 = n381 & n392;
  assign n394 = ~x108 & ~x109;
  assign n395 = n137 & n394;
  assign n396 = n394 ^ n139;
  assign n397 = ~x104 & ~x105;
  assign n398 = ~x100 & ~x101;
  assign n399 = n141 & n398;
  assign n400 = n398 ^ n143;
  assign n401 = ~x96 & ~x97;
  assign n402 = ~x92 & ~x93;
  assign n403 = n145 & n402;
  assign n404 = n402 ^ n147;
  assign n405 = ~x88 & ~x89;
  assign n406 = ~x84 & ~x85;
  assign n407 = n149 & n406;
  assign n408 = n147 & n405;
  assign n409 = n403 & n408;
  assign n410 = ~x80 & ~x81;
  assign n411 = n151 & n410;
  assign n412 = n409 & n411;
  assign n413 = n407 & n412;
  assign n414 = ~x76 & ~x77;
  assign n415 = n153 & n414;
  assign n416 = n414 ^ n155;
  assign n417 = ~x72 & ~x73;
  assign n418 = ~x68 & ~x69;
  assign n419 = n157 & n418;
  assign n420 = n418 ^ n159;
  assign n421 = n155 & n417;
  assign n422 = n415 & n421;
  assign n423 = ~x64 & ~x65;
  assign n424 = n159 & n423;
  assign n425 = n419 & n424;
  assign n426 = n422 & n425;
  assign n427 = ~x60 & ~x61;
  assign n428 = n161 & n427;
  assign n429 = ~x56 & ~x57;
  assign n430 = n163 & n429;
  assign n431 = n428 & n430;
  assign n432 = ~x52 & ~x53;
  assign n433 = n165 & n432;
  assign n434 = ~x48 & ~x49;
  assign n435 = n167 & n434;
  assign n436 = n433 & n435;
  assign n437 = n431 & n436;
  assign n438 = ~x44 & ~x45;
  assign n439 = n169 & n438;
  assign n440 = ~x40 & ~x41;
  assign n441 = n171 & n440;
  assign n442 = n439 & n441;
  assign n443 = ~x36 & ~x37;
  assign n444 = n173 & n443;
  assign n445 = ~x32 & ~x33;
  assign n446 = n175 & n445;
  assign n447 = n444 & n446;
  assign n448 = n442 & n447;
  assign n449 = n437 & n448;
  assign n450 = ~x16 & ~x17;
  assign n451 = n183 & n450;
  assign n452 = ~x28 & ~x29;
  assign n453 = n177 & n452;
  assign n454 = ~x24 & ~x25;
  assign n455 = n179 & n454;
  assign n456 = n453 & n455;
  assign n457 = ~x20 & ~x21;
  assign n458 = n181 & n457;
  assign n459 = n456 & n458;
  assign n460 = n451 & n459;
  assign n461 = ~x12 & ~x13;
  assign n462 = n185 & n461;
  assign n463 = n461 ^ n187;
  assign n464 = n139 & n397;
  assign n465 = n395 & n464;
  assign n466 = n143 & n401;
  assign n467 = n399 & n466;
  assign n468 = n465 & n467;
  assign n469 = n448 & ~n460;
  assign n470 = n437 & ~n469;
  assign n471 = n426 & ~n470;
  assign n472 = n413 & ~n471;
  assign n473 = n468 & ~n472;
  assign n474 = ~x8 & ~x9;
  assign n475 = n187 & n474;
  assign n476 = n462 & n475;
  assign n477 = ~n473 & ~n476;
  assign n478 = ~x4 & ~x5;
  assign n479 = ~n191 & n478;
  assign n480 = n189 & ~n479;
  assign n481 = ~n477 & ~n480;
  assign n482 = n481 ^ n462;
  assign n483 = n463 & n482;
  assign n484 = n483 ^ n481;
  assign n485 = n462 & n484;
  assign n486 = n485 ^ n185;
  assign n487 = n460 & ~n486;
  assign n488 = ~n181 & n455;
  assign n489 = n488 ^ n179;
  assign n490 = n453 & ~n489;
  assign n491 = ~n183 & n459;
  assign n492 = n491 ^ n177;
  assign n493 = ~n490 & n492;
  assign n494 = ~n487 & n493;
  assign n495 = n449 & ~n494;
  assign n496 = n175 & ~n495;
  assign n497 = n444 & ~n496;
  assign n498 = n173 & ~n497;
  assign n499 = n442 & ~n498;
  assign n500 = ~n171 & n438;
  assign n501 = n169 & ~n500;
  assign n502 = ~n499 & n501;
  assign n503 = n437 & ~n502;
  assign n504 = ~n167 & n432;
  assign n505 = n165 & ~n504;
  assign n506 = ~n503 & n505;
  assign n507 = n431 & ~n506;
  assign n508 = ~n163 & n427;
  assign n509 = n161 & ~n508;
  assign n510 = ~n507 & n509;
  assign n511 = n426 & ~n510;
  assign n512 = n511 ^ n419;
  assign n513 = n420 & n512;
  assign n514 = n513 ^ n511;
  assign n515 = n419 & n514;
  assign n516 = n515 ^ n157;
  assign n517 = n417 & ~n516;
  assign n518 = n517 ^ n415;
  assign n519 = n416 & n518;
  assign n520 = n519 ^ n517;
  assign n521 = n415 & n520;
  assign n522 = n521 ^ n153;
  assign n523 = n413 & ~n522;
  assign n524 = ~n151 & n406;
  assign n525 = n149 & ~n524;
  assign n526 = ~n523 & n525;
  assign n527 = n405 & ~n526;
  assign n528 = n527 ^ n403;
  assign n529 = n404 & n528;
  assign n530 = n529 ^ n527;
  assign n531 = n403 & n530;
  assign n532 = n531 ^ n145;
  assign n533 = n401 & ~n532;
  assign n534 = n533 ^ n399;
  assign n535 = n400 & n534;
  assign n536 = n535 ^ n533;
  assign n537 = n399 & n536;
  assign n538 = n537 ^ n141;
  assign n539 = n397 & ~n538;
  assign n540 = n539 ^ n395;
  assign n541 = n396 & n540;
  assign n542 = n541 ^ n539;
  assign n543 = n395 & n542;
  assign n544 = n543 ^ n137;
  assign n545 = n393 & ~n544;
  assign n546 = n135 & ~n545;
  assign n547 = n389 & ~n546;
  assign n548 = n547 ^ n381;
  assign n549 = n385 & n548;
  assign n550 = n549 ^ n547;
  assign n551 = n381 & n550;
  assign n552 = n551 ^ n129;
  assign n553 = n407 ^ n403;
  assign n554 = n189 & n478;
  assign n555 = ~n477 & ~n554;
  assign n556 = n462 & ~n555;
  assign n557 = n451 & ~n556;
  assign n558 = n458 & ~n557;
  assign n559 = n455 & ~n558;
  assign n560 = n453 & ~n559;
  assign n561 = n446 & ~n560;
  assign n562 = n444 & ~n561;
  assign n563 = n441 & ~n562;
  assign n564 = n439 & ~n563;
  assign n565 = n435 & ~n564;
  assign n566 = n433 & ~n565;
  assign n567 = n430 & ~n566;
  assign n568 = n428 & ~n567;
  assign n569 = n424 & ~n568;
  assign n570 = n419 & ~n569;
  assign n571 = n421 & ~n570;
  assign n572 = n415 & ~n571;
  assign n573 = n411 & ~n572;
  assign n574 = n573 ^ n409;
  assign n575 = n553 & n574;
  assign n576 = n575 ^ n573;
  assign n577 = n409 & n576;
  assign n578 = n577 ^ n403;
  assign n579 = n466 & ~n578;
  assign n580 = n399 & ~n579;
  assign n581 = n464 & ~n580;
  assign n582 = n395 & ~n581;
  assign n583 = n392 & ~n582;
  assign n584 = n388 & ~n583;
  assign n585 = n386 & ~n584;
  assign n586 = n381 & ~n585;
  assign n587 = n381 & n386;
  assign n588 = n413 & n426;
  assign n591 = n436 & ~n442;
  assign n592 = n431 & ~n591;
  assign n589 = n456 & ~n477;
  assign n590 = n449 & ~n589;
  assign n593 = n592 ^ n590;
  assign n594 = n588 & ~n593;
  assign n595 = n413 & ~n422;
  assign n596 = n595 ^ n409;
  assign n597 = ~n594 & n596;
  assign n598 = n467 & ~n597;
  assign n599 = n465 & ~n598;
  assign n600 = n392 & ~n599;
  assign n601 = n587 & ~n600;
  assign n602 = n393 & ~n473;
  assign n603 = n393 & n468;
  assign n604 = n588 & n603;
  assign n605 = ~n449 & n604;
  assign n606 = n605 ^ n603;
  assign n607 = ~x0 & ~x1;
  assign n608 = n449 & n607;
  assign n609 = n604 & n608;
  assign n610 = ~n471 & n609;
  assign n611 = ~n481 & n610;
  assign n612 = ~n590 & n611;
  assign n613 = ~n557 & n612;
  assign y0 = n379;
  assign y1 = ~n552;
  assign y2 = ~n586;
  assign y3 = ~n601;
  assign y4 = ~n602;
  assign y5 = ~n606;
  assign y6 = ~n604;
  assign y7 = ~n613;
endmodule
