// Benchmark "auction_BMR_2_32" written by ABC on Tue Nov 26 13:54:10 2019

module auction_BMR_2_32 ( 
    \p_input[0] , \p_input[1] , \p_input[2] , \p_input[3] , \p_input[4] ,
    \p_input[5] , \p_input[6] , \p_input[7] , \p_input[8] , \p_input[9] ,
    \p_input[10] , \p_input[11] , \p_input[12] , \p_input[13] ,
    \p_input[14] , \p_input[15] , \p_input[16] , \p_input[17] ,
    \p_input[18] , \p_input[19] , \p_input[20] , \p_input[21] ,
    \p_input[22] , \p_input[23] , \p_input[24] , \p_input[25] ,
    \p_input[26] , \p_input[27] , \p_input[28] , \p_input[29] ,
    \p_input[30] , \p_input[31] , \p_input[32] , \p_input[33] ,
    \p_input[34] , \p_input[35] , \p_input[36] , \p_input[37] ,
    \p_input[38] , \p_input[39] , \p_input[40] , \p_input[41] ,
    \p_input[42] , \p_input[43] , \p_input[44] , \p_input[45] ,
    \p_input[46] , \p_input[47] , \p_input[48] , \p_input[49] ,
    \p_input[50] , \p_input[51] , \p_input[52] , \p_input[53] ,
    \p_input[54] , \p_input[55] , \p_input[56] , \p_input[57] ,
    \p_input[58] , \p_input[59] , \p_input[60] , \p_input[61] ,
    \p_input[62] , \p_input[63] , \p_input[64] , \p_input[65] ,
    \p_input[66] , \p_input[67] , \p_input[68] , \p_input[69] ,
    \p_input[70] , \p_input[71] , \p_input[72] , \p_input[73] ,
    \p_input[74] , \p_input[75] , \p_input[76] , \p_input[77] ,
    \p_input[78] , \p_input[79] , \p_input[80] , \p_input[81] ,
    \p_input[82] , \p_input[83] , \p_input[84] , \p_input[85] ,
    \p_input[86] , \p_input[87] , \p_input[88] , \p_input[89] ,
    \p_input[90] , \p_input[91] , \p_input[92] , \p_input[93] ,
    \p_input[94] , \p_input[95] , \p_input[96] , \p_input[97] ,
    \p_input[98] , \p_input[99] , \p_input[100] , \p_input[101] ,
    \p_input[102] , \p_input[103] , \p_input[104] , \p_input[105] ,
    \p_input[106] , \p_input[107] , \p_input[108] , \p_input[109] ,
    \p_input[110] , \p_input[111] , \p_input[112] , \p_input[113] ,
    \p_input[114] , \p_input[115] , \p_input[116] , \p_input[117] ,
    \p_input[118] , \p_input[119] , \p_input[120] , \p_input[121] ,
    \p_input[122] , \p_input[123] , \p_input[124] , \p_input[125] ,
    \p_input[126] , \p_input[127] ,
    \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] , \o[8] ,
    \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] , \o[16] ,
    \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] , \o[24] ,
    \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] , \o[32] ,
    \o[33]   );
  input  \p_input[0] , \p_input[1] , \p_input[2] , \p_input[3] ,
    \p_input[4] , \p_input[5] , \p_input[6] , \p_input[7] , \p_input[8] ,
    \p_input[9] , \p_input[10] , \p_input[11] , \p_input[12] ,
    \p_input[13] , \p_input[14] , \p_input[15] , \p_input[16] ,
    \p_input[17] , \p_input[18] , \p_input[19] , \p_input[20] ,
    \p_input[21] , \p_input[22] , \p_input[23] , \p_input[24] ,
    \p_input[25] , \p_input[26] , \p_input[27] , \p_input[28] ,
    \p_input[29] , \p_input[30] , \p_input[31] , \p_input[32] ,
    \p_input[33] , \p_input[34] , \p_input[35] , \p_input[36] ,
    \p_input[37] , \p_input[38] , \p_input[39] , \p_input[40] ,
    \p_input[41] , \p_input[42] , \p_input[43] , \p_input[44] ,
    \p_input[45] , \p_input[46] , \p_input[47] , \p_input[48] ,
    \p_input[49] , \p_input[50] , \p_input[51] , \p_input[52] ,
    \p_input[53] , \p_input[54] , \p_input[55] , \p_input[56] ,
    \p_input[57] , \p_input[58] , \p_input[59] , \p_input[60] ,
    \p_input[61] , \p_input[62] , \p_input[63] , \p_input[64] ,
    \p_input[65] , \p_input[66] , \p_input[67] , \p_input[68] ,
    \p_input[69] , \p_input[70] , \p_input[71] , \p_input[72] ,
    \p_input[73] , \p_input[74] , \p_input[75] , \p_input[76] ,
    \p_input[77] , \p_input[78] , \p_input[79] , \p_input[80] ,
    \p_input[81] , \p_input[82] , \p_input[83] , \p_input[84] ,
    \p_input[85] , \p_input[86] , \p_input[87] , \p_input[88] ,
    \p_input[89] , \p_input[90] , \p_input[91] , \p_input[92] ,
    \p_input[93] , \p_input[94] , \p_input[95] , \p_input[96] ,
    \p_input[97] , \p_input[98] , \p_input[99] , \p_input[100] ,
    \p_input[101] , \p_input[102] , \p_input[103] , \p_input[104] ,
    \p_input[105] , \p_input[106] , \p_input[107] , \p_input[108] ,
    \p_input[109] , \p_input[110] , \p_input[111] , \p_input[112] ,
    \p_input[113] , \p_input[114] , \p_input[115] , \p_input[116] ,
    \p_input[117] , \p_input[118] , \p_input[119] , \p_input[120] ,
    \p_input[121] , \p_input[122] , \p_input[123] , \p_input[124] ,
    \p_input[125] , \p_input[126] , \p_input[127] ;
  output \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] ,
    \o[8] , \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] ,
    \o[16] , \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] ,
    \o[24] , \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] ,
    \o[32] , \o[33] ;
  wire new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_,
    new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_,
    new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_,
    new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_,
    new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_,
    new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_,
    new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_,
    new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_,
    new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_,
    new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_,
    new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_,
    new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_,
    new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_,
    new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_,
    new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_,
    new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_,
    new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_,
    new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_,
    new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_,
    new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_,
    new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_,
    new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_,
    new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_,
    new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_,
    new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_,
    new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_,
    new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_,
    new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_,
    new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_,
    new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_,
    new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_,
    new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_,
    new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_,
    new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_,
    new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_,
    new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_,
    new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_,
    new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_,
    new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_,
    new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n819_, new_n820_;
  assign new_n163_ = ~\p_input[95]  & \p_input[127] ;
  assign new_n164_ = \p_input[95]  & ~\p_input[127] ;
  assign new_n165_ = ~\p_input[94]  & \p_input[126] ;
  assign new_n166_ = \p_input[94]  & ~\p_input[126] ;
  assign new_n167_ = ~\p_input[93]  & \p_input[125] ;
  assign new_n168_ = \p_input[93]  & ~\p_input[125] ;
  assign new_n169_ = ~\p_input[92]  & \p_input[124] ;
  assign new_n170_ = \p_input[92]  & ~\p_input[124] ;
  assign new_n171_ = ~\p_input[91]  & \p_input[123] ;
  assign new_n172_ = \p_input[91]  & ~\p_input[123] ;
  assign new_n173_ = ~\p_input[90]  & \p_input[122] ;
  assign new_n174_ = \p_input[90]  & ~\p_input[122] ;
  assign new_n175_ = ~\p_input[89]  & \p_input[121] ;
  assign new_n176_ = \p_input[89]  & ~\p_input[121] ;
  assign new_n177_ = ~\p_input[88]  & \p_input[120] ;
  assign new_n178_ = \p_input[88]  & ~\p_input[120] ;
  assign new_n179_ = ~\p_input[87]  & \p_input[119] ;
  assign new_n180_ = \p_input[87]  & ~\p_input[119] ;
  assign new_n181_ = ~\p_input[86]  & \p_input[118] ;
  assign new_n182_ = \p_input[86]  & ~\p_input[118] ;
  assign new_n183_ = ~\p_input[85]  & \p_input[117] ;
  assign new_n184_ = \p_input[85]  & ~\p_input[117] ;
  assign new_n185_ = ~\p_input[84]  & \p_input[116] ;
  assign new_n186_ = \p_input[84]  & ~\p_input[116] ;
  assign new_n187_ = ~\p_input[83]  & \p_input[115] ;
  assign new_n188_ = \p_input[83]  & ~\p_input[115] ;
  assign new_n189_ = ~\p_input[82]  & \p_input[114] ;
  assign new_n190_ = \p_input[82]  & ~\p_input[114] ;
  assign new_n191_ = ~\p_input[81]  & \p_input[113] ;
  assign new_n192_ = \p_input[81]  & ~\p_input[113] ;
  assign new_n193_ = ~\p_input[80]  & \p_input[112] ;
  assign new_n194_ = \p_input[80]  & ~\p_input[112] ;
  assign new_n195_ = ~\p_input[79]  & \p_input[111] ;
  assign new_n196_ = \p_input[79]  & ~\p_input[111] ;
  assign new_n197_ = ~\p_input[78]  & \p_input[110] ;
  assign new_n198_ = \p_input[78]  & ~\p_input[110] ;
  assign new_n199_ = ~\p_input[77]  & \p_input[109] ;
  assign new_n200_ = \p_input[77]  & ~\p_input[109] ;
  assign new_n201_ = ~\p_input[76]  & \p_input[108] ;
  assign new_n202_ = \p_input[76]  & ~\p_input[108] ;
  assign new_n203_ = ~\p_input[75]  & \p_input[107] ;
  assign new_n204_ = \p_input[75]  & ~\p_input[107] ;
  assign new_n205_ = ~\p_input[74]  & \p_input[106] ;
  assign new_n206_ = \p_input[74]  & ~\p_input[106] ;
  assign new_n207_ = ~\p_input[73]  & \p_input[105] ;
  assign new_n208_ = \p_input[73]  & ~\p_input[105] ;
  assign new_n209_ = ~\p_input[72]  & \p_input[104] ;
  assign new_n210_ = \p_input[72]  & ~\p_input[104] ;
  assign new_n211_ = ~\p_input[71]  & \p_input[103] ;
  assign new_n212_ = \p_input[71]  & ~\p_input[103] ;
  assign new_n213_ = ~\p_input[70]  & \p_input[102] ;
  assign new_n214_ = \p_input[70]  & ~\p_input[102] ;
  assign new_n215_ = ~\p_input[69]  & \p_input[101] ;
  assign new_n216_ = \p_input[69]  & ~\p_input[101] ;
  assign new_n217_ = ~\p_input[68]  & \p_input[100] ;
  assign new_n218_ = \p_input[68]  & ~\p_input[100] ;
  assign new_n219_ = ~\p_input[67]  & \p_input[99] ;
  assign new_n220_ = \p_input[67]  & ~\p_input[99] ;
  assign new_n221_ = ~\p_input[66]  & \p_input[98] ;
  assign new_n222_ = \p_input[66]  & ~\p_input[98] ;
  assign new_n223_ = ~\p_input[65]  & \p_input[97] ;
  assign new_n224_ = \p_input[65]  & ~\p_input[97] ;
  assign new_n225_ = \p_input[64]  & ~\p_input[96] ;
  assign new_n226_ = ~new_n224_ & ~new_n225_;
  assign new_n227_ = ~new_n223_ & ~new_n226_;
  assign new_n228_ = ~new_n222_ & ~new_n227_;
  assign new_n229_ = ~new_n221_ & ~new_n228_;
  assign new_n230_ = ~new_n220_ & ~new_n229_;
  assign new_n231_ = ~new_n219_ & ~new_n230_;
  assign new_n232_ = ~new_n218_ & ~new_n231_;
  assign new_n233_ = ~new_n217_ & ~new_n232_;
  assign new_n234_ = ~new_n216_ & ~new_n233_;
  assign new_n235_ = ~new_n215_ & ~new_n234_;
  assign new_n236_ = ~new_n214_ & ~new_n235_;
  assign new_n237_ = ~new_n213_ & ~new_n236_;
  assign new_n238_ = ~new_n212_ & ~new_n237_;
  assign new_n239_ = ~new_n211_ & ~new_n238_;
  assign new_n240_ = ~new_n210_ & ~new_n239_;
  assign new_n241_ = ~new_n209_ & ~new_n240_;
  assign new_n242_ = ~new_n208_ & ~new_n241_;
  assign new_n243_ = ~new_n207_ & ~new_n242_;
  assign new_n244_ = ~new_n206_ & ~new_n243_;
  assign new_n245_ = ~new_n205_ & ~new_n244_;
  assign new_n246_ = ~new_n204_ & ~new_n245_;
  assign new_n247_ = ~new_n203_ & ~new_n246_;
  assign new_n248_ = ~new_n202_ & ~new_n247_;
  assign new_n249_ = ~new_n201_ & ~new_n248_;
  assign new_n250_ = ~new_n200_ & ~new_n249_;
  assign new_n251_ = ~new_n199_ & ~new_n250_;
  assign new_n252_ = ~new_n198_ & ~new_n251_;
  assign new_n253_ = ~new_n197_ & ~new_n252_;
  assign new_n254_ = ~new_n196_ & ~new_n253_;
  assign new_n255_ = ~new_n195_ & ~new_n254_;
  assign new_n256_ = ~new_n194_ & ~new_n255_;
  assign new_n257_ = ~new_n193_ & ~new_n256_;
  assign new_n258_ = ~new_n192_ & ~new_n257_;
  assign new_n259_ = ~new_n191_ & ~new_n258_;
  assign new_n260_ = ~new_n190_ & ~new_n259_;
  assign new_n261_ = ~new_n189_ & ~new_n260_;
  assign new_n262_ = ~new_n188_ & ~new_n261_;
  assign new_n263_ = ~new_n187_ & ~new_n262_;
  assign new_n264_ = ~new_n186_ & ~new_n263_;
  assign new_n265_ = ~new_n185_ & ~new_n264_;
  assign new_n266_ = ~new_n184_ & ~new_n265_;
  assign new_n267_ = ~new_n183_ & ~new_n266_;
  assign new_n268_ = ~new_n182_ & ~new_n267_;
  assign new_n269_ = ~new_n181_ & ~new_n268_;
  assign new_n270_ = ~new_n180_ & ~new_n269_;
  assign new_n271_ = ~new_n179_ & ~new_n270_;
  assign new_n272_ = ~new_n178_ & ~new_n271_;
  assign new_n273_ = ~new_n177_ & ~new_n272_;
  assign new_n274_ = ~new_n176_ & ~new_n273_;
  assign new_n275_ = ~new_n175_ & ~new_n274_;
  assign new_n276_ = ~new_n174_ & ~new_n275_;
  assign new_n277_ = ~new_n173_ & ~new_n276_;
  assign new_n278_ = ~new_n172_ & ~new_n277_;
  assign new_n279_ = ~new_n171_ & ~new_n278_;
  assign new_n280_ = ~new_n170_ & ~new_n279_;
  assign new_n281_ = ~new_n169_ & ~new_n280_;
  assign new_n282_ = ~new_n168_ & ~new_n281_;
  assign new_n283_ = ~new_n167_ & ~new_n282_;
  assign new_n284_ = ~new_n166_ & ~new_n283_;
  assign new_n285_ = ~new_n165_ & ~new_n284_;
  assign new_n286_ = ~new_n164_ & ~new_n285_;
  assign new_n287_ = ~new_n163_ & ~new_n286_;
  assign new_n288_ = ~\p_input[95]  & ~\p_input[127] ;
  assign new_n289_ = ~\p_input[31]  & ~\p_input[63] ;
  assign new_n290_ = ~new_n288_ & new_n289_;
  assign new_n291_ = new_n288_ & ~new_n289_;
  assign new_n292_ = \p_input[126]  & ~new_n287_;
  assign new_n293_ = \p_input[94]  & new_n287_;
  assign new_n294_ = ~new_n292_ & ~new_n293_;
  assign new_n295_ = ~\p_input[31]  & \p_input[63] ;
  assign new_n296_ = \p_input[31]  & ~\p_input[63] ;
  assign new_n297_ = ~\p_input[30]  & \p_input[62] ;
  assign new_n298_ = \p_input[30]  & ~\p_input[62] ;
  assign new_n299_ = ~\p_input[29]  & \p_input[61] ;
  assign new_n300_ = \p_input[29]  & ~\p_input[61] ;
  assign new_n301_ = ~\p_input[28]  & \p_input[60] ;
  assign new_n302_ = \p_input[28]  & ~\p_input[60] ;
  assign new_n303_ = ~\p_input[27]  & \p_input[59] ;
  assign new_n304_ = \p_input[27]  & ~\p_input[59] ;
  assign new_n305_ = ~\p_input[26]  & \p_input[58] ;
  assign new_n306_ = \p_input[26]  & ~\p_input[58] ;
  assign new_n307_ = ~\p_input[25]  & \p_input[57] ;
  assign new_n308_ = \p_input[25]  & ~\p_input[57] ;
  assign new_n309_ = ~\p_input[24]  & \p_input[56] ;
  assign new_n310_ = \p_input[24]  & ~\p_input[56] ;
  assign new_n311_ = ~\p_input[23]  & \p_input[55] ;
  assign new_n312_ = \p_input[23]  & ~\p_input[55] ;
  assign new_n313_ = ~\p_input[22]  & \p_input[54] ;
  assign new_n314_ = \p_input[22]  & ~\p_input[54] ;
  assign new_n315_ = ~\p_input[21]  & \p_input[53] ;
  assign new_n316_ = \p_input[21]  & ~\p_input[53] ;
  assign new_n317_ = ~\p_input[20]  & \p_input[52] ;
  assign new_n318_ = \p_input[20]  & ~\p_input[52] ;
  assign new_n319_ = ~\p_input[19]  & \p_input[51] ;
  assign new_n320_ = \p_input[19]  & ~\p_input[51] ;
  assign new_n321_ = ~\p_input[18]  & \p_input[50] ;
  assign new_n322_ = \p_input[18]  & ~\p_input[50] ;
  assign new_n323_ = ~\p_input[17]  & \p_input[49] ;
  assign new_n324_ = \p_input[17]  & ~\p_input[49] ;
  assign new_n325_ = ~\p_input[16]  & \p_input[48] ;
  assign new_n326_ = \p_input[16]  & ~\p_input[48] ;
  assign new_n327_ = ~\p_input[15]  & \p_input[47] ;
  assign new_n328_ = \p_input[15]  & ~\p_input[47] ;
  assign new_n329_ = ~\p_input[14]  & \p_input[46] ;
  assign new_n330_ = \p_input[14]  & ~\p_input[46] ;
  assign new_n331_ = ~\p_input[13]  & \p_input[45] ;
  assign new_n332_ = \p_input[13]  & ~\p_input[45] ;
  assign new_n333_ = ~\p_input[12]  & \p_input[44] ;
  assign new_n334_ = \p_input[12]  & ~\p_input[44] ;
  assign new_n335_ = ~\p_input[11]  & \p_input[43] ;
  assign new_n336_ = \p_input[11]  & ~\p_input[43] ;
  assign new_n337_ = ~\p_input[10]  & \p_input[42] ;
  assign new_n338_ = \p_input[10]  & ~\p_input[42] ;
  assign new_n339_ = ~\p_input[9]  & \p_input[41] ;
  assign new_n340_ = \p_input[9]  & ~\p_input[41] ;
  assign new_n341_ = ~\p_input[8]  & \p_input[40] ;
  assign new_n342_ = \p_input[8]  & ~\p_input[40] ;
  assign new_n343_ = ~\p_input[7]  & \p_input[39] ;
  assign new_n344_ = \p_input[7]  & ~\p_input[39] ;
  assign new_n345_ = ~\p_input[6]  & \p_input[38] ;
  assign new_n346_ = \p_input[6]  & ~\p_input[38] ;
  assign new_n347_ = ~\p_input[5]  & \p_input[37] ;
  assign new_n348_ = \p_input[5]  & ~\p_input[37] ;
  assign new_n349_ = ~\p_input[4]  & \p_input[36] ;
  assign new_n350_ = \p_input[4]  & ~\p_input[36] ;
  assign new_n351_ = ~\p_input[3]  & \p_input[35] ;
  assign new_n352_ = \p_input[3]  & ~\p_input[35] ;
  assign new_n353_ = ~\p_input[2]  & \p_input[34] ;
  assign new_n354_ = \p_input[2]  & ~\p_input[34] ;
  assign new_n355_ = ~\p_input[1]  & \p_input[33] ;
  assign new_n356_ = \p_input[1]  & ~\p_input[33] ;
  assign new_n357_ = \p_input[0]  & ~\p_input[32] ;
  assign new_n358_ = ~new_n356_ & ~new_n357_;
  assign new_n359_ = ~new_n355_ & ~new_n358_;
  assign new_n360_ = ~new_n354_ & ~new_n359_;
  assign new_n361_ = ~new_n353_ & ~new_n360_;
  assign new_n362_ = ~new_n352_ & ~new_n361_;
  assign new_n363_ = ~new_n351_ & ~new_n362_;
  assign new_n364_ = ~new_n350_ & ~new_n363_;
  assign new_n365_ = ~new_n349_ & ~new_n364_;
  assign new_n366_ = ~new_n348_ & ~new_n365_;
  assign new_n367_ = ~new_n347_ & ~new_n366_;
  assign new_n368_ = ~new_n346_ & ~new_n367_;
  assign new_n369_ = ~new_n345_ & ~new_n368_;
  assign new_n370_ = ~new_n344_ & ~new_n369_;
  assign new_n371_ = ~new_n343_ & ~new_n370_;
  assign new_n372_ = ~new_n342_ & ~new_n371_;
  assign new_n373_ = ~new_n341_ & ~new_n372_;
  assign new_n374_ = ~new_n340_ & ~new_n373_;
  assign new_n375_ = ~new_n339_ & ~new_n374_;
  assign new_n376_ = ~new_n338_ & ~new_n375_;
  assign new_n377_ = ~new_n337_ & ~new_n376_;
  assign new_n378_ = ~new_n336_ & ~new_n377_;
  assign new_n379_ = ~new_n335_ & ~new_n378_;
  assign new_n380_ = ~new_n334_ & ~new_n379_;
  assign new_n381_ = ~new_n333_ & ~new_n380_;
  assign new_n382_ = ~new_n332_ & ~new_n381_;
  assign new_n383_ = ~new_n331_ & ~new_n382_;
  assign new_n384_ = ~new_n330_ & ~new_n383_;
  assign new_n385_ = ~new_n329_ & ~new_n384_;
  assign new_n386_ = ~new_n328_ & ~new_n385_;
  assign new_n387_ = ~new_n327_ & ~new_n386_;
  assign new_n388_ = ~new_n326_ & ~new_n387_;
  assign new_n389_ = ~new_n325_ & ~new_n388_;
  assign new_n390_ = ~new_n324_ & ~new_n389_;
  assign new_n391_ = ~new_n323_ & ~new_n390_;
  assign new_n392_ = ~new_n322_ & ~new_n391_;
  assign new_n393_ = ~new_n321_ & ~new_n392_;
  assign new_n394_ = ~new_n320_ & ~new_n393_;
  assign new_n395_ = ~new_n319_ & ~new_n394_;
  assign new_n396_ = ~new_n318_ & ~new_n395_;
  assign new_n397_ = ~new_n317_ & ~new_n396_;
  assign new_n398_ = ~new_n316_ & ~new_n397_;
  assign new_n399_ = ~new_n315_ & ~new_n398_;
  assign new_n400_ = ~new_n314_ & ~new_n399_;
  assign new_n401_ = ~new_n313_ & ~new_n400_;
  assign new_n402_ = ~new_n312_ & ~new_n401_;
  assign new_n403_ = ~new_n311_ & ~new_n402_;
  assign new_n404_ = ~new_n310_ & ~new_n403_;
  assign new_n405_ = ~new_n309_ & ~new_n404_;
  assign new_n406_ = ~new_n308_ & ~new_n405_;
  assign new_n407_ = ~new_n307_ & ~new_n406_;
  assign new_n408_ = ~new_n306_ & ~new_n407_;
  assign new_n409_ = ~new_n305_ & ~new_n408_;
  assign new_n410_ = ~new_n304_ & ~new_n409_;
  assign new_n411_ = ~new_n303_ & ~new_n410_;
  assign new_n412_ = ~new_n302_ & ~new_n411_;
  assign new_n413_ = ~new_n301_ & ~new_n412_;
  assign new_n414_ = ~new_n300_ & ~new_n413_;
  assign new_n415_ = ~new_n299_ & ~new_n414_;
  assign new_n416_ = ~new_n298_ & ~new_n415_;
  assign new_n417_ = ~new_n297_ & ~new_n416_;
  assign new_n418_ = ~new_n296_ & ~new_n417_;
  assign new_n419_ = ~new_n295_ & ~new_n418_;
  assign new_n420_ = \p_input[62]  & ~new_n419_;
  assign new_n421_ = \p_input[30]  & new_n419_;
  assign new_n422_ = ~new_n420_ & ~new_n421_;
  assign new_n423_ = ~new_n294_ & new_n422_;
  assign new_n424_ = \p_input[97]  & ~new_n287_;
  assign new_n425_ = \p_input[65]  & new_n287_;
  assign new_n426_ = ~new_n424_ & ~new_n425_;
  assign new_n427_ = \p_input[33]  & ~new_n419_;
  assign new_n428_ = \p_input[1]  & new_n419_;
  assign new_n429_ = ~new_n427_ & ~new_n428_;
  assign new_n430_ = ~new_n426_ & new_n429_;
  assign new_n431_ = \p_input[96]  & ~new_n287_;
  assign new_n432_ = \p_input[64]  & new_n287_;
  assign new_n433_ = ~new_n431_ & ~new_n432_;
  assign new_n434_ = \p_input[32]  & ~new_n419_;
  assign new_n435_ = \p_input[0]  & new_n419_;
  assign new_n436_ = ~new_n434_ & ~new_n435_;
  assign new_n437_ = new_n433_ & ~new_n436_;
  assign new_n438_ = ~new_n430_ & new_n437_;
  assign new_n439_ = \p_input[98]  & ~new_n287_;
  assign new_n440_ = \p_input[66]  & new_n287_;
  assign new_n441_ = ~new_n439_ & ~new_n440_;
  assign new_n442_ = \p_input[34]  & ~new_n419_;
  assign new_n443_ = \p_input[2]  & new_n419_;
  assign new_n444_ = ~new_n442_ & ~new_n443_;
  assign new_n445_ = new_n441_ & ~new_n444_;
  assign new_n446_ = new_n426_ & ~new_n429_;
  assign new_n447_ = ~new_n445_ & ~new_n446_;
  assign new_n448_ = ~new_n438_ & new_n447_;
  assign new_n449_ = \p_input[99]  & ~new_n287_;
  assign new_n450_ = \p_input[67]  & new_n287_;
  assign new_n451_ = ~new_n449_ & ~new_n450_;
  assign new_n452_ = \p_input[35]  & ~new_n419_;
  assign new_n453_ = \p_input[3]  & new_n419_;
  assign new_n454_ = ~new_n452_ & ~new_n453_;
  assign new_n455_ = ~new_n451_ & new_n454_;
  assign new_n456_ = ~new_n441_ & new_n444_;
  assign new_n457_ = ~new_n455_ & ~new_n456_;
  assign new_n458_ = ~new_n448_ & new_n457_;
  assign new_n459_ = \p_input[100]  & ~new_n287_;
  assign new_n460_ = \p_input[68]  & new_n287_;
  assign new_n461_ = ~new_n459_ & ~new_n460_;
  assign new_n462_ = \p_input[36]  & ~new_n419_;
  assign new_n463_ = \p_input[4]  & new_n419_;
  assign new_n464_ = ~new_n462_ & ~new_n463_;
  assign new_n465_ = new_n461_ & ~new_n464_;
  assign new_n466_ = new_n451_ & ~new_n454_;
  assign new_n467_ = ~new_n465_ & ~new_n466_;
  assign new_n468_ = ~new_n458_ & new_n467_;
  assign new_n469_ = ~new_n461_ & new_n464_;
  assign new_n470_ = \p_input[101]  & ~new_n287_;
  assign new_n471_ = \p_input[69]  & new_n287_;
  assign new_n472_ = ~new_n470_ & ~new_n471_;
  assign new_n473_ = \p_input[37]  & ~new_n419_;
  assign new_n474_ = \p_input[5]  & new_n419_;
  assign new_n475_ = ~new_n473_ & ~new_n474_;
  assign new_n476_ = ~new_n472_ & new_n475_;
  assign new_n477_ = ~new_n469_ & ~new_n476_;
  assign new_n478_ = ~new_n468_ & new_n477_;
  assign new_n479_ = \p_input[102]  & ~new_n287_;
  assign new_n480_ = \p_input[70]  & new_n287_;
  assign new_n481_ = ~new_n479_ & ~new_n480_;
  assign new_n482_ = \p_input[38]  & ~new_n419_;
  assign new_n483_ = \p_input[6]  & new_n419_;
  assign new_n484_ = ~new_n482_ & ~new_n483_;
  assign new_n485_ = new_n481_ & ~new_n484_;
  assign new_n486_ = new_n472_ & ~new_n475_;
  assign new_n487_ = ~new_n485_ & ~new_n486_;
  assign new_n488_ = ~new_n478_ & new_n487_;
  assign new_n489_ = \p_input[39]  & ~new_n419_;
  assign new_n490_ = \p_input[7]  & new_n419_;
  assign new_n491_ = ~new_n489_ & ~new_n490_;
  assign new_n492_ = \p_input[103]  & ~new_n287_;
  assign new_n493_ = \p_input[71]  & new_n287_;
  assign new_n494_ = ~new_n492_ & ~new_n493_;
  assign new_n495_ = new_n491_ & ~new_n494_;
  assign new_n496_ = ~new_n481_ & new_n484_;
  assign new_n497_ = ~new_n495_ & ~new_n496_;
  assign new_n498_ = ~new_n488_ & new_n497_;
  assign new_n499_ = ~new_n491_ & new_n494_;
  assign new_n500_ = \p_input[104]  & ~new_n287_;
  assign new_n501_ = \p_input[72]  & new_n287_;
  assign new_n502_ = ~new_n500_ & ~new_n501_;
  assign new_n503_ = \p_input[40]  & ~new_n419_;
  assign new_n504_ = \p_input[8]  & new_n419_;
  assign new_n505_ = ~new_n503_ & ~new_n504_;
  assign new_n506_ = new_n502_ & ~new_n505_;
  assign new_n507_ = ~new_n499_ & ~new_n506_;
  assign new_n508_ = ~new_n498_ & new_n507_;
  assign new_n509_ = ~new_n502_ & new_n505_;
  assign new_n510_ = \p_input[105]  & ~new_n287_;
  assign new_n511_ = \p_input[73]  & new_n287_;
  assign new_n512_ = ~new_n510_ & ~new_n511_;
  assign new_n513_ = \p_input[41]  & ~new_n419_;
  assign new_n514_ = \p_input[9]  & new_n419_;
  assign new_n515_ = ~new_n513_ & ~new_n514_;
  assign new_n516_ = ~new_n512_ & new_n515_;
  assign new_n517_ = ~new_n509_ & ~new_n516_;
  assign new_n518_ = ~new_n508_ & new_n517_;
  assign new_n519_ = new_n512_ & ~new_n515_;
  assign new_n520_ = \p_input[42]  & ~new_n419_;
  assign new_n521_ = \p_input[10]  & new_n419_;
  assign new_n522_ = ~new_n520_ & ~new_n521_;
  assign new_n523_ = \p_input[106]  & ~new_n287_;
  assign new_n524_ = \p_input[74]  & new_n287_;
  assign new_n525_ = ~new_n523_ & ~new_n524_;
  assign new_n526_ = ~new_n522_ & new_n525_;
  assign new_n527_ = ~new_n519_ & ~new_n526_;
  assign new_n528_ = ~new_n518_ & new_n527_;
  assign new_n529_ = \p_input[43]  & ~new_n419_;
  assign new_n530_ = \p_input[11]  & new_n419_;
  assign new_n531_ = ~new_n529_ & ~new_n530_;
  assign new_n532_ = \p_input[107]  & ~new_n287_;
  assign new_n533_ = \p_input[75]  & new_n287_;
  assign new_n534_ = ~new_n532_ & ~new_n533_;
  assign new_n535_ = new_n531_ & ~new_n534_;
  assign new_n536_ = new_n522_ & ~new_n525_;
  assign new_n537_ = ~new_n535_ & ~new_n536_;
  assign new_n538_ = ~new_n528_ & new_n537_;
  assign new_n539_ = \p_input[108]  & ~new_n287_;
  assign new_n540_ = \p_input[76]  & new_n287_;
  assign new_n541_ = ~new_n539_ & ~new_n540_;
  assign new_n542_ = \p_input[44]  & ~new_n419_;
  assign new_n543_ = \p_input[12]  & new_n419_;
  assign new_n544_ = ~new_n542_ & ~new_n543_;
  assign new_n545_ = new_n541_ & ~new_n544_;
  assign new_n546_ = ~new_n531_ & new_n534_;
  assign new_n547_ = ~new_n545_ & ~new_n546_;
  assign new_n548_ = ~new_n538_ & new_n547_;
  assign new_n549_ = ~new_n541_ & new_n544_;
  assign new_n550_ = \p_input[109]  & ~new_n287_;
  assign new_n551_ = \p_input[77]  & new_n287_;
  assign new_n552_ = ~new_n550_ & ~new_n551_;
  assign new_n553_ = \p_input[45]  & ~new_n419_;
  assign new_n554_ = \p_input[13]  & new_n419_;
  assign new_n555_ = ~new_n553_ & ~new_n554_;
  assign new_n556_ = ~new_n552_ & new_n555_;
  assign new_n557_ = ~new_n549_ & ~new_n556_;
  assign new_n558_ = ~new_n548_ & new_n557_;
  assign new_n559_ = new_n552_ & ~new_n555_;
  assign new_n560_ = \p_input[46]  & ~new_n419_;
  assign new_n561_ = \p_input[14]  & new_n419_;
  assign new_n562_ = ~new_n560_ & ~new_n561_;
  assign new_n563_ = \p_input[110]  & ~new_n287_;
  assign new_n564_ = \p_input[78]  & new_n287_;
  assign new_n565_ = ~new_n563_ & ~new_n564_;
  assign new_n566_ = ~new_n562_ & new_n565_;
  assign new_n567_ = ~new_n559_ & ~new_n566_;
  assign new_n568_ = ~new_n558_ & new_n567_;
  assign new_n569_ = \p_input[47]  & ~new_n419_;
  assign new_n570_ = \p_input[15]  & new_n419_;
  assign new_n571_ = ~new_n569_ & ~new_n570_;
  assign new_n572_ = \p_input[111]  & ~new_n287_;
  assign new_n573_ = \p_input[79]  & new_n287_;
  assign new_n574_ = ~new_n572_ & ~new_n573_;
  assign new_n575_ = new_n571_ & ~new_n574_;
  assign new_n576_ = new_n562_ & ~new_n565_;
  assign new_n577_ = ~new_n575_ & ~new_n576_;
  assign new_n578_ = ~new_n568_ & new_n577_;
  assign new_n579_ = \p_input[112]  & ~new_n287_;
  assign new_n580_ = \p_input[80]  & new_n287_;
  assign new_n581_ = ~new_n579_ & ~new_n580_;
  assign new_n582_ = \p_input[48]  & ~new_n419_;
  assign new_n583_ = \p_input[16]  & new_n419_;
  assign new_n584_ = ~new_n582_ & ~new_n583_;
  assign new_n585_ = new_n581_ & ~new_n584_;
  assign new_n586_ = ~new_n571_ & new_n574_;
  assign new_n587_ = ~new_n585_ & ~new_n586_;
  assign new_n588_ = ~new_n578_ & new_n587_;
  assign new_n589_ = ~new_n581_ & new_n584_;
  assign new_n590_ = \p_input[113]  & ~new_n287_;
  assign new_n591_ = \p_input[81]  & new_n287_;
  assign new_n592_ = ~new_n590_ & ~new_n591_;
  assign new_n593_ = \p_input[49]  & ~new_n419_;
  assign new_n594_ = \p_input[17]  & new_n419_;
  assign new_n595_ = ~new_n593_ & ~new_n594_;
  assign new_n596_ = ~new_n592_ & new_n595_;
  assign new_n597_ = ~new_n589_ & ~new_n596_;
  assign new_n598_ = ~new_n588_ & new_n597_;
  assign new_n599_ = new_n592_ & ~new_n595_;
  assign new_n600_ = \p_input[50]  & ~new_n419_;
  assign new_n601_ = \p_input[18]  & new_n419_;
  assign new_n602_ = ~new_n600_ & ~new_n601_;
  assign new_n603_ = \p_input[114]  & ~new_n287_;
  assign new_n604_ = \p_input[82]  & new_n287_;
  assign new_n605_ = ~new_n603_ & ~new_n604_;
  assign new_n606_ = ~new_n602_ & new_n605_;
  assign new_n607_ = ~new_n599_ & ~new_n606_;
  assign new_n608_ = ~new_n598_ & new_n607_;
  assign new_n609_ = \p_input[51]  & ~new_n419_;
  assign new_n610_ = \p_input[19]  & new_n419_;
  assign new_n611_ = ~new_n609_ & ~new_n610_;
  assign new_n612_ = \p_input[115]  & ~new_n287_;
  assign new_n613_ = \p_input[83]  & new_n287_;
  assign new_n614_ = ~new_n612_ & ~new_n613_;
  assign new_n615_ = new_n611_ & ~new_n614_;
  assign new_n616_ = new_n602_ & ~new_n605_;
  assign new_n617_ = ~new_n615_ & ~new_n616_;
  assign new_n618_ = ~new_n608_ & new_n617_;
  assign new_n619_ = \p_input[116]  & ~new_n287_;
  assign new_n620_ = \p_input[84]  & new_n287_;
  assign new_n621_ = ~new_n619_ & ~new_n620_;
  assign new_n622_ = \p_input[52]  & ~new_n419_;
  assign new_n623_ = \p_input[20]  & new_n419_;
  assign new_n624_ = ~new_n622_ & ~new_n623_;
  assign new_n625_ = new_n621_ & ~new_n624_;
  assign new_n626_ = ~new_n611_ & new_n614_;
  assign new_n627_ = ~new_n625_ & ~new_n626_;
  assign new_n628_ = ~new_n618_ & new_n627_;
  assign new_n629_ = ~new_n621_ & new_n624_;
  assign new_n630_ = \p_input[117]  & ~new_n287_;
  assign new_n631_ = \p_input[85]  & new_n287_;
  assign new_n632_ = ~new_n630_ & ~new_n631_;
  assign new_n633_ = \p_input[53]  & ~new_n419_;
  assign new_n634_ = \p_input[21]  & new_n419_;
  assign new_n635_ = ~new_n633_ & ~new_n634_;
  assign new_n636_ = ~new_n632_ & new_n635_;
  assign new_n637_ = ~new_n629_ & ~new_n636_;
  assign new_n638_ = ~new_n628_ & new_n637_;
  assign new_n639_ = new_n632_ & ~new_n635_;
  assign new_n640_ = \p_input[54]  & ~new_n419_;
  assign new_n641_ = \p_input[22]  & new_n419_;
  assign new_n642_ = ~new_n640_ & ~new_n641_;
  assign new_n643_ = \p_input[118]  & ~new_n287_;
  assign new_n644_ = \p_input[86]  & new_n287_;
  assign new_n645_ = ~new_n643_ & ~new_n644_;
  assign new_n646_ = ~new_n642_ & new_n645_;
  assign new_n647_ = ~new_n639_ & ~new_n646_;
  assign new_n648_ = ~new_n638_ & new_n647_;
  assign new_n649_ = \p_input[55]  & ~new_n419_;
  assign new_n650_ = \p_input[23]  & new_n419_;
  assign new_n651_ = ~new_n649_ & ~new_n650_;
  assign new_n652_ = \p_input[119]  & ~new_n287_;
  assign new_n653_ = \p_input[87]  & new_n287_;
  assign new_n654_ = ~new_n652_ & ~new_n653_;
  assign new_n655_ = new_n651_ & ~new_n654_;
  assign new_n656_ = new_n642_ & ~new_n645_;
  assign new_n657_ = ~new_n655_ & ~new_n656_;
  assign new_n658_ = ~new_n648_ & new_n657_;
  assign new_n659_ = \p_input[120]  & ~new_n287_;
  assign new_n660_ = \p_input[88]  & new_n287_;
  assign new_n661_ = ~new_n659_ & ~new_n660_;
  assign new_n662_ = \p_input[56]  & ~new_n419_;
  assign new_n663_ = \p_input[24]  & new_n419_;
  assign new_n664_ = ~new_n662_ & ~new_n663_;
  assign new_n665_ = new_n661_ & ~new_n664_;
  assign new_n666_ = ~new_n651_ & new_n654_;
  assign new_n667_ = ~new_n665_ & ~new_n666_;
  assign new_n668_ = ~new_n658_ & new_n667_;
  assign new_n669_ = ~new_n661_ & new_n664_;
  assign new_n670_ = \p_input[121]  & ~new_n287_;
  assign new_n671_ = \p_input[89]  & new_n287_;
  assign new_n672_ = ~new_n670_ & ~new_n671_;
  assign new_n673_ = \p_input[57]  & ~new_n419_;
  assign new_n674_ = \p_input[25]  & new_n419_;
  assign new_n675_ = ~new_n673_ & ~new_n674_;
  assign new_n676_ = ~new_n672_ & new_n675_;
  assign new_n677_ = ~new_n669_ & ~new_n676_;
  assign new_n678_ = ~new_n668_ & new_n677_;
  assign new_n679_ = new_n672_ & ~new_n675_;
  assign new_n680_ = \p_input[58]  & ~new_n419_;
  assign new_n681_ = \p_input[26]  & new_n419_;
  assign new_n682_ = ~new_n680_ & ~new_n681_;
  assign new_n683_ = \p_input[122]  & ~new_n287_;
  assign new_n684_ = \p_input[90]  & new_n287_;
  assign new_n685_ = ~new_n683_ & ~new_n684_;
  assign new_n686_ = ~new_n682_ & new_n685_;
  assign new_n687_ = ~new_n679_ & ~new_n686_;
  assign new_n688_ = ~new_n678_ & new_n687_;
  assign new_n689_ = \p_input[59]  & ~new_n419_;
  assign new_n690_ = \p_input[27]  & new_n419_;
  assign new_n691_ = ~new_n689_ & ~new_n690_;
  assign new_n692_ = \p_input[123]  & ~new_n287_;
  assign new_n693_ = \p_input[91]  & new_n287_;
  assign new_n694_ = ~new_n692_ & ~new_n693_;
  assign new_n695_ = new_n691_ & ~new_n694_;
  assign new_n696_ = new_n682_ & ~new_n685_;
  assign new_n697_ = ~new_n695_ & ~new_n696_;
  assign new_n698_ = ~new_n688_ & new_n697_;
  assign new_n699_ = \p_input[124]  & ~new_n287_;
  assign new_n700_ = \p_input[92]  & new_n287_;
  assign new_n701_ = ~new_n699_ & ~new_n700_;
  assign new_n702_ = \p_input[60]  & ~new_n419_;
  assign new_n703_ = \p_input[28]  & new_n419_;
  assign new_n704_ = ~new_n702_ & ~new_n703_;
  assign new_n705_ = new_n701_ & ~new_n704_;
  assign new_n706_ = ~new_n691_ & new_n694_;
  assign new_n707_ = ~new_n705_ & ~new_n706_;
  assign new_n708_ = ~new_n698_ & new_n707_;
  assign new_n709_ = ~new_n701_ & new_n704_;
  assign new_n710_ = \p_input[125]  & ~new_n287_;
  assign new_n711_ = \p_input[93]  & new_n287_;
  assign new_n712_ = ~new_n710_ & ~new_n711_;
  assign new_n713_ = \p_input[61]  & ~new_n419_;
  assign new_n714_ = \p_input[29]  & new_n419_;
  assign new_n715_ = ~new_n713_ & ~new_n714_;
  assign new_n716_ = ~new_n712_ & new_n715_;
  assign new_n717_ = ~new_n709_ & ~new_n716_;
  assign new_n718_ = ~new_n708_ & new_n717_;
  assign new_n719_ = new_n294_ & ~new_n422_;
  assign new_n720_ = new_n712_ & ~new_n715_;
  assign new_n721_ = ~new_n719_ & ~new_n720_;
  assign new_n722_ = ~new_n718_ & new_n721_;
  assign new_n723_ = ~new_n423_ & ~new_n722_;
  assign new_n724_ = ~new_n291_ & ~new_n723_;
  assign \o[1]  = new_n290_ | new_n724_;
  assign new_n726_ = ~new_n287_ & \o[1] ;
  assign new_n727_ = ~new_n419_ & ~\o[1] ;
  assign \o[0]  = new_n726_ | new_n727_;
  assign new_n729_ = ~new_n436_ & ~\o[1] ;
  assign new_n730_ = ~new_n433_ & \o[1] ;
  assign \o[2]  = new_n729_ | new_n730_;
  assign new_n732_ = ~new_n429_ & ~\o[1] ;
  assign new_n733_ = ~new_n426_ & \o[1] ;
  assign \o[3]  = new_n732_ | new_n733_;
  assign new_n735_ = ~new_n444_ & ~\o[1] ;
  assign new_n736_ = ~new_n441_ & \o[1] ;
  assign \o[4]  = new_n735_ | new_n736_;
  assign new_n738_ = ~new_n454_ & ~\o[1] ;
  assign new_n739_ = ~new_n451_ & \o[1] ;
  assign \o[5]  = new_n738_ | new_n739_;
  assign new_n741_ = ~new_n464_ & ~\o[1] ;
  assign new_n742_ = ~new_n461_ & \o[1] ;
  assign \o[6]  = new_n741_ | new_n742_;
  assign new_n744_ = ~new_n475_ & ~\o[1] ;
  assign new_n745_ = ~new_n472_ & \o[1] ;
  assign \o[7]  = new_n744_ | new_n745_;
  assign new_n747_ = ~new_n484_ & ~\o[1] ;
  assign new_n748_ = ~new_n481_ & \o[1] ;
  assign \o[8]  = new_n747_ | new_n748_;
  assign new_n750_ = ~new_n491_ & ~\o[1] ;
  assign new_n751_ = ~new_n494_ & \o[1] ;
  assign \o[9]  = new_n750_ | new_n751_;
  assign new_n753_ = ~new_n505_ & ~\o[1] ;
  assign new_n754_ = ~new_n502_ & \o[1] ;
  assign \o[10]  = new_n753_ | new_n754_;
  assign new_n756_ = ~new_n515_ & ~\o[1] ;
  assign new_n757_ = ~new_n512_ & \o[1] ;
  assign \o[11]  = new_n756_ | new_n757_;
  assign new_n759_ = ~new_n522_ & ~\o[1] ;
  assign new_n760_ = ~new_n525_ & \o[1] ;
  assign \o[12]  = new_n759_ | new_n760_;
  assign new_n762_ = ~new_n531_ & ~\o[1] ;
  assign new_n763_ = ~new_n534_ & \o[1] ;
  assign \o[13]  = new_n762_ | new_n763_;
  assign new_n765_ = ~new_n544_ & ~\o[1] ;
  assign new_n766_ = ~new_n541_ & \o[1] ;
  assign \o[14]  = new_n765_ | new_n766_;
  assign new_n768_ = ~new_n555_ & ~\o[1] ;
  assign new_n769_ = ~new_n552_ & \o[1] ;
  assign \o[15]  = new_n768_ | new_n769_;
  assign new_n771_ = ~new_n562_ & ~\o[1] ;
  assign new_n772_ = ~new_n565_ & \o[1] ;
  assign \o[16]  = new_n771_ | new_n772_;
  assign new_n774_ = ~new_n571_ & ~\o[1] ;
  assign new_n775_ = ~new_n574_ & \o[1] ;
  assign \o[17]  = new_n774_ | new_n775_;
  assign new_n777_ = ~new_n584_ & ~\o[1] ;
  assign new_n778_ = ~new_n581_ & \o[1] ;
  assign \o[18]  = new_n777_ | new_n778_;
  assign new_n780_ = ~new_n595_ & ~\o[1] ;
  assign new_n781_ = ~new_n592_ & \o[1] ;
  assign \o[19]  = new_n780_ | new_n781_;
  assign new_n783_ = ~new_n602_ & ~\o[1] ;
  assign new_n784_ = ~new_n605_ & \o[1] ;
  assign \o[20]  = new_n783_ | new_n784_;
  assign new_n786_ = ~new_n611_ & ~\o[1] ;
  assign new_n787_ = ~new_n614_ & \o[1] ;
  assign \o[21]  = new_n786_ | new_n787_;
  assign new_n789_ = ~new_n624_ & ~\o[1] ;
  assign new_n790_ = ~new_n621_ & \o[1] ;
  assign \o[22]  = new_n789_ | new_n790_;
  assign new_n792_ = ~new_n635_ & ~\o[1] ;
  assign new_n793_ = ~new_n632_ & \o[1] ;
  assign \o[23]  = new_n792_ | new_n793_;
  assign new_n795_ = ~new_n642_ & ~\o[1] ;
  assign new_n796_ = ~new_n645_ & \o[1] ;
  assign \o[24]  = new_n795_ | new_n796_;
  assign new_n798_ = ~new_n651_ & ~\o[1] ;
  assign new_n799_ = ~new_n654_ & \o[1] ;
  assign \o[25]  = new_n798_ | new_n799_;
  assign new_n801_ = ~new_n664_ & ~\o[1] ;
  assign new_n802_ = ~new_n661_ & \o[1] ;
  assign \o[26]  = new_n801_ | new_n802_;
  assign new_n804_ = ~new_n675_ & ~\o[1] ;
  assign new_n805_ = ~new_n672_ & \o[1] ;
  assign \o[27]  = new_n804_ | new_n805_;
  assign new_n807_ = ~new_n682_ & ~\o[1] ;
  assign new_n808_ = ~new_n685_ & \o[1] ;
  assign \o[28]  = new_n807_ | new_n808_;
  assign new_n810_ = ~new_n691_ & ~\o[1] ;
  assign new_n811_ = ~new_n694_ & \o[1] ;
  assign \o[29]  = new_n810_ | new_n811_;
  assign new_n813_ = ~new_n704_ & ~\o[1] ;
  assign new_n814_ = ~new_n701_ & \o[1] ;
  assign \o[30]  = new_n813_ | new_n814_;
  assign new_n816_ = ~new_n715_ & ~\o[1] ;
  assign new_n817_ = ~new_n712_ & \o[1] ;
  assign \o[31]  = new_n816_ | new_n817_;
  assign new_n819_ = ~new_n422_ & ~\o[1] ;
  assign new_n820_ = ~new_n294_ & \o[1] ;
  assign \o[32]  = new_n819_ | new_n820_;
  assign \o[33]  = ~new_n288_ | ~new_n289_;
endmodule


