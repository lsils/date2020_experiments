module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614;
  assign n65 = x0 & x32;
  assign n68 = ~x32 & x33;
  assign n70 = ~x0 & n68;
  assign n69 = n68 ^ x33;
  assign n71 = n70 ^ n69;
  assign n67 = x1 & x32;
  assign n72 = n71 ^ n67;
  assign n66 = x33 & ~n65;
  assign n73 = n72 ^ n66;
  assign n78 = ~x1 & n68;
  assign n79 = n78 ^ n69;
  assign n77 = x2 & x32;
  assign n80 = n79 ^ n77;
  assign n75 = x34 ^ x33;
  assign n76 = x0 & n75;
  assign n81 = n80 ^ n76;
  assign n74 = n66 & n72;
  assign n82 = n81 ^ n74;
  assign n101 = n76 ^ n74;
  assign n102 = ~n81 & n101;
  assign n103 = n102 ^ n74;
  assign n97 = x1 & n75;
  assign n96 = x35 & n75;
  assign n98 = n97 ^ n96;
  assign n92 = x35 ^ x34;
  assign n93 = ~n75 & n92;
  assign n94 = x35 ^ x0;
  assign n95 = n93 & n94;
  assign n99 = n98 ^ n95;
  assign n88 = ~x2 & n68;
  assign n89 = n88 ^ n69;
  assign n87 = x3 & x32;
  assign n90 = n89 ^ n87;
  assign n83 = x33 ^ x0;
  assign n84 = ~n75 & n83;
  assign n85 = n84 ^ x0;
  assign n86 = x35 & ~n85;
  assign n91 = n90 ^ n86;
  assign n100 = n99 ^ n91;
  assign n104 = n103 ^ n100;
  assign n121 = n103 ^ n99;
  assign n122 = ~n100 & n121;
  assign n123 = n122 ^ n103;
  assign n116 = ~x3 & n68;
  assign n117 = n116 ^ n69;
  assign n115 = x4 & x32;
  assign n118 = n117 ^ n115;
  assign n111 = x2 & n75;
  assign n112 = n111 ^ n96;
  assign n109 = x1 & n93;
  assign n108 = x35 & n93;
  assign n110 = n109 ^ n108;
  assign n113 = n112 ^ n110;
  assign n106 = x36 ^ x35;
  assign n107 = x0 & n106;
  assign n114 = n113 ^ n107;
  assign n119 = n118 ^ n114;
  assign n105 = n86 & n90;
  assign n120 = n119 ^ n105;
  assign n124 = n123 ^ n120;
  assign n153 = n123 ^ n105;
  assign n154 = ~n120 & n153;
  assign n155 = n154 ^ n123;
  assign n148 = n118 ^ n107;
  assign n149 = n118 ^ n113;
  assign n150 = n148 & ~n149;
  assign n151 = n150 ^ n107;
  assign n143 = x1 & n106;
  assign n142 = x37 & n106;
  assign n144 = n143 ^ n142;
  assign n138 = x37 ^ x36;
  assign n139 = ~n106 & n138;
  assign n140 = x37 ^ x0;
  assign n141 = n139 & n140;
  assign n145 = n144 ^ n141;
  assign n135 = x3 & n75;
  assign n136 = n135 ^ n96;
  assign n133 = x2 & n93;
  assign n134 = n133 ^ n108;
  assign n137 = n136 ^ n134;
  assign n146 = n145 ^ n137;
  assign n129 = ~x4 & n68;
  assign n130 = n129 ^ n69;
  assign n128 = x5 & x32;
  assign n131 = n130 ^ n128;
  assign n125 = n94 & ~n106;
  assign n126 = n125 ^ x0;
  assign n127 = x37 & ~n126;
  assign n132 = n131 ^ n127;
  assign n147 = n146 ^ n132;
  assign n152 = n151 ^ n147;
  assign n156 = n155 ^ n152;
  assign n183 = n155 ^ n147;
  assign n184 = ~n152 & n183;
  assign n185 = n184 ^ n155;
  assign n179 = n145 ^ n132;
  assign n180 = n146 & ~n179;
  assign n181 = n180 ^ n137;
  assign n174 = x2 & n106;
  assign n175 = n174 ^ n142;
  assign n172 = x1 & n139;
  assign n171 = x37 & n139;
  assign n173 = n172 ^ n171;
  assign n176 = n175 ^ n173;
  assign n170 = n127 & n131;
  assign n177 = n176 ^ n170;
  assign n166 = x4 & n75;
  assign n167 = n166 ^ n96;
  assign n164 = x3 & n93;
  assign n165 = n164 ^ n108;
  assign n168 = n167 ^ n165;
  assign n160 = ~x5 & n68;
  assign n161 = n160 ^ n69;
  assign n159 = x6 & x32;
  assign n162 = n161 ^ n159;
  assign n157 = x38 ^ x37;
  assign n158 = x0 & n157;
  assign n163 = n162 ^ n158;
  assign n169 = n168 ^ n163;
  assign n178 = n177 ^ n169;
  assign n182 = n181 ^ n178;
  assign n186 = n185 ^ n182;
  assign n224 = n185 ^ n178;
  assign n225 = ~n182 & n224;
  assign n226 = n225 ^ n185;
  assign n220 = n170 ^ n169;
  assign n221 = n177 & ~n220;
  assign n222 = n221 ^ n176;
  assign n215 = n168 ^ n162;
  assign n216 = n163 & ~n215;
  assign n217 = n216 ^ n158;
  assign n211 = ~x6 & n68;
  assign n212 = n211 ^ n69;
  assign n210 = x7 & x32;
  assign n213 = n212 ^ n210;
  assign n207 = n140 & ~n157;
  assign n208 = n207 ^ x0;
  assign n209 = x39 & ~n208;
  assign n214 = n213 ^ n209;
  assign n218 = n217 ^ n214;
  assign n203 = x3 & n106;
  assign n204 = n203 ^ n142;
  assign n201 = x2 & n139;
  assign n202 = n201 ^ n171;
  assign n205 = n204 ^ n202;
  assign n197 = x5 & n75;
  assign n198 = n197 ^ n96;
  assign n195 = x4 & n93;
  assign n196 = n195 ^ n108;
  assign n199 = n198 ^ n196;
  assign n192 = x1 & n157;
  assign n191 = x39 & n157;
  assign n193 = n192 ^ n191;
  assign n187 = x39 ^ x38;
  assign n188 = ~n157 & n187;
  assign n189 = x39 ^ x0;
  assign n190 = n188 & n189;
  assign n194 = n193 ^ n190;
  assign n200 = n199 ^ n194;
  assign n206 = n205 ^ n200;
  assign n219 = n218 ^ n206;
  assign n223 = n222 ^ n219;
  assign n227 = n226 ^ n223;
  assign n266 = n226 ^ n219;
  assign n267 = ~n223 & n266;
  assign n268 = n267 ^ n226;
  assign n261 = n214 ^ n206;
  assign n262 = n217 ^ n206;
  assign n263 = n261 & ~n262;
  assign n264 = n263 ^ n214;
  assign n255 = n205 ^ n194;
  assign n256 = n205 ^ n199;
  assign n257 = n255 & ~n256;
  assign n258 = n257 ^ n194;
  assign n251 = x2 & n157;
  assign n252 = n251 ^ n191;
  assign n249 = x1 & n188;
  assign n248 = x39 & n188;
  assign n250 = n249 ^ n248;
  assign n253 = n252 ^ n250;
  assign n244 = ~x7 & n68;
  assign n245 = n244 ^ n69;
  assign n243 = x8 & x32;
  assign n246 = n245 ^ n243;
  assign n241 = x40 ^ x39;
  assign n242 = x0 & n241;
  assign n247 = n246 ^ n242;
  assign n254 = n253 ^ n247;
  assign n259 = n258 ^ n254;
  assign n236 = x4 & n106;
  assign n237 = n236 ^ n142;
  assign n234 = x3 & n139;
  assign n235 = n234 ^ n171;
  assign n238 = n237 ^ n235;
  assign n231 = x6 & n75;
  assign n232 = n231 ^ n96;
  assign n229 = x5 & n93;
  assign n230 = n229 ^ n108;
  assign n233 = n232 ^ n230;
  assign n239 = n238 ^ n233;
  assign n228 = n209 & n213;
  assign n240 = n239 ^ n228;
  assign n260 = n259 ^ n240;
  assign n265 = n264 ^ n260;
  assign n269 = n268 ^ n265;
  assign n318 = n268 ^ n260;
  assign n319 = ~n265 & n318;
  assign n320 = n319 ^ n268;
  assign n313 = n254 ^ n240;
  assign n314 = n258 ^ n240;
  assign n315 = n313 & ~n314;
  assign n316 = n315 ^ n254;
  assign n308 = n238 ^ n228;
  assign n309 = n239 & ~n308;
  assign n310 = n309 ^ n233;
  assign n304 = ~x8 & n68;
  assign n305 = n304 ^ n69;
  assign n303 = x9 & x32;
  assign n306 = n305 ^ n303;
  assign n299 = x3 & n157;
  assign n300 = n299 ^ n191;
  assign n297 = x2 & n188;
  assign n298 = n297 ^ n248;
  assign n301 = n300 ^ n298;
  assign n294 = x1 & n241;
  assign n293 = x41 & n241;
  assign n295 = n294 ^ n293;
  assign n289 = x41 ^ x40;
  assign n290 = ~n241 & n289;
  assign n291 = x41 ^ x0;
  assign n292 = n290 & n291;
  assign n296 = n295 ^ n292;
  assign n302 = n301 ^ n296;
  assign n307 = n306 ^ n302;
  assign n311 = n310 ^ n307;
  assign n285 = n253 ^ n246;
  assign n286 = n247 & ~n285;
  assign n287 = n286 ^ n242;
  assign n281 = x5 & n106;
  assign n282 = n281 ^ n142;
  assign n279 = x4 & n139;
  assign n280 = n279 ^ n171;
  assign n283 = n282 ^ n280;
  assign n275 = x7 & n75;
  assign n276 = n275 ^ n96;
  assign n273 = x6 & n93;
  assign n274 = n273 ^ n108;
  assign n277 = n276 ^ n274;
  assign n270 = n189 & ~n241;
  assign n271 = n270 ^ x0;
  assign n272 = x41 & ~n271;
  assign n278 = n277 ^ n272;
  assign n284 = n283 ^ n278;
  assign n288 = n287 ^ n284;
  assign n312 = n311 ^ n288;
  assign n317 = n316 ^ n312;
  assign n321 = n320 ^ n317;
  assign n369 = n320 ^ n312;
  assign n370 = ~n317 & n369;
  assign n371 = n370 ^ n320;
  assign n364 = n307 ^ n288;
  assign n365 = n310 ^ n288;
  assign n366 = n364 & ~n365;
  assign n367 = n366 ^ n307;
  assign n359 = n287 ^ n278;
  assign n360 = n284 & ~n359;
  assign n361 = n360 ^ n283;
  assign n355 = x6 & n106;
  assign n356 = n355 ^ n142;
  assign n353 = x5 & n139;
  assign n354 = n353 ^ n171;
  assign n357 = n356 ^ n354;
  assign n349 = ~x9 & n68;
  assign n350 = n349 ^ n69;
  assign n348 = x10 & x32;
  assign n351 = n350 ^ n348;
  assign n345 = x2 & n241;
  assign n346 = n345 ^ n293;
  assign n343 = x1 & n290;
  assign n342 = x41 & n290;
  assign n344 = n343 ^ n342;
  assign n347 = n346 ^ n344;
  assign n352 = n351 ^ n347;
  assign n358 = n357 ^ n352;
  assign n362 = n361 ^ n358;
  assign n337 = n306 ^ n296;
  assign n338 = ~n302 & n337;
  assign n339 = n338 ^ n306;
  assign n336 = n272 & n277;
  assign n340 = n339 ^ n336;
  assign n332 = x4 & n157;
  assign n333 = n332 ^ n191;
  assign n330 = x3 & n188;
  assign n331 = n330 ^ n248;
  assign n334 = n333 ^ n331;
  assign n326 = x8 & n75;
  assign n327 = n326 ^ n96;
  assign n324 = x7 & n93;
  assign n325 = n324 ^ n108;
  assign n328 = n327 ^ n325;
  assign n322 = x42 ^ x41;
  assign n323 = x0 & n322;
  assign n329 = n328 ^ n323;
  assign n335 = n334 ^ n329;
  assign n341 = n340 ^ n335;
  assign n363 = n362 ^ n341;
  assign n368 = n367 ^ n363;
  assign n372 = n371 ^ n368;
  assign n431 = n371 ^ n363;
  assign n432 = ~n368 & n431;
  assign n433 = n432 ^ n371;
  assign n426 = n358 ^ n341;
  assign n427 = n361 ^ n341;
  assign n428 = n426 & ~n427;
  assign n429 = n428 ^ n358;
  assign n422 = n336 ^ n335;
  assign n423 = ~n340 & n422;
  assign n424 = n423 ^ n335;
  assign n416 = ~x10 & n68;
  assign n417 = n416 ^ n69;
  assign n415 = x11 & x32;
  assign n418 = n417 ^ n415;
  assign n411 = x3 & n241;
  assign n412 = n411 ^ n293;
  assign n409 = x2 & n290;
  assign n410 = n409 ^ n342;
  assign n413 = n412 ^ n410;
  assign n406 = x5 & n157;
  assign n407 = n406 ^ n191;
  assign n404 = x4 & n188;
  assign n405 = n404 ^ n248;
  assign n408 = n407 ^ n405;
  assign n414 = n413 ^ n408;
  assign n419 = n418 ^ n414;
  assign n400 = n334 ^ n328;
  assign n401 = n329 & ~n400;
  assign n402 = n401 ^ n323;
  assign n397 = n357 ^ n347;
  assign n398 = n352 & ~n397;
  assign n399 = n398 ^ n351;
  assign n403 = n402 ^ n399;
  assign n420 = n419 ^ n403;
  assign n392 = x9 & n75;
  assign n393 = n392 ^ n96;
  assign n390 = x8 & n93;
  assign n391 = n390 ^ n108;
  assign n394 = n393 ^ n391;
  assign n387 = n291 & ~n322;
  assign n388 = n387 ^ x0;
  assign n389 = x43 & ~n388;
  assign n395 = n394 ^ n389;
  assign n383 = ~x1 & n322;
  assign n382 = ~x43 & n322;
  assign n384 = n383 ^ n382;
  assign n378 = x43 ^ x42;
  assign n379 = ~n322 & n378;
  assign n380 = x43 ^ x0;
  assign n381 = n379 & n380;
  assign n385 = n384 ^ n381;
  assign n375 = x7 & n106;
  assign n376 = n375 ^ n142;
  assign n373 = x6 & n139;
  assign n374 = n373 ^ n171;
  assign n377 = n376 ^ n374;
  assign n386 = n385 ^ n377;
  assign n396 = n395 ^ n386;
  assign n421 = n420 ^ n396;
  assign n425 = n424 ^ n421;
  assign n430 = n429 ^ n425;
  assign n434 = n433 ^ n430;
  assign n491 = n433 ^ n425;
  assign n492 = ~n430 & n491;
  assign n493 = n492 ^ n433;
  assign n487 = n424 ^ n420;
  assign n488 = n421 & ~n487;
  assign n489 = n488 ^ n396;
  assign n482 = n419 ^ n399;
  assign n483 = ~n403 & n482;
  assign n484 = n483 ^ n419;
  assign n478 = n418 ^ n408;
  assign n479 = ~n414 & n478;
  assign n480 = n479 ^ n418;
  assign n474 = x8 & n106;
  assign n475 = n474 ^ n142;
  assign n472 = x7 & n139;
  assign n473 = n472 ^ n171;
  assign n476 = n475 ^ n473;
  assign n471 = n389 & n394;
  assign n477 = n476 ^ n471;
  assign n481 = n480 ^ n477;
  assign n485 = n484 ^ n481;
  assign n467 = n395 ^ n385;
  assign n468 = n386 & ~n467;
  assign n469 = n468 ^ n377;
  assign n462 = ~x2 & n322;
  assign n463 = n462 ^ n382;
  assign n460 = ~x1 & n379;
  assign n459 = ~x43 & n379;
  assign n461 = n460 ^ n459;
  assign n464 = n463 ^ n461;
  assign n455 = ~x11 & n68;
  assign n456 = n455 ^ n69;
  assign n454 = x12 & x32;
  assign n457 = n456 ^ n454;
  assign n451 = x4 & n241;
  assign n452 = n451 ^ n293;
  assign n449 = x3 & n290;
  assign n450 = n449 ^ n342;
  assign n453 = n452 ^ n450;
  assign n458 = n457 ^ n453;
  assign n465 = n464 ^ n458;
  assign n445 = x6 & n157;
  assign n446 = n445 ^ n191;
  assign n443 = x5 & n188;
  assign n444 = n443 ^ n248;
  assign n447 = n446 ^ n444;
  assign n439 = x10 & n75;
  assign n440 = n439 ^ n96;
  assign n437 = x9 & n93;
  assign n438 = n437 ^ n108;
  assign n441 = n440 ^ n438;
  assign n435 = x44 ^ x43;
  assign n436 = x0 & n435;
  assign n442 = n441 ^ n436;
  assign n448 = n447 ^ n442;
  assign n466 = n465 ^ n448;
  assign n470 = n469 ^ n466;
  assign n486 = n485 ^ n470;
  assign n490 = n489 ^ n486;
  assign n494 = n493 ^ n490;
  assign n563 = n493 ^ n486;
  assign n564 = ~n490 & n563;
  assign n565 = n564 ^ n493;
  assign n559 = n481 ^ n470;
  assign n560 = ~n485 & n559;
  assign n561 = n560 ^ n470;
  assign n554 = n469 ^ n465;
  assign n555 = n466 & ~n554;
  assign n556 = n555 ^ n448;
  assign n550 = n464 ^ n453;
  assign n551 = n458 & ~n550;
  assign n552 = n551 ^ n457;
  assign n545 = n447 ^ n436;
  assign n546 = n447 ^ n441;
  assign n547 = n545 & ~n546;
  assign n548 = n547 ^ n436;
  assign n541 = ~x12 & n68;
  assign n542 = n541 ^ n69;
  assign n540 = x13 & x32;
  assign n543 = n542 ^ n540;
  assign n537 = n380 & ~n435;
  assign n538 = n537 ^ x0;
  assign n539 = x45 & ~n538;
  assign n544 = n543 ^ n539;
  assign n549 = n548 ^ n544;
  assign n553 = n552 ^ n549;
  assign n557 = n556 ^ n553;
  assign n533 = n480 ^ n471;
  assign n534 = n477 & ~n533;
  assign n535 = n534 ^ n476;
  assign n528 = x1 & n435;
  assign n527 = x45 & n435;
  assign n529 = n528 ^ n527;
  assign n523 = x45 ^ x44;
  assign n524 = ~n435 & n523;
  assign n525 = x45 ^ x0;
  assign n526 = n524 & n525;
  assign n530 = n529 ^ n526;
  assign n519 = ~x3 & n322;
  assign n520 = n519 ^ n382;
  assign n517 = ~x2 & n379;
  assign n518 = n517 ^ n459;
  assign n521 = n520 ^ n518;
  assign n514 = x9 & n106;
  assign n515 = n514 ^ n142;
  assign n512 = x8 & n139;
  assign n513 = n512 ^ n171;
  assign n516 = n515 ^ n513;
  assign n522 = n521 ^ n516;
  assign n531 = n530 ^ n522;
  assign n508 = x5 & n241;
  assign n509 = n508 ^ n293;
  assign n506 = x4 & n290;
  assign n507 = n506 ^ n342;
  assign n510 = n509 ^ n507;
  assign n502 = x11 & n75;
  assign n503 = n502 ^ n96;
  assign n500 = x10 & n93;
  assign n501 = n500 ^ n108;
  assign n504 = n503 ^ n501;
  assign n497 = x7 & n157;
  assign n498 = n497 ^ n191;
  assign n495 = x6 & n188;
  assign n496 = n495 ^ n248;
  assign n499 = n498 ^ n496;
  assign n505 = n504 ^ n499;
  assign n511 = n510 ^ n505;
  assign n532 = n531 ^ n511;
  assign n536 = n535 ^ n532;
  assign n558 = n557 ^ n536;
  assign n562 = n561 ^ n558;
  assign n566 = n565 ^ n562;
  assign n633 = n565 ^ n558;
  assign n634 = ~n562 & n633;
  assign n635 = n634 ^ n565;
  assign n629 = n556 ^ n536;
  assign n630 = n557 & ~n629;
  assign n631 = n630 ^ n553;
  assign n625 = n535 ^ n531;
  assign n626 = n532 & ~n625;
  assign n627 = n626 ^ n511;
  assign n620 = n552 ^ n548;
  assign n621 = n549 & ~n620;
  assign n622 = n621 ^ n544;
  assign n614 = x2 & n435;
  assign n615 = n614 ^ n527;
  assign n612 = x1 & n524;
  assign n611 = x45 & n524;
  assign n613 = n612 ^ n611;
  assign n616 = n615 ^ n613;
  assign n608 = ~x4 & n322;
  assign n609 = n608 ^ n382;
  assign n606 = ~x3 & n379;
  assign n607 = n606 ^ n459;
  assign n610 = n609 ^ n607;
  assign n617 = n616 ^ n610;
  assign n605 = n539 & n543;
  assign n618 = n617 ^ n605;
  assign n601 = x10 & n106;
  assign n602 = n601 ^ n142;
  assign n599 = x9 & n139;
  assign n600 = n599 ^ n171;
  assign n603 = n602 ^ n600;
  assign n595 = x6 & n241;
  assign n596 = n595 ^ n293;
  assign n593 = x5 & n290;
  assign n594 = n593 ^ n342;
  assign n597 = n596 ^ n594;
  assign n590 = x8 & n157;
  assign n591 = n590 ^ n191;
  assign n588 = x7 & n188;
  assign n589 = n588 ^ n248;
  assign n592 = n591 ^ n589;
  assign n598 = n597 ^ n592;
  assign n604 = n603 ^ n598;
  assign n619 = n618 ^ n604;
  assign n623 = n622 ^ n619;
  assign n583 = n530 ^ n521;
  assign n584 = n522 & ~n583;
  assign n585 = n584 ^ n516;
  assign n580 = n510 ^ n504;
  assign n581 = n505 & ~n580;
  assign n582 = n581 ^ n499;
  assign n586 = n585 ^ n582;
  assign n576 = x12 & n75;
  assign n577 = n576 ^ n96;
  assign n574 = x11 & n93;
  assign n575 = n574 ^ n108;
  assign n578 = n577 ^ n575;
  assign n570 = ~x13 & n68;
  assign n571 = n570 ^ n69;
  assign n569 = x14 & x32;
  assign n572 = n571 ^ n569;
  assign n567 = x46 ^ x45;
  assign n568 = x0 & n567;
  assign n573 = n572 ^ n568;
  assign n579 = n578 ^ n573;
  assign n587 = n586 ^ n579;
  assign n624 = n623 ^ n587;
  assign n628 = n627 ^ n624;
  assign n632 = n631 ^ n628;
  assign n636 = n635 ^ n632;
  assign n715 = n635 ^ n628;
  assign n716 = ~n632 & n715;
  assign n717 = n716 ^ n635;
  assign n711 = n627 ^ n623;
  assign n712 = n624 & ~n711;
  assign n713 = n712 ^ n587;
  assign n706 = n622 ^ n618;
  assign n707 = n619 & ~n706;
  assign n708 = n707 ^ n604;
  assign n700 = n603 ^ n592;
  assign n701 = n603 ^ n597;
  assign n702 = n700 & ~n701;
  assign n703 = n702 ^ n592;
  assign n696 = ~x5 & n322;
  assign n697 = n696 ^ n382;
  assign n694 = ~x4 & n379;
  assign n695 = n694 ^ n459;
  assign n698 = n697 ^ n695;
  assign n690 = x11 & n106;
  assign n691 = n690 ^ n142;
  assign n688 = x10 & n139;
  assign n689 = n688 ^ n171;
  assign n692 = n691 ^ n689;
  assign n685 = x7 & n241;
  assign n686 = n685 ^ n293;
  assign n683 = x6 & n290;
  assign n684 = n683 ^ n342;
  assign n687 = n686 ^ n684;
  assign n693 = n692 ^ n687;
  assign n699 = n698 ^ n693;
  assign n704 = n703 ^ n699;
  assign n679 = x9 & n157;
  assign n680 = n679 ^ n191;
  assign n677 = x8 & n188;
  assign n678 = n677 ^ n248;
  assign n681 = n680 ^ n678;
  assign n673 = ~x1 & n567;
  assign n672 = ~x47 & n567;
  assign n674 = n673 ^ n672;
  assign n668 = x47 ^ x46;
  assign n669 = ~n567 & n668;
  assign n670 = x47 ^ x0;
  assign n671 = n669 & n670;
  assign n675 = n674 ^ n671;
  assign n665 = x13 & n75;
  assign n666 = n665 ^ n96;
  assign n663 = x12 & n93;
  assign n664 = n663 ^ n108;
  assign n667 = n666 ^ n664;
  assign n676 = n675 ^ n667;
  assign n682 = n681 ^ n676;
  assign n705 = n704 ^ n682;
  assign n709 = n708 ^ n705;
  assign n659 = n582 ^ n579;
  assign n660 = ~n586 & n659;
  assign n661 = n660 ^ n579;
  assign n655 = n616 ^ n605;
  assign n656 = n617 & ~n655;
  assign n657 = n656 ^ n610;
  assign n651 = n578 ^ n572;
  assign n652 = n573 & ~n651;
  assign n653 = n652 ^ n568;
  assign n647 = x3 & n435;
  assign n648 = n647 ^ n527;
  assign n645 = x2 & n524;
  assign n646 = n645 ^ n611;
  assign n649 = n648 ^ n646;
  assign n641 = ~x14 & n68;
  assign n642 = n641 ^ n69;
  assign n640 = x15 & x32;
  assign n643 = n642 ^ n640;
  assign n637 = n525 & ~n567;
  assign n638 = n637 ^ x0;
  assign n639 = x47 & ~n638;
  assign n644 = n643 ^ n639;
  assign n650 = n649 ^ n644;
  assign n654 = n653 ^ n650;
  assign n658 = n657 ^ n654;
  assign n662 = n661 ^ n658;
  assign n710 = n709 ^ n662;
  assign n714 = n713 ^ n710;
  assign n718 = n717 ^ n714;
  assign n798 = n717 ^ n710;
  assign n799 = ~n714 & n798;
  assign n800 = n799 ^ n717;
  assign n793 = n705 ^ n662;
  assign n794 = n708 ^ n662;
  assign n795 = n793 & ~n794;
  assign n796 = n795 ^ n705;
  assign n788 = n661 ^ n657;
  assign n789 = n658 & ~n788;
  assign n790 = n789 ^ n654;
  assign n782 = x4 & n435;
  assign n783 = n782 ^ n527;
  assign n780 = x3 & n524;
  assign n781 = n780 ^ n611;
  assign n784 = n783 ^ n781;
  assign n776 = ~x6 & n322;
  assign n777 = n776 ^ n382;
  assign n774 = ~x5 & n379;
  assign n775 = n774 ^ n459;
  assign n778 = n777 ^ n775;
  assign n771 = x12 & n106;
  assign n772 = n771 ^ n142;
  assign n769 = x11 & n139;
  assign n770 = n769 ^ n171;
  assign n773 = n772 ^ n770;
  assign n779 = n778 ^ n773;
  assign n785 = n784 ^ n779;
  assign n765 = x14 & n75;
  assign n766 = n765 ^ n96;
  assign n763 = x13 & n93;
  assign n764 = n763 ^ n108;
  assign n767 = n766 ^ n764;
  assign n759 = ~x15 & n68;
  assign n760 = n759 ^ n69;
  assign n758 = x16 & x32;
  assign n761 = n760 ^ n758;
  assign n756 = x48 ^ x47;
  assign n757 = x0 & n756;
  assign n762 = n761 ^ n757;
  assign n768 = n767 ^ n762;
  assign n786 = n785 ^ n768;
  assign n752 = x8 & n241;
  assign n753 = n752 ^ n293;
  assign n750 = x7 & n290;
  assign n751 = n750 ^ n342;
  assign n754 = n753 ^ n751;
  assign n746 = x10 & n157;
  assign n747 = n746 ^ n191;
  assign n744 = x9 & n188;
  assign n745 = n744 ^ n248;
  assign n748 = n747 ^ n745;
  assign n741 = ~x2 & n567;
  assign n742 = n741 ^ n672;
  assign n739 = ~x1 & n669;
  assign n738 = ~x47 & n669;
  assign n740 = n739 ^ n738;
  assign n743 = n742 ^ n740;
  assign n749 = n748 ^ n743;
  assign n755 = n754 ^ n749;
  assign n787 = n786 ^ n755;
  assign n791 = n790 ^ n787;
  assign n733 = n699 ^ n682;
  assign n734 = n703 ^ n682;
  assign n735 = n733 & ~n734;
  assign n736 = n735 ^ n699;
  assign n729 = n653 ^ n644;
  assign n730 = n650 & ~n729;
  assign n731 = n730 ^ n649;
  assign n724 = n698 ^ n687;
  assign n725 = n698 ^ n692;
  assign n726 = n724 & ~n725;
  assign n727 = n726 ^ n687;
  assign n720 = n681 ^ n675;
  assign n721 = n676 & ~n720;
  assign n722 = n721 ^ n667;
  assign n719 = n639 & n643;
  assign n723 = n722 ^ n719;
  assign n728 = n727 ^ n723;
  assign n732 = n731 ^ n728;
  assign n737 = n736 ^ n732;
  assign n792 = n791 ^ n737;
  assign n797 = n796 ^ n792;
  assign n801 = n800 ^ n797;
  assign n890 = n800 ^ n792;
  assign n891 = ~n797 & n890;
  assign n892 = n891 ^ n800;
  assign n885 = n787 ^ n737;
  assign n886 = n790 ^ n737;
  assign n887 = n885 & ~n886;
  assign n888 = n887 ^ n787;
  assign n880 = n736 ^ n731;
  assign n881 = n732 & ~n880;
  assign n882 = n881 ^ n728;
  assign n874 = x1 & n756;
  assign n873 = x49 & n756;
  assign n875 = n874 ^ n873;
  assign n869 = x49 ^ x48;
  assign n870 = ~n756 & n869;
  assign n871 = x49 ^ x0;
  assign n872 = n870 & n871;
  assign n876 = n875 ^ n872;
  assign n865 = x11 & n157;
  assign n866 = n865 ^ n191;
  assign n863 = x10 & n188;
  assign n864 = n863 ^ n248;
  assign n867 = n866 ^ n864;
  assign n860 = ~x3 & n567;
  assign n861 = n860 ^ n672;
  assign n858 = ~x2 & n669;
  assign n859 = n858 ^ n738;
  assign n862 = n861 ^ n859;
  assign n868 = n867 ^ n862;
  assign n877 = n876 ^ n868;
  assign n854 = x13 & n106;
  assign n855 = n854 ^ n142;
  assign n852 = x12 & n139;
  assign n853 = n852 ^ n171;
  assign n856 = n855 ^ n853;
  assign n848 = x9 & n241;
  assign n849 = n848 ^ n293;
  assign n846 = x8 & n290;
  assign n847 = n846 ^ n342;
  assign n850 = n849 ^ n847;
  assign n843 = x15 & n75;
  assign n844 = n843 ^ n96;
  assign n841 = x14 & n93;
  assign n842 = n841 ^ n108;
  assign n845 = n844 ^ n842;
  assign n851 = n850 ^ n845;
  assign n857 = n856 ^ n851;
  assign n878 = n877 ^ n857;
  assign n836 = ~x7 & n322;
  assign n837 = n836 ^ n382;
  assign n834 = ~x6 & n379;
  assign n835 = n834 ^ n459;
  assign n838 = n837 ^ n835;
  assign n831 = x5 & n435;
  assign n832 = n831 ^ n527;
  assign n829 = x4 & n524;
  assign n830 = n829 ^ n611;
  assign n833 = n832 ^ n830;
  assign n839 = n838 ^ n833;
  assign n825 = ~x16 & n68;
  assign n826 = n825 ^ n69;
  assign n824 = x17 & x32;
  assign n827 = n826 ^ n824;
  assign n821 = n670 & ~n756;
  assign n822 = n821 ^ x0;
  assign n823 = x49 & ~n822;
  assign n828 = n827 ^ n823;
  assign n840 = n839 ^ n828;
  assign n879 = n878 ^ n840;
  assign n883 = n882 ^ n879;
  assign n817 = n785 ^ n755;
  assign n818 = n786 & ~n817;
  assign n819 = n818 ^ n768;
  assign n813 = n727 ^ n722;
  assign n814 = n723 & ~n813;
  assign n815 = n814 ^ n719;
  assign n809 = n754 ^ n748;
  assign n810 = n749 & ~n809;
  assign n811 = n810 ^ n743;
  assign n805 = n784 ^ n773;
  assign n806 = ~n779 & n805;
  assign n807 = n806 ^ n784;
  assign n802 = n767 ^ n761;
  assign n803 = n762 & ~n802;
  assign n804 = n803 ^ n757;
  assign n808 = n807 ^ n804;
  assign n812 = n811 ^ n808;
  assign n816 = n815 ^ n812;
  assign n820 = n819 ^ n816;
  assign n884 = n883 ^ n820;
  assign n889 = n888 ^ n884;
  assign n893 = n892 ^ n889;
  assign n981 = n892 ^ n884;
  assign n982 = ~n889 & n981;
  assign n983 = n982 ^ n892;
  assign n976 = n879 ^ n820;
  assign n977 = n882 ^ n820;
  assign n978 = n976 & ~n977;
  assign n979 = n978 ^ n879;
  assign n971 = n819 ^ n812;
  assign n972 = ~n816 & n971;
  assign n973 = n972 ^ n819;
  assign n966 = n838 ^ n828;
  assign n967 = n839 & ~n966;
  assign n968 = n967 ^ n833;
  assign n962 = x16 & n75;
  assign n963 = n962 ^ n96;
  assign n960 = x15 & n93;
  assign n961 = n960 ^ n108;
  assign n964 = n963 ^ n961;
  assign n956 = x2 & n756;
  assign n957 = n956 ^ n873;
  assign n954 = x1 & n870;
  assign n953 = x49 & n870;
  assign n955 = n954 ^ n953;
  assign n958 = n957 ^ n955;
  assign n950 = ~x4 & n567;
  assign n951 = n950 ^ n672;
  assign n948 = ~x3 & n669;
  assign n949 = n948 ^ n738;
  assign n952 = n951 ^ n949;
  assign n959 = n958 ^ n952;
  assign n965 = n964 ^ n959;
  assign n969 = n968 ^ n965;
  assign n944 = n876 ^ n862;
  assign n945 = ~n868 & n944;
  assign n946 = n945 ^ n876;
  assign n940 = x6 & n435;
  assign n941 = n940 ^ n527;
  assign n938 = x5 & n524;
  assign n939 = n938 ^ n611;
  assign n942 = n941 ^ n939;
  assign n937 = n823 & n827;
  assign n943 = n942 ^ n937;
  assign n947 = n946 ^ n943;
  assign n970 = n969 ^ n947;
  assign n974 = n973 ^ n970;
  assign n932 = n811 ^ n807;
  assign n933 = n808 & ~n932;
  assign n934 = n933 ^ n804;
  assign n929 = n857 ^ n840;
  assign n930 = ~n878 & n929;
  assign n931 = n930 ^ n840;
  assign n935 = n934 ^ n931;
  assign n924 = n856 ^ n850;
  assign n925 = n851 & ~n924;
  assign n926 = n925 ^ n845;
  assign n920 = ~x8 & n322;
  assign n921 = n920 ^ n382;
  assign n918 = ~x7 & n379;
  assign n919 = n918 ^ n459;
  assign n922 = n921 ^ n919;
  assign n914 = x14 & n106;
  assign n915 = n914 ^ n142;
  assign n912 = x13 & n139;
  assign n913 = n912 ^ n171;
  assign n916 = n915 ^ n913;
  assign n909 = x10 & n241;
  assign n910 = n909 ^ n293;
  assign n907 = x9 & n290;
  assign n908 = n907 ^ n342;
  assign n911 = n910 ^ n908;
  assign n917 = n916 ^ n911;
  assign n923 = n922 ^ n917;
  assign n927 = n926 ^ n923;
  assign n903 = x12 & n157;
  assign n904 = n903 ^ n191;
  assign n901 = x11 & n188;
  assign n902 = n901 ^ n248;
  assign n905 = n904 ^ n902;
  assign n897 = ~x17 & n68;
  assign n898 = n897 ^ n69;
  assign n896 = x18 & x32;
  assign n899 = n898 ^ n896;
  assign n894 = x50 ^ x49;
  assign n895 = x0 & n894;
  assign n900 = n899 ^ n895;
  assign n906 = n905 ^ n900;
  assign n928 = n927 ^ n906;
  assign n936 = n935 ^ n928;
  assign n975 = n974 ^ n936;
  assign n980 = n979 ^ n975;
  assign n984 = n983 ^ n980;
  assign n1083 = n983 ^ n975;
  assign n1084 = ~n980 & n1083;
  assign n1085 = n1084 ^ n983;
  assign n1078 = n970 ^ n936;
  assign n1079 = n973 ^ n936;
  assign n1080 = n1078 & ~n1079;
  assign n1081 = n1080 ^ n970;
  assign n1073 = n931 ^ n928;
  assign n1074 = ~n935 & n1073;
  assign n1075 = n1074 ^ n928;
  assign n1068 = n946 ^ n937;
  assign n1069 = n943 & ~n1068;
  assign n1070 = n1069 ^ n942;
  assign n1064 = x11 & n241;
  assign n1065 = n1064 ^ n293;
  assign n1062 = x10 & n290;
  assign n1063 = n1062 ^ n342;
  assign n1066 = n1065 ^ n1063;
  assign n1058 = x17 & n75;
  assign n1059 = n1058 ^ n96;
  assign n1056 = x16 & n93;
  assign n1057 = n1056 ^ n108;
  assign n1060 = n1059 ^ n1057;
  assign n1053 = ~x1 & n894;
  assign n1052 = ~x51 & n894;
  assign n1054 = n1053 ^ n1052;
  assign n1048 = x51 ^ x50;
  assign n1049 = ~n894 & n1048;
  assign n1050 = x51 ^ x0;
  assign n1051 = n1049 & n1050;
  assign n1055 = n1054 ^ n1051;
  assign n1061 = n1060 ^ n1055;
  assign n1067 = n1066 ^ n1061;
  assign n1071 = n1070 ^ n1067;
  assign n1044 = n964 ^ n952;
  assign n1045 = ~n959 & n1044;
  assign n1046 = n1045 ^ n964;
  assign n1040 = n905 ^ n899;
  assign n1041 = n900 & ~n1040;
  assign n1042 = n1041 ^ n895;
  assign n1036 = ~x18 & n68;
  assign n1037 = n1036 ^ n69;
  assign n1035 = x19 & x32;
  assign n1038 = n1037 ^ n1035;
  assign n1032 = n871 & ~n894;
  assign n1033 = n1032 ^ x0;
  assign n1034 = x51 & ~n1033;
  assign n1039 = n1038 ^ n1034;
  assign n1043 = n1042 ^ n1039;
  assign n1047 = n1046 ^ n1043;
  assign n1072 = n1071 ^ n1047;
  assign n1076 = n1075 ^ n1072;
  assign n1028 = n968 ^ n947;
  assign n1029 = n969 & ~n1028;
  assign n1030 = n1029 ^ n965;
  assign n1024 = n923 ^ n906;
  assign n1025 = ~n927 & n1024;
  assign n1026 = n1025 ^ n906;
  assign n1019 = n922 ^ n911;
  assign n1020 = ~n917 & n1019;
  assign n1021 = n1020 ^ n922;
  assign n1015 = x7 & n435;
  assign n1016 = n1015 ^ n527;
  assign n1013 = x6 & n524;
  assign n1014 = n1013 ^ n611;
  assign n1017 = n1016 ^ n1014;
  assign n1009 = ~x9 & n322;
  assign n1010 = n1009 ^ n382;
  assign n1007 = ~x8 & n379;
  assign n1008 = n1007 ^ n459;
  assign n1011 = n1010 ^ n1008;
  assign n1004 = x15 & n106;
  assign n1005 = n1004 ^ n142;
  assign n1002 = x14 & n139;
  assign n1003 = n1002 ^ n171;
  assign n1006 = n1005 ^ n1003;
  assign n1012 = n1011 ^ n1006;
  assign n1018 = n1017 ^ n1012;
  assign n1022 = n1021 ^ n1018;
  assign n998 = x3 & n756;
  assign n999 = n998 ^ n873;
  assign n996 = x2 & n870;
  assign n997 = n996 ^ n953;
  assign n1000 = n999 ^ n997;
  assign n992 = ~x5 & n567;
  assign n993 = n992 ^ n672;
  assign n990 = ~x4 & n669;
  assign n991 = n990 ^ n738;
  assign n994 = n993 ^ n991;
  assign n987 = x13 & n157;
  assign n988 = n987 ^ n191;
  assign n985 = x12 & n188;
  assign n986 = n985 ^ n248;
  assign n989 = n988 ^ n986;
  assign n995 = n994 ^ n989;
  assign n1001 = n1000 ^ n995;
  assign n1023 = n1022 ^ n1001;
  assign n1027 = n1026 ^ n1023;
  assign n1031 = n1030 ^ n1027;
  assign n1077 = n1076 ^ n1031;
  assign n1082 = n1081 ^ n1077;
  assign n1086 = n1085 ^ n1082;
  assign n1187 = n1085 ^ n1077;
  assign n1188 = ~n1082 & n1187;
  assign n1189 = n1188 ^ n1085;
  assign n1182 = n1072 ^ n1031;
  assign n1183 = n1075 ^ n1031;
  assign n1184 = n1182 & ~n1183;
  assign n1185 = n1184 ^ n1072;
  assign n1176 = n1030 ^ n1023;
  assign n1177 = n1030 ^ n1026;
  assign n1178 = n1176 & ~n1177;
  assign n1179 = n1178 ^ n1023;
  assign n1172 = n1067 ^ n1047;
  assign n1173 = n1070 ^ n1047;
  assign n1174 = n1172 & ~n1173;
  assign n1175 = n1174 ^ n1067;
  assign n1180 = n1179 ^ n1175;
  assign n1166 = n1018 ^ n1001;
  assign n1167 = n1021 ^ n1001;
  assign n1168 = n1166 & ~n1167;
  assign n1169 = n1168 ^ n1018;
  assign n1162 = n1046 ^ n1042;
  assign n1163 = n1043 & ~n1162;
  assign n1164 = n1163 ^ n1039;
  assign n1157 = x8 & n435;
  assign n1158 = n1157 ^ n527;
  assign n1155 = x7 & n524;
  assign n1156 = n1155 ^ n611;
  assign n1159 = n1158 ^ n1156;
  assign n1152 = ~x10 & n322;
  assign n1153 = n1152 ^ n382;
  assign n1150 = ~x9 & n379;
  assign n1151 = n1150 ^ n459;
  assign n1154 = n1153 ^ n1151;
  assign n1160 = n1159 ^ n1154;
  assign n1149 = n1034 & n1038;
  assign n1161 = n1160 ^ n1149;
  assign n1165 = n1164 ^ n1161;
  assign n1170 = n1169 ^ n1165;
  assign n1144 = n1066 ^ n1055;
  assign n1145 = ~n1061 & n1144;
  assign n1146 = n1145 ^ n1066;
  assign n1140 = n1000 ^ n994;
  assign n1141 = n995 & ~n1140;
  assign n1142 = n1141 ^ n989;
  assign n1137 = n1017 ^ n1011;
  assign n1138 = n1012 & ~n1137;
  assign n1139 = n1138 ^ n1006;
  assign n1143 = n1142 ^ n1139;
  assign n1147 = n1146 ^ n1143;
  assign n1131 = x18 & n75;
  assign n1132 = n1131 ^ n96;
  assign n1129 = x17 & n93;
  assign n1130 = n1129 ^ n108;
  assign n1133 = n1132 ^ n1130;
  assign n1125 = ~x6 & n567;
  assign n1126 = n1125 ^ n672;
  assign n1123 = ~x5 & n669;
  assign n1124 = n1123 ^ n738;
  assign n1127 = n1126 ^ n1124;
  assign n1120 = x4 & n756;
  assign n1121 = n1120 ^ n873;
  assign n1118 = x3 & n870;
  assign n1119 = n1118 ^ n953;
  assign n1122 = n1121 ^ n1119;
  assign n1128 = n1127 ^ n1122;
  assign n1134 = n1133 ^ n1128;
  assign n1114 = x14 & n157;
  assign n1115 = n1114 ^ n191;
  assign n1112 = x13 & n188;
  assign n1113 = n1112 ^ n248;
  assign n1116 = n1115 ^ n1113;
  assign n1108 = ~x19 & n68;
  assign n1109 = n1108 ^ n69;
  assign n1107 = x20 & x32;
  assign n1110 = n1109 ^ n1107;
  assign n1105 = x52 ^ x51;
  assign n1106 = x0 & n1105;
  assign n1111 = n1110 ^ n1106;
  assign n1117 = n1116 ^ n1111;
  assign n1135 = n1134 ^ n1117;
  assign n1101 = x16 & n106;
  assign n1102 = n1101 ^ n142;
  assign n1099 = x15 & n139;
  assign n1100 = n1099 ^ n171;
  assign n1103 = n1102 ^ n1100;
  assign n1095 = x12 & n241;
  assign n1096 = n1095 ^ n293;
  assign n1093 = x11 & n290;
  assign n1094 = n1093 ^ n342;
  assign n1097 = n1096 ^ n1094;
  assign n1090 = ~x2 & n894;
  assign n1091 = n1090 ^ n1052;
  assign n1088 = ~x1 & n1049;
  assign n1087 = ~x51 & n1049;
  assign n1089 = n1088 ^ n1087;
  assign n1092 = n1091 ^ n1089;
  assign n1098 = n1097 ^ n1092;
  assign n1104 = n1103 ^ n1098;
  assign n1136 = n1135 ^ n1104;
  assign n1148 = n1147 ^ n1136;
  assign n1171 = n1170 ^ n1148;
  assign n1181 = n1180 ^ n1171;
  assign n1186 = n1185 ^ n1181;
  assign n1190 = n1189 ^ n1186;
  assign n1300 = n1189 ^ n1181;
  assign n1301 = ~n1186 & n1300;
  assign n1302 = n1301 ^ n1189;
  assign n1296 = n1175 ^ n1171;
  assign n1297 = ~n1180 & n1296;
  assign n1298 = n1297 ^ n1171;
  assign n1292 = n1170 ^ n1147;
  assign n1293 = n1148 & ~n1292;
  assign n1294 = n1293 ^ n1136;
  assign n1287 = n1169 ^ n1161;
  assign n1288 = n1169 ^ n1164;
  assign n1289 = n1287 & ~n1288;
  assign n1290 = n1289 ^ n1161;
  assign n1281 = n1146 ^ n1142;
  assign n1282 = n1143 & ~n1281;
  assign n1283 = n1282 ^ n1139;
  assign n1276 = n1133 ^ n1122;
  assign n1277 = n1133 ^ n1127;
  assign n1278 = n1276 & ~n1277;
  assign n1279 = n1278 ^ n1122;
  assign n1272 = x9 & n435;
  assign n1273 = n1272 ^ n527;
  assign n1270 = x8 & n524;
  assign n1271 = n1270 ^ n611;
  assign n1274 = n1273 ^ n1271;
  assign n1266 = x19 & n75;
  assign n1267 = n1266 ^ n96;
  assign n1264 = x18 & n93;
  assign n1265 = n1264 ^ n108;
  assign n1268 = n1267 ^ n1265;
  assign n1261 = n1050 & ~n1105;
  assign n1262 = n1261 ^ x0;
  assign n1263 = x53 & ~n1262;
  assign n1269 = n1268 ^ n1263;
  assign n1275 = n1274 ^ n1269;
  assign n1280 = n1279 ^ n1275;
  assign n1284 = n1283 ^ n1280;
  assign n1256 = n1103 ^ n1097;
  assign n1257 = n1098 & ~n1256;
  assign n1258 = n1257 ^ n1092;
  assign n1253 = n1116 ^ n1110;
  assign n1254 = n1111 & ~n1253;
  assign n1255 = n1254 ^ n1106;
  assign n1259 = n1258 ^ n1255;
  assign n1249 = ~x11 & n322;
  assign n1250 = n1249 ^ n382;
  assign n1247 = ~x10 & n379;
  assign n1248 = n1247 ^ n459;
  assign n1251 = n1250 ^ n1248;
  assign n1243 = ~x20 & n68;
  assign n1244 = n1243 ^ n69;
  assign n1242 = x21 & x32;
  assign n1245 = n1244 ^ n1242;
  assign n1239 = x17 & n106;
  assign n1240 = n1239 ^ n142;
  assign n1237 = x16 & n139;
  assign n1238 = n1237 ^ n171;
  assign n1241 = n1240 ^ n1238;
  assign n1246 = n1245 ^ n1241;
  assign n1252 = n1251 ^ n1246;
  assign n1260 = n1259 ^ n1252;
  assign n1285 = n1284 ^ n1260;
  assign n1233 = n1134 ^ n1104;
  assign n1234 = n1135 & ~n1233;
  assign n1235 = n1234 ^ n1117;
  assign n1229 = n1159 ^ n1149;
  assign n1230 = n1160 & ~n1229;
  assign n1231 = n1230 ^ n1154;
  assign n1224 = x5 & n756;
  assign n1225 = n1224 ^ n873;
  assign n1222 = x4 & n870;
  assign n1223 = n1222 ^ n953;
  assign n1226 = n1225 ^ n1223;
  assign n1218 = x15 & n157;
  assign n1219 = n1218 ^ n191;
  assign n1216 = x14 & n188;
  assign n1217 = n1216 ^ n248;
  assign n1220 = n1219 ^ n1217;
  assign n1213 = ~x7 & n567;
  assign n1214 = n1213 ^ n672;
  assign n1211 = ~x6 & n669;
  assign n1212 = n1211 ^ n738;
  assign n1215 = n1214 ^ n1212;
  assign n1221 = n1220 ^ n1215;
  assign n1227 = n1226 ^ n1221;
  assign n1207 = x1 & n1105;
  assign n1206 = x53 & n1105;
  assign n1208 = n1207 ^ n1206;
  assign n1202 = x53 ^ x52;
  assign n1203 = ~n1105 & n1202;
  assign n1204 = x53 ^ x0;
  assign n1205 = n1203 & n1204;
  assign n1209 = n1208 ^ n1205;
  assign n1198 = ~x3 & n894;
  assign n1199 = n1198 ^ n1052;
  assign n1196 = ~x2 & n1049;
  assign n1197 = n1196 ^ n1087;
  assign n1200 = n1199 ^ n1197;
  assign n1193 = x13 & n241;
  assign n1194 = n1193 ^ n293;
  assign n1191 = x12 & n290;
  assign n1192 = n1191 ^ n342;
  assign n1195 = n1194 ^ n1192;
  assign n1201 = n1200 ^ n1195;
  assign n1210 = n1209 ^ n1201;
  assign n1228 = n1227 ^ n1210;
  assign n1232 = n1231 ^ n1228;
  assign n1236 = n1235 ^ n1232;
  assign n1286 = n1285 ^ n1236;
  assign n1291 = n1290 ^ n1286;
  assign n1295 = n1294 ^ n1291;
  assign n1299 = n1298 ^ n1295;
  assign n1303 = n1302 ^ n1299;
  assign n1412 = n1302 ^ n1295;
  assign n1413 = ~n1299 & n1412;
  assign n1414 = n1413 ^ n1302;
  assign n1407 = n1294 ^ n1286;
  assign n1408 = n1294 ^ n1290;
  assign n1409 = n1407 & ~n1408;
  assign n1410 = n1409 ^ n1286;
  assign n1403 = n1285 ^ n1232;
  assign n1404 = n1236 & ~n1403;
  assign n1405 = n1404 ^ n1235;
  assign n1397 = n1280 ^ n1260;
  assign n1398 = n1283 ^ n1260;
  assign n1399 = n1397 & ~n1398;
  assign n1400 = n1399 ^ n1280;
  assign n1392 = n1279 ^ n1269;
  assign n1393 = n1275 & ~n1392;
  assign n1394 = n1393 ^ n1274;
  assign n1387 = ~x21 & n68;
  assign n1388 = n1387 ^ n69;
  assign n1386 = x22 & x32;
  assign n1389 = n1388 ^ n1386;
  assign n1382 = x2 & n1105;
  assign n1383 = n1382 ^ n1206;
  assign n1380 = x1 & n1203;
  assign n1379 = x53 & n1203;
  assign n1381 = n1380 ^ n1379;
  assign n1384 = n1383 ^ n1381;
  assign n1376 = ~x4 & n894;
  assign n1377 = n1376 ^ n1052;
  assign n1374 = ~x3 & n1049;
  assign n1375 = n1374 ^ n1087;
  assign n1378 = n1377 ^ n1375;
  assign n1385 = n1384 ^ n1378;
  assign n1390 = n1389 ^ n1385;
  assign n1370 = x16 & n157;
  assign n1371 = n1370 ^ n191;
  assign n1368 = x15 & n188;
  assign n1369 = n1368 ^ n248;
  assign n1372 = n1371 ^ n1369;
  assign n1364 = x20 & n75;
  assign n1365 = n1364 ^ n96;
  assign n1362 = x19 & n93;
  assign n1363 = n1362 ^ n108;
  assign n1366 = n1365 ^ n1363;
  assign n1360 = x54 ^ x53;
  assign n1361 = x0 & n1360;
  assign n1367 = n1366 ^ n1361;
  assign n1373 = n1372 ^ n1367;
  assign n1391 = n1390 ^ n1373;
  assign n1395 = n1394 ^ n1391;
  assign n1355 = n1226 ^ n1220;
  assign n1356 = n1221 & ~n1355;
  assign n1357 = n1356 ^ n1215;
  assign n1351 = x10 & n435;
  assign n1352 = n1351 ^ n527;
  assign n1349 = x9 & n524;
  assign n1350 = n1349 ^ n611;
  assign n1353 = n1352 ^ n1350;
  assign n1345 = ~x12 & n322;
  assign n1346 = n1345 ^ n382;
  assign n1343 = ~x11 & n379;
  assign n1344 = n1343 ^ n459;
  assign n1347 = n1346 ^ n1344;
  assign n1340 = x18 & n106;
  assign n1341 = n1340 ^ n142;
  assign n1338 = x17 & n139;
  assign n1339 = n1338 ^ n171;
  assign n1342 = n1341 ^ n1339;
  assign n1348 = n1347 ^ n1342;
  assign n1354 = n1353 ^ n1348;
  assign n1358 = n1357 ^ n1354;
  assign n1334 = x14 & n241;
  assign n1335 = n1334 ^ n293;
  assign n1332 = x13 & n290;
  assign n1333 = n1332 ^ n342;
  assign n1336 = n1335 ^ n1333;
  assign n1328 = x6 & n756;
  assign n1329 = n1328 ^ n873;
  assign n1326 = x5 & n870;
  assign n1327 = n1326 ^ n953;
  assign n1330 = n1329 ^ n1327;
  assign n1323 = ~x8 & n567;
  assign n1324 = n1323 ^ n672;
  assign n1321 = ~x7 & n669;
  assign n1322 = n1321 ^ n738;
  assign n1325 = n1324 ^ n1322;
  assign n1331 = n1330 ^ n1325;
  assign n1337 = n1336 ^ n1331;
  assign n1359 = n1358 ^ n1337;
  assign n1396 = n1395 ^ n1359;
  assign n1401 = n1400 ^ n1396;
  assign n1317 = n1231 ^ n1227;
  assign n1318 = n1228 & ~n1317;
  assign n1319 = n1318 ^ n1210;
  assign n1313 = n1255 ^ n1252;
  assign n1314 = ~n1259 & n1313;
  assign n1315 = n1314 ^ n1252;
  assign n1309 = n1209 ^ n1195;
  assign n1310 = ~n1201 & n1309;
  assign n1311 = n1310 ^ n1209;
  assign n1305 = n1251 ^ n1241;
  assign n1306 = n1246 & ~n1305;
  assign n1307 = n1306 ^ n1245;
  assign n1304 = n1263 & n1268;
  assign n1308 = n1307 ^ n1304;
  assign n1312 = n1311 ^ n1308;
  assign n1316 = n1315 ^ n1312;
  assign n1320 = n1319 ^ n1316;
  assign n1402 = n1401 ^ n1320;
  assign n1406 = n1405 ^ n1402;
  assign n1411 = n1410 ^ n1406;
  assign n1415 = n1414 ^ n1411;
  assign n1535 = n1414 ^ n1406;
  assign n1536 = ~n1411 & n1535;
  assign n1537 = n1536 ^ n1414;
  assign n1531 = n1405 ^ n1401;
  assign n1532 = n1402 & ~n1531;
  assign n1533 = n1532 ^ n1320;
  assign n1526 = n1400 ^ n1395;
  assign n1527 = n1396 & ~n1526;
  assign n1528 = n1527 ^ n1359;
  assign n1523 = n1319 ^ n1315;
  assign n1524 = n1316 & ~n1523;
  assign n1525 = n1524 ^ n1312;
  assign n1529 = n1528 ^ n1525;
  assign n1518 = n1394 ^ n1390;
  assign n1519 = n1391 & ~n1518;
  assign n1520 = n1519 ^ n1373;
  assign n1514 = n1311 ^ n1307;
  assign n1515 = n1308 & ~n1514;
  assign n1516 = n1515 ^ n1304;
  assign n1509 = x7 & n756;
  assign n1510 = n1509 ^ n873;
  assign n1507 = x6 & n870;
  assign n1508 = n1507 ^ n953;
  assign n1511 = n1510 ^ n1508;
  assign n1503 = ~x9 & n567;
  assign n1504 = n1503 ^ n672;
  assign n1501 = ~x8 & n669;
  assign n1502 = n1501 ^ n738;
  assign n1505 = n1504 ^ n1502;
  assign n1498 = x17 & n157;
  assign n1499 = n1498 ^ n191;
  assign n1496 = x16 & n188;
  assign n1497 = n1496 ^ n248;
  assign n1500 = n1499 ^ n1497;
  assign n1506 = n1505 ^ n1500;
  assign n1512 = n1511 ^ n1506;
  assign n1491 = x21 & n75;
  assign n1492 = n1491 ^ n96;
  assign n1489 = x20 & n93;
  assign n1490 = n1489 ^ n108;
  assign n1493 = n1492 ^ n1490;
  assign n1486 = n1204 & ~n1360;
  assign n1487 = n1486 ^ x0;
  assign n1488 = x55 & ~n1487;
  assign n1494 = n1493 ^ n1488;
  assign n1482 = x11 & n435;
  assign n1483 = n1482 ^ n527;
  assign n1480 = x10 & n524;
  assign n1481 = n1480 ^ n611;
  assign n1484 = n1483 ^ n1481;
  assign n1477 = ~x13 & n322;
  assign n1478 = n1477 ^ n382;
  assign n1475 = ~x12 & n379;
  assign n1476 = n1475 ^ n459;
  assign n1479 = n1478 ^ n1476;
  assign n1485 = n1484 ^ n1479;
  assign n1495 = n1494 ^ n1485;
  assign n1513 = n1512 ^ n1495;
  assign n1517 = n1516 ^ n1513;
  assign n1521 = n1520 ^ n1517;
  assign n1469 = n1354 ^ n1337;
  assign n1470 = n1357 ^ n1337;
  assign n1471 = n1469 & ~n1470;
  assign n1472 = n1471 ^ n1354;
  assign n1464 = n1372 ^ n1361;
  assign n1465 = n1372 ^ n1366;
  assign n1466 = n1464 & ~n1465;
  assign n1467 = n1466 ^ n1361;
  assign n1460 = n1389 ^ n1378;
  assign n1461 = ~n1385 & n1460;
  assign n1462 = n1461 ^ n1389;
  assign n1457 = n1353 ^ n1347;
  assign n1458 = n1348 & ~n1457;
  assign n1459 = n1458 ^ n1342;
  assign n1463 = n1462 ^ n1459;
  assign n1468 = n1467 ^ n1463;
  assign n1473 = n1472 ^ n1468;
  assign n1452 = n1336 ^ n1325;
  assign n1453 = ~n1331 & n1452;
  assign n1454 = n1453 ^ n1336;
  assign n1448 = x1 & n1360;
  assign n1447 = x55 & n1360;
  assign n1449 = n1448 ^ n1447;
  assign n1443 = x55 ^ x54;
  assign n1444 = ~n1360 & n1443;
  assign n1445 = x55 ^ x0;
  assign n1446 = n1444 & n1445;
  assign n1450 = n1449 ^ n1446;
  assign n1439 = ~x22 & n68;
  assign n1440 = n1439 ^ n69;
  assign n1438 = x23 & x32;
  assign n1441 = n1440 ^ n1438;
  assign n1435 = x19 & n106;
  assign n1436 = n1435 ^ n142;
  assign n1433 = x18 & n139;
  assign n1434 = n1433 ^ n171;
  assign n1437 = n1436 ^ n1434;
  assign n1442 = n1441 ^ n1437;
  assign n1451 = n1450 ^ n1442;
  assign n1455 = n1454 ^ n1451;
  assign n1429 = x3 & n1105;
  assign n1430 = n1429 ^ n1206;
  assign n1427 = x2 & n1203;
  assign n1428 = n1427 ^ n1379;
  assign n1431 = n1430 ^ n1428;
  assign n1423 = ~x5 & n894;
  assign n1424 = n1423 ^ n1052;
  assign n1421 = ~x4 & n1049;
  assign n1422 = n1421 ^ n1087;
  assign n1425 = n1424 ^ n1422;
  assign n1418 = x15 & n241;
  assign n1419 = n1418 ^ n293;
  assign n1416 = x14 & n290;
  assign n1417 = n1416 ^ n342;
  assign n1420 = n1419 ^ n1417;
  assign n1426 = n1425 ^ n1420;
  assign n1432 = n1431 ^ n1426;
  assign n1456 = n1455 ^ n1432;
  assign n1474 = n1473 ^ n1456;
  assign n1522 = n1521 ^ n1474;
  assign n1530 = n1529 ^ n1522;
  assign n1534 = n1533 ^ n1530;
  assign n1538 = n1537 ^ n1534;
  assign n1656 = n1537 ^ n1530;
  assign n1657 = ~n1534 & n1656;
  assign n1658 = n1657 ^ n1537;
  assign n1652 = n1525 ^ n1522;
  assign n1653 = ~n1529 & n1652;
  assign n1654 = n1653 ^ n1522;
  assign n1647 = n1517 ^ n1474;
  assign n1648 = n1520 ^ n1474;
  assign n1649 = n1647 & ~n1648;
  assign n1650 = n1649 ^ n1517;
  assign n1642 = n1468 ^ n1456;
  assign n1643 = ~n1473 & n1642;
  assign n1644 = n1643 ^ n1456;
  assign n1638 = n1516 ^ n1512;
  assign n1639 = n1513 & ~n1638;
  assign n1640 = n1639 ^ n1495;
  assign n1633 = n1467 ^ n1459;
  assign n1634 = ~n1463 & n1633;
  assign n1635 = n1634 ^ n1467;
  assign n1630 = n1494 ^ n1484;
  assign n1631 = n1485 & ~n1630;
  assign n1632 = n1631 ^ n1479;
  assign n1636 = n1635 ^ n1632;
  assign n1626 = n1431 ^ n1420;
  assign n1627 = ~n1426 & n1626;
  assign n1628 = n1627 ^ n1431;
  assign n1622 = x12 & n435;
  assign n1623 = n1622 ^ n527;
  assign n1620 = x11 & n524;
  assign n1621 = n1620 ^ n611;
  assign n1624 = n1623 ^ n1621;
  assign n1619 = n1488 & n1493;
  assign n1625 = n1624 ^ n1619;
  assign n1629 = n1628 ^ n1625;
  assign n1637 = n1636 ^ n1629;
  assign n1641 = n1640 ^ n1637;
  assign n1645 = n1644 ^ n1641;
  assign n1614 = n1451 ^ n1432;
  assign n1615 = ~n1455 & n1614;
  assign n1616 = n1615 ^ n1432;
  assign n1609 = n1511 ^ n1500;
  assign n1610 = ~n1506 & n1609;
  assign n1611 = n1610 ^ n1511;
  assign n1606 = n1450 ^ n1437;
  assign n1607 = n1442 & ~n1606;
  assign n1608 = n1607 ^ n1441;
  assign n1612 = n1611 ^ n1608;
  assign n1602 = ~x14 & n322;
  assign n1603 = n1602 ^ n382;
  assign n1600 = ~x13 & n379;
  assign n1601 = n1600 ^ n459;
  assign n1604 = n1603 ^ n1601;
  assign n1596 = x20 & n106;
  assign n1597 = n1596 ^ n142;
  assign n1594 = x19 & n139;
  assign n1595 = n1594 ^ n171;
  assign n1598 = n1597 ^ n1595;
  assign n1591 = x2 & n1360;
  assign n1592 = n1591 ^ n1447;
  assign n1589 = x1 & n1444;
  assign n1588 = x55 & n1444;
  assign n1590 = n1589 ^ n1588;
  assign n1593 = n1592 ^ n1590;
  assign n1599 = n1598 ^ n1593;
  assign n1605 = n1604 ^ n1599;
  assign n1613 = n1612 ^ n1605;
  assign n1617 = n1616 ^ n1613;
  assign n1582 = ~x23 & n68;
  assign n1583 = n1582 ^ n69;
  assign n1581 = x24 & x32;
  assign n1584 = n1583 ^ n1581;
  assign n1577 = x4 & n1105;
  assign n1578 = n1577 ^ n1206;
  assign n1575 = x3 & n1203;
  assign n1576 = n1575 ^ n1379;
  assign n1579 = n1578 ^ n1576;
  assign n1572 = ~x6 & n894;
  assign n1573 = n1572 ^ n1052;
  assign n1570 = ~x5 & n1049;
  assign n1571 = n1570 ^ n1087;
  assign n1574 = n1573 ^ n1571;
  assign n1580 = n1579 ^ n1574;
  assign n1585 = n1584 ^ n1580;
  assign n1566 = x18 & n157;
  assign n1567 = n1566 ^ n191;
  assign n1564 = x17 & n188;
  assign n1565 = n1564 ^ n248;
  assign n1568 = n1567 ^ n1565;
  assign n1560 = x22 & n75;
  assign n1561 = n1560 ^ n96;
  assign n1558 = x21 & n93;
  assign n1559 = n1558 ^ n108;
  assign n1562 = n1561 ^ n1559;
  assign n1556 = x56 ^ x55;
  assign n1557 = x0 & n1556;
  assign n1563 = n1562 ^ n1557;
  assign n1569 = n1568 ^ n1563;
  assign n1586 = n1585 ^ n1569;
  assign n1552 = x16 & n241;
  assign n1553 = n1552 ^ n293;
  assign n1550 = x15 & n290;
  assign n1551 = n1550 ^ n342;
  assign n1554 = n1553 ^ n1551;
  assign n1546 = ~x10 & n567;
  assign n1547 = n1546 ^ n672;
  assign n1544 = ~x9 & n669;
  assign n1545 = n1544 ^ n738;
  assign n1548 = n1547 ^ n1545;
  assign n1541 = x8 & n756;
  assign n1542 = n1541 ^ n873;
  assign n1539 = x7 & n870;
  assign n1540 = n1539 ^ n953;
  assign n1543 = n1542 ^ n1540;
  assign n1549 = n1548 ^ n1543;
  assign n1555 = n1554 ^ n1549;
  assign n1587 = n1586 ^ n1555;
  assign n1618 = n1617 ^ n1587;
  assign n1646 = n1645 ^ n1618;
  assign n1651 = n1650 ^ n1646;
  assign n1655 = n1654 ^ n1651;
  assign n1659 = n1658 ^ n1655;
  assign n1791 = n1658 ^ n1651;
  assign n1792 = ~n1655 & n1791;
  assign n1793 = n1792 ^ n1658;
  assign n1787 = n1650 ^ n1645;
  assign n1788 = n1646 & ~n1787;
  assign n1789 = n1788 ^ n1618;
  assign n1782 = n1644 ^ n1640;
  assign n1783 = n1641 & ~n1782;
  assign n1784 = n1783 ^ n1637;
  assign n1777 = n1608 ^ n1605;
  assign n1778 = ~n1612 & n1777;
  assign n1779 = n1778 ^ n1605;
  assign n1773 = n1584 ^ n1574;
  assign n1774 = ~n1580 & n1773;
  assign n1775 = n1774 ^ n1584;
  assign n1768 = n1554 ^ n1543;
  assign n1769 = n1554 ^ n1548;
  assign n1770 = n1768 & ~n1769;
  assign n1771 = n1770 ^ n1543;
  assign n1764 = x23 & n75;
  assign n1765 = n1764 ^ n96;
  assign n1762 = x22 & n93;
  assign n1763 = n1762 ^ n108;
  assign n1766 = n1765 ^ n1763;
  assign n1759 = n1445 & ~n1556;
  assign n1760 = n1759 ^ x0;
  assign n1761 = x57 & ~n1760;
  assign n1767 = n1766 ^ n1761;
  assign n1772 = n1771 ^ n1767;
  assign n1776 = n1775 ^ n1772;
  assign n1780 = n1779 ^ n1776;
  assign n1753 = x5 & n1105;
  assign n1754 = n1753 ^ n1206;
  assign n1751 = x4 & n1203;
  assign n1752 = n1751 ^ n1379;
  assign n1755 = n1754 ^ n1752;
  assign n1747 = ~x7 & n894;
  assign n1748 = n1747 ^ n1052;
  assign n1745 = ~x6 & n1049;
  assign n1746 = n1745 ^ n1087;
  assign n1749 = n1748 ^ n1746;
  assign n1742 = x17 & n241;
  assign n1743 = n1742 ^ n293;
  assign n1740 = x16 & n290;
  assign n1741 = n1740 ^ n342;
  assign n1744 = n1743 ^ n1741;
  assign n1750 = n1749 ^ n1744;
  assign n1756 = n1755 ^ n1750;
  assign n1736 = x9 & n756;
  assign n1737 = n1736 ^ n873;
  assign n1734 = x8 & n870;
  assign n1735 = n1734 ^ n953;
  assign n1738 = n1737 ^ n1735;
  assign n1730 = ~x11 & n567;
  assign n1731 = n1730 ^ n672;
  assign n1728 = ~x10 & n669;
  assign n1729 = n1728 ^ n738;
  assign n1732 = n1731 ^ n1729;
  assign n1725 = x19 & n157;
  assign n1726 = n1725 ^ n191;
  assign n1723 = x18 & n188;
  assign n1724 = n1723 ^ n248;
  assign n1727 = n1726 ^ n1724;
  assign n1733 = n1732 ^ n1727;
  assign n1739 = n1738 ^ n1733;
  assign n1757 = n1756 ^ n1739;
  assign n1719 = x3 & n1360;
  assign n1720 = n1719 ^ n1447;
  assign n1717 = x2 & n1444;
  assign n1718 = n1717 ^ n1588;
  assign n1721 = n1720 ^ n1718;
  assign n1713 = ~x24 & n68;
  assign n1714 = n1713 ^ n69;
  assign n1712 = x25 & x32;
  assign n1715 = n1714 ^ n1712;
  assign n1709 = ~x15 & n322;
  assign n1710 = n1709 ^ n382;
  assign n1707 = ~x14 & n379;
  assign n1708 = n1707 ^ n459;
  assign n1711 = n1710 ^ n1708;
  assign n1716 = n1715 ^ n1711;
  assign n1722 = n1721 ^ n1716;
  assign n1758 = n1757 ^ n1722;
  assign n1781 = n1780 ^ n1758;
  assign n1785 = n1784 ^ n1781;
  assign n1701 = n1632 ^ n1629;
  assign n1702 = n1635 ^ n1629;
  assign n1703 = n1701 & ~n1702;
  assign n1704 = n1703 ^ n1632;
  assign n1698 = n1613 ^ n1587;
  assign n1699 = ~n1617 & n1698;
  assign n1700 = n1699 ^ n1587;
  assign n1705 = n1704 ^ n1700;
  assign n1693 = n1569 ^ n1555;
  assign n1694 = n1585 ^ n1555;
  assign n1695 = n1693 & ~n1694;
  assign n1696 = n1695 ^ n1569;
  assign n1689 = n1628 ^ n1619;
  assign n1690 = n1625 & ~n1689;
  assign n1691 = n1690 ^ n1624;
  assign n1683 = n1604 ^ n1593;
  assign n1684 = n1604 ^ n1598;
  assign n1685 = n1683 & ~n1684;
  assign n1686 = n1685 ^ n1593;
  assign n1680 = n1568 ^ n1562;
  assign n1681 = n1563 & ~n1680;
  assign n1682 = n1681 ^ n1557;
  assign n1687 = n1686 ^ n1682;
  assign n1676 = x13 & n435;
  assign n1677 = n1676 ^ n527;
  assign n1674 = x12 & n524;
  assign n1675 = n1674 ^ n611;
  assign n1678 = n1677 ^ n1675;
  assign n1670 = x21 & n106;
  assign n1671 = n1670 ^ n142;
  assign n1668 = x20 & n139;
  assign n1669 = n1668 ^ n171;
  assign n1672 = n1671 ^ n1669;
  assign n1665 = x1 & n1556;
  assign n1664 = x57 & n1556;
  assign n1666 = n1665 ^ n1664;
  assign n1660 = x57 ^ x56;
  assign n1661 = ~n1556 & n1660;
  assign n1662 = x57 ^ x0;
  assign n1663 = n1661 & n1662;
  assign n1667 = n1666 ^ n1663;
  assign n1673 = n1672 ^ n1667;
  assign n1679 = n1678 ^ n1673;
  assign n1688 = n1687 ^ n1679;
  assign n1692 = n1691 ^ n1688;
  assign n1697 = n1696 ^ n1692;
  assign n1706 = n1705 ^ n1697;
  assign n1786 = n1785 ^ n1706;
  assign n1790 = n1789 ^ n1786;
  assign n1794 = n1793 ^ n1790;
  assign n1925 = n1793 ^ n1786;
  assign n1926 = ~n1790 & n1925;
  assign n1927 = n1926 ^ n1793;
  assign n1920 = n1781 ^ n1706;
  assign n1921 = n1784 ^ n1706;
  assign n1922 = n1920 & ~n1921;
  assign n1923 = n1922 ^ n1781;
  assign n1915 = n1700 ^ n1697;
  assign n1916 = ~n1705 & n1915;
  assign n1917 = n1916 ^ n1697;
  assign n1908 = n1721 ^ n1715;
  assign n1909 = n1721 ^ n1711;
  assign n1910 = n1908 & ~n1909;
  assign n1911 = n1910 ^ n1715;
  assign n1903 = n1755 ^ n1744;
  assign n1904 = n1755 ^ n1749;
  assign n1905 = n1903 & ~n1904;
  assign n1906 = n1905 ^ n1744;
  assign n1900 = n1738 ^ n1732;
  assign n1901 = n1733 & ~n1900;
  assign n1902 = n1901 ^ n1727;
  assign n1907 = n1906 ^ n1902;
  assign n1912 = n1911 ^ n1907;
  assign n1897 = n1761 & n1766;
  assign n1893 = x14 & n435;
  assign n1894 = n1893 ^ n527;
  assign n1891 = x13 & n524;
  assign n1892 = n1891 ^ n611;
  assign n1895 = n1894 ^ n1892;
  assign n1888 = x22 & n106;
  assign n1889 = n1888 ^ n142;
  assign n1886 = x21 & n139;
  assign n1887 = n1886 ^ n171;
  assign n1890 = n1889 ^ n1887;
  assign n1896 = n1895 ^ n1890;
  assign n1898 = n1897 ^ n1896;
  assign n1881 = x2 & n1556;
  assign n1882 = n1881 ^ n1664;
  assign n1879 = x1 & n1661;
  assign n1878 = x57 & n1661;
  assign n1880 = n1879 ^ n1878;
  assign n1883 = n1882 ^ n1880;
  assign n1874 = ~x16 & n322;
  assign n1875 = n1874 ^ n382;
  assign n1872 = ~x15 & n379;
  assign n1873 = n1872 ^ n459;
  assign n1876 = n1875 ^ n1873;
  assign n1869 = x4 & n1360;
  assign n1870 = n1869 ^ n1447;
  assign n1867 = x3 & n1444;
  assign n1868 = n1867 ^ n1588;
  assign n1871 = n1870 ^ n1868;
  assign n1877 = n1876 ^ n1871;
  assign n1884 = n1883 ^ n1877;
  assign n1863 = x18 & n241;
  assign n1864 = n1863 ^ n293;
  assign n1861 = x17 & n290;
  assign n1862 = n1861 ^ n342;
  assign n1865 = n1864 ^ n1862;
  assign n1857 = ~x12 & n567;
  assign n1858 = n1857 ^ n672;
  assign n1855 = ~x11 & n669;
  assign n1856 = n1855 ^ n738;
  assign n1859 = n1858 ^ n1856;
  assign n1852 = x10 & n756;
  assign n1853 = n1852 ^ n873;
  assign n1850 = x9 & n870;
  assign n1851 = n1850 ^ n953;
  assign n1854 = n1853 ^ n1851;
  assign n1860 = n1859 ^ n1854;
  assign n1866 = n1865 ^ n1860;
  assign n1885 = n1884 ^ n1866;
  assign n1899 = n1898 ^ n1885;
  assign n1913 = n1912 ^ n1899;
  assign n1845 = ~x25 & n68;
  assign n1846 = n1845 ^ n69;
  assign n1844 = x26 & x32;
  assign n1847 = n1846 ^ n1844;
  assign n1840 = ~x8 & n894;
  assign n1841 = n1840 ^ n1052;
  assign n1838 = ~x7 & n1049;
  assign n1839 = n1838 ^ n1087;
  assign n1842 = n1841 ^ n1839;
  assign n1835 = x6 & n1105;
  assign n1836 = n1835 ^ n1206;
  assign n1833 = x5 & n1203;
  assign n1834 = n1833 ^ n1379;
  assign n1837 = n1836 ^ n1834;
  assign n1843 = n1842 ^ n1837;
  assign n1848 = n1847 ^ n1843;
  assign n1829 = n1678 ^ n1672;
  assign n1830 = n1673 & ~n1829;
  assign n1831 = n1830 ^ n1667;
  assign n1825 = x20 & n157;
  assign n1826 = n1825 ^ n191;
  assign n1823 = x19 & n188;
  assign n1824 = n1823 ^ n248;
  assign n1827 = n1826 ^ n1824;
  assign n1819 = x24 & n75;
  assign n1820 = n1819 ^ n96;
  assign n1817 = x23 & n93;
  assign n1818 = n1817 ^ n108;
  assign n1821 = n1820 ^ n1818;
  assign n1815 = x58 ^ x57;
  assign n1816 = x0 & n1815;
  assign n1822 = n1821 ^ n1816;
  assign n1828 = n1827 ^ n1822;
  assign n1832 = n1831 ^ n1828;
  assign n1849 = n1848 ^ n1832;
  assign n1914 = n1913 ^ n1849;
  assign n1918 = n1917 ^ n1914;
  assign n1811 = n1776 ^ n1758;
  assign n1812 = ~n1780 & n1811;
  assign n1813 = n1812 ^ n1758;
  assign n1806 = n1696 ^ n1688;
  assign n1807 = n1696 ^ n1691;
  assign n1808 = n1806 & ~n1807;
  assign n1809 = n1808 ^ n1688;
  assign n1802 = n1756 ^ n1722;
  assign n1803 = n1757 & ~n1802;
  assign n1804 = n1803 ^ n1739;
  assign n1798 = n1682 ^ n1679;
  assign n1799 = ~n1687 & n1798;
  assign n1800 = n1799 ^ n1679;
  assign n1795 = n1775 ^ n1771;
  assign n1796 = n1772 & ~n1795;
  assign n1797 = n1796 ^ n1767;
  assign n1801 = n1800 ^ n1797;
  assign n1805 = n1804 ^ n1801;
  assign n1810 = n1809 ^ n1805;
  assign n1814 = n1813 ^ n1810;
  assign n1919 = n1918 ^ n1814;
  assign n1924 = n1923 ^ n1919;
  assign n1928 = n1927 ^ n1924;
  assign n2069 = n1927 ^ n1919;
  assign n2070 = ~n1924 & n2069;
  assign n2071 = n2070 ^ n1927;
  assign n2064 = n1914 ^ n1814;
  assign n2065 = n1917 ^ n1814;
  assign n2066 = n2064 & ~n2065;
  assign n2067 = n2066 ^ n1914;
  assign n2059 = n1813 ^ n1809;
  assign n2060 = n1810 & ~n2059;
  assign n2061 = n2060 ^ n1805;
  assign n2054 = n1898 ^ n1884;
  assign n2055 = n1885 & ~n2054;
  assign n2056 = n2055 ^ n1866;
  assign n2048 = ~x1 & n1815;
  assign n2047 = ~x59 & n1815;
  assign n2049 = n2048 ^ n2047;
  assign n2043 = x59 ^ x58;
  assign n2044 = ~n1815 & n2043;
  assign n2045 = x59 ^ x0;
  assign n2046 = n2044 & n2045;
  assign n2050 = n2049 ^ n2046;
  assign n2039 = x23 & n106;
  assign n2040 = n2039 ^ n142;
  assign n2037 = x22 & n139;
  assign n2038 = n2037 ^ n171;
  assign n2041 = n2040 ^ n2038;
  assign n2034 = x3 & n1556;
  assign n2035 = n2034 ^ n1664;
  assign n2032 = x2 & n1661;
  assign n2033 = n2032 ^ n1878;
  assign n2036 = n2035 ^ n2033;
  assign n2042 = n2041 ^ n2036;
  assign n2051 = n2050 ^ n2042;
  assign n2028 = x11 & n756;
  assign n2029 = n2028 ^ n873;
  assign n2026 = x10 & n870;
  assign n2027 = n2026 ^ n953;
  assign n2030 = n2029 ^ n2027;
  assign n2022 = ~x13 & n567;
  assign n2023 = n2022 ^ n672;
  assign n2020 = ~x12 & n669;
  assign n2021 = n2020 ^ n738;
  assign n2024 = n2023 ^ n2021;
  assign n2017 = x21 & n157;
  assign n2018 = n2017 ^ n191;
  assign n2015 = x20 & n188;
  assign n2016 = n2015 ^ n248;
  assign n2019 = n2018 ^ n2016;
  assign n2025 = n2024 ^ n2019;
  assign n2031 = n2030 ^ n2025;
  assign n2052 = n2051 ^ n2031;
  assign n2011 = x5 & n1360;
  assign n2012 = n2011 ^ n1447;
  assign n2009 = x4 & n1444;
  assign n2010 = n2009 ^ n1588;
  assign n2013 = n2012 ^ n2010;
  assign n2005 = ~x26 & n68;
  assign n2006 = n2005 ^ n69;
  assign n2004 = x27 & x32;
  assign n2007 = n2006 ^ n2004;
  assign n2001 = ~x17 & n322;
  assign n2002 = n2001 ^ n382;
  assign n1999 = ~x16 & n379;
  assign n2000 = n1999 ^ n459;
  assign n2003 = n2002 ^ n2000;
  assign n2008 = n2007 ^ n2003;
  assign n2014 = n2013 ^ n2008;
  assign n2053 = n2052 ^ n2014;
  assign n2057 = n2056 ^ n2053;
  assign n1994 = n1897 ^ n1895;
  assign n1995 = n1896 & ~n1994;
  assign n1996 = n1995 ^ n1890;
  assign n1990 = x7 & n1105;
  assign n1991 = n1990 ^ n1206;
  assign n1988 = x6 & n1203;
  assign n1989 = n1988 ^ n1379;
  assign n1992 = n1991 ^ n1989;
  assign n1984 = ~x9 & n894;
  assign n1985 = n1984 ^ n1052;
  assign n1982 = ~x8 & n1049;
  assign n1983 = n1982 ^ n1087;
  assign n1986 = n1985 ^ n1983;
  assign n1979 = x19 & n241;
  assign n1980 = n1979 ^ n293;
  assign n1977 = x18 & n290;
  assign n1978 = n1977 ^ n342;
  assign n1981 = n1980 ^ n1978;
  assign n1987 = n1986 ^ n1981;
  assign n1993 = n1992 ^ n1987;
  assign n1997 = n1996 ^ n1993;
  assign n1973 = n1827 ^ n1821;
  assign n1974 = n1822 & ~n1973;
  assign n1975 = n1974 ^ n1816;
  assign n1969 = x15 & n435;
  assign n1970 = n1969 ^ n527;
  assign n1967 = x14 & n524;
  assign n1968 = n1967 ^ n611;
  assign n1971 = n1970 ^ n1968;
  assign n1963 = x25 & n75;
  assign n1964 = n1963 ^ n96;
  assign n1961 = x24 & n93;
  assign n1962 = n1961 ^ n108;
  assign n1965 = n1964 ^ n1962;
  assign n1958 = n1662 & ~n1815;
  assign n1959 = n1958 ^ x0;
  assign n1960 = x59 & ~n1959;
  assign n1966 = n1965 ^ n1960;
  assign n1972 = n1971 ^ n1966;
  assign n1976 = n1975 ^ n1972;
  assign n1998 = n1997 ^ n1976;
  assign n2058 = n2057 ^ n1998;
  assign n2062 = n2061 ^ n2058;
  assign n1953 = n1804 ^ n1797;
  assign n1954 = ~n1801 & n1953;
  assign n1955 = n1954 ^ n1804;
  assign n1949 = n1899 ^ n1849;
  assign n1950 = n1912 ^ n1849;
  assign n1951 = n1949 & ~n1950;
  assign n1952 = n1951 ^ n1899;
  assign n1956 = n1955 ^ n1952;
  assign n1944 = n1911 ^ n1906;
  assign n1945 = n1907 & ~n1944;
  assign n1946 = n1945 ^ n1902;
  assign n1941 = n1848 ^ n1828;
  assign n1942 = ~n1832 & n1941;
  assign n1943 = n1942 ^ n1848;
  assign n1947 = n1946 ^ n1943;
  assign n1937 = n1883 ^ n1876;
  assign n1938 = n1877 & ~n1937;
  assign n1939 = n1938 ^ n1871;
  assign n1933 = n1847 ^ n1837;
  assign n1934 = ~n1843 & n1933;
  assign n1935 = n1934 ^ n1847;
  assign n1929 = n1865 ^ n1854;
  assign n1930 = n1865 ^ n1859;
  assign n1931 = n1929 & ~n1930;
  assign n1932 = n1931 ^ n1854;
  assign n1936 = n1935 ^ n1932;
  assign n1940 = n1939 ^ n1936;
  assign n1948 = n1947 ^ n1940;
  assign n1957 = n1956 ^ n1948;
  assign n2063 = n2062 ^ n1957;
  assign n2068 = n2067 ^ n2063;
  assign n2072 = n2071 ^ n2068;
  assign n2212 = n2071 ^ n2063;
  assign n2213 = ~n2068 & n2212;
  assign n2214 = n2213 ^ n2071;
  assign n2207 = n2058 ^ n1957;
  assign n2208 = n2061 ^ n1957;
  assign n2209 = n2207 & ~n2208;
  assign n2210 = n2209 ^ n2058;
  assign n2201 = n1952 ^ n1948;
  assign n2202 = n1955 ^ n1948;
  assign n2203 = n2201 & ~n2202;
  assign n2204 = n2203 ^ n1952;
  assign n2197 = n1943 ^ n1940;
  assign n2198 = ~n1947 & n2197;
  assign n2199 = n2198 ^ n1940;
  assign n2193 = n1996 ^ n1976;
  assign n2194 = n1997 & ~n2193;
  assign n2195 = n2194 ^ n1993;
  assign n2188 = ~x27 & n68;
  assign n2189 = n2188 ^ n69;
  assign n2187 = x28 & x32;
  assign n2190 = n2189 ^ n2187;
  assign n2183 = x8 & n1105;
  assign n2184 = n2183 ^ n1206;
  assign n2181 = x7 & n1203;
  assign n2182 = n2181 ^ n1379;
  assign n2185 = n2184 ^ n2182;
  assign n2178 = ~x10 & n894;
  assign n2179 = n2178 ^ n1052;
  assign n2176 = ~x9 & n1049;
  assign n2177 = n2176 ^ n1087;
  assign n2180 = n2179 ^ n2177;
  assign n2186 = n2185 ^ n2180;
  assign n2191 = n2190 ^ n2186;
  assign n2171 = x16 & n435;
  assign n2172 = n2171 ^ n527;
  assign n2169 = x15 & n524;
  assign n2170 = n2169 ^ n611;
  assign n2173 = n2172 ^ n2170;
  assign n2165 = ~x2 & n1815;
  assign n2166 = n2165 ^ n2047;
  assign n2163 = ~x1 & n2044;
  assign n2162 = ~x59 & n2044;
  assign n2164 = n2163 ^ n2162;
  assign n2167 = n2166 ^ n2164;
  assign n2159 = x24 & n106;
  assign n2160 = n2159 ^ n142;
  assign n2157 = x23 & n139;
  assign n2158 = n2157 ^ n171;
  assign n2161 = n2160 ^ n2158;
  assign n2168 = n2167 ^ n2161;
  assign n2174 = n2173 ^ n2168;
  assign n2153 = x22 & n157;
  assign n2154 = n2153 ^ n191;
  assign n2151 = x21 & n188;
  assign n2152 = n2151 ^ n248;
  assign n2155 = n2154 ^ n2152;
  assign n2147 = x26 & n75;
  assign n2148 = n2147 ^ n96;
  assign n2145 = x25 & n93;
  assign n2146 = n2145 ^ n108;
  assign n2149 = n2148 ^ n2146;
  assign n2143 = x60 ^ x59;
  assign n2144 = x0 & n2143;
  assign n2150 = n2149 ^ n2144;
  assign n2156 = n2155 ^ n2150;
  assign n2175 = n2174 ^ n2156;
  assign n2192 = n2191 ^ n2175;
  assign n2196 = n2195 ^ n2192;
  assign n2200 = n2199 ^ n2196;
  assign n2205 = n2204 ^ n2200;
  assign n2138 = n2053 ^ n1998;
  assign n2139 = n2056 ^ n1998;
  assign n2140 = n2138 & ~n2139;
  assign n2141 = n2140 ^ n2053;
  assign n2133 = n1975 ^ n1966;
  assign n2134 = n1972 & ~n2133;
  assign n2135 = n2134 ^ n1971;
  assign n2129 = n1939 ^ n1932;
  assign n2130 = ~n1936 & n2129;
  assign n2131 = n2130 ^ n1939;
  assign n2125 = x4 & n1556;
  assign n2126 = n2125 ^ n1664;
  assign n2123 = x3 & n1661;
  assign n2124 = n2123 ^ n1878;
  assign n2127 = n2126 ^ n2124;
  assign n2119 = x6 & n1360;
  assign n2120 = n2119 ^ n1447;
  assign n2117 = x5 & n1444;
  assign n2118 = n2117 ^ n1588;
  assign n2121 = n2120 ^ n2118;
  assign n2114 = ~x18 & n322;
  assign n2115 = n2114 ^ n382;
  assign n2112 = ~x17 & n379;
  assign n2113 = n2112 ^ n459;
  assign n2116 = n2115 ^ n2113;
  assign n2122 = n2121 ^ n2116;
  assign n2128 = n2127 ^ n2122;
  assign n2132 = n2131 ^ n2128;
  assign n2136 = n2135 ^ n2132;
  assign n2108 = n2031 ^ n2014;
  assign n2109 = ~n2052 & n2108;
  assign n2110 = n2109 ^ n2014;
  assign n2103 = n1992 ^ n1986;
  assign n2104 = n1987 & ~n2103;
  assign n2105 = n2104 ^ n1981;
  assign n2099 = n2030 ^ n2024;
  assign n2100 = n2025 & ~n2099;
  assign n2101 = n2100 ^ n2019;
  assign n2098 = n1960 & n1965;
  assign n2102 = n2101 ^ n2098;
  assign n2106 = n2105 ^ n2102;
  assign n2093 = n2050 ^ n2041;
  assign n2094 = n2042 & ~n2093;
  assign n2095 = n2094 ^ n2036;
  assign n2090 = n2013 ^ n2003;
  assign n2091 = n2008 & ~n2090;
  assign n2092 = n2091 ^ n2007;
  assign n2096 = n2095 ^ n2092;
  assign n2086 = x20 & n241;
  assign n2087 = n2086 ^ n293;
  assign n2084 = x19 & n290;
  assign n2085 = n2084 ^ n342;
  assign n2088 = n2087 ^ n2085;
  assign n2080 = x12 & n756;
  assign n2081 = n2080 ^ n873;
  assign n2078 = x11 & n870;
  assign n2079 = n2078 ^ n953;
  assign n2082 = n2081 ^ n2079;
  assign n2075 = ~x14 & n567;
  assign n2076 = n2075 ^ n672;
  assign n2073 = ~x13 & n669;
  assign n2074 = n2073 ^ n738;
  assign n2077 = n2076 ^ n2074;
  assign n2083 = n2082 ^ n2077;
  assign n2089 = n2088 ^ n2083;
  assign n2097 = n2096 ^ n2089;
  assign n2107 = n2106 ^ n2097;
  assign n2111 = n2110 ^ n2107;
  assign n2137 = n2136 ^ n2111;
  assign n2142 = n2141 ^ n2137;
  assign n2206 = n2205 ^ n2142;
  assign n2211 = n2210 ^ n2206;
  assign n2215 = n2214 ^ n2211;
  assign n2366 = n2214 ^ n2206;
  assign n2367 = ~n2211 & n2366;
  assign n2368 = n2367 ^ n2214;
  assign n2362 = n2200 ^ n2142;
  assign n2363 = ~n2205 & n2362;
  assign n2364 = n2363 ^ n2142;
  assign n2357 = n2199 ^ n2195;
  assign n2358 = n2196 & ~n2357;
  assign n2359 = n2358 ^ n2192;
  assign n2354 = n2141 ^ n2136;
  assign n2355 = n2137 & ~n2354;
  assign n2356 = n2355 ^ n2111;
  assign n2360 = n2359 ^ n2356;
  assign n2349 = n2110 ^ n2097;
  assign n2350 = ~n2107 & n2349;
  assign n2351 = n2350 ^ n2110;
  assign n2344 = n2135 ^ n2128;
  assign n2345 = n2135 ^ n2131;
  assign n2346 = n2344 & ~n2345;
  assign n2347 = n2346 ^ n2128;
  assign n2338 = ~x11 & n894;
  assign n2339 = n2338 ^ n1052;
  assign n2336 = ~x10 & n1049;
  assign n2337 = n2336 ^ n1087;
  assign n2340 = n2339 ^ n2337;
  assign n2332 = x21 & n241;
  assign n2333 = n2332 ^ n293;
  assign n2330 = x20 & n290;
  assign n2331 = n2330 ^ n342;
  assign n2334 = n2333 ^ n2331;
  assign n2327 = x13 & n756;
  assign n2328 = n2327 ^ n873;
  assign n2325 = x12 & n870;
  assign n2326 = n2325 ^ n953;
  assign n2329 = n2328 ^ n2326;
  assign n2335 = n2334 ^ n2329;
  assign n2341 = n2340 ^ n2335;
  assign n2321 = x17 & n435;
  assign n2322 = n2321 ^ n527;
  assign n2319 = x16 & n524;
  assign n2320 = n2319 ^ n611;
  assign n2323 = n2322 ^ n2320;
  assign n2315 = x5 & n1556;
  assign n2316 = n2315 ^ n1664;
  assign n2313 = x4 & n1661;
  assign n2314 = n2313 ^ n1878;
  assign n2317 = n2316 ^ n2314;
  assign n2310 = x7 & n1360;
  assign n2311 = n2310 ^ n1447;
  assign n2308 = x6 & n1444;
  assign n2309 = n2308 ^ n1588;
  assign n2312 = n2311 ^ n2309;
  assign n2318 = n2317 ^ n2312;
  assign n2324 = n2323 ^ n2318;
  assign n2342 = n2341 ^ n2324;
  assign n2304 = ~x19 & n322;
  assign n2305 = n2304 ^ n382;
  assign n2302 = ~x18 & n379;
  assign n2303 = n2302 ^ n459;
  assign n2306 = n2305 ^ n2303;
  assign n2298 = x25 & n106;
  assign n2299 = n2298 ^ n142;
  assign n2296 = x24 & n139;
  assign n2297 = n2296 ^ n171;
  assign n2300 = n2299 ^ n2297;
  assign n2293 = x9 & n1105;
  assign n2294 = n2293 ^ n1206;
  assign n2291 = x8 & n1203;
  assign n2292 = n2291 ^ n1379;
  assign n2295 = n2294 ^ n2292;
  assign n2301 = n2300 ^ n2295;
  assign n2307 = n2306 ^ n2301;
  assign n2343 = n2342 ^ n2307;
  assign n2348 = n2347 ^ n2343;
  assign n2352 = n2351 ^ n2348;
  assign n2285 = n2191 ^ n2156;
  assign n2286 = n2191 ^ n2174;
  assign n2287 = n2285 & ~n2286;
  assign n2288 = n2287 ^ n2156;
  assign n2281 = n2105 ^ n2101;
  assign n2282 = n2102 & ~n2281;
  assign n2283 = n2282 ^ n2098;
  assign n2276 = x1 & n2143;
  assign n2275 = x61 & n2143;
  assign n2277 = n2276 ^ n2275;
  assign n2271 = x61 ^ x60;
  assign n2272 = ~n2143 & n2271;
  assign n2273 = x61 ^ x0;
  assign n2274 = n2272 & n2273;
  assign n2278 = n2277 ^ n2274;
  assign n2268 = ~x3 & n1815;
  assign n2269 = n2268 ^ n2047;
  assign n2266 = ~x2 & n2044;
  assign n2267 = n2266 ^ n2162;
  assign n2270 = n2269 ^ n2267;
  assign n2279 = n2278 ^ n2270;
  assign n2262 = ~x28 & n68;
  assign n2263 = n2262 ^ n69;
  assign n2261 = x29 & x32;
  assign n2264 = n2263 ^ n2261;
  assign n2258 = n2045 & ~n2143;
  assign n2259 = n2258 ^ x0;
  assign n2260 = x61 & ~n2259;
  assign n2265 = n2264 ^ n2260;
  assign n2280 = n2279 ^ n2265;
  assign n2284 = n2283 ^ n2280;
  assign n2289 = n2288 ^ n2284;
  assign n2253 = n2092 ^ n2089;
  assign n2254 = ~n2096 & n2253;
  assign n2255 = n2254 ^ n2089;
  assign n2249 = n2088 ^ n2082;
  assign n2250 = n2083 & ~n2249;
  assign n2251 = n2250 ^ n2077;
  assign n2245 = n2190 ^ n2180;
  assign n2246 = ~n2186 & n2245;
  assign n2247 = n2246 ^ n2190;
  assign n2241 = n2155 ^ n2144;
  assign n2242 = n2155 ^ n2149;
  assign n2243 = n2241 & ~n2242;
  assign n2244 = n2243 ^ n2144;
  assign n2248 = n2247 ^ n2244;
  assign n2252 = n2251 ^ n2248;
  assign n2256 = n2255 ^ n2252;
  assign n2236 = n2173 ^ n2161;
  assign n2237 = ~n2168 & n2236;
  assign n2238 = n2237 ^ n2173;
  assign n2233 = n2127 ^ n2116;
  assign n2234 = ~n2122 & n2233;
  assign n2235 = n2234 ^ n2127;
  assign n2239 = n2238 ^ n2235;
  assign n2229 = ~x15 & n567;
  assign n2230 = n2229 ^ n672;
  assign n2227 = ~x14 & n669;
  assign n2228 = n2227 ^ n738;
  assign n2231 = n2230 ^ n2228;
  assign n2223 = x23 & n157;
  assign n2224 = n2223 ^ n191;
  assign n2221 = x22 & n188;
  assign n2222 = n2221 ^ n248;
  assign n2225 = n2224 ^ n2222;
  assign n2218 = x27 & n75;
  assign n2219 = n2218 ^ n96;
  assign n2216 = x26 & n93;
  assign n2217 = n2216 ^ n108;
  assign n2220 = n2219 ^ n2217;
  assign n2226 = n2225 ^ n2220;
  assign n2232 = n2231 ^ n2226;
  assign n2240 = n2239 ^ n2232;
  assign n2257 = n2256 ^ n2240;
  assign n2290 = n2289 ^ n2257;
  assign n2353 = n2352 ^ n2290;
  assign n2361 = n2360 ^ n2353;
  assign n2365 = n2364 ^ n2361;
  assign n2369 = n2368 ^ n2365;
  assign n2518 = n2368 ^ n2361;
  assign n2519 = ~n2365 & n2518;
  assign n2520 = n2519 ^ n2368;
  assign n2514 = n2356 ^ n2353;
  assign n2515 = ~n2360 & n2514;
  assign n2516 = n2515 ^ n2353;
  assign n2510 = n2352 ^ n2289;
  assign n2511 = n2290 & ~n2510;
  assign n2512 = n2511 ^ n2257;
  assign n2504 = n2351 ^ n2343;
  assign n2505 = n2351 ^ n2347;
  assign n2506 = n2504 & ~n2505;
  assign n2507 = n2506 ^ n2343;
  assign n2499 = n2324 ^ n2307;
  assign n2500 = ~n2342 & n2499;
  assign n2501 = n2500 ^ n2307;
  assign n2495 = n2251 ^ n2244;
  assign n2496 = ~n2248 & n2495;
  assign n2497 = n2496 ^ n2251;
  assign n2491 = n2231 ^ n2225;
  assign n2492 = n2226 & ~n2491;
  assign n2493 = n2492 ^ n2220;
  assign n2487 = x2 & n2143;
  assign n2488 = n2487 ^ n2275;
  assign n2485 = x1 & n2272;
  assign n2484 = x61 & n2272;
  assign n2486 = n2485 ^ n2484;
  assign n2489 = n2488 ^ n2486;
  assign n2483 = n2260 & n2264;
  assign n2490 = n2489 ^ n2483;
  assign n2494 = n2493 ^ n2490;
  assign n2498 = n2497 ^ n2494;
  assign n2502 = n2501 ^ n2498;
  assign n2478 = n2235 ^ n2232;
  assign n2479 = ~n2239 & n2478;
  assign n2480 = n2479 ^ n2232;
  assign n2474 = n2323 ^ n2317;
  assign n2475 = n2318 & ~n2474;
  assign n2476 = n2475 ^ n2312;
  assign n2470 = n2340 ^ n2334;
  assign n2471 = n2335 & ~n2470;
  assign n2472 = n2471 ^ n2329;
  assign n2467 = n2306 ^ n2300;
  assign n2468 = n2301 & ~n2467;
  assign n2469 = n2468 ^ n2295;
  assign n2473 = n2472 ^ n2469;
  assign n2477 = n2476 ^ n2473;
  assign n2481 = n2480 ^ n2477;
  assign n2463 = n2278 ^ n2265;
  assign n2464 = n2279 & ~n2463;
  assign n2465 = n2464 ^ n2270;
  assign n2458 = x10 & n1105;
  assign n2459 = n2458 ^ n1206;
  assign n2456 = x9 & n1203;
  assign n2457 = n2456 ^ n1379;
  assign n2460 = n2459 ^ n2457;
  assign n2452 = ~x12 & n894;
  assign n2453 = n2452 ^ n1052;
  assign n2450 = ~x11 & n1049;
  assign n2451 = n2450 ^ n1087;
  assign n2454 = n2453 ^ n2451;
  assign n2447 = x22 & n241;
  assign n2448 = n2447 ^ n293;
  assign n2445 = x21 & n290;
  assign n2446 = n2445 ^ n342;
  assign n2449 = n2448 ^ n2446;
  assign n2455 = n2454 ^ n2449;
  assign n2461 = n2460 ^ n2455;
  assign n2441 = x14 & n756;
  assign n2442 = n2441 ^ n873;
  assign n2439 = x13 & n870;
  assign n2440 = n2439 ^ n953;
  assign n2443 = n2442 ^ n2440;
  assign n2435 = ~x16 & n567;
  assign n2436 = n2435 ^ n672;
  assign n2433 = ~x15 & n669;
  assign n2434 = n2433 ^ n738;
  assign n2437 = n2436 ^ n2434;
  assign n2430 = x24 & n157;
  assign n2431 = n2430 ^ n191;
  assign n2428 = x23 & n188;
  assign n2429 = n2428 ^ n248;
  assign n2432 = n2431 ^ n2429;
  assign n2438 = n2437 ^ n2432;
  assign n2444 = n2443 ^ n2438;
  assign n2462 = n2461 ^ n2444;
  assign n2466 = n2465 ^ n2462;
  assign n2482 = n2481 ^ n2466;
  assign n2503 = n2502 ^ n2482;
  assign n2508 = n2507 ^ n2503;
  assign n2423 = n2288 ^ n2280;
  assign n2424 = n2288 ^ n2283;
  assign n2425 = n2423 & ~n2424;
  assign n2426 = n2425 ^ n2280;
  assign n2419 = n2252 ^ n2240;
  assign n2420 = ~n2256 & n2419;
  assign n2421 = n2420 ^ n2240;
  assign n2413 = ~x4 & n1815;
  assign n2414 = n2413 ^ n2047;
  assign n2411 = ~x3 & n2044;
  assign n2412 = n2411 ^ n2162;
  assign n2415 = n2414 ^ n2412;
  assign n2407 = x18 & n435;
  assign n2408 = n2407 ^ n527;
  assign n2405 = x17 & n524;
  assign n2406 = n2405 ^ n611;
  assign n2409 = n2408 ^ n2406;
  assign n2402 = x6 & n1556;
  assign n2403 = n2402 ^ n1664;
  assign n2400 = x5 & n1661;
  assign n2401 = n2400 ^ n1878;
  assign n2404 = n2403 ^ n2401;
  assign n2410 = n2409 ^ n2404;
  assign n2416 = n2415 ^ n2410;
  assign n2396 = x28 & n75;
  assign n2397 = n2396 ^ n96;
  assign n2394 = x27 & n93;
  assign n2395 = n2394 ^ n108;
  assign n2398 = n2397 ^ n2395;
  assign n2390 = ~x29 & n68;
  assign n2391 = n2390 ^ n69;
  assign n2389 = x30 & x32;
  assign n2392 = n2391 ^ n2389;
  assign n2387 = x62 ^ x61;
  assign n2388 = x0 & n2387;
  assign n2393 = n2392 ^ n2388;
  assign n2399 = n2398 ^ n2393;
  assign n2417 = n2416 ^ n2399;
  assign n2383 = x8 & n1360;
  assign n2384 = n2383 ^ n1447;
  assign n2381 = x7 & n1444;
  assign n2382 = n2381 ^ n1588;
  assign n2385 = n2384 ^ n2382;
  assign n2377 = ~x20 & n322;
  assign n2378 = n2377 ^ n382;
  assign n2375 = ~x19 & n379;
  assign n2376 = n2375 ^ n459;
  assign n2379 = n2378 ^ n2376;
  assign n2372 = x26 & n106;
  assign n2373 = n2372 ^ n142;
  assign n2370 = x25 & n139;
  assign n2371 = n2370 ^ n171;
  assign n2374 = n2373 ^ n2371;
  assign n2380 = n2379 ^ n2374;
  assign n2386 = n2385 ^ n2380;
  assign n2418 = n2417 ^ n2386;
  assign n2422 = n2421 ^ n2418;
  assign n2427 = n2426 ^ n2422;
  assign n2509 = n2508 ^ n2427;
  assign n2513 = n2512 ^ n2509;
  assign n2517 = n2516 ^ n2513;
  assign n2521 = n2520 ^ n2517;
  assign n2683 = n2520 ^ n2513;
  assign n2684 = ~n2517 & n2683;
  assign n2685 = n2684 ^ n2520;
  assign n2678 = n2512 ^ n2427;
  assign n2679 = n2512 ^ n2508;
  assign n2680 = n2678 & ~n2679;
  assign n2681 = n2680 ^ n2427;
  assign n2674 = n2507 ^ n2502;
  assign n2675 = n2503 & ~n2674;
  assign n2676 = n2675 ^ n2482;
  assign n2669 = n2426 ^ n2421;
  assign n2670 = n2422 & ~n2669;
  assign n2671 = n2670 ^ n2418;
  assign n2663 = n2465 ^ n2461;
  assign n2664 = n2462 & ~n2663;
  assign n2665 = n2664 ^ n2444;
  assign n2659 = n2399 ^ n2386;
  assign n2660 = n2416 ^ n2386;
  assign n2661 = n2659 & ~n2660;
  assign n2662 = n2661 ^ n2399;
  assign n2666 = n2665 ^ n2662;
  assign n2653 = x3 & n2143;
  assign n2654 = n2653 ^ n2275;
  assign n2651 = x2 & n2272;
  assign n2652 = n2651 ^ n2484;
  assign n2655 = n2654 ^ n2652;
  assign n2647 = x19 & n435;
  assign n2648 = n2647 ^ n527;
  assign n2645 = x18 & n524;
  assign n2646 = n2645 ^ n611;
  assign n2649 = n2648 ^ n2646;
  assign n2642 = ~x5 & n1815;
  assign n2643 = n2642 ^ n2047;
  assign n2640 = ~x4 & n2044;
  assign n2641 = n2640 ^ n2162;
  assign n2644 = n2643 ^ n2641;
  assign n2650 = n2649 ^ n2644;
  assign n2656 = n2655 ^ n2650;
  assign n2636 = x1 & n2387;
  assign n2635 = x63 & n2387;
  assign n2637 = n2636 ^ n2635;
  assign n2630 = x63 ^ x62;
  assign n2631 = ~n2387 & n2630;
  assign n2633 = x0 & n2631;
  assign n2632 = x63 & n2631;
  assign n2634 = n2633 ^ n2632;
  assign n2638 = n2637 ^ n2634;
  assign n2626 = x25 & n157;
  assign n2627 = n2626 ^ n191;
  assign n2624 = x24 & n188;
  assign n2625 = n2624 ^ n248;
  assign n2628 = n2627 ^ n2625;
  assign n2621 = x29 & n75;
  assign n2622 = n2621 ^ n96;
  assign n2619 = x28 & n93;
  assign n2620 = n2619 ^ n108;
  assign n2623 = n2622 ^ n2620;
  assign n2629 = n2628 ^ n2623;
  assign n2639 = n2638 ^ n2629;
  assign n2657 = n2656 ^ n2639;
  assign n2615 = x23 & n241;
  assign n2616 = n2615 ^ n293;
  assign n2613 = x22 & n290;
  assign n2614 = n2613 ^ n342;
  assign n2617 = n2616 ^ n2614;
  assign n2609 = ~x17 & n567;
  assign n2610 = n2609 ^ n672;
  assign n2607 = ~x16 & n669;
  assign n2608 = n2607 ^ n738;
  assign n2611 = n2610 ^ n2608;
  assign n2604 = x15 & n756;
  assign n2605 = n2604 ^ n873;
  assign n2602 = x14 & n870;
  assign n2603 = n2602 ^ n953;
  assign n2606 = n2605 ^ n2603;
  assign n2612 = n2611 ^ n2606;
  assign n2618 = n2617 ^ n2612;
  assign n2658 = n2657 ^ n2618;
  assign n2667 = n2666 ^ n2658;
  assign n2597 = n2493 ^ n2483;
  assign n2598 = n2490 & ~n2597;
  assign n2599 = n2598 ^ n2489;
  assign n2593 = n2415 ^ n2409;
  assign n2594 = n2410 & ~n2593;
  assign n2595 = n2594 ^ n2404;
  assign n2589 = n2385 ^ n2379;
  assign n2590 = n2380 & ~n2589;
  assign n2591 = n2590 ^ n2374;
  assign n2586 = n2460 ^ n2454;
  assign n2587 = n2455 & ~n2586;
  assign n2588 = n2587 ^ n2449;
  assign n2592 = n2591 ^ n2588;
  assign n2596 = n2595 ^ n2592;
  assign n2600 = n2599 ^ n2596;
  assign n2582 = n2443 ^ n2437;
  assign n2583 = n2438 & ~n2582;
  assign n2584 = n2583 ^ n2432;
  assign n2578 = n2398 ^ n2392;
  assign n2579 = n2393 & ~n2578;
  assign n2580 = n2579 ^ n2388;
  assign n2574 = ~x30 & n68;
  assign n2575 = n2574 ^ n69;
  assign n2573 = x31 & x32;
  assign n2576 = n2575 ^ n2573;
  assign n2570 = n2273 & ~n2387;
  assign n2571 = n2570 ^ x0;
  assign n2572 = x63 & ~n2571;
  assign n2577 = n2576 ^ n2572;
  assign n2581 = n2580 ^ n2577;
  assign n2585 = n2584 ^ n2581;
  assign n2601 = n2600 ^ n2585;
  assign n2668 = n2667 ^ n2601;
  assign n2672 = n2671 ^ n2668;
  assign n2566 = n2477 ^ n2466;
  assign n2567 = ~n2481 & n2566;
  assign n2568 = n2567 ^ n2466;
  assign n2561 = n2501 ^ n2494;
  assign n2562 = n2501 ^ n2497;
  assign n2563 = n2561 & ~n2562;
  assign n2564 = n2563 ^ n2494;
  assign n2557 = n2476 ^ n2469;
  assign n2558 = ~n2473 & n2557;
  assign n2559 = n2558 ^ n2476;
  assign n2552 = x27 & n106;
  assign n2553 = n2552 ^ n142;
  assign n2550 = x26 & n139;
  assign n2551 = n2550 ^ n171;
  assign n2554 = n2553 ^ n2551;
  assign n2546 = x11 & n1105;
  assign n2547 = n2546 ^ n1206;
  assign n2544 = x10 & n1203;
  assign n2545 = n2544 ^ n1379;
  assign n2548 = n2547 ^ n2545;
  assign n2541 = ~x13 & n894;
  assign n2542 = n2541 ^ n1052;
  assign n2539 = ~x12 & n1049;
  assign n2540 = n2539 ^ n1087;
  assign n2543 = n2542 ^ n2540;
  assign n2549 = n2548 ^ n2543;
  assign n2555 = n2554 ^ n2549;
  assign n2535 = x7 & n1556;
  assign n2536 = n2535 ^ n1664;
  assign n2533 = x6 & n1661;
  assign n2534 = n2533 ^ n1878;
  assign n2537 = n2536 ^ n2534;
  assign n2529 = ~x21 & n322;
  assign n2530 = n2529 ^ n382;
  assign n2527 = ~x20 & n379;
  assign n2528 = n2527 ^ n459;
  assign n2531 = n2530 ^ n2528;
  assign n2524 = x9 & n1360;
  assign n2525 = n2524 ^ n1447;
  assign n2522 = x8 & n1444;
  assign n2523 = n2522 ^ n1588;
  assign n2526 = n2525 ^ n2523;
  assign n2532 = n2531 ^ n2526;
  assign n2538 = n2537 ^ n2532;
  assign n2556 = n2555 ^ n2538;
  assign n2560 = n2559 ^ n2556;
  assign n2565 = n2564 ^ n2560;
  assign n2569 = n2568 ^ n2565;
  assign n2673 = n2672 ^ n2569;
  assign n2677 = n2676 ^ n2673;
  assign n2682 = n2681 ^ n2677;
  assign n2686 = n2685 ^ n2682;
  assign n2840 = n2685 ^ n2677;
  assign n2841 = ~n2682 & n2840;
  assign n2842 = n2841 ^ n2685;
  assign n2836 = n2676 ^ n2672;
  assign n2837 = n2673 & ~n2836;
  assign n2838 = n2837 ^ n2569;
  assign n2831 = n2671 ^ n2667;
  assign n2832 = n2668 & ~n2831;
  assign n2833 = n2832 ^ n2601;
  assign n2828 = n2568 ^ n2564;
  assign n2829 = n2565 & ~n2828;
  assign n2830 = n2829 ^ n2560;
  assign n2834 = n2833 ^ n2830;
  assign n2823 = n2662 ^ n2658;
  assign n2824 = ~n2666 & n2823;
  assign n2825 = n2824 ^ n2658;
  assign n2819 = n2596 ^ n2585;
  assign n2820 = ~n2600 & n2819;
  assign n2821 = n2820 ^ n2585;
  assign n2815 = n2595 ^ n2591;
  assign n2816 = n2592 & ~n2815;
  assign n2817 = n2816 ^ n2588;
  assign n2810 = ~x18 & n567;
  assign n2811 = n2810 ^ n672;
  assign n2808 = ~x17 & n669;
  assign n2809 = n2808 ^ n738;
  assign n2812 = n2811 ^ n2809;
  assign n2804 = x26 & n157;
  assign n2805 = n2804 ^ n191;
  assign n2802 = x25 & n188;
  assign n2803 = n2802 ^ n248;
  assign n2806 = n2805 ^ n2803;
  assign n2799 = x2 & n2387;
  assign n2800 = n2799 ^ n2635;
  assign n2797 = x1 & n2631;
  assign n2798 = n2797 ^ n2632;
  assign n2801 = n2800 ^ n2798;
  assign n2807 = n2806 ^ n2801;
  assign n2813 = n2812 ^ n2807;
  assign n2792 = x4 & n2143;
  assign n2793 = n2792 ^ n2275;
  assign n2790 = x3 & n2272;
  assign n2791 = n2790 ^ n2484;
  assign n2794 = n2793 ^ n2791;
  assign n2787 = ~x6 & n1815;
  assign n2788 = n2787 ^ n2047;
  assign n2785 = ~x5 & n2044;
  assign n2786 = n2785 ^ n2162;
  assign n2789 = n2788 ^ n2786;
  assign n2795 = n2794 ^ n2789;
  assign n2784 = n2572 & n2576;
  assign n2796 = n2795 ^ n2784;
  assign n2814 = n2813 ^ n2796;
  assign n2818 = n2817 ^ n2814;
  assign n2822 = n2821 ^ n2818;
  assign n2826 = n2825 ^ n2822;
  assign n2779 = n2559 ^ n2555;
  assign n2780 = n2556 & ~n2779;
  assign n2781 = n2780 ^ n2538;
  assign n2773 = n2554 ^ n2543;
  assign n2774 = n2554 ^ n2548;
  assign n2775 = n2773 & ~n2774;
  assign n2776 = n2775 ^ n2543;
  assign n2769 = n2638 ^ n2628;
  assign n2770 = n2629 & ~n2769;
  assign n2771 = n2770 ^ n2623;
  assign n2766 = n2617 ^ n2606;
  assign n2767 = ~n2612 & n2766;
  assign n2768 = n2767 ^ n2617;
  assign n2772 = n2771 ^ n2768;
  assign n2777 = n2776 ^ n2772;
  assign n2760 = ~x22 & n322;
  assign n2761 = n2760 ^ n382;
  assign n2758 = ~x21 & n379;
  assign n2759 = n2758 ^ n459;
  assign n2762 = n2761 ^ n2759;
  assign n2754 = x12 & n1105;
  assign n2755 = n2754 ^ n1206;
  assign n2752 = x11 & n1203;
  assign n2753 = n2752 ^ n1379;
  assign n2756 = n2755 ^ n2753;
  assign n2749 = x28 & n106;
  assign n2750 = n2749 ^ n142;
  assign n2747 = x27 & n139;
  assign n2748 = n2747 ^ n171;
  assign n2751 = n2750 ^ n2748;
  assign n2757 = n2756 ^ n2751;
  assign n2763 = n2762 ^ n2757;
  assign n2743 = ~x14 & n894;
  assign n2744 = n2743 ^ n1052;
  assign n2741 = ~x13 & n1049;
  assign n2742 = n2741 ^ n1087;
  assign n2745 = n2744 ^ n2742;
  assign n2737 = x16 & n756;
  assign n2738 = n2737 ^ n873;
  assign n2735 = x15 & n870;
  assign n2736 = n2735 ^ n953;
  assign n2739 = n2738 ^ n2736;
  assign n2732 = x24 & n241;
  assign n2733 = n2732 ^ n293;
  assign n2730 = x23 & n290;
  assign n2731 = n2730 ^ n342;
  assign n2734 = n2733 ^ n2731;
  assign n2740 = n2739 ^ n2734;
  assign n2746 = n2745 ^ n2740;
  assign n2764 = n2763 ^ n2746;
  assign n2726 = x20 & n435;
  assign n2727 = n2726 ^ n527;
  assign n2724 = x19 & n524;
  assign n2725 = n2724 ^ n611;
  assign n2728 = n2727 ^ n2725;
  assign n2720 = x8 & n1556;
  assign n2721 = n2720 ^ n1664;
  assign n2718 = x7 & n1661;
  assign n2719 = n2718 ^ n1878;
  assign n2722 = n2721 ^ n2719;
  assign n2715 = x10 & n1360;
  assign n2716 = n2715 ^ n1447;
  assign n2713 = x9 & n1444;
  assign n2714 = n2713 ^ n1588;
  assign n2717 = n2716 ^ n2714;
  assign n2723 = n2722 ^ n2717;
  assign n2729 = n2728 ^ n2723;
  assign n2765 = n2764 ^ n2729;
  assign n2778 = n2777 ^ n2765;
  assign n2782 = n2781 ^ n2778;
  assign n2708 = n2584 ^ n2580;
  assign n2709 = n2581 & ~n2708;
  assign n2710 = n2709 ^ n2577;
  assign n2705 = n2639 ^ n2618;
  assign n2706 = ~n2657 & n2705;
  assign n2707 = n2706 ^ n2618;
  assign n2711 = n2710 ^ n2707;
  assign n2700 = n2655 ^ n2644;
  assign n2701 = ~n2650 & n2700;
  assign n2702 = n2701 ^ n2655;
  assign n2697 = n2537 ^ n2526;
  assign n2698 = ~n2532 & n2697;
  assign n2699 = n2698 ^ n2537;
  assign n2703 = n2702 ^ n2699;
  assign n2693 = x30 & n75;
  assign n2694 = n2693 ^ n96;
  assign n2691 = x29 & n93;
  assign n2692 = n2691 ^ n108;
  assign n2695 = n2694 ^ n2692;
  assign n2688 = x31 & n68;
  assign n2689 = n2688 ^ x33;
  assign n2687 = x0 & x63;
  assign n2690 = n2689 ^ n2687;
  assign n2696 = n2695 ^ n2690;
  assign n2704 = n2703 ^ n2696;
  assign n2712 = n2711 ^ n2704;
  assign n2783 = n2782 ^ n2712;
  assign n2827 = n2826 ^ n2783;
  assign n2835 = n2834 ^ n2827;
  assign n2839 = n2838 ^ n2835;
  assign n2843 = n2842 ^ n2839;
  assign n3000 = n2842 ^ n2835;
  assign n3001 = ~n2839 & n3000;
  assign n3002 = n3001 ^ n2842;
  assign n2996 = n2830 ^ n2827;
  assign n2997 = ~n2834 & n2996;
  assign n2998 = n2997 ^ n2827;
  assign n2992 = n2826 ^ n2782;
  assign n2993 = n2783 & ~n2992;
  assign n2994 = n2993 ^ n2712;
  assign n2987 = n2825 ^ n2821;
  assign n2988 = n2822 & ~n2987;
  assign n2989 = n2988 ^ n2818;
  assign n2983 = n2781 ^ n2777;
  assign n2984 = n2778 & ~n2983;
  assign n2985 = n2984 ^ n2765;
  assign n2979 = n2817 ^ n2813;
  assign n2980 = n2814 & ~n2979;
  assign n2981 = n2980 ^ n2796;
  assign n2972 = n2762 ^ n2751;
  assign n2973 = n2762 ^ n2756;
  assign n2974 = n2972 & ~n2973;
  assign n2975 = n2974 ^ n2751;
  assign n2967 = x3 & n2387;
  assign n2968 = n2967 ^ n2635;
  assign n2965 = x2 & n2631;
  assign n2966 = n2965 ^ n2632;
  assign n2969 = n2968 ^ n2966;
  assign n2962 = ~x19 & n567;
  assign n2963 = n2962 ^ n672;
  assign n2960 = ~x18 & n669;
  assign n2961 = n2960 ^ n738;
  assign n2964 = n2963 ^ n2961;
  assign n2970 = n2969 ^ n2964;
  assign n2959 = x1 & x63;
  assign n2971 = n2970 ^ n2959;
  assign n2976 = n2975 ^ n2971;
  assign n2955 = ~x7 & n1815;
  assign n2956 = n2955 ^ n2047;
  assign n2953 = ~x6 & n2044;
  assign n2954 = n2953 ^ n2162;
  assign n2957 = n2956 ^ n2954;
  assign n2949 = x9 & n1556;
  assign n2950 = n2949 ^ n1664;
  assign n2947 = x8 & n1661;
  assign n2948 = n2947 ^ n1878;
  assign n2951 = n2950 ^ n2948;
  assign n2944 = x21 & n435;
  assign n2945 = n2944 ^ n527;
  assign n2942 = x20 & n524;
  assign n2943 = n2942 ^ n611;
  assign n2946 = n2945 ^ n2943;
  assign n2952 = n2951 ^ n2946;
  assign n2958 = n2957 ^ n2952;
  assign n2977 = n2976 ^ n2958;
  assign n2936 = x27 & n157;
  assign n2937 = n2936 ^ n191;
  assign n2934 = x26 & n188;
  assign n2935 = n2934 ^ n248;
  assign n2938 = n2937 ^ n2935;
  assign n2930 = x17 & n756;
  assign n2931 = n2930 ^ n873;
  assign n2928 = x16 & n870;
  assign n2929 = n2928 ^ n953;
  assign n2932 = n2931 ^ n2929;
  assign n2925 = x31 & n75;
  assign n2926 = n2925 ^ n96;
  assign n2923 = x30 & n93;
  assign n2924 = n2923 ^ n108;
  assign n2927 = n2926 ^ n2924;
  assign n2933 = n2932 ^ n2927;
  assign n2939 = n2938 ^ n2933;
  assign n2919 = x11 & n1360;
  assign n2920 = n2919 ^ n1447;
  assign n2917 = x10 & n1444;
  assign n2918 = n2917 ^ n1588;
  assign n2921 = n2920 ^ n2918;
  assign n2913 = ~x23 & n322;
  assign n2914 = n2913 ^ n382;
  assign n2911 = ~x22 & n379;
  assign n2912 = n2911 ^ n459;
  assign n2915 = n2914 ^ n2912;
  assign n2908 = x29 & n106;
  assign n2909 = n2908 ^ n142;
  assign n2906 = x28 & n139;
  assign n2907 = n2906 ^ n171;
  assign n2910 = n2909 ^ n2907;
  assign n2916 = n2915 ^ n2910;
  assign n2922 = n2921 ^ n2916;
  assign n2940 = n2939 ^ n2922;
  assign n2902 = x13 & n1105;
  assign n2903 = n2902 ^ n1206;
  assign n2900 = x12 & n1203;
  assign n2901 = n2900 ^ n1379;
  assign n2904 = n2903 ^ n2901;
  assign n2896 = x25 & n241;
  assign n2897 = n2896 ^ n293;
  assign n2894 = x24 & n290;
  assign n2895 = n2894 ^ n342;
  assign n2898 = n2897 ^ n2895;
  assign n2891 = ~x15 & n894;
  assign n2892 = n2891 ^ n1052;
  assign n2889 = ~x14 & n1049;
  assign n2890 = n2889 ^ n1087;
  assign n2893 = n2892 ^ n2890;
  assign n2899 = n2898 ^ n2893;
  assign n2905 = n2904 ^ n2899;
  assign n2941 = n2940 ^ n2905;
  assign n2978 = n2977 ^ n2941;
  assign n2982 = n2981 ^ n2978;
  assign n2986 = n2985 ^ n2982;
  assign n2990 = n2989 ^ n2986;
  assign n2883 = n2707 ^ n2704;
  assign n2884 = n2710 ^ n2704;
  assign n2885 = n2883 & ~n2884;
  assign n2886 = n2885 ^ n2707;
  assign n2879 = n2699 ^ n2696;
  assign n2880 = ~n2703 & n2879;
  assign n2881 = n2880 ^ n2696;
  assign n2875 = n2776 ^ n2771;
  assign n2876 = n2772 & ~n2875;
  assign n2877 = n2876 ^ n2768;
  assign n2872 = n2794 ^ n2784;
  assign n2873 = n2795 & ~n2872;
  assign n2874 = n2873 ^ n2789;
  assign n2878 = n2877 ^ n2874;
  assign n2882 = n2881 ^ n2878;
  assign n2887 = n2886 ^ n2882;
  assign n2868 = n2763 ^ n2729;
  assign n2869 = n2764 & ~n2868;
  assign n2870 = n2869 ^ n2746;
  assign n2862 = n2728 ^ n2717;
  assign n2863 = n2728 ^ n2722;
  assign n2864 = n2862 & ~n2863;
  assign n2865 = n2864 ^ n2717;
  assign n2858 = n2745 ^ n2739;
  assign n2859 = n2740 & ~n2858;
  assign n2860 = n2859 ^ n2734;
  assign n2854 = n2812 ^ n2801;
  assign n2855 = n2812 ^ n2806;
  assign n2856 = n2854 & ~n2855;
  assign n2857 = n2856 ^ n2801;
  assign n2861 = n2860 ^ n2857;
  assign n2866 = n2865 ^ n2861;
  assign n2850 = n2695 ^ n2689;
  assign n2851 = n2690 & ~n2850;
  assign n2852 = n2851 ^ n2687;
  assign n2846 = x5 & n2143;
  assign n2847 = n2846 ^ n2275;
  assign n2844 = x4 & n2272;
  assign n2845 = n2844 ^ n2484;
  assign n2848 = n2847 ^ n2845;
  assign n2849 = n2848 ^ x33;
  assign n2853 = n2852 ^ n2849;
  assign n2867 = n2866 ^ n2853;
  assign n2871 = n2870 ^ n2867;
  assign n2888 = n2887 ^ n2871;
  assign n2991 = n2990 ^ n2888;
  assign n2995 = n2994 ^ n2991;
  assign n2999 = n2998 ^ n2995;
  assign n3003 = n3002 ^ n2999;
  assign n3158 = n3002 ^ n2995;
  assign n3159 = ~n2999 & n3158;
  assign n3160 = n3159 ^ n3002;
  assign n3154 = n2994 ^ n2990;
  assign n3155 = n2991 & ~n3154;
  assign n3156 = n3155 ^ n2888;
  assign n3150 = n2989 ^ n2985;
  assign n3151 = n2986 & ~n3150;
  assign n3152 = n3151 ^ n2982;
  assign n3145 = n2882 ^ n2871;
  assign n3146 = ~n2887 & n3145;
  assign n3147 = n3146 ^ n2871;
  assign n3141 = n2981 ^ n2977;
  assign n3142 = n2978 & ~n3141;
  assign n3143 = n3142 ^ n2941;
  assign n3136 = n2870 ^ n2853;
  assign n3137 = n2870 ^ n2866;
  assign n3138 = n3136 & ~n3137;
  assign n3139 = n3138 ^ n2853;
  assign n3129 = n2957 ^ n2946;
  assign n3130 = n2957 ^ n2951;
  assign n3131 = n3129 & ~n3130;
  assign n3132 = n3131 ^ n2946;
  assign n3125 = x4 & n2387;
  assign n3126 = n3125 ^ n2635;
  assign n3123 = x3 & n2631;
  assign n3124 = n3123 ^ n2632;
  assign n3127 = n3126 ^ n3124;
  assign n3119 = ~x20 & n567;
  assign n3120 = n3119 ^ n672;
  assign n3117 = ~x19 & n669;
  assign n3118 = n3117 ^ n738;
  assign n3121 = n3120 ^ n3118;
  assign n3114 = x6 & n2143;
  assign n3115 = n3114 ^ n2275;
  assign n3112 = x5 & n2272;
  assign n3113 = n3112 ^ n2484;
  assign n3116 = n3115 ^ n3113;
  assign n3122 = n3121 ^ n3116;
  assign n3128 = n3127 ^ n3122;
  assign n3133 = n3132 ^ n3128;
  assign n3108 = ~x24 & n322;
  assign n3109 = n3108 ^ n382;
  assign n3106 = ~x23 & n379;
  assign n3107 = n3106 ^ n459;
  assign n3110 = n3109 ^ n3107;
  assign n3102 = ~x16 & n894;
  assign n3103 = n3102 ^ n1052;
  assign n3100 = ~x15 & n1049;
  assign n3101 = n3100 ^ n1087;
  assign n3104 = n3103 ^ n3101;
  assign n3097 = x18 & n756;
  assign n3098 = n3097 ^ n873;
  assign n3095 = x17 & n870;
  assign n3096 = n3095 ^ n953;
  assign n3099 = n3098 ^ n3096;
  assign n3105 = n3104 ^ n3099;
  assign n3111 = n3110 ^ n3105;
  assign n3134 = n3133 ^ n3111;
  assign n3089 = x28 & n157;
  assign n3090 = n3089 ^ n191;
  assign n3087 = x27 & n188;
  assign n3088 = n3087 ^ n248;
  assign n3091 = n3090 ^ n3088;
  assign n3083 = x14 & n1105;
  assign n3084 = n3083 ^ n1206;
  assign n3081 = x13 & n1203;
  assign n3082 = n3081 ^ n1379;
  assign n3085 = n3084 ^ n3082;
  assign n3078 = x12 & n1360;
  assign n3079 = n3078 ^ n1447;
  assign n3076 = x11 & n1444;
  assign n3077 = n3076 ^ n1588;
  assign n3080 = n3079 ^ n3077;
  assign n3086 = n3085 ^ n3080;
  assign n3092 = n3091 ^ n3086;
  assign n3071 = x30 & n106;
  assign n3072 = n3071 ^ n142;
  assign n3069 = x29 & n139;
  assign n3070 = n3069 ^ n171;
  assign n3073 = n3072 ^ n3070;
  assign n3066 = x26 & n241;
  assign n3067 = n3066 ^ n293;
  assign n3064 = x25 & n290;
  assign n3065 = n3064 ^ n342;
  assign n3068 = n3067 ^ n3065;
  assign n3074 = n3073 ^ n3068;
  assign n3063 = x2 & x63;
  assign n3075 = n3074 ^ n3063;
  assign n3093 = n3092 ^ n3075;
  assign n3059 = ~x8 & n1815;
  assign n3060 = n3059 ^ n2047;
  assign n3057 = ~x7 & n2044;
  assign n3058 = n3057 ^ n2162;
  assign n3061 = n3060 ^ n3058;
  assign n3053 = x10 & n1556;
  assign n3054 = n3053 ^ n1664;
  assign n3051 = x9 & n1661;
  assign n3052 = n3051 ^ n1878;
  assign n3055 = n3054 ^ n3052;
  assign n3048 = x22 & n435;
  assign n3049 = n3048 ^ n527;
  assign n3046 = x21 & n524;
  assign n3047 = n3046 ^ n611;
  assign n3050 = n3049 ^ n3047;
  assign n3056 = n3055 ^ n3050;
  assign n3062 = n3061 ^ n3056;
  assign n3094 = n3093 ^ n3062;
  assign n3135 = n3134 ^ n3094;
  assign n3140 = n3139 ^ n3135;
  assign n3144 = n3143 ^ n3140;
  assign n3148 = n3147 ^ n3144;
  assign n3040 = n2881 ^ n2874;
  assign n3041 = n2881 ^ n2877;
  assign n3042 = n3040 & ~n3041;
  assign n3043 = n3042 ^ n2874;
  assign n3035 = n2865 ^ n2857;
  assign n3036 = ~n2861 & n3035;
  assign n3037 = n3036 ^ n2865;
  assign n3032 = n2852 ^ n2848;
  assign n3033 = n2849 & ~n3032;
  assign n3034 = n3033 ^ x33;
  assign n3038 = n3037 ^ n3034;
  assign n3028 = n2921 ^ n2910;
  assign n3029 = ~n2916 & n3028;
  assign n3030 = n3029 ^ n2921;
  assign n3024 = n2938 ^ n2927;
  assign n3025 = ~n2933 & n3024;
  assign n3026 = n3025 ^ n2938;
  assign n3021 = n2904 ^ n2898;
  assign n3022 = n2899 & ~n3021;
  assign n3023 = n3022 ^ n2893;
  assign n3027 = n3026 ^ n3023;
  assign n3031 = n3030 ^ n3027;
  assign n3039 = n3038 ^ n3031;
  assign n3044 = n3043 ^ n3039;
  assign n3016 = n2922 ^ n2905;
  assign n3017 = n2939 ^ n2905;
  assign n3018 = n3016 & ~n3017;
  assign n3019 = n3018 ^ n2922;
  assign n3012 = n2971 ^ n2958;
  assign n3013 = ~n2976 & n3012;
  assign n3014 = n3013 ^ n2958;
  assign n3008 = n2964 ^ n2959;
  assign n3009 = ~n2970 & n3008;
  assign n3010 = n3009 ^ n2959;
  assign n3004 = x31 & n93;
  assign n3005 = n3004 ^ n96;
  assign n3006 = n3005 ^ n108;
  assign n3007 = n3006 ^ x33;
  assign n3011 = n3010 ^ n3007;
  assign n3015 = n3014 ^ n3011;
  assign n3020 = n3019 ^ n3015;
  assign n3045 = n3044 ^ n3020;
  assign n3149 = n3148 ^ n3045;
  assign n3153 = n3152 ^ n3149;
  assign n3157 = n3156 ^ n3153;
  assign n3161 = n3160 ^ n3157;
  assign n3314 = n3160 ^ n3153;
  assign n3315 = ~n3157 & n3314;
  assign n3316 = n3315 ^ n3160;
  assign n3310 = n3152 ^ n3148;
  assign n3311 = n3149 & ~n3310;
  assign n3312 = n3311 ^ n3045;
  assign n3305 = n3147 ^ n3140;
  assign n3306 = n3147 ^ n3143;
  assign n3307 = n3305 & ~n3306;
  assign n3308 = n3307 ^ n3140;
  assign n3300 = n3039 ^ n3020;
  assign n3301 = ~n3044 & n3300;
  assign n3302 = n3301 ^ n3020;
  assign n3296 = n3139 ^ n3134;
  assign n3297 = n3135 & ~n3296;
  assign n3298 = n3297 ^ n3094;
  assign n3291 = n3010 ^ n3006;
  assign n3292 = n3007 & n3291;
  assign n3293 = n3292 ^ x33;
  assign n3287 = n3030 ^ n3026;
  assign n3288 = n3027 & ~n3287;
  assign n3289 = n3288 ^ n3023;
  assign n3283 = n3068 ^ n3063;
  assign n3284 = ~n3074 & n3283;
  assign n3285 = n3284 ^ n3063;
  assign n3279 = x5 & n2387;
  assign n3280 = n3279 ^ n2635;
  assign n3277 = x4 & n2631;
  assign n3278 = n3277 ^ n2632;
  assign n3281 = n3280 ^ n3278;
  assign n3282 = n3281 ^ n3006;
  assign n3286 = n3285 ^ n3282;
  assign n3290 = n3289 ^ n3286;
  assign n3294 = n3293 ^ n3290;
  assign n3271 = n3127 ^ n3116;
  assign n3272 = ~n3122 & n3271;
  assign n3273 = n3272 ^ n3127;
  assign n3267 = ~x17 & n894;
  assign n3268 = n3267 ^ n1052;
  assign n3265 = ~x16 & n1049;
  assign n3266 = n3265 ^ n1087;
  assign n3269 = n3268 ^ n3266;
  assign n3261 = x19 & n756;
  assign n3262 = n3261 ^ n873;
  assign n3259 = x18 & n870;
  assign n3260 = n3259 ^ n953;
  assign n3263 = n3262 ^ n3260;
  assign n3258 = x3 & x63;
  assign n3264 = n3263 ^ n3258;
  assign n3270 = n3269 ^ n3264;
  assign n3274 = n3273 ^ n3270;
  assign n3254 = x27 & n241;
  assign n3255 = n3254 ^ n293;
  assign n3252 = x26 & n290;
  assign n3253 = n3252 ^ n342;
  assign n3256 = n3255 ^ n3253;
  assign n3248 = x31 & n106;
  assign n3249 = n3248 ^ n142;
  assign n3246 = x30 & n139;
  assign n3247 = n3246 ^ n171;
  assign n3250 = n3249 ^ n3247;
  assign n3245 = n108 ^ n96;
  assign n3251 = n3250 ^ n3245;
  assign n3257 = n3256 ^ n3251;
  assign n3275 = n3274 ^ n3257;
  assign n3239 = x13 & n1360;
  assign n3240 = n3239 ^ n1447;
  assign n3237 = x12 & n1444;
  assign n3238 = n3237 ^ n1588;
  assign n3241 = n3240 ^ n3238;
  assign n3233 = x15 & n1105;
  assign n3234 = n3233 ^ n1206;
  assign n3231 = x14 & n1203;
  assign n3232 = n3231 ^ n1379;
  assign n3235 = n3234 ^ n3232;
  assign n3228 = ~x25 & n322;
  assign n3229 = n3228 ^ n382;
  assign n3226 = ~x24 & n379;
  assign n3227 = n3226 ^ n459;
  assign n3230 = n3229 ^ n3227;
  assign n3236 = n3235 ^ n3230;
  assign n3242 = n3241 ^ n3236;
  assign n3222 = x7 & n2143;
  assign n3223 = n3222 ^ n2275;
  assign n3220 = x6 & n2272;
  assign n3221 = n3220 ^ n2484;
  assign n3224 = n3223 ^ n3221;
  assign n3216 = ~x9 & n1815;
  assign n3217 = n3216 ^ n2047;
  assign n3214 = ~x8 & n2044;
  assign n3215 = n3214 ^ n2162;
  assign n3218 = n3217 ^ n3215;
  assign n3211 = ~x21 & n567;
  assign n3212 = n3211 ^ n672;
  assign n3209 = ~x20 & n669;
  assign n3210 = n3209 ^ n738;
  assign n3213 = n3212 ^ n3210;
  assign n3219 = n3218 ^ n3213;
  assign n3225 = n3224 ^ n3219;
  assign n3243 = n3242 ^ n3225;
  assign n3205 = x11 & n1556;
  assign n3206 = n3205 ^ n1664;
  assign n3203 = x10 & n1661;
  assign n3204 = n3203 ^ n1878;
  assign n3207 = n3206 ^ n3204;
  assign n3199 = x23 & n435;
  assign n3200 = n3199 ^ n527;
  assign n3197 = x22 & n524;
  assign n3198 = n3197 ^ n611;
  assign n3201 = n3200 ^ n3198;
  assign n3194 = x29 & n157;
  assign n3195 = n3194 ^ n191;
  assign n3192 = x28 & n188;
  assign n3193 = n3192 ^ n248;
  assign n3196 = n3195 ^ n3193;
  assign n3202 = n3201 ^ n3196;
  assign n3208 = n3207 ^ n3202;
  assign n3244 = n3243 ^ n3208;
  assign n3276 = n3275 ^ n3244;
  assign n3295 = n3294 ^ n3276;
  assign n3299 = n3298 ^ n3295;
  assign n3303 = n3302 ^ n3299;
  assign n3187 = n3034 ^ n3031;
  assign n3188 = ~n3038 & n3187;
  assign n3189 = n3188 ^ n3031;
  assign n3183 = n3019 ^ n3011;
  assign n3184 = n3019 ^ n3014;
  assign n3185 = n3183 & ~n3184;
  assign n3186 = n3185 ^ n3011;
  assign n3190 = n3189 ^ n3186;
  assign n3178 = n3128 ^ n3111;
  assign n3179 = n3132 ^ n3111;
  assign n3180 = n3178 & ~n3179;
  assign n3181 = n3180 ^ n3128;
  assign n3173 = n3075 ^ n3062;
  assign n3174 = n3092 ^ n3062;
  assign n3175 = n3173 & ~n3174;
  assign n3176 = n3175 ^ n3075;
  assign n3169 = n3061 ^ n3055;
  assign n3170 = n3056 & ~n3169;
  assign n3171 = n3170 ^ n3050;
  assign n3165 = n3110 ^ n3104;
  assign n3166 = n3105 & ~n3165;
  assign n3167 = n3166 ^ n3099;
  assign n3162 = n3091 ^ n3080;
  assign n3163 = ~n3086 & n3162;
  assign n3164 = n3163 ^ n3091;
  assign n3168 = n3167 ^ n3164;
  assign n3172 = n3171 ^ n3168;
  assign n3177 = n3176 ^ n3172;
  assign n3182 = n3181 ^ n3177;
  assign n3191 = n3190 ^ n3182;
  assign n3304 = n3303 ^ n3191;
  assign n3309 = n3308 ^ n3304;
  assign n3313 = n3312 ^ n3309;
  assign n3317 = n3316 ^ n3313;
  assign n3468 = n3316 ^ n3309;
  assign n3469 = ~n3313 & n3468;
  assign n3470 = n3469 ^ n3316;
  assign n3464 = n3308 ^ n3303;
  assign n3465 = n3304 & ~n3464;
  assign n3466 = n3465 ^ n3191;
  assign n3460 = n3302 ^ n3298;
  assign n3461 = n3299 & ~n3460;
  assign n3462 = n3461 ^ n3295;
  assign n3455 = n3186 ^ n3182;
  assign n3456 = ~n3190 & n3455;
  assign n3457 = n3456 ^ n3182;
  assign n3451 = n3294 ^ n3275;
  assign n3452 = ~n3276 & ~n3451;
  assign n3453 = n3452 ^ n3244;
  assign n3446 = n3293 ^ n3286;
  assign n3447 = n3293 ^ n3289;
  assign n3448 = ~n3446 & n3447;
  assign n3449 = n3448 ^ n3286;
  assign n3442 = n3225 ^ n3208;
  assign n3443 = ~n3243 & n3442;
  assign n3444 = n3443 ^ n3208;
  assign n3436 = x14 & n1360;
  assign n3437 = n3436 ^ n1447;
  assign n3434 = x13 & n1444;
  assign n3435 = n3434 ^ n1588;
  assign n3438 = n3437 ^ n3435;
  assign n3430 = x24 & n435;
  assign n3431 = n3430 ^ n527;
  assign n3428 = x23 & n524;
  assign n3429 = n3428 ^ n611;
  assign n3432 = n3431 ^ n3429;
  assign n3425 = x16 & n1105;
  assign n3426 = n3425 ^ n1206;
  assign n3423 = x15 & n1203;
  assign n3424 = n3423 ^ n1379;
  assign n3427 = n3426 ^ n3424;
  assign n3433 = n3432 ^ n3427;
  assign n3439 = n3438 ^ n3433;
  assign n3419 = x20 & n756;
  assign n3420 = n3419 ^ n873;
  assign n3417 = x19 & n870;
  assign n3418 = n3417 ^ n953;
  assign n3421 = n3420 ^ n3418;
  assign n3413 = x8 & n2143;
  assign n3414 = n3413 ^ n2275;
  assign n3411 = x7 & n2272;
  assign n3412 = n3411 ^ n2484;
  assign n3415 = n3414 ^ n3412;
  assign n3408 = ~x10 & n1815;
  assign n3409 = n3408 ^ n2047;
  assign n3406 = ~x9 & n2044;
  assign n3407 = n3406 ^ n2162;
  assign n3410 = n3409 ^ n3407;
  assign n3416 = n3415 ^ n3410;
  assign n3422 = n3421 ^ n3416;
  assign n3440 = n3439 ^ n3422;
  assign n3402 = ~x22 & n567;
  assign n3403 = n3402 ^ n672;
  assign n3400 = ~x21 & n669;
  assign n3401 = n3400 ^ n738;
  assign n3404 = n3403 ^ n3401;
  assign n3396 = x12 & n1556;
  assign n3397 = n3396 ^ n1664;
  assign n3394 = x11 & n1661;
  assign n3395 = n3394 ^ n1878;
  assign n3398 = n3397 ^ n3395;
  assign n3391 = x28 & n241;
  assign n3392 = n3391 ^ n293;
  assign n3389 = x27 & n290;
  assign n3390 = n3389 ^ n342;
  assign n3393 = n3392 ^ n3390;
  assign n3399 = n3398 ^ n3393;
  assign n3405 = n3404 ^ n3399;
  assign n3441 = n3440 ^ n3405;
  assign n3445 = n3444 ^ n3441;
  assign n3450 = n3449 ^ n3445;
  assign n3454 = n3453 ^ n3450;
  assign n3458 = n3457 ^ n3454;
  assign n3384 = n3181 ^ n3176;
  assign n3385 = n3177 & ~n3384;
  assign n3386 = n3385 ^ n3172;
  assign n3380 = n3285 ^ n3281;
  assign n3381 = n3282 & ~n3380;
  assign n3382 = n3381 ^ n3006;
  assign n3375 = n3171 ^ n3164;
  assign n3376 = n3171 ^ n3167;
  assign n3377 = n3375 & ~n3376;
  assign n3378 = n3377 ^ n3164;
  assign n3371 = x31 & n139;
  assign n3372 = n3371 ^ n142;
  assign n3373 = n3372 ^ n171;
  assign n3367 = x6 & n2387;
  assign n3368 = n3367 ^ n2635;
  assign n3365 = x5 & n2631;
  assign n3366 = n3365 ^ n2632;
  assign n3369 = n3368 ^ n3366;
  assign n3364 = x4 & x63;
  assign n3370 = n3369 ^ n3364;
  assign n3374 = n3373 ^ n3370;
  assign n3379 = n3378 ^ n3374;
  assign n3383 = n3382 ^ n3379;
  assign n3387 = n3386 ^ n3383;
  assign n3358 = n3270 ^ n3257;
  assign n3359 = n3273 ^ n3257;
  assign n3360 = ~n3358 & n3359;
  assign n3361 = n3360 ^ n3270;
  assign n3353 = n3241 ^ n3230;
  assign n3354 = n3241 ^ n3235;
  assign n3355 = n3353 & ~n3354;
  assign n3356 = n3355 ^ n3230;
  assign n3348 = n3269 ^ n3258;
  assign n3349 = n3269 ^ n3263;
  assign n3350 = n3348 & ~n3349;
  assign n3351 = n3350 ^ n3258;
  assign n3344 = n3256 ^ n3245;
  assign n3345 = n3256 ^ n3250;
  assign n3346 = ~n3344 & ~n3345;
  assign n3347 = n3346 ^ n3245;
  assign n3352 = n3351 ^ n3347;
  assign n3357 = n3356 ^ n3352;
  assign n3362 = n3361 ^ n3357;
  assign n3338 = n3224 ^ n3213;
  assign n3339 = n3224 ^ n3218;
  assign n3340 = n3338 & ~n3339;
  assign n3341 = n3340 ^ n3213;
  assign n3335 = n3207 ^ n3201;
  assign n3336 = n3202 & ~n3335;
  assign n3337 = n3336 ^ n3196;
  assign n3342 = n3341 ^ n3337;
  assign n3331 = ~x18 & n894;
  assign n3332 = n3331 ^ n1052;
  assign n3329 = ~x17 & n1049;
  assign n3330 = n3329 ^ n1087;
  assign n3333 = n3332 ^ n3330;
  assign n3325 = x30 & n157;
  assign n3326 = n3325 ^ n191;
  assign n3323 = x29 & n188;
  assign n3324 = n3323 ^ n248;
  assign n3327 = n3326 ^ n3324;
  assign n3320 = ~x26 & n322;
  assign n3321 = n3320 ^ n382;
  assign n3318 = ~x25 & n379;
  assign n3319 = n3318 ^ n459;
  assign n3322 = n3321 ^ n3319;
  assign n3328 = n3327 ^ n3322;
  assign n3334 = n3333 ^ n3328;
  assign n3343 = n3342 ^ n3334;
  assign n3363 = n3362 ^ n3343;
  assign n3388 = n3387 ^ n3363;
  assign n3459 = n3458 ^ n3388;
  assign n3463 = n3462 ^ n3459;
  assign n3467 = n3466 ^ n3463;
  assign n3471 = n3470 ^ n3467;
  assign n3616 = n3470 ^ n3463;
  assign n3617 = ~n3467 & n3616;
  assign n3618 = n3617 ^ n3470;
  assign n3612 = n3462 ^ n3458;
  assign n3613 = n3459 & ~n3612;
  assign n3614 = n3613 ^ n3388;
  assign n3608 = n3457 ^ n3453;
  assign n3609 = n3454 & ~n3608;
  assign n3610 = n3609 ^ n3450;
  assign n3602 = n3383 ^ n3363;
  assign n3603 = n3386 ^ n3363;
  assign n3604 = n3602 & n3603;
  assign n3605 = n3604 ^ n3383;
  assign n3598 = n3449 ^ n3444;
  assign n3599 = n3445 & ~n3598;
  assign n3600 = n3599 ^ n3441;
  assign n3592 = n3356 ^ n3347;
  assign n3593 = n3356 ^ n3351;
  assign n3594 = ~n3592 & ~n3593;
  assign n3595 = n3594 ^ n3347;
  assign n3587 = n3373 ^ n3364;
  assign n3588 = n3373 ^ n3369;
  assign n3589 = ~n3587 & n3588;
  assign n3590 = n3589 ^ n3364;
  assign n3583 = x29 & n241;
  assign n3584 = n3583 ^ n293;
  assign n3581 = x28 & n290;
  assign n3582 = n3581 ^ n342;
  assign n3585 = n3584 ^ n3582;
  assign n3577 = x13 & n1556;
  assign n3578 = n3577 ^ n1664;
  assign n3575 = x12 & n1661;
  assign n3576 = n3575 ^ n1878;
  assign n3579 = n3578 ^ n3576;
  assign n3572 = x15 & n1360;
  assign n3573 = n3572 ^ n1447;
  assign n3570 = x14 & n1444;
  assign n3571 = n3570 ^ n1588;
  assign n3574 = n3573 ^ n3571;
  assign n3580 = n3579 ^ n3574;
  assign n3586 = n3585 ^ n3580;
  assign n3591 = n3590 ^ n3586;
  assign n3596 = n3595 ^ n3591;
  assign n3565 = n3422 ^ n3405;
  assign n3566 = n3439 ^ n3405;
  assign n3567 = n3565 & ~n3566;
  assign n3568 = n3567 ^ n3422;
  assign n3558 = x7 & n2387;
  assign n3559 = n3558 ^ n2635;
  assign n3556 = x6 & n2631;
  assign n3557 = n3556 ^ n2632;
  assign n3560 = n3559 ^ n3557;
  assign n3553 = x21 & n756;
  assign n3554 = n3553 ^ n873;
  assign n3551 = x20 & n870;
  assign n3552 = n3551 ^ n953;
  assign n3555 = n3554 ^ n3552;
  assign n3561 = n3560 ^ n3555;
  assign n3550 = x5 & x63;
  assign n3562 = n3561 ^ n3550;
  assign n3546 = ~x27 & n322;
  assign n3547 = n3546 ^ n382;
  assign n3544 = ~x26 & n379;
  assign n3545 = n3544 ^ n459;
  assign n3548 = n3547 ^ n3545;
  assign n3540 = x31 & n157;
  assign n3541 = n3540 ^ n191;
  assign n3538 = x30 & n188;
  assign n3539 = n3538 ^ n248;
  assign n3542 = n3541 ^ n3539;
  assign n3537 = n171 ^ n142;
  assign n3543 = n3542 ^ n3537;
  assign n3549 = n3548 ^ n3543;
  assign n3563 = n3562 ^ n3549;
  assign n3533 = x9 & n2143;
  assign n3534 = n3533 ^ n2275;
  assign n3531 = x8 & n2272;
  assign n3532 = n3531 ^ n2484;
  assign n3535 = n3534 ^ n3532;
  assign n3527 = ~x11 & n1815;
  assign n3528 = n3527 ^ n2047;
  assign n3525 = ~x10 & n2044;
  assign n3526 = n3525 ^ n2162;
  assign n3529 = n3528 ^ n3526;
  assign n3522 = ~x23 & n567;
  assign n3523 = n3522 ^ n672;
  assign n3520 = ~x22 & n669;
  assign n3521 = n3520 ^ n738;
  assign n3524 = n3523 ^ n3521;
  assign n3530 = n3529 ^ n3524;
  assign n3536 = n3535 ^ n3530;
  assign n3564 = n3563 ^ n3536;
  assign n3569 = n3568 ^ n3564;
  assign n3597 = n3596 ^ n3569;
  assign n3601 = n3600 ^ n3597;
  assign n3606 = n3605 ^ n3601;
  assign n3515 = n3357 ^ n3343;
  assign n3516 = n3362 & ~n3515;
  assign n3517 = n3516 ^ n3343;
  assign n3511 = n3382 ^ n3374;
  assign n3512 = n3382 ^ n3378;
  assign n3513 = ~n3511 & ~n3512;
  assign n3514 = n3513 ^ n3374;
  assign n3518 = n3517 ^ n3514;
  assign n3507 = n3337 ^ n3334;
  assign n3508 = ~n3342 & n3507;
  assign n3509 = n3508 ^ n3334;
  assign n3502 = n3438 ^ n3432;
  assign n3503 = n3433 & ~n3502;
  assign n3504 = n3503 ^ n3427;
  assign n3498 = n3333 ^ n3327;
  assign n3499 = n3328 & ~n3498;
  assign n3500 = n3499 ^ n3322;
  assign n3501 = n3500 ^ n3373;
  assign n3505 = n3504 ^ n3501;
  assign n3492 = n3404 ^ n3393;
  assign n3493 = n3404 ^ n3398;
  assign n3494 = n3492 & ~n3493;
  assign n3495 = n3494 ^ n3393;
  assign n3489 = n3421 ^ n3410;
  assign n3490 = ~n3416 & n3489;
  assign n3491 = n3490 ^ n3421;
  assign n3496 = n3495 ^ n3491;
  assign n3485 = x25 & n435;
  assign n3486 = n3485 ^ n527;
  assign n3483 = x24 & n524;
  assign n3484 = n3483 ^ n611;
  assign n3487 = n3486 ^ n3484;
  assign n3479 = x17 & n1105;
  assign n3480 = n3479 ^ n1206;
  assign n3477 = x16 & n1203;
  assign n3478 = n3477 ^ n1379;
  assign n3481 = n3480 ^ n3478;
  assign n3474 = ~x19 & n894;
  assign n3475 = n3474 ^ n1052;
  assign n3472 = ~x18 & n1049;
  assign n3473 = n3472 ^ n1087;
  assign n3476 = n3475 ^ n3473;
  assign n3482 = n3481 ^ n3476;
  assign n3488 = n3487 ^ n3482;
  assign n3497 = n3496 ^ n3488;
  assign n3506 = n3505 ^ n3497;
  assign n3510 = n3509 ^ n3506;
  assign n3519 = n3518 ^ n3510;
  assign n3607 = n3606 ^ n3519;
  assign n3611 = n3610 ^ n3607;
  assign n3615 = n3614 ^ n3611;
  assign n3619 = n3618 ^ n3615;
  assign n3755 = n3618 ^ n3611;
  assign n3756 = ~n3615 & n3755;
  assign n3757 = n3756 ^ n3618;
  assign n3751 = n3610 ^ n3606;
  assign n3752 = n3607 & n3751;
  assign n3753 = n3752 ^ n3519;
  assign n3747 = n3605 ^ n3600;
  assign n3748 = n3601 & n3747;
  assign n3749 = n3748 ^ n3597;
  assign n3743 = n3514 ^ n3510;
  assign n3744 = n3518 & ~n3743;
  assign n3745 = n3744 ^ n3510;
  assign n3738 = n3596 ^ n3568;
  assign n3739 = ~n3569 & n3738;
  assign n3740 = n3739 ^ n3564;
  assign n3734 = n3595 ^ n3590;
  assign n3735 = n3591 & n3734;
  assign n3736 = n3735 ^ n3586;
  assign n3729 = n3549 ^ n3536;
  assign n3730 = n3562 ^ n3536;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = n3731 ^ n3549;
  assign n3724 = n3555 ^ n3550;
  assign n3725 = ~n3561 & n3724;
  assign n3726 = n3725 ^ n3550;
  assign n3719 = x8 & n2387;
  assign n3720 = n3719 ^ n2635;
  assign n3717 = x7 & n2631;
  assign n3718 = n3717 ^ n2632;
  assign n3721 = n3720 ^ n3718;
  assign n3714 = ~x28 & n322;
  assign n3715 = n3714 ^ n382;
  assign n3712 = ~x27 & n379;
  assign n3713 = n3712 ^ n459;
  assign n3716 = n3715 ^ n3713;
  assign n3722 = n3721 ^ n3716;
  assign n3711 = x6 & x63;
  assign n3723 = n3722 ^ n3711;
  assign n3727 = n3726 ^ n3723;
  assign n3707 = x16 & n1360;
  assign n3708 = n3707 ^ n1447;
  assign n3705 = x15 & n1444;
  assign n3706 = n3705 ^ n1588;
  assign n3709 = n3708 ^ n3706;
  assign n3701 = x18 & n1105;
  assign n3702 = n3701 ^ n1206;
  assign n3699 = x17 & n1203;
  assign n3700 = n3699 ^ n1379;
  assign n3703 = n3702 ^ n3700;
  assign n3696 = x26 & n435;
  assign n3697 = n3696 ^ n527;
  assign n3694 = x25 & n524;
  assign n3695 = n3694 ^ n611;
  assign n3698 = n3697 ^ n3695;
  assign n3704 = n3703 ^ n3698;
  assign n3710 = n3709 ^ n3704;
  assign n3728 = n3727 ^ n3710;
  assign n3733 = n3732 ^ n3728;
  assign n3737 = n3736 ^ n3733;
  assign n3741 = n3740 ^ n3737;
  assign n3689 = n3509 ^ n3505;
  assign n3690 = n3506 & ~n3689;
  assign n3691 = n3690 ^ n3497;
  assign n3684 = n3535 ^ n3524;
  assign n3685 = ~n3530 & n3684;
  assign n3686 = n3685 ^ n3535;
  assign n3680 = ~x20 & n894;
  assign n3681 = n3680 ^ n1052;
  assign n3678 = ~x19 & n1049;
  assign n3679 = n3678 ^ n1087;
  assign n3682 = n3681 ^ n3679;
  assign n3675 = x30 & n241;
  assign n3676 = n3675 ^ n293;
  assign n3673 = x29 & n290;
  assign n3674 = n3673 ^ n342;
  assign n3677 = n3676 ^ n3674;
  assign n3683 = n3682 ^ n3677;
  assign n3687 = n3686 ^ n3683;
  assign n3668 = ~x12 & n1815;
  assign n3669 = n3668 ^ n2047;
  assign n3666 = ~x11 & n2044;
  assign n3667 = n3666 ^ n2162;
  assign n3670 = n3669 ^ n3667;
  assign n3662 = x14 & n1556;
  assign n3663 = n3662 ^ n1664;
  assign n3660 = x13 & n1661;
  assign n3661 = n3660 ^ n1878;
  assign n3664 = n3663 ^ n3661;
  assign n3657 = ~x24 & n567;
  assign n3658 = n3657 ^ n672;
  assign n3655 = ~x23 & n669;
  assign n3656 = n3655 ^ n738;
  assign n3659 = n3658 ^ n3656;
  assign n3665 = n3664 ^ n3659;
  assign n3671 = n3670 ^ n3665;
  assign n3651 = x10 & n2143;
  assign n3652 = n3651 ^ n2275;
  assign n3649 = x9 & n2272;
  assign n3650 = n3649 ^ n2484;
  assign n3653 = n3652 ^ n3650;
  assign n3645 = x22 & n756;
  assign n3646 = n3645 ^ n873;
  assign n3643 = x21 & n870;
  assign n3644 = n3643 ^ n953;
  assign n3647 = n3646 ^ n3644;
  assign n3640 = x31 & n188;
  assign n3641 = n3640 ^ n191;
  assign n3642 = n3641 ^ n248;
  assign n3648 = n3647 ^ n3642;
  assign n3654 = n3653 ^ n3648;
  assign n3672 = n3671 ^ n3654;
  assign n3688 = n3687 ^ n3672;
  assign n3692 = n3691 ^ n3688;
  assign n3636 = n3491 ^ n3488;
  assign n3637 = ~n3496 & n3636;
  assign n3638 = n3637 ^ n3488;
  assign n3632 = n3504 ^ n3500;
  assign n3633 = n3501 & ~n3632;
  assign n3634 = n3633 ^ n3373;
  assign n3628 = n3585 ^ n3579;
  assign n3629 = n3580 & ~n3628;
  assign n3630 = n3629 ^ n3574;
  assign n3624 = n3487 ^ n3476;
  assign n3625 = ~n3482 & n3624;
  assign n3626 = n3625 ^ n3487;
  assign n3620 = n3548 ^ n3537;
  assign n3621 = n3548 ^ n3542;
  assign n3622 = ~n3620 & ~n3621;
  assign n3623 = n3622 ^ n3537;
  assign n3627 = n3626 ^ n3623;
  assign n3631 = n3630 ^ n3627;
  assign n3635 = n3634 ^ n3631;
  assign n3639 = n3638 ^ n3635;
  assign n3693 = n3692 ^ n3639;
  assign n3742 = n3741 ^ n3693;
  assign n3746 = n3745 ^ n3742;
  assign n3750 = n3749 ^ n3746;
  assign n3754 = n3753 ^ n3750;
  assign n3758 = n3757 ^ n3754;
  assign n3890 = n3757 ^ n3750;
  assign n3891 = n3754 & n3890;
  assign n3892 = n3891 ^ n3757;
  assign n3886 = n3749 ^ n3745;
  assign n3887 = n3746 & ~n3886;
  assign n3888 = n3887 ^ n3742;
  assign n3881 = n3737 ^ n3693;
  assign n3882 = n3740 ^ n3693;
  assign n3883 = ~n3881 & n3882;
  assign n3884 = n3883 ^ n3737;
  assign n3876 = n3688 ^ n3639;
  assign n3877 = n3691 ^ n3639;
  assign n3878 = n3876 & n3877;
  assign n3879 = n3878 ^ n3688;
  assign n3871 = n3736 ^ n3732;
  assign n3872 = ~n3733 & n3871;
  assign n3873 = n3872 ^ n3728;
  assign n3866 = n3723 ^ n3710;
  assign n3867 = ~n3727 & n3866;
  assign n3868 = n3867 ^ n3710;
  assign n3861 = n3716 ^ n3711;
  assign n3862 = ~n3722 & n3861;
  assign n3863 = n3862 ^ n3711;
  assign n3857 = ~x25 & n567;
  assign n3858 = n3857 ^ n672;
  assign n3855 = ~x24 & n669;
  assign n3856 = n3855 ^ n738;
  assign n3859 = n3858 ^ n3856;
  assign n3851 = x17 & n1360;
  assign n3852 = n3851 ^ n1447;
  assign n3849 = x16 & n1444;
  assign n3850 = n3849 ^ n1588;
  assign n3853 = n3852 ^ n3850;
  assign n3846 = x19 & n1105;
  assign n3847 = n3846 ^ n1206;
  assign n3844 = x18 & n1203;
  assign n3845 = n3844 ^ n1379;
  assign n3848 = n3847 ^ n3845;
  assign n3854 = n3853 ^ n3848;
  assign n3860 = n3859 ^ n3854;
  assign n3864 = n3863 ^ n3860;
  assign n3840 = x27 & n435;
  assign n3841 = n3840 ^ n527;
  assign n3838 = x26 & n524;
  assign n3839 = n3838 ^ n611;
  assign n3842 = n3841 ^ n3839;
  assign n3834 = x31 & n241;
  assign n3835 = n3834 ^ n293;
  assign n3832 = x30 & n290;
  assign n3833 = n3832 ^ n342;
  assign n3836 = n3835 ^ n3833;
  assign n3831 = n248 ^ n191;
  assign n3837 = n3836 ^ n3831;
  assign n3843 = n3842 ^ n3837;
  assign n3865 = n3864 ^ n3843;
  assign n3869 = n3868 ^ n3865;
  assign n3825 = ~x29 & n322;
  assign n3826 = n3825 ^ n382;
  assign n3823 = ~x28 & n379;
  assign n3824 = n3823 ^ n459;
  assign n3827 = n3826 ^ n3824;
  assign n3819 = ~x13 & n1815;
  assign n3820 = n3819 ^ n2047;
  assign n3817 = ~x12 & n2044;
  assign n3818 = n3817 ^ n2162;
  assign n3821 = n3820 ^ n3818;
  assign n3814 = x15 & n1556;
  assign n3815 = n3814 ^ n1664;
  assign n3812 = x14 & n1661;
  assign n3813 = n3812 ^ n1878;
  assign n3816 = n3815 ^ n3813;
  assign n3822 = n3821 ^ n3816;
  assign n3828 = n3827 ^ n3822;
  assign n3808 = x9 & n2387;
  assign n3809 = n3808 ^ n2635;
  assign n3806 = x8 & n2631;
  assign n3807 = n3806 ^ n2632;
  assign n3810 = n3809 ^ n3807;
  assign n3802 = x11 & n2143;
  assign n3803 = n3802 ^ n2275;
  assign n3800 = x10 & n2272;
  assign n3801 = n3800 ^ n2484;
  assign n3804 = n3803 ^ n3801;
  assign n3797 = x23 & n756;
  assign n3798 = n3797 ^ n873;
  assign n3795 = x22 & n870;
  assign n3796 = n3795 ^ n953;
  assign n3799 = n3798 ^ n3796;
  assign n3805 = n3804 ^ n3799;
  assign n3811 = n3810 ^ n3805;
  assign n3829 = n3828 ^ n3811;
  assign n3790 = ~x21 & n894;
  assign n3791 = n3790 ^ n1052;
  assign n3788 = ~x20 & n1049;
  assign n3789 = n3788 ^ n1087;
  assign n3792 = n3791 ^ n3789;
  assign n3787 = x7 & x63;
  assign n3793 = n3792 ^ n3787;
  assign n3794 = n3793 ^ n3677;
  assign n3830 = n3829 ^ n3794;
  assign n3870 = n3869 ^ n3830;
  assign n3874 = n3873 ^ n3870;
  assign n3782 = n3638 ^ n3631;
  assign n3783 = n3638 ^ n3634;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = n3784 ^ n3631;
  assign n3778 = n3687 ^ n3671;
  assign n3779 = n3672 & n3778;
  assign n3780 = n3779 ^ n3654;
  assign n3773 = n3630 ^ n3626;
  assign n3774 = ~n3627 & ~n3773;
  assign n3775 = n3774 ^ n3623;
  assign n3770 = n3686 ^ n3682;
  assign n3771 = ~n3683 & ~n3770;
  assign n3772 = n3771 ^ n3677;
  assign n3776 = n3775 ^ n3772;
  assign n3766 = n3653 ^ n3647;
  assign n3767 = n3648 & ~n3766;
  assign n3768 = n3767 ^ n3642;
  assign n3762 = n3709 ^ n3698;
  assign n3763 = ~n3704 & n3762;
  assign n3764 = n3763 ^ n3709;
  assign n3759 = n3670 ^ n3659;
  assign n3760 = ~n3665 & n3759;
  assign n3761 = n3760 ^ n3670;
  assign n3765 = n3764 ^ n3761;
  assign n3769 = n3768 ^ n3765;
  assign n3777 = n3776 ^ n3769;
  assign n3781 = n3780 ^ n3777;
  assign n3786 = n3785 ^ n3781;
  assign n3875 = n3874 ^ n3786;
  assign n3880 = n3879 ^ n3875;
  assign n3885 = n3884 ^ n3880;
  assign n3889 = n3888 ^ n3885;
  assign n3893 = n3892 ^ n3889;
  assign n4020 = n3892 ^ n3885;
  assign n4021 = ~n3889 & n4020;
  assign n4022 = n4021 ^ n3892;
  assign n4015 = n3884 ^ n3879;
  assign n4016 = n3884 ^ n3875;
  assign n4017 = n4015 & n4016;
  assign n4018 = n4017 ^ n3879;
  assign n4010 = n3870 ^ n3786;
  assign n4011 = n3873 ^ n3786;
  assign n4012 = n4010 & n4011;
  assign n4013 = n4012 ^ n3870;
  assign n4005 = n3785 ^ n3777;
  assign n4006 = n3781 & n4005;
  assign n4007 = n4006 ^ n3780;
  assign n4001 = n3865 ^ n3830;
  assign n4002 = n3869 & ~n4001;
  assign n4003 = n4002 ^ n3830;
  assign n3997 = n3811 ^ n3794;
  assign n3998 = ~n3829 & n3997;
  assign n3999 = n3998 ^ n3794;
  assign n3993 = n3860 ^ n3843;
  assign n3994 = ~n3864 & ~n3993;
  assign n3995 = n3994 ^ n3843;
  assign n3988 = n3810 ^ n3804;
  assign n3989 = n3805 & ~n3988;
  assign n3990 = n3989 ^ n3799;
  assign n3984 = n3842 ^ n3831;
  assign n3985 = n3842 ^ n3836;
  assign n3986 = ~n3984 & ~n3985;
  assign n3987 = n3986 ^ n3831;
  assign n3991 = n3990 ^ n3987;
  assign n3980 = x20 & n1105;
  assign n3981 = n3980 ^ n1206;
  assign n3978 = x19 & n1203;
  assign n3979 = n3978 ^ n1379;
  assign n3982 = n3981 ^ n3979;
  assign n3974 = x28 & n435;
  assign n3975 = n3974 ^ n527;
  assign n3972 = x27 & n524;
  assign n3973 = n3972 ^ n611;
  assign n3976 = n3975 ^ n3973;
  assign n3971 = x8 & x63;
  assign n3977 = n3976 ^ n3971;
  assign n3983 = n3982 ^ n3977;
  assign n3992 = n3991 ^ n3983;
  assign n3996 = n3995 ^ n3992;
  assign n4000 = n3999 ^ n3996;
  assign n4004 = n4003 ^ n4000;
  assign n4008 = n4007 ^ n4004;
  assign n3966 = n3772 ^ n3769;
  assign n3967 = ~n3776 & ~n3966;
  assign n3968 = n3967 ^ n3769;
  assign n3960 = x10 & n2387;
  assign n3961 = n3960 ^ n2635;
  assign n3958 = x9 & n2631;
  assign n3959 = n3958 ^ n2632;
  assign n3962 = n3961 ^ n3959;
  assign n3954 = ~x22 & n894;
  assign n3955 = n3954 ^ n1052;
  assign n3952 = ~x21 & n1049;
  assign n3953 = n3952 ^ n1087;
  assign n3956 = n3955 ^ n3953;
  assign n3949 = x31 & n290;
  assign n3950 = n3949 ^ n293;
  assign n3951 = n3950 ^ n342;
  assign n3957 = n3956 ^ n3951;
  assign n3963 = n3962 ^ n3957;
  assign n3945 = x16 & n1556;
  assign n3946 = n3945 ^ n1664;
  assign n3943 = x15 & n1661;
  assign n3944 = n3943 ^ n1878;
  assign n3947 = n3946 ^ n3944;
  assign n3939 = ~x26 & n567;
  assign n3940 = n3939 ^ n672;
  assign n3937 = ~x25 & n669;
  assign n3938 = n3937 ^ n738;
  assign n3941 = n3940 ^ n3938;
  assign n3934 = x18 & n1360;
  assign n3935 = n3934 ^ n1447;
  assign n3932 = x17 & n1444;
  assign n3933 = n3932 ^ n1588;
  assign n3936 = n3935 ^ n3933;
  assign n3942 = n3941 ^ n3936;
  assign n3948 = n3947 ^ n3942;
  assign n3964 = n3963 ^ n3948;
  assign n3928 = x12 & n2143;
  assign n3929 = n3928 ^ n2275;
  assign n3926 = x11 & n2272;
  assign n3927 = n3926 ^ n2484;
  assign n3930 = n3929 ^ n3927;
  assign n3922 = ~x14 & n1815;
  assign n3923 = n3922 ^ n2047;
  assign n3920 = ~x13 & n2044;
  assign n3921 = n3920 ^ n2162;
  assign n3924 = n3923 ^ n3921;
  assign n3917 = x24 & n756;
  assign n3918 = n3917 ^ n873;
  assign n3915 = x23 & n870;
  assign n3916 = n3915 ^ n953;
  assign n3919 = n3918 ^ n3916;
  assign n3925 = n3924 ^ n3919;
  assign n3931 = n3930 ^ n3925;
  assign n3965 = n3964 ^ n3931;
  assign n3969 = n3968 ^ n3965;
  assign n3910 = n3768 ^ n3764;
  assign n3911 = n3765 & ~n3910;
  assign n3912 = n3911 ^ n3761;
  assign n3907 = n3792 ^ n3677;
  assign n3908 = n3793 & ~n3907;
  assign n3909 = n3908 ^ n3787;
  assign n3913 = n3912 ^ n3909;
  assign n3903 = n3827 ^ n3816;
  assign n3904 = ~n3822 & n3903;
  assign n3905 = n3904 ^ n3827;
  assign n3899 = ~x30 & n322;
  assign n3900 = n3899 ^ n382;
  assign n3897 = ~x29 & n379;
  assign n3898 = n3897 ^ n459;
  assign n3901 = n3900 ^ n3898;
  assign n3894 = n3859 ^ n3848;
  assign n3895 = ~n3854 & n3894;
  assign n3896 = n3895 ^ n3859;
  assign n3902 = n3901 ^ n3896;
  assign n3906 = n3905 ^ n3902;
  assign n3914 = n3913 ^ n3906;
  assign n3970 = n3969 ^ n3914;
  assign n4009 = n4008 ^ n3970;
  assign n4014 = n4013 ^ n4009;
  assign n4019 = n4018 ^ n4014;
  assign n4023 = n4022 ^ n4019;
  assign n4148 = n4022 ^ n4014;
  assign n4149 = n4019 & n4148;
  assign n4150 = n4149 ^ n4022;
  assign n4144 = n4013 ^ n4008;
  assign n4145 = ~n4009 & n4144;
  assign n4146 = n4145 ^ n3970;
  assign n4140 = n4007 ^ n4003;
  assign n4141 = n4004 & ~n4140;
  assign n4142 = n4141 ^ n4000;
  assign n4134 = n3965 ^ n3914;
  assign n4135 = n3968 ^ n3914;
  assign n4136 = ~n4134 & n4135;
  assign n4137 = n4136 ^ n3965;
  assign n4129 = n3999 ^ n3992;
  assign n4130 = n3999 ^ n3995;
  assign n4131 = ~n4129 & n4130;
  assign n4132 = n4131 ^ n3992;
  assign n4124 = n3948 ^ n3931;
  assign n4125 = n3963 ^ n3931;
  assign n4126 = n4124 & ~n4125;
  assign n4127 = n4126 ^ n3948;
  assign n4120 = n3987 ^ n3983;
  assign n4121 = n3991 & ~n4120;
  assign n4122 = n4121 ^ n3983;
  assign n4115 = n3947 ^ n3936;
  assign n4116 = n3947 ^ n3941;
  assign n4117 = n4115 & ~n4116;
  assign n4118 = n4117 ^ n3936;
  assign n4110 = n3962 ^ n3951;
  assign n4111 = n3962 ^ n3956;
  assign n4112 = n4110 & ~n4111;
  assign n4113 = n4112 ^ n3951;
  assign n4107 = n3982 ^ n3976;
  assign n4108 = n3977 & ~n4107;
  assign n4109 = n4108 ^ n3971;
  assign n4114 = n4113 ^ n4109;
  assign n4119 = n4118 ^ n4114;
  assign n4123 = n4122 ^ n4119;
  assign n4128 = n4127 ^ n4123;
  assign n4133 = n4132 ^ n4128;
  assign n4138 = n4137 ^ n4133;
  assign n4101 = n3909 ^ n3906;
  assign n4102 = n3912 ^ n3906;
  assign n4103 = ~n4101 & n4102;
  assign n4104 = n4103 ^ n3909;
  assign n4095 = x29 & n435;
  assign n4096 = n4095 ^ n527;
  assign n4093 = x28 & n524;
  assign n4094 = n4093 ^ n611;
  assign n4097 = n4096 ^ n4094;
  assign n4089 = x13 & n2143;
  assign n4090 = n4089 ^ n2275;
  assign n4087 = x12 & n2272;
  assign n4088 = n4087 ^ n2484;
  assign n4091 = n4090 ^ n4088;
  assign n4084 = ~x15 & n1815;
  assign n4085 = n4084 ^ n2047;
  assign n4082 = ~x14 & n2044;
  assign n4083 = n4082 ^ n2162;
  assign n4086 = n4085 ^ n4083;
  assign n4092 = n4091 ^ n4086;
  assign n4098 = n4097 ^ n4092;
  assign n4078 = ~x27 & n567;
  assign n4079 = n4078 ^ n672;
  assign n4076 = ~x26 & n669;
  assign n4077 = n4076 ^ n738;
  assign n4080 = n4079 ^ n4077;
  assign n4072 = ~x31 & n322;
  assign n4073 = n4072 ^ n382;
  assign n4070 = ~x30 & n379;
  assign n4071 = n4070 ^ n459;
  assign n4074 = n4073 ^ n4071;
  assign n4069 = n342 ^ n293;
  assign n4075 = n4074 ^ n4069;
  assign n4081 = n4080 ^ n4075;
  assign n4099 = n4098 ^ n4081;
  assign n4065 = x25 & n756;
  assign n4066 = n4065 ^ n873;
  assign n4063 = x24 & n870;
  assign n4064 = n4063 ^ n953;
  assign n4067 = n4066 ^ n4064;
  assign n4059 = x17 & n1556;
  assign n4060 = n4059 ^ n1664;
  assign n4057 = x16 & n1661;
  assign n4058 = n4057 ^ n1878;
  assign n4061 = n4060 ^ n4058;
  assign n4054 = x19 & n1360;
  assign n4055 = n4054 ^ n1447;
  assign n4052 = x18 & n1444;
  assign n4053 = n4052 ^ n1588;
  assign n4056 = n4055 ^ n4053;
  assign n4062 = n4061 ^ n4056;
  assign n4068 = n4067 ^ n4062;
  assign n4100 = n4099 ^ n4068;
  assign n4105 = n4104 ^ n4100;
  assign n4048 = n3905 ^ n3896;
  assign n4049 = ~n3902 & ~n4048;
  assign n4050 = n4049 ^ n3901;
  assign n4043 = n3930 ^ n3919;
  assign n4044 = ~n3925 & n4043;
  assign n4045 = n4044 ^ n3930;
  assign n4039 = x21 & n1105;
  assign n4040 = n4039 ^ n1206;
  assign n4037 = x20 & n1203;
  assign n4038 = n4037 ^ n1379;
  assign n4041 = n4040 ^ n4038;
  assign n4042 = n4041 ^ n3901;
  assign n4046 = n4045 ^ n4042;
  assign n4032 = x11 & n2387;
  assign n4033 = n4032 ^ n2635;
  assign n4030 = x10 & n2631;
  assign n4031 = n4030 ^ n2632;
  assign n4034 = n4033 ^ n4031;
  assign n4027 = ~x23 & n894;
  assign n4028 = n4027 ^ n1052;
  assign n4025 = ~x22 & n1049;
  assign n4026 = n4025 ^ n1087;
  assign n4029 = n4028 ^ n4026;
  assign n4035 = n4034 ^ n4029;
  assign n4024 = x9 & x63;
  assign n4036 = n4035 ^ n4024;
  assign n4047 = n4046 ^ n4036;
  assign n4051 = n4050 ^ n4047;
  assign n4106 = n4105 ^ n4051;
  assign n4139 = n4138 ^ n4106;
  assign n4143 = n4142 ^ n4139;
  assign n4147 = n4146 ^ n4143;
  assign n4151 = n4150 ^ n4147;
  assign n4269 = n4150 ^ n4143;
  assign n4270 = ~n4147 & ~n4269;
  assign n4271 = n4270 ^ n4150;
  assign n4265 = n4142 ^ n4138;
  assign n4266 = ~n4139 & n4265;
  assign n4267 = n4266 ^ n4106;
  assign n4261 = n4137 ^ n4132;
  assign n4262 = ~n4133 & n4261;
  assign n4263 = n4262 ^ n4128;
  assign n4255 = n4100 ^ n4051;
  assign n4256 = n4104 ^ n4051;
  assign n4257 = n4255 & n4256;
  assign n4258 = n4257 ^ n4100;
  assign n4251 = n4127 ^ n4119;
  assign n4252 = ~n4123 & n4251;
  assign n4253 = n4252 ^ n4127;
  assign n4247 = n4098 ^ n4068;
  assign n4248 = ~n4099 & ~n4247;
  assign n4249 = n4248 ^ n4081;
  assign n4243 = n4045 ^ n4041;
  assign n4244 = n4042 & ~n4243;
  assign n4245 = n4244 ^ n3901;
  assign n4239 = n4080 ^ n4074;
  assign n4240 = ~n4075 & ~n4239;
  assign n4241 = n4240 ^ n4069;
  assign n4235 = n4029 ^ n4024;
  assign n4236 = ~n4035 & n4235;
  assign n4237 = n4236 ^ n4024;
  assign n4232 = n4097 ^ n4086;
  assign n4233 = ~n4092 & n4232;
  assign n4234 = n4233 ^ n4097;
  assign n4238 = n4237 ^ n4234;
  assign n4242 = n4241 ^ n4238;
  assign n4246 = n4245 ^ n4242;
  assign n4250 = n4249 ^ n4246;
  assign n4254 = n4253 ^ n4250;
  assign n4259 = n4258 ^ n4254;
  assign n4227 = n4050 ^ n4046;
  assign n4228 = n4047 & n4227;
  assign n4229 = n4228 ^ n4036;
  assign n4222 = n4067 ^ n4061;
  assign n4223 = n4062 & ~n4222;
  assign n4224 = n4223 ^ n4056;
  assign n4217 = ~x28 & n567;
  assign n4218 = n4217 ^ n672;
  assign n4215 = ~x27 & n669;
  assign n4216 = n4215 ^ n738;
  assign n4219 = n4218 ^ n4216;
  assign n4212 = x31 & n379;
  assign n4211 = n382 ^ n322;
  assign n4213 = n4212 ^ n4211;
  assign n4210 = n459 ^ n379;
  assign n4214 = n4213 ^ n4210;
  assign n4220 = n4219 ^ n4214;
  assign n4209 = x10 & x63;
  assign n4221 = n4220 ^ n4209;
  assign n4225 = n4224 ^ n4221;
  assign n4205 = ~x16 & n1815;
  assign n4206 = n4205 ^ n2047;
  assign n4203 = ~x15 & n2044;
  assign n4204 = n4203 ^ n2162;
  assign n4207 = n4206 ^ n4204;
  assign n4199 = x26 & n756;
  assign n4200 = n4199 ^ n873;
  assign n4197 = x25 & n870;
  assign n4198 = n4197 ^ n953;
  assign n4201 = n4200 ^ n4198;
  assign n4194 = x18 & n1556;
  assign n4195 = n4194 ^ n1664;
  assign n4192 = x17 & n1661;
  assign n4193 = n4192 ^ n1878;
  assign n4196 = n4195 ^ n4193;
  assign n4202 = n4201 ^ n4196;
  assign n4208 = n4207 ^ n4202;
  assign n4226 = n4225 ^ n4208;
  assign n4230 = n4229 ^ n4226;
  assign n4187 = n4118 ^ n4109;
  assign n4188 = n4118 ^ n4113;
  assign n4189 = n4187 & ~n4188;
  assign n4190 = n4189 ^ n4109;
  assign n4182 = x12 & n2387;
  assign n4183 = n4182 ^ n2635;
  assign n4180 = x11 & n2631;
  assign n4181 = n4180 ^ n2632;
  assign n4184 = n4183 ^ n4181;
  assign n4176 = ~x24 & n894;
  assign n4177 = n4176 ^ n1052;
  assign n4174 = ~x23 & n1049;
  assign n4175 = n4174 ^ n1087;
  assign n4178 = n4177 ^ n4175;
  assign n4171 = x14 & n2143;
  assign n4172 = n4171 ^ n2275;
  assign n4169 = x13 & n2272;
  assign n4170 = n4169 ^ n2484;
  assign n4173 = n4172 ^ n4170;
  assign n4179 = n4178 ^ n4173;
  assign n4185 = n4184 ^ n4179;
  assign n4165 = x30 & n435;
  assign n4166 = n4165 ^ n527;
  assign n4163 = x29 & n524;
  assign n4164 = n4163 ^ n611;
  assign n4167 = n4166 ^ n4164;
  assign n4159 = x22 & n1105;
  assign n4160 = n4159 ^ n1206;
  assign n4157 = x21 & n1203;
  assign n4158 = n4157 ^ n1379;
  assign n4161 = n4160 ^ n4158;
  assign n4154 = x20 & n1360;
  assign n4155 = n4154 ^ n1447;
  assign n4152 = x19 & n1444;
  assign n4153 = n4152 ^ n1588;
  assign n4156 = n4155 ^ n4153;
  assign n4162 = n4161 ^ n4156;
  assign n4168 = n4167 ^ n4162;
  assign n4186 = n4185 ^ n4168;
  assign n4191 = n4190 ^ n4186;
  assign n4231 = n4230 ^ n4191;
  assign n4260 = n4259 ^ n4231;
  assign n4264 = n4263 ^ n4260;
  assign n4268 = n4267 ^ n4264;
  assign n4272 = n4271 ^ n4268;
  assign n4387 = n4271 ^ n4264;
  assign n4388 = ~n4268 & n4387;
  assign n4389 = n4388 ^ n4271;
  assign n4383 = n4263 ^ n4259;
  assign n4384 = n4260 & n4383;
  assign n4385 = n4384 ^ n4231;
  assign n4379 = n4258 ^ n4253;
  assign n4380 = n4254 & n4379;
  assign n4381 = n4380 ^ n4250;
  assign n4373 = n4226 ^ n4191;
  assign n4374 = n4229 ^ n4191;
  assign n4375 = ~n4373 & n4374;
  assign n4376 = n4375 ^ n4226;
  assign n4368 = n4249 ^ n4242;
  assign n4369 = n4249 ^ n4245;
  assign n4370 = n4368 & n4369;
  assign n4371 = n4370 ^ n4242;
  assign n4362 = n4241 ^ n4234;
  assign n4363 = n4241 ^ n4237;
  assign n4364 = ~n4362 & n4363;
  assign n4365 = n4364 ^ n4234;
  assign n4358 = n4221 ^ n4208;
  assign n4359 = n4224 ^ n4208;
  assign n4360 = n4358 & ~n4359;
  assign n4361 = n4360 ^ n4221;
  assign n4366 = n4365 ^ n4361;
  assign n4354 = n4207 ^ n4201;
  assign n4355 = n4202 & ~n4354;
  assign n4356 = n4355 ^ n4196;
  assign n4350 = n4214 ^ n4209;
  assign n4351 = ~n4220 & n4350;
  assign n4352 = n4351 ^ n4209;
  assign n4353 = n4352 ^ n4167;
  assign n4357 = n4356 ^ n4353;
  assign n4367 = n4366 ^ n4357;
  assign n4372 = n4371 ^ n4367;
  assign n4377 = n4376 ^ n4372;
  assign n4346 = n4190 ^ n4185;
  assign n4347 = ~n4186 & ~n4346;
  assign n4348 = n4347 ^ n4168;
  assign n4340 = n4167 ^ n4156;
  assign n4341 = n4167 ^ n4161;
  assign n4342 = ~n4340 & n4341;
  assign n4343 = n4342 ^ n4156;
  assign n4335 = ~x25 & n894;
  assign n4336 = n4335 ^ n1052;
  assign n4333 = ~x24 & n1049;
  assign n4334 = n4333 ^ n1087;
  assign n4337 = n4336 ^ n4334;
  assign n4329 = ~x17 & n1815;
  assign n4330 = n4329 ^ n2047;
  assign n4327 = ~x16 & n2044;
  assign n4328 = n4327 ^ n2162;
  assign n4331 = n4330 ^ n4328;
  assign n4324 = x19 & n1556;
  assign n4325 = n4324 ^ n1664;
  assign n4322 = x18 & n1661;
  assign n4323 = n4322 ^ n1878;
  assign n4326 = n4325 ^ n4323;
  assign n4332 = n4331 ^ n4326;
  assign n4338 = n4337 ^ n4332;
  assign n4318 = x27 & n756;
  assign n4319 = n4318 ^ n873;
  assign n4316 = x26 & n870;
  assign n4317 = n4316 ^ n953;
  assign n4320 = n4319 ^ n4317;
  assign n4312 = x31 & n435;
  assign n4313 = n4312 ^ n527;
  assign n4310 = x30 & n524;
  assign n4311 = n4310 ^ n611;
  assign n4314 = n4313 ^ n4311;
  assign n4309 = n4211 ^ n4210;
  assign n4315 = n4314 ^ n4309;
  assign n4321 = n4320 ^ n4315;
  assign n4339 = n4338 ^ n4321;
  assign n4344 = n4343 ^ n4339;
  assign n4303 = n4184 ^ n4173;
  assign n4304 = n4184 ^ n4178;
  assign n4305 = n4303 & ~n4304;
  assign n4306 = n4305 ^ n4173;
  assign n4299 = ~x29 & n567;
  assign n4300 = n4299 ^ n672;
  assign n4297 = ~x28 & n669;
  assign n4298 = n4297 ^ n738;
  assign n4301 = n4300 ^ n4298;
  assign n4293 = x13 & n2387;
  assign n4294 = n4293 ^ n2635;
  assign n4291 = x12 & n2631;
  assign n4292 = n4291 ^ n2632;
  assign n4295 = n4294 ^ n4292;
  assign n4288 = x15 & n2143;
  assign n4289 = n4288 ^ n2275;
  assign n4286 = x14 & n2272;
  assign n4287 = n4286 ^ n2484;
  assign n4290 = n4289 ^ n4287;
  assign n4296 = n4295 ^ n4290;
  assign n4302 = n4301 ^ n4296;
  assign n4307 = n4306 ^ n4302;
  assign n4282 = x21 & n1360;
  assign n4283 = n4282 ^ n1447;
  assign n4280 = x20 & n1444;
  assign n4281 = n4280 ^ n1588;
  assign n4284 = n4283 ^ n4281;
  assign n4276 = x23 & n1105;
  assign n4277 = n4276 ^ n1206;
  assign n4274 = x22 & n1203;
  assign n4275 = n4274 ^ n1379;
  assign n4278 = n4277 ^ n4275;
  assign n4273 = x11 & x63;
  assign n4279 = n4278 ^ n4273;
  assign n4285 = n4284 ^ n4279;
  assign n4308 = n4307 ^ n4285;
  assign n4345 = n4344 ^ n4308;
  assign n4349 = n4348 ^ n4345;
  assign n4378 = n4377 ^ n4349;
  assign n4382 = n4381 ^ n4378;
  assign n4386 = n4385 ^ n4382;
  assign n4390 = n4389 ^ n4386;
  assign n4495 = n4389 ^ n4382;
  assign n4496 = ~n4386 & ~n4495;
  assign n4497 = n4496 ^ n4389;
  assign n4491 = n4381 ^ n4377;
  assign n4492 = ~n4378 & n4491;
  assign n4493 = n4492 ^ n4349;
  assign n4487 = n4376 ^ n4371;
  assign n4488 = ~n4372 & n4487;
  assign n4489 = n4488 ^ n4367;
  assign n4482 = n4348 ^ n4344;
  assign n4483 = ~n4345 & ~n4482;
  assign n4484 = n4483 ^ n4308;
  assign n4478 = n4361 ^ n4357;
  assign n4479 = ~n4366 & n4478;
  assign n4480 = n4479 ^ n4357;
  assign n4473 = n4356 ^ n4352;
  assign n4474 = n4353 & ~n4473;
  assign n4475 = n4474 ^ n4167;
  assign n4468 = n4301 ^ n4290;
  assign n4469 = n4301 ^ n4295;
  assign n4470 = n4468 & ~n4469;
  assign n4471 = n4470 ^ n4290;
  assign n4464 = x20 & n1556;
  assign n4465 = n4464 ^ n1664;
  assign n4462 = x19 & n1661;
  assign n4463 = n4462 ^ n1878;
  assign n4466 = n4465 ^ n4463;
  assign n4459 = ~x30 & n567;
  assign n4460 = n4459 ^ n672;
  assign n4457 = ~x29 & n669;
  assign n4458 = n4457 ^ n738;
  assign n4461 = n4460 ^ n4458;
  assign n4467 = n4466 ^ n4461;
  assign n4472 = n4471 ^ n4467;
  assign n4476 = n4475 ^ n4472;
  assign n4453 = n4337 ^ n4331;
  assign n4454 = n4332 & ~n4453;
  assign n4455 = n4454 ^ n4326;
  assign n4449 = n4320 ^ n4314;
  assign n4450 = ~n4315 & ~n4449;
  assign n4451 = n4450 ^ n4309;
  assign n4446 = n4284 ^ n4278;
  assign n4447 = n4279 & ~n4446;
  assign n4448 = n4447 ^ n4273;
  assign n4452 = n4451 ^ n4448;
  assign n4456 = n4455 ^ n4452;
  assign n4477 = n4476 ^ n4456;
  assign n4481 = n4480 ^ n4477;
  assign n4485 = n4484 ^ n4481;
  assign n4441 = n4343 ^ n4338;
  assign n4442 = ~n4339 & ~n4441;
  assign n4443 = n4442 ^ n4321;
  assign n4438 = n4302 ^ n4285;
  assign n4439 = ~n4307 & n4438;
  assign n4440 = n4439 ^ n4285;
  assign n4444 = n4443 ^ n4440;
  assign n4431 = x14 & n2387;
  assign n4432 = n4431 ^ n2635;
  assign n4429 = x13 & n2631;
  assign n4430 = n4429 ^ n2632;
  assign n4433 = n4432 ^ n4430;
  assign n4426 = x24 & n1105;
  assign n4427 = n4426 ^ n1206;
  assign n4424 = x23 & n1203;
  assign n4425 = n4424 ^ n1379;
  assign n4428 = n4427 ^ n4425;
  assign n4434 = n4433 ^ n4428;
  assign n4423 = x12 & x63;
  assign n4435 = n4434 ^ n4423;
  assign n4419 = x22 & n1360;
  assign n4420 = n4419 ^ n1447;
  assign n4417 = x21 & n1444;
  assign n4418 = n4417 ^ n1588;
  assign n4421 = n4420 ^ n4418;
  assign n4413 = x28 & n756;
  assign n4414 = n4413 ^ n873;
  assign n4411 = x27 & n870;
  assign n4412 = n4411 ^ n953;
  assign n4415 = n4414 ^ n4412;
  assign n4408 = x31 & n524;
  assign n4409 = n4408 ^ n527;
  assign n4410 = n4409 ^ n611;
  assign n4416 = n4415 ^ n4410;
  assign n4422 = n4421 ^ n4416;
  assign n4436 = n4435 ^ n4422;
  assign n4404 = x16 & n2143;
  assign n4405 = n4404 ^ n2275;
  assign n4402 = x15 & n2272;
  assign n4403 = n4402 ^ n2484;
  assign n4406 = n4405 ^ n4403;
  assign n4398 = ~x26 & n894;
  assign n4399 = n4398 ^ n1052;
  assign n4396 = ~x25 & n1049;
  assign n4397 = n4396 ^ n1087;
  assign n4400 = n4399 ^ n4397;
  assign n4393 = ~x18 & n1815;
  assign n4394 = n4393 ^ n2047;
  assign n4391 = ~x17 & n2044;
  assign n4392 = n4391 ^ n2162;
  assign n4395 = n4394 ^ n4392;
  assign n4401 = n4400 ^ n4395;
  assign n4407 = n4406 ^ n4401;
  assign n4437 = n4436 ^ n4407;
  assign n4445 = n4444 ^ n4437;
  assign n4486 = n4485 ^ n4445;
  assign n4490 = n4489 ^ n4486;
  assign n4494 = n4493 ^ n4490;
  assign n4498 = n4497 ^ n4494;
  assign n4602 = n4497 ^ n4490;
  assign n4603 = n4494 & ~n4602;
  assign n4604 = n4603 ^ n4497;
  assign n4598 = n4489 ^ n4485;
  assign n4599 = ~n4486 & ~n4598;
  assign n4600 = n4599 ^ n4445;
  assign n4594 = n4484 ^ n4480;
  assign n4595 = n4481 & ~n4594;
  assign n4596 = n4595 ^ n4477;
  assign n4590 = n4440 ^ n4437;
  assign n4591 = n4444 & n4590;
  assign n4592 = n4591 ^ n4437;
  assign n4584 = n4472 ^ n4456;
  assign n4585 = n4475 ^ n4456;
  assign n4586 = n4584 & n4585;
  assign n4587 = n4586 ^ n4472;
  assign n4580 = n4471 ^ n4466;
  assign n4581 = ~n4467 & ~n4580;
  assign n4582 = n4581 ^ n4461;
  assign n4575 = n4455 ^ n4448;
  assign n4576 = n4455 ^ n4451;
  assign n4577 = n4575 & n4576;
  assign n4578 = n4577 ^ n4448;
  assign n4570 = x23 & n1360;
  assign n4571 = n4570 ^ n1447;
  assign n4568 = x22 & n1444;
  assign n4569 = n4568 ^ n1588;
  assign n4572 = n4571 ^ n4569;
  assign n4565 = x21 & n1556;
  assign n4566 = n4565 ^ n1664;
  assign n4563 = x20 & n1661;
  assign n4564 = n4563 ^ n1878;
  assign n4567 = n4566 ^ n4564;
  assign n4573 = n4572 ^ n4567;
  assign n4574 = n4573 ^ n4461;
  assign n4579 = n4578 ^ n4574;
  assign n4583 = n4582 ^ n4579;
  assign n4588 = n4587 ^ n4583;
  assign n4557 = n4422 ^ n4407;
  assign n4558 = n4435 ^ n4407;
  assign n4559 = n4557 & ~n4558;
  assign n4560 = n4559 ^ n4422;
  assign n4553 = n4428 ^ n4423;
  assign n4554 = ~n4434 & n4553;
  assign n4555 = n4554 ^ n4423;
  assign n4548 = n4406 ^ n4395;
  assign n4549 = n4406 ^ n4400;
  assign n4550 = n4548 & ~n4549;
  assign n4551 = n4550 ^ n4395;
  assign n4544 = n4421 ^ n4410;
  assign n4545 = n4421 ^ n4415;
  assign n4546 = n4544 & ~n4545;
  assign n4547 = n4546 ^ n4410;
  assign n4552 = n4551 ^ n4547;
  assign n4556 = n4555 ^ n4552;
  assign n4561 = n4560 ^ n4556;
  assign n4538 = x29 & n756;
  assign n4539 = n4538 ^ n873;
  assign n4536 = x28 & n870;
  assign n4537 = n4536 ^ n953;
  assign n4540 = n4539 ^ n4537;
  assign n4532 = x15 & n2387;
  assign n4533 = n4532 ^ n2635;
  assign n4530 = x14 & n2631;
  assign n4531 = n4530 ^ n2632;
  assign n4534 = n4533 ^ n4531;
  assign n4529 = x13 & x63;
  assign n4535 = n4534 ^ n4529;
  assign n4541 = n4540 ^ n4535;
  assign n4525 = x25 & n1105;
  assign n4526 = n4525 ^ n1206;
  assign n4523 = x24 & n1203;
  assign n4524 = n4523 ^ n1379;
  assign n4527 = n4526 ^ n4524;
  assign n4519 = x17 & n2143;
  assign n4520 = n4519 ^ n2275;
  assign n4517 = x16 & n2272;
  assign n4518 = n4517 ^ n2484;
  assign n4521 = n4520 ^ n4518;
  assign n4514 = ~x19 & n1815;
  assign n4515 = n4514 ^ n2047;
  assign n4512 = ~x18 & n2044;
  assign n4513 = n4512 ^ n2162;
  assign n4516 = n4515 ^ n4513;
  assign n4522 = n4521 ^ n4516;
  assign n4528 = n4527 ^ n4522;
  assign n4542 = n4541 ^ n4528;
  assign n4508 = ~x27 & n894;
  assign n4509 = n4508 ^ n1052;
  assign n4506 = ~x26 & n1049;
  assign n4507 = n4506 ^ n1087;
  assign n4510 = n4509 ^ n4507;
  assign n4502 = ~x31 & n567;
  assign n4503 = n4502 ^ n672;
  assign n4500 = ~x30 & n669;
  assign n4501 = n4500 ^ n738;
  assign n4504 = n4503 ^ n4501;
  assign n4499 = n611 ^ n527;
  assign n4505 = n4504 ^ n4499;
  assign n4511 = n4510 ^ n4505;
  assign n4543 = n4542 ^ n4511;
  assign n4562 = n4561 ^ n4543;
  assign n4589 = n4588 ^ n4562;
  assign n4593 = n4592 ^ n4589;
  assign n4597 = n4596 ^ n4593;
  assign n4601 = n4600 ^ n4597;
  assign n4605 = n4604 ^ n4601;
  assign n4704 = n4604 ^ n4597;
  assign n4705 = ~n4601 & ~n4704;
  assign n4706 = n4705 ^ n4604;
  assign n4700 = n4596 ^ n4592;
  assign n4701 = ~n4593 & ~n4700;
  assign n4702 = n4701 ^ n4589;
  assign n4696 = n4583 ^ n4562;
  assign n4697 = ~n4588 & n4696;
  assign n4698 = n4697 ^ n4562;
  assign n4691 = n4560 ^ n4543;
  assign n4692 = ~n4561 & ~n4691;
  assign n4693 = n4692 ^ n4543;
  assign n4686 = n4582 ^ n4574;
  assign n4687 = n4582 ^ n4578;
  assign n4688 = ~n4686 & n4687;
  assign n4689 = n4688 ^ n4574;
  assign n4682 = n4555 ^ n4551;
  assign n4683 = n4552 & ~n4682;
  assign n4684 = n4683 ^ n4547;
  assign n4677 = n4567 ^ n4461;
  assign n4678 = n4572 ^ n4461;
  assign n4679 = n4677 & ~n4678;
  assign n4680 = n4679 ^ n4567;
  assign n4673 = ~x20 & n1815;
  assign n4674 = n4673 ^ n2047;
  assign n4671 = ~x19 & n2044;
  assign n4672 = n4671 ^ n2162;
  assign n4675 = n4674 ^ n4672;
  assign n4667 = ~x28 & n894;
  assign n4668 = n4667 ^ n1052;
  assign n4665 = ~x27 & n1049;
  assign n4666 = n4665 ^ n1087;
  assign n4669 = n4668 ^ n4666;
  assign n4662 = x22 & n1556;
  assign n4663 = n4662 ^ n1664;
  assign n4660 = x21 & n1661;
  assign n4661 = n4660 ^ n1878;
  assign n4664 = n4663 ^ n4661;
  assign n4670 = n4669 ^ n4664;
  assign n4676 = n4675 ^ n4670;
  assign n4681 = n4680 ^ n4676;
  assign n4685 = n4684 ^ n4681;
  assign n4690 = n4689 ^ n4685;
  assign n4694 = n4693 ^ n4690;
  assign n4655 = n4528 ^ n4511;
  assign n4656 = ~n4542 & ~n4655;
  assign n4657 = n4656 ^ n4511;
  assign n4651 = n4527 ^ n4516;
  assign n4652 = ~n4522 & n4651;
  assign n4653 = n4652 ^ n4527;
  assign n4647 = x31 & n669;
  assign n4646 = n672 ^ n567;
  assign n4648 = n4647 ^ n4646;
  assign n4645 = n738 ^ n669;
  assign n4649 = n4648 ^ n4645;
  assign n4642 = n4510 ^ n4504;
  assign n4643 = ~n4505 & ~n4642;
  assign n4644 = n4643 ^ n4499;
  assign n4650 = n4649 ^ n4644;
  assign n4654 = n4653 ^ n4650;
  assign n4658 = n4657 ^ n4654;
  assign n4636 = n4540 ^ n4529;
  assign n4637 = n4540 ^ n4534;
  assign n4638 = n4636 & ~n4637;
  assign n4639 = n4638 ^ n4529;
  assign n4632 = x16 & n2387;
  assign n4633 = n4632 ^ n2635;
  assign n4630 = x15 & n2631;
  assign n4631 = n4630 ^ n2632;
  assign n4634 = n4633 ^ n4631;
  assign n4626 = x18 & n2143;
  assign n4627 = n4626 ^ n2275;
  assign n4624 = x17 & n2272;
  assign n4625 = n4624 ^ n2484;
  assign n4628 = n4627 ^ n4625;
  assign n4621 = x26 & n1105;
  assign n4622 = n4621 ^ n1206;
  assign n4619 = x25 & n1203;
  assign n4620 = n4619 ^ n1379;
  assign n4623 = n4622 ^ n4620;
  assign n4629 = n4628 ^ n4623;
  assign n4635 = n4634 ^ n4629;
  assign n4640 = n4639 ^ n4635;
  assign n4615 = x24 & n1360;
  assign n4616 = n4615 ^ n1447;
  assign n4613 = x23 & n1444;
  assign n4614 = n4613 ^ n1588;
  assign n4617 = n4616 ^ n4614;
  assign n4609 = x30 & n756;
  assign n4610 = n4609 ^ n873;
  assign n4607 = x29 & n870;
  assign n4608 = n4607 ^ n953;
  assign n4611 = n4610 ^ n4608;
  assign n4606 = x14 & x63;
  assign n4612 = n4611 ^ n4606;
  assign n4618 = n4617 ^ n4612;
  assign n4641 = n4640 ^ n4618;
  assign n4659 = n4658 ^ n4641;
  assign n4695 = n4694 ^ n4659;
  assign n4699 = n4698 ^ n4695;
  assign n4703 = n4702 ^ n4699;
  assign n4707 = n4706 ^ n4703;
  assign n4799 = n4706 ^ n4699;
  assign n4800 = ~n4703 & ~n4799;
  assign n4801 = n4800 ^ n4706;
  assign n4795 = n4698 ^ n4694;
  assign n4796 = n4695 & ~n4795;
  assign n4797 = n4796 ^ n4659;
  assign n4790 = n4693 ^ n4685;
  assign n4791 = n4693 ^ n4689;
  assign n4792 = ~n4790 & n4791;
  assign n4793 = n4792 ^ n4685;
  assign n4785 = n4654 ^ n4641;
  assign n4786 = n4658 & n4785;
  assign n4787 = n4786 ^ n4641;
  assign n4781 = n4684 ^ n4680;
  assign n4782 = n4681 & ~n4781;
  assign n4783 = n4782 ^ n4676;
  assign n4776 = n4634 ^ n4628;
  assign n4777 = n4629 & ~n4776;
  assign n4778 = n4777 ^ n4623;
  assign n4772 = ~x21 & n1815;
  assign n4773 = n4772 ^ n2047;
  assign n4770 = ~x20 & n2044;
  assign n4771 = n4770 ^ n2162;
  assign n4774 = n4773 ^ n4771;
  assign n4775 = n4774 ^ n4649;
  assign n4779 = n4778 ^ n4775;
  assign n4765 = x25 & n1360;
  assign n4766 = n4765 ^ n1447;
  assign n4763 = x24 & n1444;
  assign n4764 = n4763 ^ n1588;
  assign n4767 = n4766 ^ n4764;
  assign n4759 = x17 & n2387;
  assign n4760 = n4759 ^ n2635;
  assign n4757 = x16 & n2631;
  assign n4758 = n4757 ^ n2632;
  assign n4761 = n4760 ^ n4758;
  assign n4754 = x19 & n2143;
  assign n4755 = n4754 ^ n2275;
  assign n4752 = x18 & n2272;
  assign n4753 = n4752 ^ n2484;
  assign n4756 = n4755 ^ n4753;
  assign n4762 = n4761 ^ n4756;
  assign n4768 = n4767 ^ n4762;
  assign n4748 = x27 & n1105;
  assign n4749 = n4748 ^ n1206;
  assign n4746 = x26 & n1203;
  assign n4747 = n4746 ^ n1379;
  assign n4750 = n4749 ^ n4747;
  assign n4742 = x31 & n756;
  assign n4743 = n4742 ^ n873;
  assign n4740 = x30 & n870;
  assign n4741 = n4740 ^ n953;
  assign n4744 = n4743 ^ n4741;
  assign n4739 = n4646 ^ n4645;
  assign n4745 = n4744 ^ n4739;
  assign n4751 = n4750 ^ n4745;
  assign n4769 = n4768 ^ n4751;
  assign n4780 = n4779 ^ n4769;
  assign n4784 = n4783 ^ n4780;
  assign n4788 = n4787 ^ n4784;
  assign n4733 = n4653 ^ n4649;
  assign n4734 = n4653 ^ n4644;
  assign n4735 = ~n4733 & n4734;
  assign n4736 = n4735 ^ n4649;
  assign n4730 = n4635 ^ n4618;
  assign n4731 = ~n4640 & n4730;
  assign n4732 = n4731 ^ n4618;
  assign n4737 = n4736 ^ n4732;
  assign n4724 = n4675 ^ n4664;
  assign n4725 = n4675 ^ n4669;
  assign n4726 = n4724 & ~n4725;
  assign n4727 = n4726 ^ n4664;
  assign n4721 = n4617 ^ n4611;
  assign n4722 = n4612 & ~n4721;
  assign n4723 = n4722 ^ n4606;
  assign n4728 = n4727 ^ n4723;
  assign n4717 = x23 & n1556;
  assign n4718 = n4717 ^ n1664;
  assign n4715 = x22 & n1661;
  assign n4716 = n4715 ^ n1878;
  assign n4719 = n4718 ^ n4716;
  assign n4711 = ~x29 & n894;
  assign n4712 = n4711 ^ n1052;
  assign n4709 = ~x28 & n1049;
  assign n4710 = n4709 ^ n1087;
  assign n4713 = n4712 ^ n4710;
  assign n4708 = x15 & x63;
  assign n4714 = n4713 ^ n4708;
  assign n4720 = n4719 ^ n4714;
  assign n4729 = n4728 ^ n4720;
  assign n4738 = n4737 ^ n4729;
  assign n4789 = n4788 ^ n4738;
  assign n4794 = n4793 ^ n4789;
  assign n4798 = n4797 ^ n4794;
  assign n4802 = n4801 ^ n4798;
  assign n4887 = n4801 ^ n4794;
  assign n4888 = n4798 & n4887;
  assign n4889 = n4888 ^ n4801;
  assign n4883 = n4793 ^ n4788;
  assign n4884 = n4789 & n4883;
  assign n4885 = n4884 ^ n4738;
  assign n4878 = n4787 ^ n4780;
  assign n4879 = n4787 ^ n4783;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = n4880 ^ n4780;
  assign n4873 = n4732 ^ n4729;
  assign n4874 = n4737 & n4873;
  assign n4875 = n4874 ^ n4729;
  assign n4869 = n4779 ^ n4768;
  assign n4870 = ~n4769 & ~n4869;
  assign n4871 = n4870 ^ n4751;
  assign n4862 = x26 & n1360;
  assign n4863 = n4862 ^ n1447;
  assign n4860 = x25 & n1444;
  assign n4861 = n4860 ^ n1588;
  assign n4864 = n4863 ^ n4861;
  assign n4857 = x18 & n2387;
  assign n4858 = n4857 ^ n2635;
  assign n4855 = x17 & n2631;
  assign n4856 = n4855 ^ n2632;
  assign n4859 = n4858 ^ n4856;
  assign n4865 = n4864 ^ n4859;
  assign n4854 = x16 & x63;
  assign n4866 = n4865 ^ n4854;
  assign n4850 = x28 & n1105;
  assign n4851 = n4850 ^ n1206;
  assign n4848 = x27 & n1203;
  assign n4849 = n4848 ^ n1379;
  assign n4852 = n4851 ^ n4849;
  assign n4844 = ~x30 & n894;
  assign n4845 = n4844 ^ n1052;
  assign n4842 = ~x29 & n1049;
  assign n4843 = n4842 ^ n1087;
  assign n4846 = n4845 ^ n4843;
  assign n4839 = x24 & n1556;
  assign n4840 = n4839 ^ n1664;
  assign n4837 = x23 & n1661;
  assign n4838 = n4837 ^ n1878;
  assign n4841 = n4840 ^ n4838;
  assign n4847 = n4846 ^ n4841;
  assign n4853 = n4852 ^ n4847;
  assign n4867 = n4866 ^ n4853;
  assign n4833 = x31 & n870;
  assign n4834 = n4833 ^ n873;
  assign n4835 = n4834 ^ n953;
  assign n4829 = ~x22 & n1815;
  assign n4830 = n4829 ^ n2047;
  assign n4827 = ~x21 & n2044;
  assign n4828 = n4827 ^ n2162;
  assign n4831 = n4830 ^ n4828;
  assign n4824 = x20 & n2143;
  assign n4825 = n4824 ^ n2275;
  assign n4822 = x19 & n2272;
  assign n4823 = n4822 ^ n2484;
  assign n4826 = n4825 ^ n4823;
  assign n4832 = n4831 ^ n4826;
  assign n4836 = n4835 ^ n4832;
  assign n4868 = n4867 ^ n4836;
  assign n4872 = n4871 ^ n4868;
  assign n4876 = n4875 ^ n4872;
  assign n4817 = n4723 ^ n4720;
  assign n4818 = ~n4728 & n4817;
  assign n4819 = n4818 ^ n4720;
  assign n4814 = n4778 ^ n4774;
  assign n4815 = n4775 & ~n4814;
  assign n4816 = n4815 ^ n4649;
  assign n4820 = n4819 ^ n4816;
  assign n4810 = n4719 ^ n4713;
  assign n4811 = n4714 & ~n4810;
  assign n4812 = n4811 ^ n4708;
  assign n4806 = n4767 ^ n4761;
  assign n4807 = n4762 & ~n4806;
  assign n4808 = n4807 ^ n4756;
  assign n4803 = n4750 ^ n4744;
  assign n4804 = ~n4745 & ~n4803;
  assign n4805 = n4804 ^ n4739;
  assign n4809 = n4808 ^ n4805;
  assign n4813 = n4812 ^ n4809;
  assign n4821 = n4820 ^ n4813;
  assign n4877 = n4876 ^ n4821;
  assign n4882 = n4881 ^ n4877;
  assign n4886 = n4885 ^ n4882;
  assign n4890 = n4889 ^ n4886;
  assign n4969 = n4889 ^ n4882;
  assign n4970 = n4886 & n4969;
  assign n4971 = n4970 ^ n4889;
  assign n4965 = n4881 ^ n4876;
  assign n4966 = ~n4877 & n4965;
  assign n4967 = n4966 ^ n4821;
  assign n4961 = n4875 ^ n4871;
  assign n4962 = n4872 & n4961;
  assign n4963 = n4962 ^ n4868;
  assign n4956 = n4816 ^ n4813;
  assign n4957 = ~n4820 & ~n4956;
  assign n4958 = n4957 ^ n4813;
  assign n4952 = n4853 ^ n4836;
  assign n4953 = ~n4867 & ~n4952;
  assign n4954 = n4953 ^ n4836;
  assign n4946 = x27 & n1360;
  assign n4947 = n4946 ^ n1447;
  assign n4944 = x26 & n1444;
  assign n4945 = n4944 ^ n1588;
  assign n4948 = n4947 ^ n4945;
  assign n4940 = ~x31 & n894;
  assign n4941 = n4940 ^ n1052;
  assign n4938 = ~x30 & n1049;
  assign n4939 = n4938 ^ n1087;
  assign n4942 = n4941 ^ n4939;
  assign n4937 = n953 ^ n873;
  assign n4943 = n4942 ^ n4937;
  assign n4949 = n4948 ^ n4943;
  assign n4933 = x21 & n2143;
  assign n4934 = n4933 ^ n2275;
  assign n4931 = x20 & n2272;
  assign n4932 = n4931 ^ n2484;
  assign n4935 = n4934 ^ n4932;
  assign n4927 = ~x23 & n1815;
  assign n4928 = n4927 ^ n2047;
  assign n4925 = ~x22 & n2044;
  assign n4926 = n4925 ^ n2162;
  assign n4929 = n4928 ^ n4926;
  assign n4922 = x29 & n1105;
  assign n4923 = n4922 ^ n1206;
  assign n4920 = x28 & n1203;
  assign n4921 = n4920 ^ n1379;
  assign n4924 = n4923 ^ n4921;
  assign n4930 = n4929 ^ n4924;
  assign n4936 = n4935 ^ n4930;
  assign n4950 = n4949 ^ n4936;
  assign n4916 = x25 & n1556;
  assign n4917 = n4916 ^ n1664;
  assign n4914 = x24 & n1661;
  assign n4915 = n4914 ^ n1878;
  assign n4918 = n4917 ^ n4915;
  assign n4910 = x19 & n2387;
  assign n4911 = n4910 ^ n2635;
  assign n4908 = x18 & n2631;
  assign n4909 = n4908 ^ n2632;
  assign n4912 = n4911 ^ n4909;
  assign n4907 = x17 & x63;
  assign n4913 = n4912 ^ n4907;
  assign n4919 = n4918 ^ n4913;
  assign n4951 = n4950 ^ n4919;
  assign n4955 = n4954 ^ n4951;
  assign n4959 = n4958 ^ n4955;
  assign n4902 = n4812 ^ n4805;
  assign n4903 = n4809 & ~n4902;
  assign n4904 = n4903 ^ n4812;
  assign n4899 = n4835 ^ n4826;
  assign n4900 = ~n4832 & ~n4899;
  assign n4901 = n4900 ^ n4835;
  assign n4905 = n4904 ^ n4901;
  assign n4895 = n4852 ^ n4846;
  assign n4896 = n4847 & ~n4895;
  assign n4897 = n4896 ^ n4841;
  assign n4891 = n4859 ^ n4854;
  assign n4892 = ~n4865 & n4891;
  assign n4893 = n4892 ^ n4854;
  assign n4894 = n4893 ^ n4835;
  assign n4898 = n4897 ^ n4894;
  assign n4906 = n4905 ^ n4898;
  assign n4960 = n4959 ^ n4906;
  assign n4964 = n4963 ^ n4960;
  assign n4968 = n4967 ^ n4964;
  assign n4972 = n4971 ^ n4968;
  assign n5051 = n4971 ^ n4964;
  assign n5052 = ~n4968 & ~n5051;
  assign n5053 = n5052 ^ n4971;
  assign n5047 = n4963 ^ n4959;
  assign n5048 = n4960 & ~n5047;
  assign n5049 = n5048 ^ n4906;
  assign n5043 = n4958 ^ n4954;
  assign n5044 = n4955 & ~n5043;
  assign n5045 = n5044 ^ n4951;
  assign n5038 = n4901 ^ n4898;
  assign n5039 = n4904 ^ n4898;
  assign n5040 = ~n5038 & ~n5039;
  assign n5041 = n5040 ^ n4901;
  assign n5033 = n4897 ^ n4893;
  assign n5034 = n4894 & ~n5033;
  assign n5035 = n5034 ^ n4835;
  assign n5027 = n4948 ^ n4937;
  assign n5028 = n4948 ^ n4942;
  assign n5029 = ~n5027 & ~n5028;
  assign n5030 = n5029 ^ n4937;
  assign n5023 = x20 & n2387;
  assign n5024 = n5023 ^ n2635;
  assign n5021 = x19 & n2631;
  assign n5022 = n5021 ^ n2632;
  assign n5025 = n5024 ^ n5022;
  assign n5018 = x31 & n1049;
  assign n5017 = n1052 ^ n894;
  assign n5019 = n5018 ^ n5017;
  assign n5016 = n1087 ^ n1049;
  assign n5020 = n5019 ^ n5016;
  assign n5026 = n5025 ^ n5020;
  assign n5031 = n5030 ^ n5026;
  assign n5012 = x26 & n1556;
  assign n5013 = n5012 ^ n1664;
  assign n5010 = x25 & n1661;
  assign n5011 = n5010 ^ n1878;
  assign n5014 = n5013 ^ n5011;
  assign n5006 = x30 & n1105;
  assign n5007 = n5006 ^ n1206;
  assign n5004 = x29 & n1203;
  assign n5005 = n5004 ^ n1379;
  assign n5008 = n5007 ^ n5005;
  assign n5003 = x18 & x63;
  assign n5009 = n5008 ^ n5003;
  assign n5015 = n5014 ^ n5009;
  assign n5032 = n5031 ^ n5015;
  assign n5036 = n5035 ^ n5032;
  assign n4999 = n4949 ^ n4919;
  assign n5000 = ~n4950 & n4999;
  assign n5001 = n5000 ^ n4936;
  assign n4994 = n4935 ^ n4929;
  assign n4995 = n4930 & ~n4994;
  assign n4996 = n4995 ^ n4924;
  assign n4990 = n4918 ^ n4907;
  assign n4991 = n4918 ^ n4912;
  assign n4992 = n4990 & ~n4991;
  assign n4993 = n4992 ^ n4907;
  assign n4997 = n4996 ^ n4993;
  assign n4986 = x22 & n2143;
  assign n4987 = n4986 ^ n2275;
  assign n4984 = x21 & n2272;
  assign n4985 = n4984 ^ n2484;
  assign n4988 = n4987 ^ n4985;
  assign n4980 = x28 & n1360;
  assign n4981 = n4980 ^ n1447;
  assign n4978 = x27 & n1444;
  assign n4979 = n4978 ^ n1588;
  assign n4982 = n4981 ^ n4979;
  assign n4975 = ~x24 & n1815;
  assign n4976 = n4975 ^ n2047;
  assign n4973 = ~x23 & n2044;
  assign n4974 = n4973 ^ n2162;
  assign n4977 = n4976 ^ n4974;
  assign n4983 = n4982 ^ n4977;
  assign n4989 = n4988 ^ n4983;
  assign n4998 = n4997 ^ n4989;
  assign n5002 = n5001 ^ n4998;
  assign n5037 = n5036 ^ n5002;
  assign n5042 = n5041 ^ n5037;
  assign n5046 = n5045 ^ n5042;
  assign n5050 = n5049 ^ n5046;
  assign n5054 = n5053 ^ n5050;
  assign n5123 = n5053 ^ n5046;
  assign n5124 = n5050 & n5123;
  assign n5125 = n5124 ^ n5053;
  assign n5119 = n5045 ^ n5041;
  assign n5120 = ~n5042 & ~n5119;
  assign n5121 = n5120 ^ n5037;
  assign n5115 = n5036 ^ n5001;
  assign n5116 = n5002 & ~n5115;
  assign n5117 = n5116 ^ n4998;
  assign n5110 = n5035 ^ n5031;
  assign n5111 = n5032 & ~n5110;
  assign n5112 = n5111 ^ n5015;
  assign n5106 = n4993 ^ n4989;
  assign n5107 = ~n4997 & n5106;
  assign n5108 = n5107 ^ n4989;
  assign n5101 = n4988 ^ n4977;
  assign n5102 = ~n4983 & n5101;
  assign n5103 = n5102 ^ n4988;
  assign n5098 = n5014 ^ n5008;
  assign n5099 = n5009 & ~n5098;
  assign n5100 = n5099 ^ n5003;
  assign n5104 = n5103 ^ n5100;
  assign n5094 = x27 & n1556;
  assign n5095 = n5094 ^ n1664;
  assign n5092 = x26 & n1661;
  assign n5093 = n5092 ^ n1878;
  assign n5096 = n5095 ^ n5093;
  assign n5088 = x31 & n1105;
  assign n5089 = n5088 ^ n1206;
  assign n5086 = x30 & n1203;
  assign n5087 = n5086 ^ n1379;
  assign n5090 = n5089 ^ n5087;
  assign n5085 = n5017 ^ n5016;
  assign n5091 = n5090 ^ n5085;
  assign n5097 = n5096 ^ n5091;
  assign n5105 = n5104 ^ n5097;
  assign n5109 = n5108 ^ n5105;
  assign n5113 = n5112 ^ n5109;
  assign n5081 = n5030 ^ n5025;
  assign n5082 = ~n5026 & n5081;
  assign n5083 = n5082 ^ n5020;
  assign n5076 = x29 & n1360;
  assign n5077 = n5076 ^ n1447;
  assign n5074 = x28 & n1444;
  assign n5075 = n5074 ^ n1588;
  assign n5078 = n5077 ^ n5075;
  assign n5070 = ~x25 & n1815;
  assign n5071 = n5070 ^ n2047;
  assign n5068 = ~x24 & n2044;
  assign n5069 = n5068 ^ n2162;
  assign n5072 = n5071 ^ n5069;
  assign n5067 = x19 & x63;
  assign n5073 = n5072 ^ n5067;
  assign n5079 = n5078 ^ n5073;
  assign n5062 = x21 & n2387;
  assign n5063 = n5062 ^ n2635;
  assign n5060 = x20 & n2631;
  assign n5061 = n5060 ^ n2632;
  assign n5064 = n5063 ^ n5061;
  assign n5057 = x23 & n2143;
  assign n5058 = n5057 ^ n2275;
  assign n5055 = x22 & n2272;
  assign n5056 = n5055 ^ n2484;
  assign n5059 = n5058 ^ n5056;
  assign n5065 = n5064 ^ n5059;
  assign n5066 = n5065 ^ n5020;
  assign n5080 = n5079 ^ n5066;
  assign n5084 = n5083 ^ n5080;
  assign n5114 = n5113 ^ n5084;
  assign n5118 = n5117 ^ n5114;
  assign n5122 = n5121 ^ n5118;
  assign n5126 = n5125 ^ n5122;
  assign n5191 = n5125 ^ n5118;
  assign n5192 = ~n5122 & n5191;
  assign n5193 = n5192 ^ n5125;
  assign n5186 = n5117 ^ n5084;
  assign n5187 = n5117 ^ n5113;
  assign n5188 = ~n5186 & n5187;
  assign n5189 = n5188 ^ n5084;
  assign n5182 = n5112 ^ n5108;
  assign n5183 = ~n5109 & ~n5182;
  assign n5184 = n5183 ^ n5105;
  assign n5178 = n5083 ^ n5079;
  assign n5179 = n5080 & n5178;
  assign n5180 = n5179 ^ n5066;
  assign n5173 = n5100 ^ n5097;
  assign n5174 = ~n5104 & ~n5173;
  assign n5175 = n5174 ^ n5097;
  assign n5169 = n5078 ^ n5072;
  assign n5170 = n5073 & ~n5169;
  assign n5171 = n5170 ^ n5067;
  assign n5165 = x31 & n1203;
  assign n5166 = n5165 ^ n1206;
  assign n5167 = n5166 ^ n1379;
  assign n5162 = n5096 ^ n5090;
  assign n5163 = ~n5091 & ~n5162;
  assign n5164 = n5163 ^ n5085;
  assign n5168 = n5167 ^ n5164;
  assign n5172 = n5171 ^ n5168;
  assign n5176 = n5175 ^ n5172;
  assign n5158 = n5059 ^ n5020;
  assign n5159 = ~n5065 & n5158;
  assign n5160 = n5159 ^ n5020;
  assign n5153 = x24 & n2143;
  assign n5154 = n5153 ^ n2275;
  assign n5151 = x23 & n2272;
  assign n5152 = n5151 ^ n2484;
  assign n5155 = n5154 ^ n5152;
  assign n5147 = ~x26 & n1815;
  assign n5148 = n5147 ^ n2047;
  assign n5145 = ~x25 & n2044;
  assign n5146 = n5145 ^ n2162;
  assign n5149 = n5148 ^ n5146;
  assign n5142 = x30 & n1360;
  assign n5143 = n5142 ^ n1447;
  assign n5140 = x29 & n1444;
  assign n5141 = n5140 ^ n1588;
  assign n5144 = n5143 ^ n5141;
  assign n5150 = n5149 ^ n5144;
  assign n5156 = n5155 ^ n5150;
  assign n5135 = x22 & n2387;
  assign n5136 = n5135 ^ n2635;
  assign n5133 = x21 & n2631;
  assign n5134 = n5133 ^ n2632;
  assign n5137 = n5136 ^ n5134;
  assign n5130 = x28 & n1556;
  assign n5131 = n5130 ^ n1664;
  assign n5128 = x27 & n1661;
  assign n5129 = n5128 ^ n1878;
  assign n5132 = n5131 ^ n5129;
  assign n5138 = n5137 ^ n5132;
  assign n5127 = x20 & x63;
  assign n5139 = n5138 ^ n5127;
  assign n5157 = n5156 ^ n5139;
  assign n5161 = n5160 ^ n5157;
  assign n5177 = n5176 ^ n5161;
  assign n5181 = n5180 ^ n5177;
  assign n5185 = n5184 ^ n5181;
  assign n5190 = n5189 ^ n5185;
  assign n5194 = n5193 ^ n5190;
  assign n5254 = n5193 ^ n5185;
  assign n5255 = n5190 & n5254;
  assign n5256 = n5255 ^ n5193;
  assign n5250 = n5184 ^ n5180;
  assign n5251 = ~n5181 & n5250;
  assign n5252 = n5251 ^ n5177;
  assign n5246 = n5172 ^ n5161;
  assign n5247 = n5176 & n5246;
  assign n5248 = n5247 ^ n5161;
  assign n5241 = n5160 ^ n5156;
  assign n5242 = n5157 & ~n5241;
  assign n5243 = n5242 ^ n5139;
  assign n5236 = n5171 ^ n5167;
  assign n5237 = n5171 ^ n5164;
  assign n5238 = ~n5236 & n5237;
  assign n5239 = n5238 ^ n5167;
  assign n5232 = n5155 ^ n5149;
  assign n5233 = n5150 & ~n5232;
  assign n5234 = n5233 ^ n5144;
  assign n5230 = x21 & x63;
  assign n5231 = n5230 ^ n5167;
  assign n5235 = n5234 ^ n5231;
  assign n5240 = n5239 ^ n5235;
  assign n5244 = n5243 ^ n5240;
  assign n5225 = n5132 ^ n5127;
  assign n5226 = ~n5138 & n5225;
  assign n5227 = n5226 ^ n5127;
  assign n5221 = x23 & n2387;
  assign n5222 = n5221 ^ n2635;
  assign n5219 = x22 & n2631;
  assign n5220 = n5219 ^ n2632;
  assign n5223 = n5222 ^ n5220;
  assign n5215 = x29 & n1556;
  assign n5216 = n5215 ^ n1664;
  assign n5213 = x28 & n1661;
  assign n5214 = n5213 ^ n1878;
  assign n5217 = n5216 ^ n5214;
  assign n5210 = x25 & n2143;
  assign n5211 = n5210 ^ n2275;
  assign n5208 = x24 & n2272;
  assign n5209 = n5208 ^ n2484;
  assign n5212 = n5211 ^ n5209;
  assign n5218 = n5217 ^ n5212;
  assign n5224 = n5223 ^ n5218;
  assign n5228 = n5227 ^ n5224;
  assign n5204 = ~x27 & n1815;
  assign n5205 = n5204 ^ n2047;
  assign n5202 = ~x26 & n2044;
  assign n5203 = n5202 ^ n2162;
  assign n5206 = n5205 ^ n5203;
  assign n5198 = x31 & n1360;
  assign n5199 = n5198 ^ n1447;
  assign n5196 = x30 & n1444;
  assign n5197 = n5196 ^ n1588;
  assign n5200 = n5199 ^ n5197;
  assign n5195 = n1379 ^ n1206;
  assign n5201 = n5200 ^ n5195;
  assign n5207 = n5206 ^ n5201;
  assign n5229 = n5228 ^ n5207;
  assign n5245 = n5244 ^ n5229;
  assign n5249 = n5248 ^ n5245;
  assign n5253 = n5252 ^ n5249;
  assign n5257 = n5256 ^ n5253;
  assign n5314 = n5256 ^ n5249;
  assign n5315 = n5253 & n5314;
  assign n5316 = n5315 ^ n5256;
  assign n5310 = n5248 ^ n5244;
  assign n5311 = n5245 & n5310;
  assign n5312 = n5311 ^ n5229;
  assign n5305 = n5243 ^ n5235;
  assign n5306 = n5243 ^ n5239;
  assign n5307 = n5305 & n5306;
  assign n5308 = n5307 ^ n5235;
  assign n5299 = n5224 ^ n5207;
  assign n5300 = n5227 ^ n5207;
  assign n5301 = ~n5299 & n5300;
  assign n5302 = n5301 ^ n5224;
  assign n5295 = n5234 ^ n5167;
  assign n5296 = n5231 & ~n5295;
  assign n5297 = n5296 ^ n5230;
  assign n5291 = x30 & n1556;
  assign n5292 = n5291 ^ n1664;
  assign n5289 = x29 & n1661;
  assign n5290 = n5289 ^ n1878;
  assign n5293 = n5292 ^ n5290;
  assign n5285 = ~x28 & n1815;
  assign n5286 = n5285 ^ n2047;
  assign n5283 = ~x27 & n2044;
  assign n5284 = n5283 ^ n2162;
  assign n5287 = n5286 ^ n5284;
  assign n5282 = x22 & x63;
  assign n5288 = n5287 ^ n5282;
  assign n5294 = n5293 ^ n5288;
  assign n5298 = n5297 ^ n5294;
  assign n5303 = n5302 ^ n5298;
  assign n5276 = n5223 ^ n5212;
  assign n5277 = n5223 ^ n5217;
  assign n5278 = n5276 & ~n5277;
  assign n5279 = n5278 ^ n5212;
  assign n5273 = n5206 ^ n5200;
  assign n5274 = ~n5201 & ~n5273;
  assign n5275 = n5274 ^ n5195;
  assign n5280 = n5279 ^ n5275;
  assign n5269 = x31 & n1444;
  assign n5270 = n5269 ^ n1447;
  assign n5271 = n5270 ^ n1588;
  assign n5265 = x26 & n2143;
  assign n5266 = n5265 ^ n2275;
  assign n5263 = x25 & n2272;
  assign n5264 = n5263 ^ n2484;
  assign n5267 = n5266 ^ n5264;
  assign n5260 = x24 & n2387;
  assign n5261 = n5260 ^ n2635;
  assign n5258 = x23 & n2631;
  assign n5259 = n5258 ^ n2632;
  assign n5262 = n5261 ^ n5259;
  assign n5268 = n5267 ^ n5262;
  assign n5272 = n5271 ^ n5268;
  assign n5281 = n5280 ^ n5272;
  assign n5304 = n5303 ^ n5281;
  assign n5309 = n5308 ^ n5304;
  assign n5313 = n5312 ^ n5309;
  assign n5317 = n5316 ^ n5313;
  assign n5367 = n5316 ^ n5309;
  assign n5368 = n5313 & n5367;
  assign n5369 = n5368 ^ n5316;
  assign n5363 = n5308 ^ n5303;
  assign n5364 = n5304 & n5363;
  assign n5365 = n5364 ^ n5281;
  assign n5359 = n5302 ^ n5297;
  assign n5360 = ~n5298 & ~n5359;
  assign n5361 = n5360 ^ n5294;
  assign n5355 = n5275 ^ n5272;
  assign n5356 = n5280 & ~n5355;
  assign n5357 = n5356 ^ n5272;
  assign n5349 = n5293 ^ n5282;
  assign n5350 = n5293 ^ n5287;
  assign n5351 = ~n5349 & n5350;
  assign n5352 = n5351 ^ n5282;
  assign n5345 = x27 & n2143;
  assign n5346 = n5345 ^ n2275;
  assign n5343 = x26 & n2272;
  assign n5344 = n5343 ^ n2484;
  assign n5347 = n5346 ^ n5344;
  assign n5339 = x31 & n1556;
  assign n5340 = n5339 ^ n1664;
  assign n5337 = x30 & n1661;
  assign n5338 = n5337 ^ n1878;
  assign n5341 = n5340 ^ n5338;
  assign n5336 = n1588 ^ n1447;
  assign n5342 = n5341 ^ n5336;
  assign n5348 = n5347 ^ n5342;
  assign n5353 = n5352 ^ n5348;
  assign n5331 = n5271 ^ n5262;
  assign n5332 = ~n5268 & n5331;
  assign n5333 = n5332 ^ n5271;
  assign n5334 = n5333 ^ n5293;
  assign n5326 = x25 & n2387;
  assign n5327 = n5326 ^ n2635;
  assign n5324 = x24 & n2631;
  assign n5325 = n5324 ^ n2632;
  assign n5328 = n5327 ^ n5325;
  assign n5321 = ~x29 & n1815;
  assign n5322 = n5321 ^ n2047;
  assign n5319 = ~x28 & n2044;
  assign n5320 = n5319 ^ n2162;
  assign n5323 = n5322 ^ n5320;
  assign n5329 = n5328 ^ n5323;
  assign n5318 = x23 & x63;
  assign n5330 = n5329 ^ n5318;
  assign n5335 = n5334 ^ n5330;
  assign n5354 = n5353 ^ n5335;
  assign n5358 = n5357 ^ n5354;
  assign n5362 = n5361 ^ n5358;
  assign n5366 = n5365 ^ n5362;
  assign n5370 = n5369 ^ n5366;
  assign n5415 = n5369 ^ n5362;
  assign n5416 = n5366 & n5415;
  assign n5417 = n5416 ^ n5369;
  assign n5411 = n5361 ^ n5357;
  assign n5412 = ~n5358 & n5411;
  assign n5413 = n5412 ^ n5354;
  assign n5407 = n5352 ^ n5335;
  assign n5408 = ~n5353 & ~n5407;
  assign n5409 = n5408 ^ n5348;
  assign n5402 = n5330 ^ n5293;
  assign n5403 = n5333 ^ n5330;
  assign n5404 = n5402 & ~n5403;
  assign n5405 = n5404 ^ n5293;
  assign n5397 = n5347 ^ n5341;
  assign n5398 = ~n5342 & ~n5397;
  assign n5399 = n5398 ^ n5336;
  assign n5393 = x31 & n1661;
  assign n5394 = n5393 ^ n1664;
  assign n5395 = n5394 ^ n1878;
  assign n5389 = x26 & n2387;
  assign n5390 = n5389 ^ n2635;
  assign n5387 = x25 & n2631;
  assign n5388 = n5387 ^ n2632;
  assign n5391 = n5390 ^ n5388;
  assign n5386 = x24 & x63;
  assign n5392 = n5391 ^ n5386;
  assign n5396 = n5395 ^ n5392;
  assign n5400 = n5399 ^ n5396;
  assign n5382 = n5323 ^ n5318;
  assign n5383 = ~n5329 & n5382;
  assign n5384 = n5383 ^ n5318;
  assign n5378 = x28 & n2143;
  assign n5379 = n5378 ^ n2275;
  assign n5376 = x27 & n2272;
  assign n5377 = n5376 ^ n2484;
  assign n5380 = n5379 ^ n5377;
  assign n5373 = ~x30 & n1815;
  assign n5374 = n5373 ^ n2047;
  assign n5371 = ~x29 & n2044;
  assign n5372 = n5371 ^ n2162;
  assign n5375 = n5374 ^ n5372;
  assign n5381 = n5380 ^ n5375;
  assign n5385 = n5384 ^ n5381;
  assign n5401 = n5400 ^ n5385;
  assign n5406 = n5405 ^ n5401;
  assign n5410 = n5409 ^ n5406;
  assign n5414 = n5413 ^ n5410;
  assign n5418 = n5417 ^ n5414;
  assign n5458 = n5417 ^ n5410;
  assign n5459 = ~n5414 & ~n5458;
  assign n5460 = n5459 ^ n5417;
  assign n5454 = n5409 ^ n5405;
  assign n5455 = n5406 & n5454;
  assign n5456 = n5455 ^ n5401;
  assign n5450 = n5399 ^ n5385;
  assign n5451 = ~n5400 & ~n5450;
  assign n5452 = n5451 ^ n5396;
  assign n5446 = n5384 ^ n5380;
  assign n5447 = ~n5381 & ~n5446;
  assign n5448 = n5447 ^ n5375;
  assign n5440 = n5395 ^ n5386;
  assign n5441 = n5395 ^ n5391;
  assign n5442 = n5440 & ~n5441;
  assign n5443 = n5442 ^ n5386;
  assign n5436 = x27 & n2387;
  assign n5437 = n5436 ^ n2635;
  assign n5434 = x26 & n2631;
  assign n5435 = n5434 ^ n2632;
  assign n5438 = n5437 ^ n5435;
  assign n5430 = ~x31 & n1815;
  assign n5431 = n5430 ^ n2047;
  assign n5428 = ~x30 & n2044;
  assign n5429 = n5428 ^ n2162;
  assign n5432 = n5431 ^ n5429;
  assign n5427 = n1878 ^ n1664;
  assign n5433 = n5432 ^ n5427;
  assign n5439 = n5438 ^ n5433;
  assign n5444 = n5443 ^ n5439;
  assign n5422 = x29 & n2143;
  assign n5423 = n5422 ^ n2275;
  assign n5420 = x28 & n2272;
  assign n5421 = n5420 ^ n2484;
  assign n5424 = n5423 ^ n5421;
  assign n5419 = x25 & x63;
  assign n5425 = n5424 ^ n5419;
  assign n5426 = n5425 ^ n5375;
  assign n5445 = n5444 ^ n5426;
  assign n5449 = n5448 ^ n5445;
  assign n5453 = n5452 ^ n5449;
  assign n5457 = n5456 ^ n5453;
  assign n5461 = n5460 ^ n5457;
  assign n5499 = n5460 ^ n5453;
  assign n5500 = ~n5457 & n5499;
  assign n5501 = n5500 ^ n5460;
  assign n5495 = n5452 ^ n5448;
  assign n5496 = n5449 & n5495;
  assign n5497 = n5496 ^ n5445;
  assign n5491 = n5439 ^ n5426;
  assign n5492 = n5444 & ~n5491;
  assign n5493 = n5492 ^ n5426;
  assign n5486 = n5419 ^ n5375;
  assign n5487 = n5424 ^ n5375;
  assign n5488 = n5486 & ~n5487;
  assign n5489 = n5488 ^ n5419;
  assign n5481 = x31 & n2044;
  assign n5480 = n2047 ^ n1815;
  assign n5482 = n5481 ^ n5480;
  assign n5479 = n2162 ^ n2044;
  assign n5483 = n5482 ^ n5479;
  assign n5475 = n5438 ^ n5427;
  assign n5476 = n5438 ^ n5432;
  assign n5477 = ~n5475 & ~n5476;
  assign n5478 = n5477 ^ n5427;
  assign n5484 = n5483 ^ n5478;
  assign n5471 = x28 & n2387;
  assign n5472 = n5471 ^ n2635;
  assign n5469 = x27 & n2631;
  assign n5470 = n5469 ^ n2632;
  assign n5473 = n5472 ^ n5470;
  assign n5465 = x30 & n2143;
  assign n5466 = n5465 ^ n2275;
  assign n5463 = x29 & n2272;
  assign n5464 = n5463 ^ n2484;
  assign n5467 = n5466 ^ n5464;
  assign n5462 = x26 & x63;
  assign n5468 = n5467 ^ n5462;
  assign n5474 = n5473 ^ n5468;
  assign n5485 = n5484 ^ n5474;
  assign n5490 = n5489 ^ n5485;
  assign n5494 = n5493 ^ n5490;
  assign n5498 = n5497 ^ n5494;
  assign n5502 = n5501 ^ n5498;
  assign n5532 = n5501 ^ n5494;
  assign n5533 = n5498 & n5532;
  assign n5534 = n5533 ^ n5501;
  assign n5528 = n5493 ^ n5485;
  assign n5529 = n5490 & ~n5528;
  assign n5530 = n5529 ^ n5489;
  assign n5523 = n5483 ^ n5474;
  assign n5524 = n5478 ^ n5474;
  assign n5525 = ~n5523 & n5524;
  assign n5526 = n5525 ^ n5483;
  assign n5518 = n5473 ^ n5467;
  assign n5519 = n5468 & ~n5518;
  assign n5520 = n5519 ^ n5462;
  assign n5514 = x29 & n2387;
  assign n5515 = n5514 ^ n2635;
  assign n5512 = x28 & n2631;
  assign n5513 = n5512 ^ n2632;
  assign n5516 = n5515 ^ n5513;
  assign n5517 = n5516 ^ n5483;
  assign n5521 = n5520 ^ n5517;
  assign n5507 = x31 & n2143;
  assign n5508 = n5507 ^ n2275;
  assign n5505 = x30 & n2272;
  assign n5506 = n5505 ^ n2484;
  assign n5509 = n5508 ^ n5506;
  assign n5504 = n5480 ^ n5479;
  assign n5510 = n5509 ^ n5504;
  assign n5503 = x27 & x63;
  assign n5511 = n5510 ^ n5503;
  assign n5522 = n5521 ^ n5511;
  assign n5527 = n5526 ^ n5522;
  assign n5531 = n5530 ^ n5527;
  assign n5535 = n5534 ^ n5531;
  assign n5559 = n5534 ^ n5527;
  assign n5560 = ~n5531 & n5559;
  assign n5561 = n5560 ^ n5534;
  assign n5555 = n5526 ^ n5521;
  assign n5556 = ~n5522 & n5555;
  assign n5557 = n5556 ^ n5511;
  assign n5551 = n5520 ^ n5516;
  assign n5552 = n5517 & ~n5551;
  assign n5553 = n5552 ^ n5483;
  assign n5547 = n5504 ^ n5503;
  assign n5548 = n5510 & ~n5547;
  assign n5549 = n5548 ^ n5503;
  assign n5543 = x31 & n2272;
  assign n5544 = n5543 ^ n2275;
  assign n5545 = n5544 ^ n2484;
  assign n5539 = x30 & n2387;
  assign n5540 = n5539 ^ n2635;
  assign n5537 = x29 & n2631;
  assign n5538 = n5537 ^ n2632;
  assign n5541 = n5540 ^ n5538;
  assign n5536 = x28 & x63;
  assign n5542 = n5541 ^ n5536;
  assign n5546 = n5545 ^ n5542;
  assign n5550 = n5549 ^ n5546;
  assign n5554 = n5553 ^ n5550;
  assign n5558 = n5557 ^ n5554;
  assign n5562 = n5561 ^ n5558;
  assign n5582 = n5561 ^ n5554;
  assign n5583 = ~n5558 & ~n5582;
  assign n5584 = n5583 ^ n5561;
  assign n5578 = n5553 ^ n5549;
  assign n5579 = ~n5550 & ~n5578;
  assign n5580 = n5579 ^ n5546;
  assign n5573 = n5545 ^ n5536;
  assign n5574 = n5545 ^ n5541;
  assign n5575 = ~n5573 & n5574;
  assign n5576 = n5575 ^ n5536;
  assign n5567 = x31 & n2387;
  assign n5568 = n5567 ^ n2635;
  assign n5565 = x30 & n2631;
  assign n5566 = n5565 ^ n2632;
  assign n5569 = n5568 ^ n5566;
  assign n5564 = n2484 ^ n2275;
  assign n5570 = n5569 ^ n5564;
  assign n5563 = x29 & x63;
  assign n5571 = n5570 ^ n5563;
  assign n5572 = n5571 ^ n5545;
  assign n5577 = n5576 ^ n5572;
  assign n5581 = n5580 ^ n5577;
  assign n5585 = n5584 ^ n5581;
  assign n5599 = n5584 ^ n5577;
  assign n5600 = ~n5581 & ~n5599;
  assign n5601 = n5600 ^ n5584;
  assign n5595 = n5576 ^ n5571;
  assign n5596 = ~n5572 & n5595;
  assign n5597 = n5596 ^ n5545;
  assign n5591 = n5564 ^ n5563;
  assign n5592 = n5570 & ~n5591;
  assign n5593 = n5592 ^ n5563;
  assign n5587 = x31 & n2631;
  assign n5588 = n5587 ^ n2635;
  assign n5589 = n5588 ^ n2632;
  assign n5586 = x30 & x63;
  assign n5590 = n5589 ^ n5586;
  assign n5594 = n5593 ^ n5590;
  assign n5598 = n5597 ^ n5594;
  assign n5602 = n5601 ^ n5598;
  assign n5611 = n5601 ^ n5594;
  assign n5612 = n5598 & ~n5611;
  assign n5613 = n5612 ^ n5601;
  assign n5607 = n5593 ^ n5589;
  assign n5608 = ~n5590 & ~n5607;
  assign n5609 = n5608 ^ n5586;
  assign n5603 = n2631 ^ n2387;
  assign n5604 = n5603 ^ x31;
  assign n5605 = x63 & n5604;
  assign n5606 = n5605 ^ n5586;
  assign n5610 = n5609 ^ n5606;
  assign n5614 = n5613 ^ n5610;
  assign y0 = n65;
  assign y1 = n73;
  assign y2 = n82;
  assign y3 = n104;
  assign y4 = n124;
  assign y5 = n156;
  assign y6 = n186;
  assign y7 = n227;
  assign y8 = n269;
  assign y9 = n321;
  assign y10 = n372;
  assign y11 = n434;
  assign y12 = n494;
  assign y13 = n566;
  assign y14 = n636;
  assign y15 = n718;
  assign y16 = n801;
  assign y17 = n893;
  assign y18 = n984;
  assign y19 = n1086;
  assign y20 = n1190;
  assign y21 = n1303;
  assign y22 = n1415;
  assign y23 = n1538;
  assign y24 = n1659;
  assign y25 = n1794;
  assign y26 = n1928;
  assign y27 = n2072;
  assign y28 = n2215;
  assign y29 = n2369;
  assign y30 = n2521;
  assign y31 = n2686;
  assign y32 = n2843;
  assign y33 = n3003;
  assign y34 = n3161;
  assign y35 = n3317;
  assign y36 = n3471;
  assign y37 = n3619;
  assign y38 = ~n3758;
  assign y39 = n3893;
  assign y40 = ~n4023;
  assign y41 = n4151;
  assign y42 = n4272;
  assign y43 = n4390;
  assign y44 = ~n4498;
  assign y45 = n4605;
  assign y46 = n4707;
  assign y47 = ~n4802;
  assign y48 = ~n4890;
  assign y49 = n4972;
  assign y50 = ~n5054;
  assign y51 = n5126;
  assign y52 = ~n5194;
  assign y53 = ~n5257;
  assign y54 = ~n5317;
  assign y55 = ~n5370;
  assign y56 = n5418;
  assign y57 = n5461;
  assign y58 = ~n5502;
  assign y59 = n5535;
  assign y60 = n5562;
  assign y61 = n5585;
  assign y62 = ~n5602;
  assign y63 = n5614;
endmodule
